Offentlig tandvård
Du kan använda de kommunala tandläkartjänsterna om du har hemkommun i Esbo.
I nödfall kan du använda kommunala tjänster även om Esbo inte är din hemkommun.
Du kan boka tid hos en tandläkare på Esbo tandklinikers gemensamma nummer.
Tandklinikernas tidsbeställning
Tfn (09) 816 30300
Du kan ringa numret på vardagar.
Om du behöver besöka tandläkaren snabbt, ta kontakt med social- och hälsostationen i Kilo.
Social- och hälsostationen i Kilo
Trillagatan 5
Tfn (09) 816 35900
Tidsbeställning på vardagar.
Om du behöver akut tandläkarvård kvällstid eller under veckoslut, kan du kontakta Haartmanska sjukhuset i Helsingfors.
Jourmottagningen vid Haartmanska sjukhuset har öppet vardagar kl. 14–21 och lö-sö kl. 8–21.
Tfn (09) 310 49999.
linkkiEsbo stad:
Mun- och tandhälsovårdenfinska _ svenska _ engelska
Privat tandvård
I Esbo finns också privata tandläkare.
Du kan gå till en privat tandläkare även om du inte har rätt att använda den offentliga hälsovårdens tjänster.
Privat tandvård är dyrare än offentlig tandvård.
Läs mer: Tandvård.
Sök tandläkarefinska
Mental hälsa
Om du behöver hjälp eller stöd i mental- och/eller missbruksfrågor, boka tid till en psykiatriskötare.
Du kan boka tid vardagar kl. 8–16 på numret 09 816 31300.
linkkiEsbo stad:
Information om mentalvårdstjänsternafinska _ svenska _ engelska
Psykiatriskötarna har mottagning på hälsostationerna.
Mottagning för unga finns vid Nupoli.
Du kan även besöka mottagningen vid Kliniken för mental- och missbruksvård på servicetorget i Iso Omena utan tidsbokning måndag till fredag kl. 8.30–10.30 och dessutom måndag till torsdag kl. 13–14.30.
Adress: Finnviksvägen 1, Köpcentret Iso Omena.
Om du behöver krishjälp snabbt, ta kontakt med Esbo social- och krisjour (Espoon sosiaali- ja kriisipäivystys).
Social- och krisjouren
Åbovägen 150
Tfn (09) 816 42439
Öppet alla dagar dygnet runt.
linkkiEsbo stad:
Social- och krisjourenfinska _ svenska _ engelska
Läs mer: Mental hälsa.
linkkiFöreningen för mental hälsa i Finland:
Krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Information om mentalvårdstjänsternafinska _ svenska _ engelska
Sexuell hälsa
Vid hälsostationernas preventivrådgivning (ehkäisyneuvola) får du hjälp med graviditetsprevention och familjeplanering.
Ungdomar kan diskutera frågor kring sexuell hälsa med hälsovårdaren vid sin egen skola.
linkkiEsbo stad:
Preventivrådgivningsbyråerfinska _ svenska _ engelska
Om du behöver en gynekologisk undersökning, ta kontakt med hälsostationen.
Du kan också boka tid vid hälsostationen om du behöver ett recept för preventivmedel eller om du överväger abort.
Hälsostationernas kontaktuppgifter finns på Esbo stads webbplats.
linkkiEsbo stad:
Hälsostationernafinska _ svenska _ engelska
Könssjukdomar behandlas i huvudstadsregionen på polikliniken för könssjukdomar i Helsingfors.
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Polikliniken för könssjukdomarfinska _ svenska _ engelska
När du väntar barn
Kontakta rådgivningen (neuvola) när du upptäcker att du är gravid.
Vid rådgivningen följs moderns, fostrets och hela familjens hälsotillstånd under graviditeten.
I Esbo finns flera rådgivningsbyråer på olika håll i staden.
Du kan boka tid vid alla rådgivningsbyråer på samma nummer.
Rådgivning och tidsbeställning vid rådgivningsbyrån
Tfn (09) 816 22800
Läs mer: När du väntar barn.
linkkiEsbo stad:
Rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
Förlossning
I Esbo finns Jorv sjukhus där man kan föda barn.
Om du vill kan du även föda barnet på något annat sjukhus inom samkommunen Helsingfors och Nylands sjukvårdsdistrikt (HNS).
Mer information hittar du på HNS webbplats.
Läs mer: Förlossning.
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Förlossningfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Handikappade personer
Esbo stad ordnar olika tjänster för handikappade, till exempel dagverksamhet och färdtjänster.
Personer som har sin hemkommun i Esbo har rätt till dessa tjänster.
Du kan ansöka om tjänster och stödfunktioner hos stadens socialarbetare.
Mer information om tjänsterna för handikappade hittar du på Esbo stads handikappservice.
Esbo handikappservice
Kamrersvägen 2 A, vån. 4
Tfn (09) 816 45285
Läs mer: Handikappade personer
linkkiEsbo stad:
Kontaktuppgifter till socialarbetarefinska _ svenska _ engelska
linkkiEsbo stad:
Stödtjänster för handikappadefinska _ svenska _ engelska
Ett handikappat barn
Om du har ett handikappat barn kan du kontakta socialarbetaren vid handikappservicen för ditt eget område vammaispalvelut(at)espoo.fi.
Frågor som rör skolgången för ett handikappat barn kan du ställa till skolväsendet (opetustoimi) samt till servicehandledaren för skolelever (koululaisten palveluohjaaja).
Läs mer: Ett handikappat barn
linkkiEsbo stad:
Kontaktuppgifter till utbildningsväsendetfinska _ engelska
Hälsovårdstjänsterna i Esbo
Tandvården
Mental hälsa
Sexuell hälsa
När du väntar barn
Handikappade personer
Ring nödnumret 112 om det är fråga om en brådskande nödsituation.
Ring nödnumret till exempel vid en allvarlig olycka eller när någon drabbas av en sjukdomsattack.
Ring inte nödnumret om det inte är en nödsituation.
Om du har din hemkommun i Esbo kan du utnyttja de offentliga hälsovårdstjänsterna.
Offentliga hälsovårdstjänster tillhandahålls vid hälsostationer, tandkliniker, rådgivningsbyråer och sjukhus.
Om du inte har rätt till de offentliga hälsovårdstjänsterna, kan du söka hjälp på en privat läkarstation.
På en privat läkarstation måste du betala samtliga kostnader själv.
Läs mer: Hälsa.
Hälsovårdstjänsterna i Esbo
Offentliga hälsovårdstjänster tillhandahålls av hälsostationerna (terveysasema).
Hälsostationerna har öppet vardagar klockan 8–16.
På hälsostationerna finns vanligtvis läkarens, sjukskötarens och hälsovårdarens mottagningar.
Du kan boka tid på hälsostationen per telefon.
På Esbo stads webbplats finns kontaktuppgifterna och telefonnumren till hälsostationerna.
När du ringer hälsostationen, besvaras ditt samtal inte nödvändigtvis omedelbart.
Ditt nummer sparas dock i en automat och du blir uppringd.
Kom i tid till mottagningen.
Om du inte kan komma till mottagningen, kom ihåg att avboka din tid senast föregående vardag före klockan 14.
Om du behöver första hjälpen snabbt, kan du komma till hälsostationen utan tidsbeställning.
linkkiEsbo stad:
Hälsostationernafinska _ svenska _ engelska
linkkiEsbo stad:
Hälsovårdscentralsavgifterfinska _ svenska
Privata hälsovårdstjänster
Vem som helst kan gå till en privat hälsostation.
Också de personer som inte har rätt till den offentliga hälsovården i Finland kan besöka privata hälsostationer.
På en privat hälsostation måste kunden själv betala samtliga kostnader.
I Esbo finns flera privata läkarstationer.
Kontaktuppgifter till privata läkare hittar du till exempel på Internet.
linkkietsilaakari.fi:
Privata hälsovårdstjänsterfinska
Privat läkarstationfinska _ svenska _ engelska
Privat läkarstationfinska _ svenska _ engelska
Läkemedel
Information om köp av läkemedel hittar du på InfoFinlands sida Läkemedel.
Hälsovård för papperslösa
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärhälsovård.
Tjänsterna vid Global Clinic är avgiftsfria för kunderna.
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter.
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
Telefonnumret till Global Clinic i Helsingfors är 044 977 4547.
Samtalet besvaras av en sjukskötare eller en läkare.
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Läs mer: Hälsovårdstjänster i Finland
Kvällstid och under veckoslut har hälsostationen stängt.
Då vårdas akuta sjukfall och olycksfall på jourmottagningen (päivystys).
Den närmaste jourmottagningen för vuxna finns vid Jorv sjukhus.
Ring den kostnadsfria Jourhjälpen på tfn 116 117 innan du kommer till jourmottagningen.
Jourmottagningen vid Jorv sjukhus
Åbovägen 150
Tfn (09) 4711
Jourmottagningar för barn under 16 år finns i Jorv och på Barnkliniken i Helsingfors.
Du behöver inte boka tid på jourmottagningen.
linkkiEsbo stad:
Jourmottagningarfinska _ svenska _ engelska
Läs mer: Hälsovårdstjänster i Finland
Barns hälsa
I hälsovården av 1–6-åriga barn får man hjälp av rådgivningsbyråns (neuvola) hälsovårdare och läkare.
Dem kan du fråga om råd och få hjälp med fostran av barn.
På rådgivningsbyrån följs att barnet är friskt och växer som det ska.
I Esbo finns flera rådgivningsbyråer på olika håll i staden.
Rådgivningsbyråernas kontaktuppgifter finns på Esbo stads webbplats.
Du kan boka tid vid alla rådgivningsbyråer på samma nummer.
Om ett barn blir sjukt och behöver snabbt vård, ta kontakt med hälsostationen (terveysasema).
Skolhälsovårdaren har hand om skolbarns hälsa.
Under kvällar och veckoslut finns jourmottagningen för barn under 16 år vid Jorv sjukhus och på Barnkliniken i Helsingfors.
Du kan också ta ditt barn till en privat läkarstation.
Läs mer: Barns hälsa.
linkkiEsbo stad:
Barnrådgivningsbyråernas tjänsterfinska _ svenska _ engelska
linkkiEsbo stad:
Rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
linkkiEsbo stad:
Hälsostationernafinska _ svenska _ engelska
linkkiEsbo stad:
Information om hälsovården för skolbarnfinska _ svenska _ engelska
linkkiEsbo stad:
Jourmottagningarfinska _ svenska _ engelska
Tandvården
Offentlig tandvård
Du kan använda de kommunala tandläkartjänsterna om du har hemkommun i Esbo.
I nödfall kan du använda kommunala tjänster även om Esbo inte är din hemkommun.
Du kan boka tid hos en tandläkare på Esbo tandklinikers gemensamma nummer.
Tandklinikernas tidsbeställning
Tfn (09) 816 30300
Du kan ringa numret på vardagar.
Om du behöver besöka tandläkaren snabbt, ta kontakt med social- och hälsostationen i Kilo.
Social- och hälsostationen i Kilo
Trillagatan 5
Tfn (09) 816 35900
Tidsbeställning på vardagar.
Om du behöver akut tandläkarvård kvällstid eller under veckoslut, kan du kontakta Haartmanska sjukhuset i Helsingfors.
Jourmottagningen vid Haartmanska sjukhuset har öppet vardagar kl. 14–21 och lö-sö kl. 8–21.
Tfn (09) 310 49999.
linkkiEsbo stad:
Mun- och tandhälsovårdenfinska _ svenska _ engelska
Privat tandvård
I Esbo finns också privata tandläkare.
Du kan gå till en privat tandläkare även om du inte har rätt att använda den offentliga hälsovårdens tjänster.
Privat tandvård är dyrare än offentlig tandvård.
Läs mer: Tandvård.
Sök tandläkarefinska
Mental hälsa
Om du behöver hjälp eller stöd i mental- och/eller missbruksfrågor, boka tid till en psykiatriskötare.
Du kan boka tid vardagar kl. 8–16 på numret 09 816 31300.
linkkiEsbo stad:
Information om mentalvårdstjänsternafinska _ svenska _ engelska
Psykiatriskötarna har mottagning på hälsostationerna.
Mottagning för unga finns vid Nupoli.
Du kan även besöka mottagningen vid Kliniken för mental- och missbruksvård på servicetorget i Iso Omena utan tidsbokning måndag till fredag kl. 8.30–10.30 och dessutom måndag till torsdag kl. 13–14.30.
Adress: Finnviksvägen 1, Köpcentret Iso Omena.
Om du behöver krishjälp snabbt, ta kontakt med Esbo social- och krisjour (Espoon sosiaali- ja kriisipäivystys).
Social- och krisjouren
Åbovägen 150
Tfn (09) 816 42439
Öppet alla dagar dygnet runt.
linkkiEsbo stad:
Social- och krisjourenfinska _ svenska _ engelska
Läs mer: Mental hälsa.
linkkiFöreningen för mental hälsa i Finland:
Krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Information om mentalvårdstjänsternafinska _ svenska _ engelska
Sexuell hälsa
Vid hälsostationernas preventivrådgivning (ehkäisyneuvola) får du hjälp med graviditetsprevention och familjeplanering.
Ungdomar kan diskutera frågor kring sexuell hälsa med hälsovårdaren vid sin egen skola.
linkkiEsbo stad:
Preventivrådgivningsbyråerfinska _ svenska _ engelska
Om du behöver en gynekologisk undersökning, ta kontakt med hälsostationen.
Du kan också boka tid vid hälsostationen om du behöver ett recept för preventivmedel eller om du överväger abort.
Hälsostationernas kontaktuppgifter finns på Esbo stads webbplats.
linkkiEsbo stad:
Hälsostationernafinska _ svenska _ engelska
Könssjukdomar behandlas i huvudstadsregionen på polikliniken för könssjukdomar i Helsingfors.
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Polikliniken för könssjukdomarfinska _ svenska _ engelska
När du väntar barn
Kontakta rådgivningen (neuvola) när du upptäcker att du är gravid.
Vid rådgivningen följs moderns, fostrets och hela familjens hälsotillstånd under graviditeten.
I Esbo finns flera rådgivningsbyråer på olika håll i staden.
Du kan boka tid vid alla rådgivningsbyråer på samma nummer.
Rådgivning och tidsbeställning vid rådgivningsbyrån
Tfn (09) 816 22800
Läs mer: När du väntar barn.
linkkiEsbo stad:
Rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
Förlossning
I Esbo finns Jorv sjukhus där man kan föda barn.
Om du vill kan du även föda barnet på något annat sjukhus inom samkommunen Helsingfors och Nylands sjukvårdsdistrikt (HNS).
Mer information hittar du på HNS webbplats.
Läs mer: Förlossning.
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Förlossningfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Handikappade personer
Esbo stad ordnar olika tjänster för handikappade, till exempel dagverksamhet och färdtjänster.
Personer som har sin hemkommun i Esbo har rätt till dessa tjänster.
Du kan ansöka om tjänster och stödfunktioner hos stadens socialarbetare.
Mer information om tjänsterna för handikappade hittar du på Esbo stads handikappservice.
Esbo handikappservice
Kamrersvägen 2 A, vån. 4
Tfn (09) 816 45285
Handikappade personerlinkkiEsbo stad:
linkkiEsbo stad:
Stödtjänster för handikappadefinska _ svenska _ engelska
Ett handikappat barn
Om du har ett handikappat barn kan du kontakta socialarbetaren vid handikappservicen för ditt eget område vammaispalvelut(at)espoo.fi.
Frågor som rör skolgången för ett handikappat barn kan du ställa till skolväsendet (opetustoimi) samt till servicehandledaren för skolelever (koululaisten palveluohjaaja).
Läs mer: Ett handikappat barn
linkkiEsbo stad:
Kontaktuppgifter till utbildningsväsendetfinska _ engelska
Hälsovårdstjänsterna i Esbo
Tandvården
Mental hälsa
Sexuell hälsa
När du väntar barn
Handikappade personer
Ring nödnumret 112 om det är fråga om en brådskande nödsituation.
Ring nödnumret till exempel vid en allvarlig olycka eller när någon drabbas av en sjukdomsattack.
Ring inte nödnumret om det inte är en nödsituation.
Om du har din hemkommun i Esbo kan du utnyttja de offentliga hälsovårdstjänsterna.
Offentliga hälsovårdstjänster tillhandahålls vid hälsostationer, tandkliniker, rådgivningsbyråer och sjukhus.
Om du inte har rätt till de offentliga hälsovårdstjänsterna, kan du söka hjälp på en privat läkarstation.
På en privat läkarstation måste du betala samtliga kostnader själv.
Läs mer: Hälsa.
Hälsovårdstjänsterna i Esbo
Offentliga hälsovårdstjänster tillhandahålls av hälsostationerna (terveysasema).
Hälsostationerna har öppet vardagar klockan 8–16.
På hälsostationerna finns vanligtvis läkarens, sjukskötarens och hälsovårdarens mottagningar.
Du kan boka tid på hälsostationen per telefon.
På Esbo stads webbplats finns kontaktuppgifterna och telefonnumren till hälsostationerna.
När du ringer hälsostationen, besvaras ditt samtal inte nödvändigtvis omedelbart.
Ditt nummer sparas dock i en automat och du blir uppringd.
Kom i tid till mottagningen.
Om du inte kan komma till mottagningen, kom ihåg att avboka din tid senast föregående vardag före klockan 14.
Om du behöver första hjälpen snabbt, kan du komma till hälsostationen utan tidsbeställning.
linkkiEsbo stad:
Hälsostationernafinska _ svenska _ engelska
linkkiEsbo stad:
Hälsovårdscentralsavgifterfinska _ svenska
Privata hälsovårdstjänster
Vem som helst kan gå till en privat hälsostation.
Också de personer som inte har rätt till den offentliga hälsovården i Finland kan besöka privata hälsostationer.
På en privat hälsostation måste kunden själv betala samtliga kostnader.
I Esbo finns flera privata läkarstationer.
Kontaktuppgifter till privata läkare hittar du till exempel på Internet.
linkkietsilaakari.fi:
Privata hälsovårdstjänsterfinska
Privat läkarstationfinska _ svenska _ engelska
Privat läkarstationfinska _ svenska _ engelska
Läkemedel
Information om köp av läkemedel hittar du på InfoFinlands sida Läkemedel.
Hälsovård för papperslösa
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärhälsovård.
Tjänsterna vid Global Clinic är avgiftsfria för kunderna.
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter.
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
Telefonnumret till Global Clinic i Helsingfors är 044 977 4547.
Samtalet besvaras av en sjukskötare eller en läkare.
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Läs mer: Hälsovårdstjänster i Finland
Kvällstid och under veckoslut har hälsostationen stängt.
Då vårdas akuta sjukfall och olycksfall på jourmottagningen (päivystys).
Den närmaste jourmottagningen för vuxna finns vid Jorv sjukhus.
Ring den kostnadsfria Jourhjälpen på tfn 116 117 innan du kommer till jourmottagningen.
Jourmottagningen vid Jorv sjukhus
Åbovägen 150
Tfn (09) 4711
Jourmottagningar för barn under 16 år finns i Jorv och på Barnkliniken i Helsingfors.
Du behöver inte boka tid på jourmottagningen.
linkkiEsbo stad:
Jourmottagningarfinska _ svenska _ engelska
Läs mer: Hälsovårdstjänster i Finland
Barns hälsa
I hälsovården av 1–6-åriga barn får man hjälp av rådgivningsbyråns (neuvola) hälsovårdare och läkare.
Dem kan du fråga om råd och få hjälp med fostran av barn.
På rådgivningsbyrån följs att barnet är friskt och växer som det ska.
I Esbo finns flera rådgivningsbyråer på olika håll i staden.
Rådgivningsbyråernas kontaktuppgifter finns på Esbo stads webbplats.
Du kan boka tid vid alla rådgivningsbyråer på samma nummer.
Om ett barn blir sjukt och behöver snabbt vård, ta kontakt med hälsostationen (terveysasema).
Skolhälsovårdaren har hand om skolbarns hälsa.
Under kvällar och veckoslut finns jourmottagningen för barn under 16 år vid Jorv sjukhus och på Barnkliniken i Helsingfors.
Du kan också ta ditt barn till en privat läkarstation.
Läs mer: Barns hälsa.
linkkiEsbo stad:
Barnrådgivningsbyråernas tjänsterfinska _ svenska _ engelska
linkkiEsbo stad:
Rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
linkkiEsbo stad:
Hälsostationernafinska _ svenska _ engelska
linkkiEsbo stad:
Information om hälsovården för skolbarnfinska _ svenska _ engelska
linkkiEsbo stad:
Jourmottagningarfinska _ svenska _ engelska
Tandvården
Offentlig tandvård
Du kan använda de kommunala tandläkartjänsterna om du har hemkommun i Esbo.
I nödfall kan du använda kommunala tjänster även om Esbo inte är din hemkommun.
Du kan boka tid hos en tandläkare på Esbo tandklinikers gemensamma nummer.
Tandklinikernas tidsbeställning
Tfn (09) 816 30300
Du kan ringa numret på vardagar.
Om du behöver besöka tandläkaren snabbt, ta kontakt med social- och hälsostationen i Kilo.
Social- och hälsostationen i Kilo
Trillagatan 5
Tfn (09) 816 35900
Tidsbeställning på vardagar.
Om du behöver akut tandläkarvård kvällstid eller under veckoslut, kan du kontakta Haartmanska sjukhuset i Helsingfors.
Jourmottagningen vid Haartmanska sjukhuset har öppet vardagar kl. 14–21 och lö-sö kl. 8–21.
Tfn (09) 310 49999.
linkkiEsbo stad:
Mun- och tandhälsovårdenfinska _ svenska _ engelska
Privat tandvård
I Esbo finns också privata tandläkare.
Du kan gå till en privat tandläkare även om du inte har rätt att använda den offentliga hälsovårdens tjänster.
Privat tandvård är dyrare än offentlig tandvård.
Läs mer: Tandvård.
Sök tandläkarefinska
Mental hälsa
Om du behöver hjälp eller stöd i mental- och/eller missbruksfrågor, boka tid till en psykiatriskötare.
Du kan boka tid vardagar kl. 8–16 på numret 09 816 31300.
linkkiEsbo stad:
Information om mentalvårdstjänsternafinska _ svenska _ engelska
Psykiatriskötarna har mottagning på hälsostationerna.
Mottagning för unga finns vid Nupoli.
Du kan även besöka mottagningen vid Kliniken för mental- och missbruksvård på servicetorget i Iso Omena utan tidsbokning måndag till fredag kl. 8.30–10.30 och dessutom måndag till torsdag kl. 13–14.30.
Adress: Finnviksvägen 1, Köpcentret Iso Omena.
Om du behöver krishjälp snabbt, ta kontakt med Esbo social- och krisjour (Espoon sosiaali- ja kriisipäivystys).
Social- och krisjouren
Åbovägen 150
Tfn (09) 816 42439
Öppet alla dagar dygnet runt.
linkkiEsbo stad:
Social- och krisjourenfinska _ svenska _ engelska
Läs mer: Mental hälsa.
linkkiFöreningen för mental hälsa i Finland:
Krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Information om mentalvårdstjänsternafinska _ svenska _ engelska
Sexuell hälsa
Vid hälsostationernas preventivrådgivning (ehkäisyneuvola) får du hjälp med graviditetsprevention och familjeplanering.
Ungdomar kan diskutera frågor kring sexuell hälsa med hälsovårdaren vid sin egen skola.
linkkiEsbo stad:
Preventivrådgivningsbyråerfinska _ svenska _ engelska
Om du behöver en gynekologisk undersökning, ta kontakt med hälsostationen.
Du kan också boka tid vid hälsostationen om du behöver ett recept för preventivmedel eller om du överväger abort.
Hälsostationernas kontaktuppgifter finns på Esbo stads webbplats.
linkkiEsbo stad:
Hälsostationernafinska _ svenska _ engelska
Könssjukdomar behandlas i huvudstadsregionen på polikliniken för könssjukdomar i Helsingfors.
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Polikliniken för könssjukdomarfinska _ svenska _ engelska
Läs mer: Sexualhälsa
När du väntar barn
Kontakta rådgivningen (neuvola) när du upptäcker att du är gravid.
Vid rådgivningen följs moderns, fostrets och hela familjens hälsotillstånd under graviditeten.
I Esbo finns flera rådgivningsbyråer på olika håll i staden.
Du kan boka tid vid alla rådgivningsbyråer på samma nummer.
Rådgivning och tidsbeställning vid rådgivningsbyrån
Tfn (09) 816 22800
Läs mer: Graviditet och förlossning.
linkkiEsbo stad:
Rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
Förlossning
I Esbo finns Jorv sjukhus där man kan föda barn.
Om du vill kan du även föda barnet på något annat sjukhus inom samkommunen Helsingfors och Nylands sjukvårdsdistrikt (HNS).
Mer information hittar du på HNS webbplats.
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Förlossningfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Handikappade personer
Esbo stad ordnar olika tjänster för handikappade, till exempel dagverksamhet och färdtjänster.
Personer som har sin hemkommun i Esbo har rätt till dessa tjänster.
Du kan ansöka om tjänster och stödfunktioner hos stadens socialarbetare.
Mer information om tjänsterna för handikappade hittar du på Esbo stads handikappservice.
Esbo handikappservice
Kamrersvägen 2 A, vån. 4
Tfn (09) 816 45285
Läs mer: Handikappade personer
linkkiEsbo stad:
Stödtjänster för handikappadefinska _ svenska _ engelska
Ett handikappat barn
Om du har ett handikappat barn kan du kontakta socialarbetaren vid handikappservicen för ditt eget område vammaispalvelut(at)espoo.fi.
Frågor som rör skolgången för ett handikappat barn kan du ställa till skolväsendet (opetustoimi) samt till servicehandledaren för skolelever (koululaisten palveluohjaaja).
Läs mer: Ett handikappat barn
linkkiEsbo stad:
Kontaktuppgifter till utbildningsväsendetfinska _ engelska
Detta innehåll finns inte på det språk som du har valt.
Välj något annat språk.
Finska
Detta innehåll finns inte på det språk som du har valt.
Välj något annat språk.
Finska
Detta innehåll finns inte på det språk som du har valt.
Välj något annat språk.
Finska
Dagvård
Förskoleundervisning
Grundläggande utbildning
Hemspråksundervisning för invandrare
Yrkesutbildning
Gymnasium
Stöd och handledning för unga
Högskoleutbildning
Andra studiemöjligheter
Dagvård
I Esbo finns både kommunala och privata daghem.
I Esbo finns dessutom familjedagvårdare.
Dagvård fås på finska och på svenska.
Ansök om dagvårdsplats minst fyra månader innan barnet ska börja i dagvården.
Om du till exempel oväntat får arbete eller en studieplats kan du ansöka om vårdplats senare.
När du ansöker om vårdplats ska du fylla i en ansökningsblankett.
Du kan också söka dagvårdsplats via Internet.
Familjer som bor i Esbo kan också söka dagvårdsplats till sitt barn i Helsingfors, Vanda eller Grankulla.
Du ska ändå lämna in din ansökan i Esbo.
Mer information får du via tjänsten Helsingforsregionen.fi.
Läs mer: Dagvård.
linkkiEsbo stad:
Dagvårdfinska _ svenska _ engelska
linkkiEsbo stad:
Ansökan om dagvårdsplatsfinska
linkkiEsbo stad:
Servicepunktfinska _ svenska _ engelska
linkkiEsbo stad:
Dagvårdens samanvändningsområdefinska _ svenska _ engelska
Förskoleundervisning
I Esbo anordnas förskoleundervisningen (esiopetus) i daghemmen.
Förskoleundervisning ges på finska och på svenska.
Till förskoleundervisningen anmäler man sig via Esbo stads webbplats.
Förskoleundervisningen börjar i augusti.
Ansökningstiden är vanligtvis i januari.
I frågor kring barndagvård och förskoleundervisning kan du också kontakta daghemsföreståndarna eller stadens chef för småbarnsfostran (varhaiskasvatuspäällikkö).
Kontaktuppgifterna finns på stadens webbplats.
Läs mer: Förskoleundervisning.
linkkiEsbo stad:
Förskoleundervisningfinska _ svenska _ engelska
linkkiEsbo stad:
Ansökan till förskoleundervisningfinska _ svenska _ engelska
Grundläggande utbildning
