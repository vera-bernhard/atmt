��&      ]�(�numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i4�����R�(K�<�NNNJ����J����K t�b�CT   �       �  �      (  G   �     ~  �      �  �  �  �            �t�bhhK ��h��R�(KK!��h�C�      �   A      8      �   `     �   �     ,   \   Q   B         �      #  �         !     �   8   �  	         �t�bhhK ��h��R�(KK;��h�C�          �  D     �      �           J  �   s   �  �     O           X     �                 t   �   _   a     �   X         #   6           �    y         *   �      �     n   �         �t�bhhK ��h��R�(KK��h�C`�	  c  ]      �      
   �  "           K  
      	   p     6         4   	      �t�bhhK ��h��R�(KK��h�C`   f   �
  p   _  9      d   "     ,      W   "   �           f      d           �t�bhhK ��h��R�(KK��h�CP      "      e            "             M   �         s           �t�bhhK ��h��R�(KK$��h�C�   +               �      #   �     �     F             T     u     g	        �              >  �   C   �         �t�bhhK ��h��R�(KK��h�CH         �  [              D           y     �        �t�bhhK ��h��R�(KK��h�CD   I     �         �         �  �  �         �        �t�bhhK ��h��R�(KK��h�Cd    �  �   �     �        ?     t        1   �   @  �   �  +   
   J   .   �        �t�bhhK ��h��R�(KK��h�C4      �              0   c  #   v         �t�bhhK ��h��R�(KKB��h�B     -            |   .         �      *   �               �   v   5     �         �   !   �   �  �  ;      5   �      q   E  �                     %  ;              X      l            �  �         \   Q   �             �t�bhhK ��h��R�(KK��h�C@   �           �     U       �   /      �         �t�bhhK ��h��R�(KK��h�Ct      �      �  #   ?          �         6      +            �   b        ^   |   \  k        �t�bhhK ��h��R�(KK&��h�C�   `   5  �  �     !   g
  V      l        	   >   A   t  �            L      �  �     2   A   B   �   3         �   �   4   	      �t�bhhK ��h��R�(KK��h�C|      L            L   :  �     0      �
              ?        �                    3            �t�bhhK ��h��R�(KKG��h�B     c   ]                 <   `   #          N            c   �   �            W     �     	        �   �  �   �     s  "   k        
      U   d                 x           %   (   �        
      U      >        
  	         �t�bhhK ��h��R�(KK7��h�C�   -   <   *      �     &   S     �           	     }         v         �  t   h   H   	            �        �        �        �  =  E   �     �        }              �  �     �t�bhhK ��h��R�(KK+��h�C�         �        '           ^   �               0   T      +               �
        *     #   �        0   �  T   >     #   G            �t�bhhK ��h��R�(KK��h�C|              �                                Q        �     �      
   �   �  �     n        �t�bhhK ��h��R�(KK	��h�C$�  0   �        �           �t�bhhK ��h��R�(KK��h�C8D        k   x     <
  �         k   x        �t�bhhK ��h��R�(KK,��h�C�   �  �         \   V      	   M   �         �  �
  	   �   `   0  p   \     �  Y         '      \   V   4            (  )   �         �     �
  4      �t�bhhK ��h��R�(KK��h�C\    4  }     '   p   �     6         �         �   E     �  %     �        �t�bhhK ��h��R�(KK+��h�C�      n   �   P      �         �      %   _      �      �        �            �        �      V     ?  �              S   
      M  �         �t�bhhK ��h��R�(KK'��h�C�A        V  )      �  �            %   �         #                        '      r   �  2      n               B   �   �        �t�bhhK ��h��R�(KK��h�C@        �           �      �        M            �t�bhhK ��h��R�(KK��h�CT      <         .   �     j   P      	      �      �         	         �t�bhhK ��h��R�(KK��h�CD       f      3   U           G  �   Y   �     �      �t�bhhK ��h��R�(KK��h�Cx
               .   5  C     i            L   0      �   `   
   �   �  �   �      L   I         4      �t�bhhK ��h��R�(KK8��h�C�         a      �  �         h     5           &      [   �      	         t   <  �   	   �            �      `              f  �  �   0      a   ?   ]   >   �  8           �          �t�bhhK ��h��R�(KK��h�CD2   !   *   1  �      *   \   Q      0   �  �   I   �        �t�bhhK ��h��R�(KK��h�CD   B        �              t   s        E   �        �t�bhhK ��h��R�(KK(��h�C�            D     �            L      !      �   /         
      �  L      +  �           s      #   J   k     �   �              �t�bhhK ��h��R�(KK/��h�C�          �     +            �  M   �   
      Z  B     ,      D  �        �      �       �     2   !      �                  >   �         !   F	        �t�bhhK ��h��R�(KK��h�CP   �  �  H   .   �   ;   .  �            �  9        .  Z         �t�bhhK ��h��R�(KK��h�CT   �   9  x   y   M   �      �  �     w	        y      �               �t�bhhK ��h��R�(KK$��h�C�               �   �  �        �      *  K      �     �     ?     �            f        N      �     �  �        �t�bhhK ��h��R�(KK��h�Ch   <  A       �     �        F                     �   �  F         �           �t�bhhK ��h��R�(KK(��h�C��   &   
      	   �     	         -   
   *   �        &   
      \   �      	        �   	         �  
   �   S     j   �  
   9         �t�bhhK ��h��R�(KK��h�C8   @  y    �  ;   %                       �t�bhhK ��h��R�(KK��h�Cp   �   q   �   �  
   j   �               
   �   *            0      �         �   
   �         �t�bhhK ��h��R�(KK��h�CP�                  b     �            �  �     D      a        �t�bhhK ��h��R�(KK$��h�C�     �         �     %   _         O         `  O   *        O           O   u     H     �      I         0         �t�bhhK ��h��R�(KK��h�C\j   �   I   s   �     +            [          �   6  %         z	  [   �        �t�bhhK ��h��R�(KK��h�CPD      w     
   �         [   T            
   �      �  �        �t�bhhK ��h��R�(KK,��h�C�   
      {  e  [
     �	  �   8   �   T         >         D              D   �           �  >   �   �   �
    G   L        �   �  #      �        �t�bhhK ��h��R�(KK��h�C\n        n        n        o   l      �     <  Z      +   U     #         �t�bhhK ��h��R�(KK��h�Cx-      f   q   �            #   X  �        �     ,      u  �        ^            �	     �
        �t�bhhK ��h��R�(KK��h�C<   �   w             �               Z         �t�bhhK ��h��R�(KK��h�CX   &  �     �  �      �  X   [   w     �  �         �   =              �t�bhhK ��h��R�(KK,��h�C�  �  %  N      u   �            ]       &      	         {   C  	          
               �
           �   �      �      �     
   +   A        �t�bhhK ��h��R�(KK#��h�C�,         !            �  )   9   u   .  Z                  Y   )   /         r   '   3   Y   #     ,         �        �t�bhhK ��h��R�(KK��h�C\         k           =  Z     �  J   I      ?      I      ?               �t�bhhK ��h��R�(KK��h�C        �         �t�bhhK ��h��R�(KK��h�CL�     "               �   $   j     �     �  W     �        �t�bhhK ��h��R�(KK$��h�C�%   _      X     "         ]  
   H   2         �              <   x  E  �  7     �        �           �
  9         �t�bhhK ��h��R�(KK��h�C|   d  �        i  
      �                       
   �            1      v     K     �  �         �t�bhhK ��h��R�(KK&��h�C�   
   3   `  �     4     �   
   K   �   �      B        ^  �        m     (        �  H   �     4     ,      l            �t�bhhK ��h��R�(KK#��h�C�  P      )           �                  �               >   �   {                    �      >   U           �t�bhhK ��h��R�(KK��h�Cl+            �  .        
                  '   �     t         �  �         #         �t�bhhK ��h��R�(KK,��h�C�       �     '   )   8   H     �     '      �        �      '      �     M  y     '   U     	   �  L   �      n     ,        �   A   G  	         �t�bhhK ��h��R�(KK(��h�C�              �      9                  *   �  2            x	  2   1              �      .   b     .   �     �      �   J        �t�bhhK ��h��R�(KK��h�C4   n   �                                �t�bhhK ��h��R�(KK��h�C\%      !                       �            `   (      �  a   u            �t�bhhK ��h��R�(KK��h�C<      �  6           �          �  �         �t�bhhK ��h��R�(KK��h�C<   �   �
        �      c	  �      �   C   �         �t�bhhK ��h��R�(KK��h�CHj      *     #              j  X      �        Z        �t�bhhK ��h��R�(KK��h�C\@   �            �     s   �   �      �        �  ]   �      ^              �t�bhhK ��h��R�(KK"��h�C�!      �  �     
   �   �      +     �  
   .   �   a   ]                 �            �          _   ^        �t�bhhK ��h��R�(KK)��h�C�%      �                      �      I        �         �  $      G     ,            �             n   �     �        M        �t�bhhK ��h��R�(KK	��h�C$                          �t�bhhK ��h��R�(KK��h�CpK      @   a  �  �   p   �                     �        �   d	     e      d	     E   l        �t�bhhK ��h��R�(KK��h�Cx&        
         )   �     A	     �   )   �   @      w      #         O   ~     '         ;        �t�bhhK ��h��R�(KK,��h�C�    �         6   b   �   2         Y     8   !               �  9               i           �   M   �   >      �      B   �              T        �t�bhhK ��h��R�(KK'��h�C�      2     �     
     3   2   �     �  �     i        V              5            N            �  =            �        �t�bhhK ��h��R�(KK��h�Cl,   !   /            R     !   !       V     
            �   �         /     s        �t�bhhK ��h��R�(KK(��h�C�K      
  >   h      P   !               �      �     �  8   �      
      =  2   �      B   �        
      �  �      I     �         �t�bhhK ��h��R�(KK!��h�C�   �	  #      �   G        
  G   �         �  v      c      &      	   S   7   �      �   �      ?  �  �   	      �t�bhhK ��h��R�(KK*��h�C�         ^         1   C  T      �         \   �           	  �   >      0   B         >      �   Y   �   T         �   Y   �     �   5        �t�bhhK ��h��R�(KK!��h�C�      �  �  �  H            �   o        :  �   X   �  �  u   �   W     u      W     u   T  W     �         �t�bhhK ��h��R�(KK(��h�C�   0      u   0   (      >   �             %   R  U   �        >      Z     8   0            '   r              !         [        �t�bhhK ��h��R�(KK#��h�C�,   c   *      5        Z                g  �  >  �   w      �     �      #        F                          �t�bhhK ��h��R�(KK��h�CD�   7   w  0    
  $      B        $	  "   d   v        �t�bhhK ��h��R�(KK#��h�C�   ^        n         �  |   p   '  
     m  �        w     .   I        m        O     N  ?     .   �        �t�bhhK ��h��R�(KK!��h�C��      �   `      �   m   $              M   "      	  4   G         G      J   Z     G         
   |	           �t�bhhK ��h��R�(KK/��h�C�   &   
      D   �      	           �  ?      1   �  J   0     R                  
          3   �           �  	               �
  �                 �t�bhhK ��h��R�(KK��h�CD   $     w        B           5   �  0     
        �t�bhhK ��h��R�(KK��h�Cl          .   F   �        0   D   �   %        �             F   �  +   �   �            �t�bhhK ��h��R�(KK��h�C`      �     �         
      U   B                  �     
      U            �t�bhhK ��h��R�(KK��h�C0   7   s    #      /      7            �t�bhhK ��h��R�(KK��h�Cp   W   A      �  J   �   9     A     �      A   W   �  y   �         O  A   W   �     y        �t�bhhK ��h��R�(KK��h�C`   �   
   �      �  u        �   �   �  �   *   �               0   �  #         �t�bhhK ��h��R�(KK.��h�C�   q   �      #   ;   �     ,      *            I   [   �            �  !      q   .           
   �   #   �              
   �      m   $     0   A        �t�bhhK ��h��R�(KK3��h�C�   S           -   "  �     M   �               
      [     �                    @   �      !         [                 "  [                 �        	         �t�bhhK ��h��R�(KK3��h�C�j   �         7   �  �                  ]   !           �            	               ;   �  a     -      �   �  �        >   m
     �     �   D      

  �   	      �t�bhhK ��h��R�(KK��h�C0      "              �   d   "        �t�bhhK ��h��R�(KK��h�Cx�   $   S      �  _      �  .   F   O   *  a   X        O         #        O      O      O            �t�bhhK ��h��R�(KK��h�CX       I         )        L     ,   	                �  	         �t�bhhK ��h��R�(KK��h�Cl   2   
         L         �            �   �   P     7   8           �  �      	         �t�bhhK ��h��R�(KK��h�Cd2   ~   �      �  /         �  N   ~   �  P  �  W     :   �  �      �     I        �t�bhhK ��h��R�(KK&��h�C�   S   3      R     �     �   �  y   M   �         \   �      �  H         
  C      C  �        2   <            %  	         �t�bhhK ��h��R�(KK-��h�C�   �       �   !  %  N   �   �     g         *   �     M   �     
   �  q  <   �   s      ]  �   <         s   S
  G     !   *   �     �   �   s         �t�bhhK ��h��R�(KK��h�C`
   �         �     (      >         K        �      
   �  X   {   w  �        �t�bhhK ��h��R�(KK��h�CT   @      �  %   s     :  �   >   ,  ]      �   M   �         �        �t�bhhK ��h��R�(KK1��h�C�   &      	   %         �       d   �      �        S   �   a      L      ,   �         1      T             f   �     L   �   �     �     �   L      :   �  	         �t�bhhK ��h��R�(KK(��h�C�         ;   )   h   I   �                �      �   y      �       P     =         =   	       (      '      e  9     �        �t�bhhK ��h��R�(KK��h�CpK            [     �    $            �  $      E     +  $         8           4        �t�bhhK ��h��R�(KK'��h�C�         �     K  
        �  ?   M   V         �   ?   d        Y        �  %     �  ;   n   �        0   �	  >   �  �         �t�bhhK ��h��R�(KK��h�C<               -   E   �    �  e     e        �t�bhhK ��h��R�(KK:��h�C�     O  j      �       �   +   �      +            +   	     �     �            $      !      :   /      �            Y      �     R   T   �      e            Y      U  ;   R   T   �   	         �t�bhhK ��h��R�(KK��h�C\A   Y  $      �  /      A   Y  $      ~   �      L         <      d   |         �t�bhhK ��h��R�(KK��h�CX�   �  
   #         $     �                   (   3     �   T         �t�bhhK ��h��R�(KK��h�CP�   z      	         [  �               D  h   �   ~   �   	         �t�bhhK ��h��R�(KK��h�CP
      +         {   �                         /   2   1   2        �t�bhhK ��h��R�(KK!��h�C�          �     �   3   6      �     $      +      �	  2   @   �  d     �  :   �     �  6      !  $   	         �t�bhhK ��h��R�(KK7��h�C�   
   �   �  8                 `            �        �   �   *   �     H   u   h        
         	   �          n   �  m     @   	      j   �   
   l     �  #         <  �        �t�bhhK ��h��R�(KK��h�Ct%  A            �  2   �     -   
     L   4   j      
   �   N   �  6   
   �      �     L         �t�bhhK ��h��R�(KK%��h�C�j   6     M  �  �      �   v   5   �       ;   �     �         o     �  F            �        I   6      *               �t�bhhK ��h��R�(KK,��h�C�   <   �   ]   �   K     �   �     �   �        N   �   D     �     
        Y        �         
     :  �      �        r  @      M   �        �t�bhhK ��h��R�(KK��h�Cl�   �  �  2   �  �  �   K     1   �     �      >
           {   V      c      I   s         �t�bhhK ��h��R�(KK��h�CX                  �           �         �           �     _        �t�bhhK ��h��R�(KK��h�C`�   �           #     B   �              �   {   "     �  �     �   	         �t�bhhK ��h��R�(KK��h�Cp      �   �     9      �                       ^                       Z               �t�bhhK ��h��R�(KK��h�CD      y     X        �   �      |     
   2  �        �t�bhhK ��h��R�(KK)��h�C�%   
   �   �  $   .            �   
   (       e         �
  ?                 /      $               �	  8         �     :   �        �t�bhhK ��h��R�(KK��h�CT         u   [   x	  �   C   �  2      �           �	  `      �         �t�bhhK ��h��R�(KK��h�Ch   K   3         ,   !        $      (  1   V      Y     +   �
     a      �  	         �t�bhhK ��h��R�(KK*��h�C�   8  +   [       X        +           �  �     �   k            �  l      �  �     C            !   *   �
  �   *   �   `  ^   8        �t�bhhK ��h��R�(KK��h�C@    "  Y     <     *     .     �     
            �t�bhhK ��h��R�(KK��h�ClD  �         c      &      	           �   "      �  	                    c         �t�bhhK ��h��R�(KK��h�C@o   �  #      `        ^  �           n   Y        �t�bhhK ��h��R�(KK��h�C@�   B      D   �      �   E     �  %     �  �         �t�bhhK ��h��R�(KK ��h�C�   �     p   \               "      p   	     p   �        �      >        #   �        �  .   �        �t�bhhK ��h��R�(KK��h�C                     �t�bhhK ��h��R�(KK'��h�C�   !      :   /            o   W     $          �                    b  m   s                 �
     S   3  #      :   a        �t�bhhK ��h��R�(KK&��h�C��   D  �  %         ]            (  #      9   �  %   t  �         �   �           (  #   9         ~
  �  #   j   G            �t�bhhK ��h��R�(KK ��h�C�      N       (   �      �               
         ;   [   V         I   6   
   �  1  
      (           �t�bhhK ��h��R�(KK"��h�C�   %   
   �  1          I  C   I     1             1        6        S   
   �   �     �  �   �  	         �t�bhhK ��h��R�(KK��h�C`,      P   )            �         �   �     �     �      `     {   �  	         �t�bhhK ��h��R�(KK��h�Ct   z   
         	   �           N      ^   $                           $        �  %         �t�bhhK ��h��R�(KK3��h�C�f  +      T           �        *               �     S   3   �   �     ,   t         W     R   �  �   �   "   �            �      �      ,   #     s        $   	         �t�bhhK ��h��R�(KK#��h�C�       �  3  D     X   E   �     n     #   �           �      �   �   _            �  %         �   k  �        �t�bhhK ��h��R�(KK��h�CX       �     =      H  *   �  �      h     �  6      +         �        �t�bhhK ��h��R�(KK��h�Cp         �   :   �  U   2   #     �      �   _   `  #     �            N   :   �  �   +        �t�bhhK ��h��R�(KK,��h�C�        A  G   f        
   �  �            &      f     	         �
  p   �  �     $   �        K               �  3   �   S  `           �t�bhhK ��h��R�(KK��h�Cx   
   U        
   �              
  a         �	  E	  9      Z     t     
   J  �      �         �t�bhhK ��h��R�(KK9��h�C�%      <   �     �   Q        ?     �   �      e      %   (   �  P  �      �          (   u          #   �     (   t        %   
      P  i            P            �   
      1               �t�bhhK ��h��R�(KK��h�CL   M  (                 (                        �        �t�bhhK ��h��R�(KK��h�C,   �  X               �          �t�bhhK ��h��R�(KK+��h�C�   +            )   S   �   [         c  �  �        j   ,  [      ]   �   M   �      �   �   ]           �      �  �  N   �   +   [      	         �t�bhhK ��h��R�(KK'��h�C�   �   &            	   ~     �  ;   ~   �     ,   :   5  �        G   $                  &      =         �  M   �     =   	      �t�bhhK ��h��R�(KK!��h�C�   �  �	  �   #   �         �                         k  Q  �   �      ;                  %     |   o         �t�bhhK ��h��R�(KK&��h�C�     �                       �        "         7   h  �   %        "         "            7   5  �          �        �t�bhhK ��h��R�(KK(��h�C�   �     �     4     "      �        �   )   u  ?        f   �     )   1   �  �        '   r   �  :                G  �         �t�bhhK ��h��R�(KK��h�C4d   	  �         I        d   �           �t�bhhK ��h��R�(KK��h�Cx   �      �  �   0   o   |   �   }         !      �  �            
      �  \   Q   H   u   [   Z         �t�bhhK ��h��R�(KK��h�C`   -   '   4  }      _   $  ?   <   �  �   )         |  6      �  ]   8   )         �t�bhhK ��h��R�(KK��h�Ct         P   M   �     e         k   a     g         �   �   !      F     !      F  �   *        �t�bhhK ��h��R�(KK��h�Ct   &   3   /           	   @      Y            �              e  "      I   �     �   	         �t�bhhK ��h��R�(KK��h�Cd    -      5   �  �  #   H               �      �  *   �         �                 �t�bhhK ��h��R�(KK��h�CX   P   !      K            8  G   �     G      �      a        s        �t�bhhK ��h��R�(KK��h�C@g         V     u  �  �      )      �              �t�bhhK ��h��R�(KK��h�CP   j   
  *   �       �  
     �      �        �      �        �t�bhhK ��h��R�(KK/��h�C��      j  '      �              �        4      �  �   %   .   �     	   
         �   "   	   4   O         �   %                     	   
   p  �   	   4      �t�bhhK ��h��R�(KK=��h�C�      �   7   >  a   ;   $               &     ]   G   $         >         $                      U   �      $   >   �          <      +  x   d   �      �        6      �   �      $                    �t�bhhK ��h��R�(KK��h�CD          #            
   &          n   �           �t�bhhK ��h��R�(KK��h�CP                    �t�bhhK ��h��R�(KK.��h�C�        �  Y   �                                  �            X   L	        X   W           �                        Z        �   n  �   �      �t�bhhK ��h��R�(KK��h�Cl-      *   �     �                       �   v  5            n   v        K   �        �t�bhhK ��h��R�(KK��h�C|A   B   �     �            <           �  �   0   �     q   �           
         6                 �t�bhhK ��h��R�(KK��h�C|  2               0   �     "   C   0         �  7   5        i                     >   U   M	        �t�bhhK ��h��R�(KK,��h�C�   �   l   �     �         �  �     D   �      �  �               2                  �  �      �  �   !      ^   �  �         M     (   �         �t�bhhK ��h��R�(KK"��h�C�        +               �     !        !  �  N            0        +            �  0     �  �  @        �t�bhhK ��h��R�(KK��h�Cx&     p   �  �        _           �  �     B  �     �   '   �     �  �              �         �t�bhhK ��h��R�(KK2��h�C�   -      3      �        *   �   "   ?     �     "      �                     �             �                    A   `      �   j           �               �t�bhhK ��h��R�(KK;��h�C�   !   &            	   @         Z            .     G  8   �     ,                   &      =   8   :   �        �         =         3   `  $   K         d   �          �           h   	         �t�bhhK ��h��R�(KK)��h�C�-   �  �   Y        F      t     �      �   C            (   $  �           (   �   �        *              +   *        �            �t�bhhK ��h��R�(KK"��h�C�<      '     +            .      �      e      <         �	  .   	  �      <      �   $   .   o     .   �  *        �t�bhhK ��h��R�(KK��h�CH   M      w      "      
   &         �     {              �t�bhhK ��h��R�(KK��h�C0   �   �  #                  {        �t�bhhK ��h��R�(KK"��h�C�i      8     !      )   /      �  �  _      �   �        ?   �  [   �      �     r   '   
     �         a         �t�bhhK ��h��R�(KK,��h�C�e                     R   V   �   /   4   
      �         "   1   �  �           �           e      �     
   �   :  �     �  (  9   8   "         �t�bhhK ��h��R�(KK.��h�C��  '               �     >   m   {   �     �  4   �
     �     z  W  �   O      O         z        �   �  #      �  G      O           u  f  �        �t�bhhK ��h��R�(KK-��h�C�   
   �   �  0  9   #            M   V           e     d     2   �                       "  Y  *   1     ,        +   V     !   X   (   �        �t�bhhK ��h��R�(KK��h�CH            �   '   �        '   �     �  �               �t�bhhK ��h��R�(KK��h�C|c   K     	         
   4   	      z   c      	   
      3              	     V         �      	         �t�bhhK ��h��R�(KK��h�Cd                     >   h         s  :           �        0  9      '        �t�bhhK ��h��R�(KK��h�Cx�            O         �           O   u     �         <      q     0   j  '   1      �   �         �t�bhhK ��h��R�(KK��h�CL   W             /                 
         I      0         �t�bhhK ��h��R�(KK.��h�C�	     j      E   �  9               x         -         �   �  r           ~   �                  �  �      ,      �   $      1   �     \   V   	         �t�bhhK ��h��R�(KK��h�CP   &         7   �      =       %   3   �     f   �     "   4   =      �t�bhhK ��h��R�(KK��h�C@I   2   !   *   1  �         
            �  �        �t�bhhK ��h��R�(KK��h�CT(   �     c  +   C  2   ~  �     2   >        (   �   l   2            �t�bhhK ��h��R�(KK.��h�C�    �  �      �               �   /  .         �   �   H                  ]  �         �      q   m  �      �     ,  -      �   9           �   a         �t�bhhK ��h��R�(KK/��h�C�	   o   l      �   5            �  9   u      �	     _     �      *   �              c      �           6  �      �         �      +            .   $        �t�bhhK ��h��R�(KK��h�CH�            �  .   �      4   -   
   �  #   C   ~            �t�bhhK ��h��R�(KK��h�C<         q     
   #  6   �  P        	         �t�bhhK ��h��R�(KK(��h�C�   �  *  w   v      �        �        �        �  �     -   b   3   �   K                 b   .     �      �   #        #         �t�bhhK ��h��R�(KK��h�C\0   o   n     H      �  �     v     �  )        R  n     ~
  �  �         �t�bhhK ��h��R�(KK+��h�C�        I      T      
   *   �   #   �  #      �           ?   �     K         �  *   	  [     G      �              �   �      *   �        �t�bhhK ��h��R�(KK��h�Cp,         �	  %      z  �  O   �      z  �  O         z  �      3      O   �         h         �t�bhhK ��h��R�(KK-��h�C�   S   Y           %      �      2   (   �        +     %      �      2   (   �      %      B   h        �     �   �   �   >            &  (   �  �      �t�bhhK ��h��R�(KK"��h�C�g   P   !      %      �            �   C   ~   �      �      	   m        M   �      %         f   G     �   �   	      �t�bhhK ��h��R�(KK��h�Cdj   �     ]            &      	      $         �  �   �   	      �        �        �t�bhhK ��h��R�(KK-��h�C�8   �         �         ?   <   �  �  c  }   s          �	        4     �     y             +   c	  8   �          $
        N      8   �        �t�bhhK ��h��R�(KK��h�C|e      0   n   T   /  �     1      .      �          A     /     M      �   {      �      �     �        �t�bhhK ��h��R�(KK��h�CX-   8  J  @      �     #      &      	   �     �        b     4   	      �t�bhhK ��h��R�(KK.��h�C�   �     Q  �      >   �  ]      ,         !      :   /              ^   �  �               M     M   �         2      !  >   0         0               �t�bhhK ��h��R�(KK��h�C@     L  *         �        h        9   �         �t�bhhK ��h��R�(KK��h�C8J   E   �     �     {     0                 �t�bhhK ��h��R�(KK��h�CD   �  +   1   �   �  �   �     -   
   t     �          �t�bhhK ��h��R�(KK��h�Cl   	    �   R  �
  ]      &            	      $   �   x   2     ,   �  f   �  $   	         �t�bhhK ��h��R�(KK��h�CL   
   �   ]            �     (   �   i  D   _        �        �t�bhhK ��h��R�(KK&��h�C�   �           [  ]            *   Y  E         �	     
   *         �      �   K        	   �        �     0      4   	      �t�bhhK ��h��R�(KK,��h�C��   '   X        �   �      �        .              �  �   j           �         �  9           
      �  %   5   .     �      �  [   �         �t�bhhK ��h��R�(KK��h�C\    �  �   5   /               L      #   �   X   �      �   8   L      V	        �t�bhhK ��h��R�(KK!��h�C�       D  )   �   �  5   n   0  �     �      /  �      q   �  Z            �   (   �           �      ,        �t�bhhK ��h��R�(KK��h�C@   }  �        D   �         r        r           �t�bhhK ��h��R�(KK&��h�C�   3   �   7     
   *            &   
            	              y   {   �  	      j      #   t      D  0  _   �              �t�bhhK ��h��R�(KK��h�CD   &      	   �      7   �   �              �  	         �t�bhhK ��h��R�(KK ��h�C�   z   I   s         �     &      	   I   6   !      [    A   ^   	         �   �   �      !      y  �        �t�bhhK ��h��R�(KK��h�Cl   %   ~        1   �                          Y        �     �                   �t�bhhK ��h��R�(KK��h�CH                    .   �                 .   �        �t�bhhK ��h��R�(KK'��h�C�%   
   f   ,  ]   1   �                 
   p  �   1   $  �     �     +     ]      �  '           
   S   U   
  �   M   �         �t�bhhK ��h��R�(KK)��h�C�   	  X  *   
   �      �  Q                          
         |                    "  #      E   Z      ?        �      �         �t�bhhK ��h��R�(KK<��h�C�   "     �     �  F      �   D   Q               `   n  y           �            �      �   n        y           G   .   �  "         �         �       [     )         '   �   �         "         �t�bhhK ��h��R�(KK%��h�C�   *            A   /  C      "  
      �      e      @               '   r   /          �  6   '   �   Y  5   �        �t�bhhK ��h��R�(KK��h�CLb   �   N      X   $     [   .     X      }     I   P  �        �t�bhhK ��h��R�(KK��h�C<'  g   x        )            �   �  U            �t�bhhK ��h��R�(KK2��h�C�    ?   +   N      <  �         �   j           �        K         �   �  3         D   7        5   �  ?      +     	     D      G               
   `               �t�bhhK ��h��R�(KK!��h�C�   f   �   6   /      !      �     K      
   �  �     [   T         D   �     S      �     H  �      �        �t�bhhK ��h��R�(KK��h�C0               +            F         �t�bhhK ��h��R�(KK��h�C|,      j           B   P           ^   6   �           W   o      i      B   P     #   �      P        �t�bhhK ��h��R�(KK-��h�C�   �   �   &      q        	   7   F   �     L     /              �                   e     ,   �   &                 |     i      !   /         �t�bhhK ��h��R�(KK&��h�C�   3   �   7     
   *            &   
            	              y   {   �  	      j      #   t      D  0  _   �              �t�bhhK ��h��R�(KK��h�CH   �      �     (   �         D   _     �     �   
        �t�bhhK ��h��R�(KK"��h�C�	          P      )               �   }         X   �     i   D  }   _   <  �      
         >                 �t�bhhK ��h��R�(KK��h�C\            m   \     
   �      =         \  �     �   �  �              �t�bhhK ��h��R�(KK&��h�C�(   o  +   1   R     1   �   @       H              %   q       C   �  H     M  ?       �     �             �        �t�bhhK ��h��R�(KK��h�CDX      �               W  .                         �t�bhhK ��h��R�(KK2��h�C�         �     m    �         P   �      !   %   0  Q      %   E   �     {     1        e      1                             +        Z                       �t�bhhK ��h��R�(KK)��h�C�g      E   �   U         2         i     �        >         m
  �      �     ,      f   �   =  @        -   E         �      P   !         �t�bhhK ��h��R�(KK0��h�C��  M  �	  (  �  P  c        -   c          f      �            =      ,  E                             �
  9            j   }         7         =   	      �t�bhhK ��h��R�(KK��h�CH       ]     !      .   �        
         u   E   t        �t�bhhK ��h��R�(KK��h�C<            �        k  �   �   �  �            �t�bhhK ��h��R�(KK��h�CT         '      r   �      i         )   /	  @        �      )         �t�bhhK ��h��R�(KK+��h�C�   !   7  L      ^   C   :  o           �  !      �   /               �  `   a   L   �               
      L   J   �      2   N         �        �t�bhhK ��h��R�(KK1��h�C�   /   >        /   &            	     �        )            �      	     |   )            ;   �     Z     ;      |   �      ;   0   �     �  #      �   	         �t�bhhK ��h��R�(KK��h�CLd   #  �   B   �      �     �     �      �     �      `        �t�bhhK ��h��R�(KK��h�CX   
   �   L   h   �     �   L   @   Z      1   Z      I     _     �        �t�bhhK ��h��R�(KK��h�Ch%   3   �  f  H   �           
   �      �     #   �      �   �      (   �  B   |  4      �t�bhhK ��h��R�(KK��h�C4   /     �  ^	  �   <           T         �t�bhhK ��h��R�(KK��h�Cd   6      �                        :   {   V         S      �      u              �t�bhhK ��h��R�(KK��h�C4�  !      �     4  �   (   �      R        �t�bhhK ��h��R�(KK$��h�C�   u            �  >          �   M   �      �   
         $                       i  @               �           �t�bhhK ��h��R�(KK��h�Ct   �                k     x  �               n            +   ]  @       \  @  f        �t�bhhK ��h��R�(KK��h�C\e         

        �  Z            �  k   �          �      k   �        �t�bhhK ��h��R�(KK.��h�C�i         a         8     �      :   /      �       8   [   �         ?         +     %   5     -   �  �   v      �      �            (  H   u           �t�bhhK ��h��R�(KK��h�CL,      <  �  �   t   c     �                  5  �   �         �t�bhhK ��h��R�(KK��h�Cd   t   <  �  �  '   ^   8   )            �      Y      �        Y   $      !         �t�bhhK ��h��R�(KK(��h�C�   <  �         �   I            \   �   �  #   �      5        .   p     |  G   @         J      �      �  �   v   �   
   9   '        �t�bhhK ��h��R�(KK��h�C\�        �     '      �  h      J     3     V         /        	         �t�bhhK ��h��R�(KK��h�Cx   z   �         	      B            �  �  B   v	         +     t   8  ?   
   �   h  [   �  	         �t�bhhK ��h��R�(KK��h�CL1   �	  �  �                        	     
   �      =        �t�bhhK ��h��R�(KK.��h�C�!  �     3   �   o   �                        �      )   �           �   �     B   �   9	       ,      2      �     �         f      '   r   Y   �        �t�bhhK ��h��R�(KK��h�CLF	        7   �         �  
            �         �            �t�bhhK ��h��R�(KK)��h�C�   ;   �  �     E   {   \           <   ^        c  �         E              k   �  *   �   �        j   `   <   [        E          �t�bhhK ��h��R�(KK.��h�C�c   K     	   �   t   �         V      G   �      �   �  �     2   /      �  4   	      z   c      	   �   �   �      F      �                    K  	         �t�bhhK ��h��R�(KK��h�C\
   �  5  %  �        $    �   .  �     ,   
   *   .   �                 �t�bhhK ��h��R�(KK��h�C\,      J        f           I  �     e      
      �        ;   #         �t�bhhK ��h��R�(KK��h�CX      �  !      
   �     t               �	        
   �      \        �t�bhhK ��h��R�(KK��h�CH�        �      
         �   �
     �           �        �t�bhhK ��h��R�(KK#��h�C�?      
   #      �   k     -   
   j   �     l              
      �   �     �   W  G            ^      X            �t�bhhK ��h��R�(KK��h�Cl      M
                �  �   �    
            n        "  \     �	  =   F         �t�bhhK ��h��R�(KK��h�Cd         ^   ]                E        L                 �     1   ?        �t�bhhK ��h��R�(KK��h�Ch   &      	      r   '   �      =   (   3  �   %   m        x         >  A         =      �t�bhhK ��h��R�(KK"��h�C�         >   h   �               c     U   1      T            !      -   '                   b  �  @         �t�bhhK ��h��R�(KK��h�Cd      �     &      	   �            D    �     X  L   �      o   �              �t�bhhK ��h��R�(KK��h�C,7  
   �     �  M   �     &         �t�bhhK ��h��R�(KK��h�C<'  g   x        )            �   �  U            �t�bhhK ��h��R�(KK��h�CX,   �                  <   f   �  �        �  H         q      �        �t�bhhK ��h��R�(KK'��h�C�   +               �   C   :   {   P       P     ;         K              �   #      �  O         O         O      :  	         �t�bhhK ��h��R�(KK��h�C@e      p     �                 k   )  ;   �   4      �t�bhhK ��h��R�(KK ��h�C�       )  �     +            .   8     x  �   �        �  0      �     O  �     �      �     r        �t�bhhK ��h��R�(KK��h�CTS   E   >       U         �        1   �     -     a   ?            �t�bhhK ��h��R�(KK��h�CX      �   ~   �     �  �               $   9   G   "      +   :   F        �t�bhhK ��h��R�(KK��h�Ct    �     �  ,     +   �
     
   +      �        <               F      +      �     �         �t�bhhK ��h��R�(KK��h�CT   k  Q         �              F         I              F         �t�bhhK ��h��R�(KK&��h�C��   
   (
        �  <            �     �           �         
   �   {  9   8         r     �        �  ?         �         �t�bhhK ��h��R�(KK&��h�C�            F            _  G            F         �        '     �      �      (   +                 	        H        �t�bhhK ��h��R�(KK��h�Cl    h  �   k  c               9                  j   q   (   �   *   �           #         �t�bhhK ��h��R�(KK��h�Cp,   +            �     
   �               �     
   �                       Z           �t�bhhK ��h��R�(KK+��h�C�         $         q            <  <      W  �   �            (  1   V             m     *           B
     �            m   l
  k   �        �t�bhhK ��h��R�(KK.��h�C�%      3                  �  '         
      7         7   
     �  �        %         {
  %   n   �   �         �  '            W         %  V        �t�bhhK ��h��R�(KK#��h�C��            A     p   �         y                 "      g   !     �      �     $      T      �     ~   �         �t�bhhK ��h��R�(KK��h�CPp   �	  r   '   �            7   �  r   '   B   J           !         �t�bhhK ��h��R�(KK��h�C|j  �   B   N  �  /      (      �            N   �     	   �  f      �  $   �   j     u
  ~   �   	         �t�bhhK ��h��R�(KK��h�C8~      v     V  f            d      �        �t�bhhK ��h��R�(KK��h�Ch       �     �  �           �  9           �   �                      	         �t�bhhK ��h��R�(KK��h�CH    -   
   �   @      �   
   �	        ,   
   +   �   �        �t�bhhK ��h��R�(KK��h�Cp6      �   '         �  @   �     \   Z      	      �                  �  U      ~  	   4      �t�bhhK ��h��R�(KK��h�CT     �     �  �  �   �        q           
  �      
   �        �t�bhhK ��h��R�(KK��h�Cx   
   w   �      �      &      	            �  �      p  P   s            t         �   ?   	         �t�bhhK ��h��R�(KK2��h�C�      �      "      �   �     �      '   3      �   �            �           '   �   S	  c     R   �     �      '        �   �  �         '        �     ^   �         �t�bhhK ��h��R�(KK��h�CX   =   �   l   G                                �   l         f        �t�bhhK ��h��R�(KK��h�C8!     �  a  b      J   E     ?               �t�bhhK ��h��R�(KK��h�C\%   _      f   X  #            
   [        .   �     
      �      �        �t�bhhK ��h��R�(KK"��h�C�{  &      .   �      	            �      C       7   �   4   M  �   "      7   �   	         {  u  H      �        �t�bhhK ��h��R�(KK��h�CD!      [   �  k        1      �	     
      .   �        �t�bhhK ��h��R�(KK.��h�C�   
   ;  �   m   �  �  %   �   �        �     �   
   �   �   �               7  }     q   �        h   �     j   �   
   +  �  J	     :     �            �t�bhhK ��h��R�(KK��h�C\%         *     #   X               b   .   �      b      �
  9              �t�bhhK ��h��R�(KK��h�Cp  b         �     &      	      �   "   	          
   1  �     �   �      �     w   H         �t�bhhK ��h��R�(KK3��h�C�   &   
            	   �                  M        g      1       v   $      -      �   y   "   	         -   
   �   .   �   y         w   1     �         �  v            �t�bhhK ��h��R�(KK��h�CT�   �            ~   V   B   �   i  �  �   ?     1   $     1   �        �t�bhhK ��h��R�(KK"��h�C�s           ?      �   @      &         	      +   1      	      n   &      	      +      �             	         �t�bhhK ��h��R�(KK��h�CP�  �         k
  #         �   �  �  #      d      �      B        �t�bhhK ��h��R�(KK"��h�C��   Q  #      �        �  %   m        <           ?      ~        &      	   �  ;            F  L   	         �t�bhhK ��h��R�(KK/��h�C�9      0   '      j        4  �     a  �         '        �  �      4  �        �     |     e      4  �        �  i   �        �      y     _        �t�bhhK ��h��R�(KK��h�Cx!     7   /      8     r  9     C   o   (   -        N                  n   l     �   <  "   �      �t�bhhK ��h��R�(KK/��h�C�          �   �  �   $            �   $   R     �   d  J      �     (      t    �   
   `   c     �     \   Q               `   �   �  5         �  "        �t�bhhK ��h��R�(KK5��h�C�   3   L     �   I   6   
   *            s      &   
      	   6         I                  s   4   �   �     �      �	  �	  |         I   s   �   �   �   $   5   �  �      5  4   	      �t�bhhK ��h��R�(KK��h�C,   ~        p  �         (        �t�bhhK ��h��R�(KK��h�C<,   E   B  �   �      4        �   �   %  4   	      �t�bhhK ��h��R�(KK��h�CL   m  �      h  �   D           (   F   I  �   �   C            �t�bhhK ��h��R�(KK*��h�C�         r   '   �      =            R   �       4   /      "   3      t     %            :  :   �      U      �   "      h
  +     =   	      �t�bhhK ��h��R�(KK��h�Ct         �      !   7  [     ;     (   D          |   (   v              C     �          �t�bhhK ��h��R�(KK��h�C|,   o   i  0   �      [   i         b   i  �      [      I   6   b   *         �      �     �   :  	         �t�bhhK ��h��R�(KK2��h�C�        �      *   �   �         .
  �     9      �   �     z              
        N            �
        |             J   �     
       �  �      �        �t�bhhK ��h��R�(KK��h�CD   �     g  i   P         -      w      �     �         �t�bhhK ��h��R�(KK��h�C\A   Y        '  �         X     L               Y      L      f  �         �t�bhhK ��h��R�(KK-��h�C�@      6              p     "  �    5   �         �     �   �  �      H	           �     l     I   s              *   �  x   y   �      �        �t�bhhK ��h��R�(KK��h�C|   +     @       @	  @  x     5  J         �   <     �        J      )             +   �        �t�bhhK ��h��R�(KK��h�C\-         D    5   �
        �      5   �
        �        r  �  �        �t�bhhK ��h��R�(KK��h�C\   "                     �  �     �   "               �      �   >        �t�bhhK ��h��R�(KK��h�Cl,      �  `   ?        
   *   �      	                  �   "              _   	         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CP         
   *      e       N      F      �   �   
   �  �        �t�bhhK ��h��R�(KK��h�CT         �   1   y  O   1                  �   k  H   �  G   "   4      �t�bhhK ��h��R�(KK ��h�C��   �  $      �            7   u  �   �  #   y   $                  �   $         `        1      Z         �t�bhhK ��h��R�(KK#��h�C�   �              &      	   6   f               ^   $   4   	         z         	         �   "   m   7   �  	         �t�bhhK ��h��R�(KK(��h�C�  �         �	     7     
   *   y  F      �        �     7     
   *   N              �          I  �   �      -              �t�bhhK ��h��R�(KK��h�Cd         Y  !      :   /         I   ~   �         :  :   u        :  :   w        �t�bhhK ��h��R�(KK��h�Ct     &      D   �     	      E  �  	            z  �     �   1         n  �  ?               �t�bhhK ��h��R�(KK-��h�C�%     _      d     [   T              �         i   �   �  .   5                [   T           �   .      *  v  2   b            �   �   �         �t�bhhK ��h��R�(KK-��h�C�            A     �   D   T     �     I   [   c     �  #      �         �   
   �     �   j   a   }      �     �      
   b  l  [   �     �   
        �t�bhhK ��h��R�(KK"��h�C�              �  �  2      8   !   �                   \                       <
           �           �t�bhhK ��h��R�(KK��h�CT     *   T                   %   D   V     �     
	              �t�bhhK ��h��R�(KK%��h�C�?  $      
     M   V         �  ?   @         {     �  M         '   0      �           }   X   o   g        �  !         �t�bhhK ��h��R�(KK1��h�C�-     3   *   �  �  ;   �      �     �   
     G   0   D   �  x  �      G   �     G   0  Q      G   �     G              G   �        �  
   6  #      
            �t�bhhK ��h��R�(KK��h�Ct      t     -   
   +   1   �   U  �   �        <               
                             �t�bhhK ��h��R�(KK��h�Ch   �   #                           �  9   D   Q        8                  �        �t�bhhK ��h��R�(KK��h�Ct   T  #      [              �  %   �      >   c  H           �      	   �   `   K   L   4   	      �t�bhhK ��h��R�(KK��h�Cx�  _      <   �
        C  
  <            *   �  Q      �      �                 O   �           �t�bhhK ��h��R�(KK��h�CX      H
                            �   �  �   �  �      E   �        �t�bhhK ��h��R�(KK ��h�C�_  �      )      n     d    �      )         ,         '      �         e         R  3      '            �t�bhhK ��h��R�(KK!��h�C�g   P   �      !         �   �       �     �   	  W   	     K      g         h   ;   )      P   �      !         �t�bhhK ��h��R�(KK��h�C@   M   �   �   t  ?      �  Z      2   !   *   �         �t�bhhK ��h��R�(KK��h�C<,   �  �       I   6   �	     I     K           �t�bhhK ��h��R�(KK'��h�C�   -   s   �         ^     �  .   f     &      	   �   f     �   �   ?     �   �            T  Z      �     �      L   �  	         �t�bhhK ��h��R�(KK*��h�C�-      �   @      �     /            &            	      �     �       �   �   �   �           B   �      ;        0            �        �t�bhhK ��h��R�(KK��h�C8�	  �           �           e  �  �         �t�bhhK ��h��R�(KK4��h�Cе     I   @   N  �   %   #      Y   	   U  	      �   *  �  1            1   i  	      	         �            �  �  *  	      �	     	         �  �                  �        �t�bhhK ��h��R�(KK��h�Ct   z        &      �     	      ;     $      ,      �        `      O  �   d   �  y   "         �t�bhhK ��h��R�(KK��h�C4   (  �   G  H   5   �        q   �         �t�bhhK ��h��R�(KK��h�CH!      �   �     :   /      �     5   d     d       �      �t�bhhK ��h��R�(KK+��h�C�    �      I   6   *        �     �  8   !      �            m   ?       0      W        �   V      g      b   �           A   *   �  �         �t�bhhK ��h��R�(KK��h�C<   �      X  W          �  b  �     �         �t�bhhK ��h��R�(KK=��h�C�    ;   �  V      ;     �        ~              s              K   9      "         K   �      B               >   �   �	  C         2   <   �  �	  C   L  �        >   z  �        2   <      .   r        �t�bhhK ��h��R�(KK#��h�C��     �            &      	         �             �  "      
      e     /     �     i      B   M    	         �t�bhhK ��h��R�(KK��h�CL  g   y      (   �        ?     8               U           �t�bhhK ��h��R�(KK��h�CPO      /   �   �  /   4      
      N   �  4   v     e  �   �        �t�bhhK ��h��R�(KK��h�CX   �  +   
         X      *   �  �             �  �                    �t�bhhK ��h��R�(KK.��h�C�   �  L   �    !      e      �  L   &  C      �          (            �	              
      h   ;   L   �  1   �     �  1               �   	         �t�bhhK ��h��R�(KK��h�Cd8   �   �      B  �  1   �     &            	   {  �            
   �  %   	         �t�bhhK ��h��R�(KK��h�C<   �      |  W          �     �   9  �         �t�bhhK ��h��R�(KK��h�CL    9   5   (            5   (   �          5            �t�bhhK ��h��R�(KK��h�CL�  D      -  �      �          m              �  �        �t�bhhK ��h��R�(KK��h�Cx   �  �         �         �   �            
   �   �                �      Z           6        �t�bhhK ��h��R�(KK��h�C<�  �  �         |     +  �   ]   �      K	        �t�bhhK ��h��R�(KK!��h�C�     '   '  )   �  -  	         &            	   A   W            �     A   B   /      �      t   <  	         �t�bhhK ��h��R�(KK��h�C\         k           =  Z     �  J   I      ?      I      ?               �t�bhhK ��h��R�(KK%��h�C�g      %   3      �  �  %   j        �   <   ,     -            �      `       
         �     !      K     �  	         �t�bhhK ��h��R�(KK��h�C|   �   P
  >   Z        �                     )         U   �           �   U   �  �   �   �  H        �t�bhhK ��h��R�(KK��h�CP           (   F   +         (   F   +         (   F   +            �t�bhhK ��h��R�(KK��h�Cl%   _   �  �   .            >      M  �     �        B   W              �  J            �t�bhhK ��h��R�(KK2��h�C�   &      R   �      	   K            U
  "   �   U                                        �  "   B      ;   �      e      U     r     R   �            ?  	         �t�bhhK ��h��R�(KK��h�C`    -   �  w      
     �     �  9   G         ,   
   *                       �t�bhhK ��h��R�(KK#��h�C�           8   !   I         �  �     I      �  �              �   :   M        %         �     �   !            �t�bhhK ��h��R�(KK&��h�C�      �  �  >   V  "                  g         �  �   5          �                 R   T      7         �   m   n        �t�bhhK ��h��R�(KK��h�Cd?   �  5           J   �                     F     N  �        �  �            �t�bhhK ��h��R�(KK��h�CP      "      /      1   �  �         q  "      ;     �
  s        �t�bhhK ��h��R�(KK��h�CT   �   �         @         3           �  �        �     *        �t�bhhK ��h��R�(KK��h�C<,   0               {   @        W   {   Q         �t�bhhK ��h��R�(KK'��h�C��   �      �   �   X      �           =   !   &      7   �      X  $      7   �  �        k         �  d   �  $         �
     =      �t�bhhK ��h��R�(KK)��h�C�%         @      �        �     $   2      �  %  �  �            �   �  :         L        t                                      �t�bhhK ��h��R�(KK��h�C4      )   %      �  �     X              �t�bhhK ��h��R�(KK��h�Cpl  �      ]   f
  G   #        <
  �            �         D              g  #               �t�bhhK ��h��R�(KK��h�CL   -   /     9      K           �  0   �     �      �        �t�bhhK ��h��R�(KK��h�Cl      �   <   �         #  �       e      0                *   �   	     �   	         �t�bhhK ��h��R�(KK,��h�C�-   
   j   �   T  W  a   ]   C   k   �               �     �  o       +	  =   F         �         -         �  C           
         W        �t�bhhK ��h��R�(KK��h�C8   �  �   �   "  A   B   �   )   X   �   �         �t�bhhK ��h��R�(KK��h�CH�      �        (      4   �      #   }   e  (      I  4      �t�bhhK ��h��R�(KK��h�Cx?   S     �     "  Y  �        �   ;   �      j   r   '   m
     �     �     =   Y
  �   �  �   =      �t�bhhK ��h��R�(KK��h�Ch      �              -      *      9            x      �         ?   *   _            �t�bhhK ��h��R�(KK��h�CD   �   L      1         �   �	        �   �     L         �t�bhhK ��h��R�(KK��h�CD  �      )      �  y   /      A        �   �   �         �t�bhhK ��h��R�(KK��h�Cd      U      �   2   �     
         2               2      �     
   _           �t�bhhK ��h��R�(KK*��h�C�g   P   !      %   c      R     
         h   }      �   $        _  _      �     
         G      +  ]   _   R  O   �  9   _      G            �t�bhhK ��h��R�(KK��h�CHq  "      7   F      ~   �         �   p   \  
  d   �         �t�bhhK ��h��R�(KK��h�Cdf        F               N      \   Q             n         %  �              �t�bhhK ��h��R�(KK+��h�C�g   P   �      !   7        �        R   T            1     �        �     -   
   �  $               .   1  G   $      2   <   �              �t�bhhK ��h��R�(KK&��h�C�-      �  w   }      �     &   �           	                  [  	      A   ^   2   
      �   4   �           �      	         �t�bhhK ��h��R�(KK+��h�C��      �  R   T   �     �  Z      	   �         !      �  4        �      �   ?   4   	   e      �   B         "      D   �	        D   p  H  4      �t�bhhK ��h��R�(KK,��h�C�      :   �           ^   _                        :   �              9            V  @   �   8           8              !      )   /         �t�bhhK ��h��R�(KK��h�C0   <   ^  |   D   �  0   �     �         �t�bhhK ��h��R�(KK#��h�C�   �   r      �  �     @      a     '   r   6  v   E   P
     =       '   �      �  �   7        6   �   '   �   �   �      �t�bhhK ��h��R�(KK��h�CH      �  w   H               (   �      �      �  �        �t�bhhK ��h��R�(KK��h�C`   �     L                 �           "           B  V     �   �        �t�bhhK ��h��R�(KK��h�Cx   -   S  w   }   X   
     ]  b      	   I   a  �   �                           �  :   �   4   	      �t�bhhK ��h��R�(KK ��h�C�   !         �   Y  $   �        f   Y   (         2   
      �      $               f   �   0   (   "        �t�bhhK ��h��R�(KK��h�C4j   �  
   #   �                  �        �t�bhhK ��h��R�(KK��h�C|   9  �   .         �       (   �     (        &      	   K      !         $      U  ;   .   �        �t�bhhK ��h��R�(KK��h�C<              
     -   
   +      �   �        �t�bhhK ��h��R�(KK!��h�C�(     W                    h     B                K         2      K   �           
   2               �t�bhhK ��h��R�(KK��h�C<,   E         -     
      �  E   �  G   $         �t�bhhK ��h��R�(KK��h�Ct   �     �     $
             �        s   ~
           q   �      "  #      D   �   	         �t�bhhK ��h��R�(KK��h�C@!   �  �   [         �                 M  �        �t�bhhK ��h��R�(KK,��h�C�      &      D   �      	               /      e  K      )         +  )   9   5   @   Z         Z      
      .     G  8   �     ,       	         �t�bhhK ��h��R�(KK��h�C@  �     �   u                                   �t�bhhK ��h��R�(KK��h�Ct�   &      .   �     	        7   �   �  �   "     �        `   �           5   (     �   	      �t�bhhK ��h��R�(KK��h�CD   �         9   X            _  7  �  1      �        �t�bhhK ��h��R�(KK*��h�C�  
  �   l   (   3  �   �           +      �            w   �      >  �  l              R   �           &      	   �  �      )   �   	      �t�bhhK ��h��R�(KK��h�Cl         �  :   F      	   A   l   �  �                 -  �   �   !   L   H   u           �t�bhhK ��h��R�(KK��h�Ct               �   K         ?   
   h  J   �  :  J           &      	   �   �   +               �t�bhhK ��h��R�(KK��h�Cp      <      �  z         	   �           �     $   7   F                        s        �t�bhhK ��h��R�(KK��h�Cx    %      �     �            ;   �         �     _   C        �         �   �   �  �  �            �t�bhhK ��h��R�(KK��h�CD6   <   3   &  �  �   ;           f  S      Y   �        �t�bhhK ��h��R�(KK��h�CH7   r  f      #     y         8   7   �  f      �  �         �t�bhhK ��h��R�(KK'��h�C��  '      �        �  �   �  6   �   �         �   '      j     �     i      "   �   �           H   u   �     g   �  �  )         �t�bhhK ��h��R�(KK#��h�C�{     �   M            �   �         �     �  �     �            d   �      ~   T      '        }   X   o   g        �t�bhhK ��h��R�(KK��h�Cp   
   w         �     &   e        z   �      &      =   e      �   =          
   �            �t�b��      hhK ��h��R�(KK��h�C|   &   b      	   K      :         t  �      [   T         .   f     |  N      �         :      	         �t�bhhK ��h��R�(KK��h�Ch   I   s      q   �            c   t   �  *   Y        w        F      *   �   �	        �t�bhhK ��h��R�(KK%��h�C�   �   &      	         K        �   �     �                    K   >   Z                       K   >   Z  N  	         �t�bhhK ��h��R�(KK��h�C0   @      �  %               �
        �t�bhhK ��h��R�(KK%��h�C�         +  �   �      (   "
        
      m   a   �     �
                   X  �        7     
   m   �   #   �        �t�bhhK ��h��R�(KK��h�C<"     (   V              �  %   0   (   |         �t�bhhK ��h��R�(KK$��h�C�O            
      -   
         �            p     �	  �	     _   �     6      3   S   Y      �     |  �      #         �t�bhhK ��h��R�(KK��h�C<         �       <   ^         0   o   �        �t�bhhK ��h��R�(KK��h�C8   >      %   M   \     ,   M   V     �         �t�bhhK ��h��R�(KK��h�Cl                                 0   �                               0   �        �t�bhhK ��h��R�(KK��h�CP-   �     @      �         v      +
          l  D              �t�bhhK ��h��R�(KK��h�C\      j   E     L        C  1              U         1      :   �         �t�bhhK ��h��R�(KK1��h�Cď   z      &            	   %      �   �  %   "   �         �  �   R   |     ,      J  �        �         �     �          '   �     �     �      O   �     �         �t�bhhK ��h��R�(KK��h�C �  �      �     L         �t�bhhK ��h��R�(KK��h�CL    �  :
  �         <   m                 �   N     |        �t�bhhK ��h��R�(KK��h�Cd�   O     B           �     i         �   �  �   $   ;   O     i         D  4      �t�bhhK ��h��R�(KK��h�Cx   &   
            	   5               5         w      	          |   �   
          �           �t�bhhK ��h��R�(KK��h�C`   %      q     .   �  V   �   1   =     O      .     #            �   -        �t�bhhK ��h��R�(KK
��h�C(M                           �t�bhhK ��h��R�(KK$��h�C�    �    H            0   \   �     �   �      	   -   '   �     

        �     =   3      �  �   �      4     =   	      �t�bhhK ��h��R�(KK��h�C|!   w   2      ?     
  �      
   
  0   k   ?	     
   }  k   �           
   ;   �  �   �     �        �t�bhhK ��h��R�(KK#��h�C�t         �     �  O         h   }      M   2        R           4  L             f     h   }      M   2        �t�bhhK ��h��R�(KK��h�CD�        u     �  �   x         
                    �t�bhhK ��h��R�(KKA��h�B     !   &      9     	   �   O  �     �  ;     4         �   *        ,      f      E     
      Y   �   ;   �         ~   �          a   �      f   [  $               ,         (   �         4  8   "      �   	         �t�bhhK ��h��R�(KK��h�CP   0      �                 J                 #      �         �t�bhhK ��h��R�(KK��h�Ch         z  �   (   �    �  #                       �      J   �  �   �   �	        �t�bhhK ��h��R�(KK��h�C|8      �   
     �     8      <  �      8      >  1   �     8   +         C   (            �           �t�bhhK ��h��R�(KK&��h�C�-      &  6  "            U           �  �   ,   6   �      �   ^         h   C   c      �  �   7     <   �  �     �   4   �      �t�bhhK ��h��R�(KK��h�Ch   E   Q        z     �   ,   Z          �   �  �   O   N   �         n   �  r        �t�bhhK ��h��R�(KK��h�C ,   �   W         �        �t�bhhK ��h��R�(KK��h�Cx
   �      ]   ;   �  �     �      �      �  �     
   �         �  u           u         s        �t�bhhK ��h��R�(KK��h�CX-      j     l     ~               �  ]  `   �         %   	  �        �t�bhhK ��h��R�(KK��h�CX   
         m      .   J                          t   �      �         �t�bhhK ��h��R�(KK#��h�C�   !   �   "        ?   
                 	   !   �   !   �   �      /      �                �            �        �t�bhhK ��h��R�(KK��h�CX   
   &            	   �   9      a   d   o     :   ;     B  $   	         �t�bhhK ��h��R�(KK��h�C4g         �      �  �  �      i           �t�bhhK ��h��R�(KK'��h�C�              +         �      �   @         -      *   Y     �        �     v         �  �      �     (      Q  "   @         �t�bhhK ��h��R�(KK ��h�C�%     �   m   �         �           
   `  C   @      #      �        `  �     #   C   
     D   �         �t�bhhK ��h��R�(KK��h�CT   &   
      "      a         f   [  $   �     x      j     =   	      �t�bhhK ��h��R�(KK��h�C<      �  #      �      >  �     9     H        �t�bhhK ��h��R�(KK��h�C<1      �  E  A         1         �   �  �         �t�bhhK ��h��R�(KK��h�CPe      S   :   �   Y   3  ;   d   �        S   0   d   �  U   $  �      �t�bhhK ��h��R�(KK��h�C`   
   &            	         �
        �   @         )      �  R   z  C        �t�bhhK ��h��R�(KK!��h�C�,   �  �     �      2   A   ;        $        �     �  �     N   /   X   �   +        W   �  ]              �t�bhhK ��h��R�(KK$��h�C�   -   b      �        F	  b   E  D               P      =   B     "      ,         �              *      x      =      �t�bhhK ��h��R�(KK��h�CL      i  �        �   b      9            �  �  |            �t�bhhK ��h��R�(KK��h�C`   0   #  �     \   Q   �   2      �     �      ,  ]           >   �  �         �t�bhhK ��h��R�(KK6��h�C�j   �  �  �     #      &            	   6         �   G   L   �   �           "   G   $      �         �  h   "      R   �     �        �   �  4         X          G   "   	         �t�bhhK ��h��R�(KK=��h�C�,      J     '   C   7   �  r   �   )         6   �           �     y      �            1  )   a      g      =  L  )      K  
     -   '   '  6   2        M   �            '         X   �     �  	         �t�bhhK ��h��R�(KK��h�CD            s                    �                 �t�bhhK ��h��R�(KK��h�CT    o      �   C   R   �        i           >   &  v      �  �        �t�bhhK ��h��R�(KK��h�C4   �   �  �   �                  &         �t�bhhK ��h��R�(KK#��h�C�      `   +  �                 	     �   c            
   `   �   �     �  K   �         ,   b   +         W        �t�bhhK ��h��R�(KK��h�C`e      7        Y   �                  Y   E   /            >   Y   R   T         �t�bhhK ��h��R�(KK��h�Cd,   K            B   �  x   y   $   >   �        Y  +                  5   $         �t�bhhK ��h��R�(KK��h�C8         +  ]   (   �      k                 �t�bhhK ��h��R�(KK��h�Cx            <   *   h  9   ;                  6   
   +            *   �         	   �  �   	         �t�bhhK ��h��R�(KK'��h�C�
   `   N   U      �            5     �        �   W         i   N   /              ;     �   �   �  *      >  
   �   +   *        �t�be.