i Esbo finns finskspråkiga och svenskspråkiga grundskolor ( peruskoulu ) .
undervisning kan även fås på engelska .
skolan börjar vanligtvis det året då barnet fyller sju år .
anmälan till grundskolan ska göras på förhand .
Anmälningstiden är vanligtvis i januari .
på stadens webbplats hittar du kontaktuppgifterna till skolorna och mer information om anmälan .
om du har frågor om den grundläggande utbildningen kan du kontakta Resultatenheten för den finskspråkiga undervisningen ( Suomenkielisen opetuksen tulosyksikkö ) .
Resultatenheten för den finskspråkiga undervisningen
Kamrersvägen 3 B
tfn ( 09 ) 816.52044 och ( 09 ) 816.52043
grundläggande utbildning .
linkkiEsbo stad :
grundläggande utbildningfinska _ svenska _ engelska
linkkiEsbo stad :
anmälan till skolanfinska _ svenska _ engelska
linkkiEsbo stad :
Espoo International Schoolfinska _ engelska
internationella skolor i huvudstadsregionenfinska
linkkiExpatFinland.fi :
internationella skolor i huvudstadsregionenengelska
linkkiEsbo stad :
Eftermiddagsverksamhetfinska _ engelska
hemspråksundervisning för invandrare
barn med invandrarbakgrund och barn från tvåspråkiga familjer kan få hemspråksundervisning ( oman äidinkielen opetus ) om tillräckligt många barn anmäler sig till gruppen för det egna språket .
undervisning ges två timmar i veckan .
anmälan till hemspråksundervisning görs varje år i mars .
mer information hittar du på Esbo stads webbplats .
linkkiEsbo stad :
förberedande undervisning för barn i förskoleåldern ( pdf , 100 kb ) finska _ engelska _ ryska _ estniska _ somaliska _ kinesiska _ arabiska _ kurdiska _ albanska
linkkiEsbo stad :
förberedande undervisning för barn i förskoleåldernfinska _ engelska
linkkiEsbo stad :
hemspråksundervisningfinska _ engelska
yrkesutbildning
på Omnia kan man studera många olika yrken .
på Omnia ordnas för invandrare utbildning som förbereder dem på yrkesutbildning .
den förberedande utbildningen är avsedd för unga och vuxna , som är intresserade av yrkesstudier och vill förbättra sina kunskaper i finska ..
Esbobor kan också ansöka till yrkesskolorna i Helsingfors och Vanda .
Läs mer : yrkesutbildning
yrkesutbildningfinska _ engelska
linkkiEsbo stad :
Yrkesläroanstalterfinska _ engelska
Yrkesläroanstalterfinska _ svenska _ engelska
linkkiVanda stad :
yrkesutbildningfinska _ svenska
gymnasium
i Esbo finns elva finskspråkiga och ett svenskspråkigt gymnasium ( lukio ) .
i två av gymnasierna i Esbo finns en engelskspråkig IB @-@ linje .
ungdomar från Esbo kan också söka till gymnasier i andra städer .
i Esbo finns ett vuxengymnasium ( aikuislukio ) där vuxna kan avlägga gymnasie- och studentexamen .
på gymnasiet kan man även höja vitsorden i sitt avgångsbetyg eller studera enskilda ämnen .
invandrarungdomar kan dessutom studera finska och avlägga grundskolans lärokurs .
i gymnasiet Leppävaaran lukio ordnas för invandrare och utlänningar utbildning som förbereder dem på gymnasiet .
utbildningen är avsedd för unga som vill studera på gymnasiet , men vars språkkunskaper inte är tillräckliga för gymnasiestudier .
Läs mer : gymnasium
linkkiEsbo stad :
Gymnasierfinska _ svenska _ engelska
linkkiEsbo stad :
Vuxengymnasietfinska
linkkiEsbo stad :
Gymnasieförberedande utbildning för invandrarefinska _ engelska
linkkiEsbo vuxengymnasium Omnia :
grundläggande utbildning för invandrarefinska
om du är under 30 år gammal kan du få råd och handledning via Ohjaamo @-@ tjänsten .
Ohjaamos personal hjälper dig om du inte har ett arbete eller en studieplats .
du kan även fråga om andra saker , som till exempel boende eller ekonomiska frågor .
kontaktuppgifter :
Fågelbergavägen 2 A
Puh . 040.126.7513
linkkiEsbo stad :
Ohjaamofinska _ svenska _ engelska
Högskoleutbildning
i Esbo finns tre högskolor :
yrkeshögskolan Laurea
yrkeshögskolan Metropolia .
vid högskolorna kan du avlägga högskoleexamen .
mer information finns på Aalto @-@ universitetets , Laureas och Metropolias webbplatser .
också i Helsingfors finns det universitet och yrkeshögskolor där man kan studera inom många områden .
mer information hittar du på Helsingfors stads webbplats .
Läs mer : Högskoleutbildning
universitet inom teknik , konst och ekonomifinska _ svenska _ engelska
yrkeshögskolafinska _ engelska
linkkiMetropolia :
yrkeshögskolafinska _ engelska
Högskolorfinska
andra studiemöjligheter
vid Esbo arbetarinstitut ( Espoon työväenopisto ) kan du studera till exempel språk , handarbete och matlagning eller delta i ledd motion .
kurserna är avgiftsbelagda . kurser anordnas både dagtid och kvällstid .
vid arbetarinstitutet kan vem som helst studera .
vid Esbo bildkonstskola ( Espoon kuvataidekoulu ) kan barn och unga studera bildkonst .
studierna är avgiftsbelagda .
vid Esbo musikinstitut ( Espoon musiikkiopisto ) kan barn och vuxna studera musik .
Läs mer : andra studiemöjligheter
linkkiEsbo stad :
Arbetarinstitutetfinska _ svenska _ engelska
linkkiEsbo biIdkonstskola :
bildkonst för barn och ungafinska _ svenska _ engelska
linkkiEsbo musikinstitut :
Musikundervisning för barn och vuxnafinska _ engelska
dagvård
förskoleundervisning
grundläggande utbildning
hemspråksundervisning för invandrare
yrkesutbildning
gymnasium
stöd och handledning för unga
Högskoleutbildning
andra studiemöjligheter
dagvård
i Esbo finns både kommunala och privata daghem .
i Esbo finns dessutom familjedagvårdare .
dagvård fås på finska och på svenska .
Ansök om dagvårdsplats minst fyra månader innan barnet ska börja i dagvården .
om du till exempel oväntat får arbete eller en studieplats kan du ansöka om vårdplats senare .
när du ansöker om vårdplats ska du fylla i en ansökningsblankett .
du kan också söka dagvårdsplats via Internet .
familjer som bor i Esbo kan också söka dagvårdsplats till sitt barn i Helsingfors , Vanda eller Grankulla .
du ska ändå lämna in din ansökan i Esbo .
mer information får du via tjänsten Helsingforsregionen.fi .
Läs mer : dagvård .
linkkiEsbo stad :
dagvårdfinska _ svenska _ engelska
linkkiEsbo stad :
ansökan om dagvårdsplatsfinska
linkkiEsbo stad :
Servicepunktfinska _ svenska _ engelska
linkkiEsbo stad :
Dagvårdens samanvändningsområdefinska _ svenska _ engelska
förskoleundervisning
i Esbo anordnas förskoleundervisningen ( esiopetus ) i daghemmen .
förskoleundervisning ges på finska och på svenska .
till förskoleundervisningen anmäler man sig via Esbo stads webbplats .
förskoleundervisningen börjar i augusti .
ansökningstiden är vanligtvis i januari .
i frågor kring barndagvård och förskoleundervisning kan du också kontakta daghemsföreståndarna eller stadens chef för småbarnsfostran ( varhaiskasvatuspäällikkö ) .
kontaktuppgifterna finns på stadens webbplats .
Läs mer : förskoleundervisning .
linkkiEsbo stad :
förskoleundervisningfinska _ svenska _ engelska
linkkiEsbo stad :
ansökan till förskoleundervisningfinska _ engelska
grundläggande utbildning
i Esbo finns finskspråkiga och svenskspråkiga grundskolor ( peruskoulu ) .
undervisning kan även fås på engelska .
skolan börjar vanligtvis det året då barnet fyller sju år .
anmälan till grundskolan ska göras på förhand .
Anmälningstiden är vanligtvis i januari .
på stadens webbplats hittar du kontaktuppgifterna till skolorna och mer information om anmälan .
om du har frågor om den grundläggande utbildningen kan du kontakta Resultatenheten för den finskspråkiga undervisningen ( Suomenkielisen opetuksen tulosyksikkö ) .
Resultatenheten för den finskspråkiga undervisningen
Kamrersvägen 3 B
tfn ( 09 ) 816.52044 och ( 09 ) 816.52043
grundläggande utbildning .
linkkiEsbo stad :
grundläggande utbildningfinska _ svenska _ engelska
linkkiEsbo stad :
anmälan till skolanfinska _ svenska _ engelska
linkkiEsbo stad :
Espoo International Schoolfinska _ engelska
internationella skolor i huvudstadsregionenfinska
linkkiExpatFinland.fi :
internationella skolor i huvudstadsregionenengelska
linkkiEsbo stad :
Eftermiddagsverksamhetfinska _ engelska
hemspråksundervisning för invandrare
barn med invandrarbakgrund och barn från tvåspråkiga familjer kan få hemspråksundervisning ( oman äidinkielen opetus ) om tillräckligt många barn anmäler sig till gruppen för det egna språket .
undervisning ges två timmar i veckan .
anmälan till hemspråksundervisning görs varje år i mars .
mer information hittar du på Esbo stads webbplats .
linkkiEsbo stad :
förberedande undervisning för barn i förskoleåldern ( pdf , 100 kb ) finska _ engelska _ ryska _ estniska _ somaliska _ kinesiska _ arabiska _ kurdiska _ albanska
linkkiEsbo stad :
förberedande undervisning för barn i förskoleåldernfinska _ engelska
linkkiEsbo stad :
hemspråksundervisningfinska _ engelska
yrkesutbildning
på Omnia kan man studera många olika yrken .
på Omnia ordnas för invandrare utbildning som förbereder dem på yrkesutbildning .
den förberedande utbildningen är avsedd för unga och vuxna , som är intresserade av yrkesstudier och vill förbättra sina kunskaper i finska ..
Esbobor kan också ansöka till yrkesskolorna i Helsingfors och Vanda .
Läs mer : yrkesutbildning
yrkesutbildningfinska _ engelska
linkkiEsbo stad :
Yrkesläroanstalterfinska _ engelska
Yrkesläroanstalterfinska _ svenska _ engelska
linkkiVanda stad :
yrkesutbildningfinska _ svenska
gymnasium
i Esbo finns elva finskspråkiga och ett svenskspråkigt gymnasium ( lukio ) .
i två av gymnasierna i Esbo finns en engelskspråkig IB @-@ linje .
ungdomar från Esbo kan också söka till gymnasier i andra städer .
i Esbo finns ett vuxengymnasium ( aikuislukio ) där vuxna kan avlägga gymnasie- och studentexamen .
på gymnasiet kan man även höja vitsorden i sitt avgångsbetyg eller studera enskilda ämnen .
invandrarungdomar kan dessutom studera finska och avlägga grundskolans lärokurs .
i gymnasiet Leppävaaran lukio ordnas för invandrare och utlänningar utbildning som förbereder dem på gymnasiet .
utbildningen är avsedd för unga som vill studera på gymnasiet , men vars språkkunskaper inte är tillräckliga för gymnasiestudier .
Läs mer : gymnasium
linkkiEsbo stad :
Gymnasierfinska _ svenska _ engelska
linkkiEsbo stad :
Vuxengymnasietfinska
linkkiEsbo stad :
Gymnasieförberedande utbildning för invandrarefinska _ engelska
linkkiEsbo vuxengymnasium Omnia :
grundläggande utbildning för invandrarefinska
om du är under 30 år gammal kan du få råd och handledning via Ohjaamo @-@ tjänsten .
Ohjaamos personal hjälper dig om du inte har ett arbete eller en studieplats .
du kan även fråga om andra saker , som till exempel boende eller ekonomiska frågor .
kontaktuppgifter :
Fågelbergavägen 2 A
Puh . 040.126.7513
linkkiEsbo stad :
Ohjaamofinska _ svenska _ engelska
Högskoleutbildning
i Esbo finns tre högskolor :
yrkeshögskolan Laurea
yrkeshögskolan Metropolia .
vid högskolorna kan du avlägga högskoleexamen .
mer information finns på Aalto @-@ universitetets , Laureas och Metropolias webbplatser .
också i Helsingfors finns det universitet och yrkeshögskolor där man kan studera inom många områden .
mer information hittar du på Helsingfors stads webbplats .
Läs mer : Högskoleutbildning
universitet inom teknik , konst och ekonomifinska _ svenska _ engelska
yrkeshögskolafinska _ engelska
linkkiMetropolia :
yrkeshögskolafinska _ engelska
Högskolorfinska
andra studiemöjligheter
vid Esbo arbetarinstitut ( Espoon työväenopisto ) kan du studera till exempel språk , handarbete och matlagning eller delta i ledd motion .
kurserna är avgiftsbelagda . kurser anordnas både dagtid och kvällstid .
vid arbetarinstitutet kan vem som helst studera .
vid Esbo bildkonstskola ( Espoon kuvataidekoulu ) kan barn och unga studera bildkonst .
studierna är avgiftsbelagda .
vid Esbo musikinstitut ( Espoon musiikkiopisto ) kan barn och vuxna studera musik .
Läs mer : andra studiemöjligheter
linkkiEsbo stad :
Arbetarinstitutetfinska _ svenska _ engelska
linkkiEsbo biIdkonstskola :
bildkonst för barn och ungafinska _ svenska _ engelska
linkkiEsbo musikinstitut :
Musikundervisning för barn och vuxnafinska _ engelska
dagvård
förskoleundervisning
grundläggande utbildning
hemspråksundervisning för invandrare
yrkesutbildning
gymnasium
stöd och handledning för unga
Högskoleutbildning
andra studiemöjligheter
dagvård
i Esbo finns både kommunala och privata daghem .
i Esbo finns dessutom familjedagvårdare .
dagvård fås på finska och på svenska .
Ansök om dagvårdsplats minst fyra månader innan barnet ska börja i dagvården .
om du till exempel oväntat får arbete eller en studieplats kan du ansöka om vårdplats senare .
när du ansöker om vårdplats ska du fylla i en ansökningsblankett .
du kan också söka dagvårdsplats via Internet .
familjer som bor i Esbo kan också söka dagvårdsplats till sitt barn i Helsingfors , Vanda eller Grankulla .
du ska ändå lämna in din ansökan i Esbo .
mer information får du via tjänsten Helsingforsregionen.fi .
Läs mer : småbarnspedagogik
linkkiEsbo stad :
dagvårdfinska _ svenska _ engelska
linkkiEsbo stad :
ansökan om dagvårdsplatsfinska _ engelska
linkkiEsbo stad :
Servicepunktfinska _ svenska _ engelska
linkkiEsbo stad :
Dagvårdens samanvändningsområdefinska _ svenska _ engelska
förskoleundervisning
i Esbo anordnas förskoleundervisningen ( esiopetus ) i daghemmen .
förskoleundervisning ges på finska och på svenska .
till förskoleundervisningen anmäler man sig via Esbo stads webbplats .
förskoleundervisningen börjar i augusti .
ansökningstiden är vanligtvis i januari .
i frågor kring barndagvård och förskoleundervisning kan du också kontakta daghemsföreståndarna eller stadens chef för småbarnsfostran ( varhaiskasvatuspäällikkö ) .
kontaktuppgifterna finns på stadens webbplats .
Läs mer : förskoleundervisning .
linkkiEsbo stad :
förskoleundervisningfinska _ svenska _ engelska
linkkiEsbo stad :
ansökan till förskoleundervisningfinska _ engelska
grundläggande utbildning
i Esbo finns finskspråkiga och svenskspråkiga grundskolor ( peruskoulu ) .
undervisning kan även fås på engelska .
skolan börjar vanligtvis det året då barnet fyller sju år .
anmälan till grundskolan ska göras på förhand .
Anmälningstiden är vanligtvis i januari .
på stadens webbplats hittar du kontaktuppgifterna till skolorna och mer information om anmälan .
om du har frågor om den grundläggande utbildningen kan du kontakta Resultatenheten för den finskspråkiga undervisningen ( Suomenkielisen opetuksen tulosyksikkö ) .
Resultatenheten för den finskspråkiga undervisningen
Kamrersvägen 3 B
tfn ( 09 ) 816.52044 och ( 09 ) 816.52043
grundläggande utbildning .
linkkiEsbo stad :
grundläggande utbildningfinska _ svenska _ engelska
linkkiEsbo stad :
anmälan till skolanfinska _ svenska _ engelska
linkkiEsbo stad :
Espoo International Schoolfinska _ engelska
internationella skolor i huvudstadsregionenfinska
linkkiExpatFinland.fi :
internationella skolor i huvudstadsregionenengelska
linkkiEsbo stad :
Eftermiddagsverksamhetfinska _ engelska
hemspråksundervisning för invandrare
barn med invandrarbakgrund och barn från tvåspråkiga familjer kan få hemspråksundervisning ( oman äidinkielen opetus ) om tillräckligt många barn anmäler sig till gruppen för det egna språket .
undervisning ges två timmar i veckan .
anmälan till hemspråksundervisning görs varje år i mars .
mer information hittar du på Esbo stads webbplats .
linkkiEsbo stad :
förberedande undervisning för barn i förskoleåldern ( pdf , 100 kb ) finska _ engelska _ ryska _ estniska _ somaliska _ kinesiska _ arabiska _ kurdiska _ albanska
linkkiEsbo stad :
förberedande undervisning för barn i förskoleåldernfinska _ engelska
linkkiEsbo stad :
hemspråksundervisningfinska _ engelska
yrkesutbildning
på Omnia kan man studera många olika yrken .
på Omnia ordnas för invandrare utbildning som förbereder dem på yrkesutbildning .
den förberedande utbildningen är avsedd för unga och vuxna , som är intresserade av yrkesstudier och vill förbättra sina kunskaper i finska ..
Esbobor kan också ansöka till yrkesskolorna i Helsingfors och Vanda .
Läs mer : yrkesutbildning
yrkesutbildningfinska _ engelska
linkkiEsbo stad :
Yrkesläroanstalterfinska _ engelska
Yrkesläroanstalterfinska _ svenska _ engelska
linkkiVanda stad :
yrkesutbildningfinska _ svenska
gymnasium
i Esbo finns elva finskspråkiga och ett svenskspråkigt gymnasium ( lukio ) .
i två av gymnasierna i Esbo finns en engelskspråkig IB @-@ linje .
ungdomar från Esbo kan också söka till gymnasier i andra städer .
i Esbo finns ett vuxengymnasium ( aikuislukio ) där vuxna kan avlägga gymnasie- och studentexamen .
på gymnasiet kan man även höja vitsorden i sitt avgångsbetyg eller studera enskilda ämnen .
invandrarungdomar kan dessutom studera finska och avlägga grundskolans lärokurs .
i gymnasiet Leppävaaran lukio ordnas för invandrare och utlänningar utbildning som förbereder dem på gymnasiet .
utbildningen är avsedd för unga som vill studera på gymnasiet , men vars språkkunskaper inte är tillräckliga för gymnasiestudier .
Läs mer : gymnasium
linkkiEsbo stad :
Gymnasierfinska _ svenska _ engelska
linkkiEsbo stad :
Vuxengymnasietfinska
linkkiEsbo stad :
Gymnasieförberedande utbildning för invandrarefinska _ engelska
linkkiEsbo vuxengymnasium Omnia :
grundläggande utbildning för invandrarefinska
om du är under 30 år gammal kan du få råd och handledning via Ohjaamo @-@ tjänsten .
Ohjaamos personal hjälper dig om du inte har ett arbete eller en studieplats .
du kan även fråga om andra saker , som till exempel boende eller ekonomiska frågor .
kontaktuppgifter :
Fågelbergavägen 2 A
Puh . 040.126.7513
linkkiEsbo stad :
Ohjaamofinska _ svenska _ engelska
Högskoleutbildning
i Esbo finns tre högskolor :
yrkeshögskolan Laurea
yrkeshögskolan Metropolia .
vid högskolorna kan du avlägga högskoleexamen .
mer information finns på Aalto @-@ universitetets , Laureas och Metropolias webbplatser .
också i Helsingfors finns det universitet och yrkeshögskolor där man kan studera inom många områden .
mer information hittar du på Helsingfors stads webbplats .
Läs mer : yrkeshögskolor
universitet inom teknik , konst och ekonomifinska _ svenska _ engelska
yrkeshögskolafinska _ engelska
linkkiMetropolia :
yrkeshögskolafinska _ engelska
Högskolorfinska
andra studiemöjligheter
vid Esbo arbetarinstitut ( Espoon työväenopisto ) kan du studera till exempel språk , handarbete och matlagning eller delta i ledd motion .
kurserna är avgiftsbelagda . kurser anordnas både dagtid och kvällstid .
vid arbetarinstitutet kan vem som helst studera .
vid Esbo bildkonstskola ( Espoon kuvataidekoulu ) kan barn och unga studera bildkonst .
studierna är avgiftsbelagda .
vid Esbo musikinstitut ( Espoon musiikkiopisto ) kan barn och vuxna studera musik .
Läs mer : studier som hobby
linkkiEsbo stad :
Arbetarinstitutetfinska _ svenska _ engelska
linkkiEsbo biIdkonstskola :
bildkonst för barn och ungafinska _ svenska _ engelska
linkkiEsbo musikinstitut :
Musikundervisning för barn och vuxnafinska _ engelska
hyresbostad
Ägarbostad
Bostadsrättsbostad
Delägarbostad
tillfälligt boende
boende i en krissituation
Stöd- och serviceboende
Bostadslöshet
avfallshantering och återvinning
hyresbostad
i Esbo och huvudstadsregionen är hyrorna ofta högre än i resten av Finland .
det kan vara svårt att hitta en bostad med lämplig hyra .
det lönar sig att avsätta tid för bostadssökandet och undersöka olika alternativ .
privata hyresbostäder
hos en privat hyresvärd kan det gå snabbt att få en bostad , men hyran kan vara högre än i stadens hyresbostäder .
du kan söka privata hyresbostäder i Esbo via hyresvärdarnas webbplatser :
Sökning av hyresbostäderfinska
Sökning av hyresbostäderfinska _ engelska
hyresbostäder för ungafinska _ engelska
hyresbostäder för ungafinska _ engelska
om du är studerande kan du få en hyresbostad för studerande i Esbo .
hyresbostäder för studerande erbjuds av Helsingforsregionens studentbostadsstiftelse HOAS och Aalto @-@ universitets studentkår AUS .
linkkiHOAS :
hyresbostäder för studerandefinska _ svenska _ engelska
hyresbostäder för studerandefinska _ svenska _ engelska
stadens hyresbostäder
stadens hyresbostäder är ofta billigare än bostäder som man hyr av företag eller privatpersoner .
det är dock många som ansöker om stadens bostäder och endast en liten del av de sökande får en bostad .
Störst är bristen på små bostäder .
stadens hyresbostäder förvaltas av Espoon Asunnot Oy ( Espoon Asunnot Oy ) .
om du vill ansöka om en hyresbostad , fyll i en ansökningsblankett för hyresbostad på Espoon Asunnot Oy:s webbplats .
du kan även fylla i ansökningsblanketten på Espoon Asunnot Oy:s kontor .
du kan också få blanketten hemskickad per post .
dina möjligheter att få en bostad påverkas av ditt bostadsbehov och dina tillgångar och inkomster .
för att kunna ansöka om en hyresbostad hos staden , måste du ha uppehållstillstånd för minst ett år .
tfn ( 09 ) 816.5800
ansökan är giltig i tre månader .
efter det måste du förnya din ansökan om du fortfarande letar efter bostad .
Läs mer : hyresbostad
linkkiEsbo bostäder Ab :
ansökan om hyresbostad i stadenfinska _ engelska
linkkiEsbo stad :
stadens hyresbostäderfinska _ svenska _ engelska
linkkiEsbo stad :
Seniorbostäderfinska _ svenska
Ägarbostad
på internet finns många bostadsförsäljningsannonser . bostäderna i Esbo är tämligen dyra .
information om köp av bostad hittar du på InfoFinlands sida Ägarbostad .
Bostadsrättsbostad
om du ansöker om en bostadsrättsbostad , behöver du ett ordningsnummer . du ansöker om ordningsnumret vid Esbo eller Helsingfors stad .
Läs mer : Bostadsrättsbostad .
linkkiEsbo stad :
Bostadsrättsbostäderfinska _ svenska _ engelska
Delägarbostad
asuntosäätiö har delägarbostäder i Esbo .
mer information hittar du på Asuntosäätiös webbplats .
Läs mer : Delägarbostad .
Delägarbostadfinska
tillfälligt boende
i Esbo finns många olika hotell där man kan bo tillfälligt .
Läs mer : tillfälligt boende .
linkkiVisitEspoo.fi :
Hotellfinska _ svenska _ engelska _ ryska _ kinesiska
brand eller vattenskada
om din bostad har skadats till exempel till följd av brand eller vattenskada kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna .
kontakta ditt försäkringsbolag direkt när skadan har inträffat .
våld i hemmet
om någon i din familj utövar våld mot dig eller hotar dig med våld , kan du kontakta tjänsten Omatila ( Omatila ) .
Omatila ordnar vid behov boende för dig och dina barn .
Omatila @-@ tjänsten
Kamrersvägen 6 A
tfn 043.825.0535
öppet
Lördag @-@ söndag kl . 9 @-@ 16
social- och krisjouren 24 h
tfn 09.816.42439
linkkiEsbo stad :
hjälp till offer för familjevåldfinska _ svenska _ engelska
om du är ung och har problem hemma , kan du kontakta Finlands Röda Kors De ungas skyddshus .
skyddshuset finns i Alberga .
de ungas skyddshus
tfn ( 09 ) 8195.5360
linkkiFinlands Röda Kors :
de ungas skyddshusfinska _ svenska _ engelska
Stöd- och serviceboende
en del människor , till exempel åldringar och handikappade , har svårt att klara av de dagliga sysslorna utan hjälp .
personer som har sin hemkommun i Esbo kan få hemvårdens stödtjänster av Esbo stad , till exempel måltidstjänster eller färdtjänst .
dessa tjänster hjälper människorna att klara sig bättre hemma .
åldringar och handikappade som inte klarar av att bo självständigt , kan bo i ett servicehus eller på en vårdinrättning .
Läs mer : Stöd- och serviceboende
om du har frågor kring stödtjänsterna för handikappade , kontakta handikappservicen vid Esbo stad .
Esbo stads handikappservice
telefonrådgivning : ( 09 ) 816.45285
linkkiEsbo stad :
stödtjänster för handikappadefinska _ svenska _ engelska
om du har frågor kring stödtjänsterna för äldre , kontakta Esbo stads rådgivning för seniorer .
Esbo stads rådgivning för seniorer
tfn ( 09 ) 816.33333
linkkiEsbo stad :
stödtjänster för äldrefinska _ svenska _ engelska
linkkiEsbo stad :
information om hemvårdens stödtjänsterfinska _ svenska
linkkiEsbo stad :
information om boende i servicehusfinska _ svenska
Bostadslöshet
om du blir bostadslös , kontakta Esbo stads verksamhetsställe för vuxensocialarbete .
linkkiEsbo stad :
kontaktuppgifter till vuxensocialarbetetfinska _ svenska _ engelska
om läget är akut , kan du även kontakta social- och krisjouren i Esbo .
social- och krisjouren
Jorvs sjukhus
Åbovägen 150
tfn ( 09 ) 816.42439
linkkiEsbo stad :
social- och krisjourenfinska _ svenska _ engelska
Läs mer : Bostadslöshet
avfallshantering och återvinning
