Grundläggande information
Historia
Trafik
Religion
Beslutsfattande och påverkan
Grundläggande information
Karleby finns i Mellersta Österbotten invid Bottniska viken.
Karleby stad är grundad 1620 och hette då Gamlakarleby.
Senare blev Kokkola stadens finska namn.
Vid Karleby centrum finns en av landets mest omfattande historiska trästadshelheter.
Stadsplanen är från 1650-talet.
Den omfattar 12 kvarter med hundratals trähus och gårdsbyggnader.
De äldsta av dessa är från 1600-talet.
Karleby är en kulturstad med mycket att se och uppleva.
Karleby hamn ligger i stadsdelen Yxpila och är en av Finlands mest trafikerade godshamnar.
Grunden för näringslivet i Karleby är den internationella storindustrin.
I Karleby är den kemiska industrin och industri i anslutning till denna särskilt viktig.
Karleby är även en betydande handelsstad.
Information om Karlebyfinska _ svenska _ engelska
Historia
Redan under medeltiden fanns det hamn, båtbygge och handelsplats i Karleby.
Landhöjningen har varit en central faktor i Karlebys historia.
Den har format omgivningen i hög grad och bland annat påverkat utvecklingen av hamnverksamheten och handeln.
Handel bedrevs längs med Bottniska vikens kust och jordbruk, jakt, fiske och sälfångst var även viktiga näringar.
Exporten av tjära, som blev mycket viktig för Karlebys historia, inleddes redan på 1500-talet.
Den sjunde september 1620 undertecknade Sveriges kung Gustav II Adolf en handling som gav den lilla jordbruks- och fiskebyn vid Ristrand status som stad.
Dagens stadssund var då en smal havsvik som sträckte sig ända till Kyrkbacken.
Sakta men säkert blev Karleby en viktig stad för sjöfart och skeppsbygge.
Skeppsvarv fanns bland annat i Kaustarviken, Svartskär och Soldatskär.
Inledningsvis seglade man endast till Åbo och Stockholm, eftersom Karleby som s.k. uppstad inte fick bedriva utrikeshandel.
År 1765 erhöll staden stapelrättigheter, dvs. rätt till fri utrikeshandel, främst tack vare den aktiva kyrkoherden och lantdagsmannen Anders Chydenius.
Karleby blev snabbt en förmögen stad i början av 1800-talet tack vare just handeln med tjära och rederiverksamheten.
Stadens borgare köpte tjära av bönder och exporterade den, ofta till hamnar vid Medelhavet och i England.
Karleby handelsflotta var under perioder Finlands största.
Den snabba ekonomiska utvecklingen avtog i mitten av 1800-talet, men tog ny fart i slutet av århundradet tack vare industrialiseringen.
Karleby blev en viktig industristad främst tack vare läder- och metallindustrin.
Karlebys historiafinska _ svenska _ engelska
Trafik
Karleby har goda trafikförbindelser.
Via Karleby löper riksväg 8 och 13.
Järnvägsstationen finns i stadens centrum.
Restiden med tåg till Helsingfors är cirka fyra timmar.
Flygplatsen finns i Kronoby på endast 22 kilometers avstånd från Karleby centrum.
Stadsborna erbjuds även ett tryggt, omfattande, fungerande och trivsamt nätverk för den lätta trafiken.
Karleby har satsat på att förbättra förhållandena för cyklister.
Lokalbussarna trafikerar de olika delarna av staden på vardagar.
Läs mer: Trafik.
Gator och trafikfinska _ svenska
Kollektivtrafikfinska _ svenska
linkkiVR:
Tågtidtabellerfinska _ svenska _ engelska _ ryska
Busstidtabellerfinska _ svenska _ engelska
Flyg från Karleby-Jakobstad flygplatsfinska _ svenska _ engelska
Religion
I Karleby finns flera olika religiösa samfund.
I tjänsten Uskonnot Suomessa (Religioner i Finland) finns information om religiösa samfund enligt ort.
Den evangelisk-lutherska kyrkan har fyra finskspråkiga församlingar och en svenskspråkig församling i Karleby.
Läs mer på Karleby kyrkliga samfällighets webbplats.
I Karleby finns en ortodox kyrka.
Mer information om den ortodoxa församlingens verksamhet i Karleby finns på Vasa ortodoxa församlings webbplats.
Läs mer: Kulturer och religioner i Finland.
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiVasa ortodoxa församling:
Vasa ortodoxa församlingfinska _ engelska _ ryska
Beslutsfattande och påverkan
Den högsta beslutsfattande makten i Karleby stad innehas av stadsfullmäktige.
Fullmäktigeledamöterna och deras suppleanter väljs vid kommunalval vart fjärde år.
På stadens webbplats finns information om stadsfullmäktige och dess beslut.
Invånarna kan påverka stadens beslutsfattande redan då beslut bereds.
Information om olika sätt att delta och påverka finns på stadens webbplats.
Kommunens invånare har enligt kommunallagen rätt att lämna in motioner till kommunen i ärenden som gäller dess verksamhet.
I Karleby finns ungdomsfullmäktige, äldre- och handikappråd samt ett råd för kulturell mångfald.
Läs mer: Finlands förvaltning, Val och röstning i Finland
Beslutsfattandefinska _ svenska _ engelska
Grundläggande information
Historia
Trafik
Religion
Beslutsfattande och påverkan
Grundläggande information
Karleby finns i Mellersta Österbotten invid Bottniska viken.
Karleby stad är grundad 1620 och hette då Gamlakarleby.
Senare blev Kokkola stadens finska namn.
Vid Karleby centrum finns en av landets mest omfattande historiska trästadshelheter.
Stadsplanen är från 1650-talet.
Den omfattar 12 kvarter med hundratals trähus och gårdsbyggnader.
De äldsta av dessa är från 1600-talet.
Karleby är en kulturstad med mycket att se och uppleva.
Karleby hamn ligger i stadsdelen Yxpila och är en av Finlands mest trafikerade godshamnar.
Grunden för näringslivet i Karleby är den internationella storindustrin.
I Karleby är den kemiska industrin och industri i anslutning till denna särskilt viktig.
Karleby är även en betydande handelsstad.
Information om Karlebyfinska _ svenska _ engelska
Historia
Redan under medeltiden fanns det hamn, båtbygge och handelsplats i Karleby.
Landhöjningen har varit en central faktor i Karlebys historia.
Den har format omgivningen i hög grad och bland annat påverkat utvecklingen av hamnverksamheten och handeln.
Handel bedrevs längs med Bottniska vikens kust och jordbruk, jakt, fiske och sälfångst var även viktiga näringar.
Exporten av tjära, som blev mycket viktig för Karlebys historia, inleddes redan på 1500-talet.
Den sjunde september 1620 undertecknade Sveriges kung Gustav II Adolf en handling som gav den lilla jordbruks- och fiskebyn vid Ristrand status som stad.
Dagens stadssund var då en smal havsvik som sträckte sig ända till Kyrkbacken.
Sakta men säkert blev Karleby en viktig stad för sjöfart och skeppsbygge.
Skeppsvarv fanns bland annat i Kaustarviken, Svartskär och Soldatskär.
Inledningsvis seglade man endast till Åbo och Stockholm, eftersom Karleby som s.k. uppstad inte fick bedriva utrikeshandel.
År 1765 erhöll staden stapelrättigheter, dvs. rätt till fri utrikeshandel, främst tack vare den aktiva kyrkoherden och lantdagsmannen Anders Chydenius.
Karleby blev snabbt en förmögen stad i början av 1800-talet tack vare just handeln med tjära och rederiverksamheten.
Stadens borgare köpte tjära av bönder och exporterade den, ofta till hamnar vid Medelhavet och i England.
Karleby handelsflotta var under perioder Finlands största.
Den snabba ekonomiska utvecklingen avtog i mitten av 1800-talet, men tog ny fart i slutet av århundradet tack vare industrialiseringen.
Karleby blev en viktig industristad främst tack vare läder- och metallindustrin.
Karlebys historiafinska _ svenska _ engelska
Trafik
Karleby har goda trafikförbindelser.
Via Karleby löper riksväg 8 och 13.
Järnvägsstationen finns i stadens centrum.
Restiden med tåg till Helsingfors är cirka fyra timmar.
Flygplatsen finns i Kronoby på endast 22 kilometers avstånd från Karleby centrum.
Stadsborna erbjuds även ett tryggt, omfattande, fungerande och trivsamt nätverk för den lätta trafiken.
Karleby har satsat på att förbättra förhållandena för cyklister.
Lokalbussarna trafikerar de olika delarna av staden på vardagar.
Läs mer: Trafik.
Gator och trafikfinska _ svenska
Kollektivtrafikfinska _ svenska
linkkiVR:
Tågtidtabellerfinska _ svenska _ engelska _ ryska
Busstidtabellerfinska _ svenska _ engelska
Flyg från Karleby-Jakobstad flygplatsfinska _ svenska _ engelska
Religion
I Karleby finns flera olika religiösa samfund.
I tjänsten Uskonnot Suomessa (Religioner i Finland) finns information om religiösa samfund enligt ort.
Den evangelisk-lutherska kyrkan har fyra finskspråkiga församlingar och en svenskspråkig församling i Karleby.
Läs mer på Karleby kyrkliga samfällighets webbplats.
I Karleby finns en ortodox kyrka.
Mer information om den ortodoxa församlingens verksamhet i Karleby finns på Vasa ortodoxa församlings webbplats.
Läs mer: Kulturer och religioner i Finland.
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiVasa ortodoxa församling:
Vasa ortodoxa församlingfinska _ engelska _ ryska
Beslutsfattande och påverkan
Den högsta beslutsfattande makten i Karleby stad innehas av stadsfullmäktige.
Fullmäktigeledamöterna och deras suppleanter väljs vid kommunalval vart fjärde år.
På stadens webbplats finns information om stadsfullmäktige och dess beslut.
Invånarna kan påverka stadens beslutsfattande redan då beslut bereds.
Information om olika sätt att delta och påverka finns på stadens webbplats.
Kommunens invånare har enligt kommunallagen rätt att lämna in motioner till kommunen i ärenden som gäller dess verksamhet.
I Karleby finns ungdomsfullmäktige, äldre- och handikappråd samt ett råd för kulturell mångfald.
Läs mer: Finlands förvaltning, Val och röstning i Finland
Beslutsfattandefinska _ svenska _ engelska
Grundläggande information
Historia
Trafik
Religion
Beslutsfattande och påverkan
Grundläggande information
Karleby finns i Mellersta Österbotten invid Bottniska viken.
Karleby stad är grundad 1620 och hette då Gamlakarleby.
Senare blev Kokkola stadens finska namn.
Vid Karleby centrum finns en av landets mest omfattande historiska trästadshelheter.
Stadsplanen är från 1650-talet.
Den omfattar 12 kvarter med hundratals trähus och gårdsbyggnader.
De äldsta av dessa är från 1600-talet.
Karleby är en kulturstad med mycket att se och uppleva.
Karleby hamn ligger i stadsdelen Yxpila och är en av Finlands mest trafikerade godshamnar.
Grunden för näringslivet i Karleby är den internationella storindustrin.
I Karleby är den kemiska industrin och industri i anslutning till denna särskilt viktig.
Karleby är även en betydande handelsstad.
Information om Karlebyfinska _ svenska _ engelska
Historia
Redan under medeltiden fanns det hamn, båtbygge och handelsplats i Karleby.
Landhöjningen har varit en central faktor i Karlebys historia.
Den har format omgivningen i hög grad och bland annat påverkat utvecklingen av hamnverksamheten och handeln.
Handel bedrevs längs med Bottniska vikens kust och jordbruk, jakt, fiske och sälfångst var även viktiga näringar.
Exporten av tjära, som blev mycket viktig för Karlebys historia, inleddes redan på 1500-talet.
Den sjunde september 1620 undertecknade Sveriges kung Gustav II Adolf en handling som gav den lilla jordbruks- och fiskebyn vid Ristrand status som stad.
Dagens stadssund var då en smal havsvik som sträckte sig ända till Kyrkbacken.
Sakta men säkert blev Karleby en viktig stad för sjöfart och skeppsbygge.
Skeppsvarv fanns bland annat i Kaustarviken, Svartskär och Soldatskär.
Inledningsvis seglade man endast till Åbo och Stockholm, eftersom Karleby som s.k. uppstad inte fick bedriva utrikeshandel.
År 1765 erhöll staden stapelrättigheter, dvs. rätt till fri utrikeshandel, främst tack vare den aktiva kyrkoherden och lantdagsmannen Anders Chydenius.
Karleby blev snabbt en förmögen stad i början av 1800-talet tack vare just handeln med tjära och rederiverksamheten.
Stadens borgare köpte tjära av bönder och exporterade den, ofta till hamnar vid Medelhavet och i England.
Karleby handelsflotta var under perioder Finlands största.
Den snabba ekonomiska utvecklingen avtog i mitten av 1800-talet, men tog ny fart i slutet av århundradet tack vare industrialiseringen.
Karleby blev en viktig industristad främst tack vare läder- och metallindustrin.
Karlebys historiafinska _ svenska _ engelska
Trafik
Karleby har goda trafikförbindelser.
Via Karleby löper riksväg 8 och 13.
Järnvägsstationen finns i stadens centrum.
Restiden med tåg till Helsingfors är cirka fyra timmar.
Flygplatsen finns i Kronoby på endast 22 kilometers avstånd från Karleby centrum.
Stadsborna erbjuds även ett tryggt, omfattande, fungerande och trivsamt nätverk för den lätta trafiken.
Karleby har satsat på att förbättra förhållandena för cyklister.
Lokalbussarna trafikerar de olika delarna av staden på vardagar.
Läs mer: Trafik.
Gator och trafikfinska _ svenska
Kollektivtrafikfinska _ svenska
linkkiVR:
Tågtidtabellerfinska _ svenska _ engelska _ ryska
Busstidtabellerfinska _ svenska _ engelska
Flyg från Karleby-Jakobstad flygplatsfinska _ svenska _ engelska
Religion
I Karleby finns flera olika religiösa samfund.
I tjänsten Uskonnot Suomessa (Religioner i Finland) finns information om religiösa samfund enligt ort.
Den evangelisk-lutherska kyrkan har fyra finskspråkiga församlingar och en svenskspråkig församling i Karleby.
Läs mer på Karleby kyrkliga samfällighets webbplats.
I Karleby finns en ortodox kyrka.
Mer information om den ortodoxa församlingens verksamhet i Karleby finns på Vasa ortodoxa församlings webbplats.
Läs mer: Kulturer och religioner i Finland.
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiVasa ortodoxa församling:
Vasa ortodoxa församlingfinska _ engelska _ ryska
Beslutsfattande och påverkan
Den högsta beslutsfattande makten i Karleby stad innehas av stadsfullmäktige.
Fullmäktigeledamöterna och deras suppleanter väljs vid kommunalval vart fjärde år.
På stadens webbplats finns information om stadsfullmäktige och dess beslut.
Invånarna kan påverka stadens beslutsfattande redan då beslut bereds.
Information om olika sätt att delta och påverka finns på stadens webbplats.
Kommunens invånare har enligt kommunallagen rätt att lämna in motioner till kommunen i ärenden som gäller dess verksamhet.
I Karleby finns ungdomsfullmäktige, äldre- och handikappråd samt ett råd för kulturell mångfald.
Läs mer: Finlands förvaltning, Val och röstning i Finland
Beslutsfattandefinska _ svenska _ engelska
Detta innehåll finns inte på det språk som du har valt.
Välj något annat språk.
Finska
Detta innehåll finns inte på det språk som du har valt.
Välj något annat språk.
Finska
Detta innehåll finns inte på det språk som du har valt.
Välj något annat språk.
Finska
Bibliotek
Motion
Att röra sig i naturen
Teater och film
Museer
Hobbyer för barn och unga
Föreningar
Karleby är en gammal sjöstad som erbjuder mångsidiga möjligheter för utfärder och friluftsliv.
Personer ntresserad av friluftsliv bör läsa mer om allemansrätten under rubriken ”Att röra sig i naturen” i denna tjänst.
Flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet.
Föreningar och organisationer samt hobbygrupper och kommunala institut erbjuder kurser i idrott och kultur samt bl.a. språk och hantverk.
I Snellman-salen och i stadens övriga kulturlokaler erbjuds kulturevenemang av varierande slag.
Årliga evenemang i Karleby är bland annat Veneziansk afton i slutet av sommaren, Kokkola Cup för fotbollsjuniorer, Stadsfestivalen Karleby sommarveckor, Lochteå kyrkomusikfest samt Vinterdans i Karleby och festivalen Karleby Vinterharmonika.
Mer information om fritidstjänsterna i Karleby finns på Karleby stads webbplats.
På stadens webbplats finns även en länk till Evenemangskalendern med daglig information om stadens kultur- och motionsevenemang.
Läs mer: Fritid.
Evenemangskalenderfinska
Kulturtjänsterfinska _ svenska _ engelska
Idrottstjänsterfinska _ svenska _ engelska
Bibliotek
Karleby stadsbibliotek finns i stadens centrum.
Närbiblioteken finns i Björkhagen, Kelviå, Lochteå samt Ullava kyrkby och Rahkonen.
Information om bibliotekets öppettider och tjänster finns på dess webbplats.
Biblioteket finns även på nätet.
Där kan kunderna bläddra i bibliotekets samlingar, reservera material, förnya sina lån, beställa fjärrlån och låna e-böcker under alla tider på dygnet.
Tack vare det effektiva biblioteksnätverket i Finland är nästan alla finländska biblioteks samlingar tillgängliga för bibliotekskunderna i Karleby.
Karleby stadsbibliotek/huvudbiblioteket
Storgatan 3, 67100 Karleby
Telefon: 040 806 5124, 040 806 5133
Läs mer: Bibliotek.
Bibliotekstjänsterfinska _ svenska _ engelska
Motion
I Karleby finns mångsidiga motionsmöjligheter året runt.
Staden anordnar ledda aktiviteter i Simcentret VesiVeijari och motionshallarna.
Dessutom finns det gym av flera olika slag.
Gym anpassade för äldre finns i Furuåsens aktivitetscenter och Kuusikumpu servicehus.
Staden underhåller cykelvägar, motionsrutter, joggingbanor, skidspår, badstränder, bollplaner och skridskobanor samt platser för närmotion.
I Karlebynejdens instituts nättjänst finns information om institutets mångsidiga motionsutbud.
I Karleby finns nära på hundra idrottsföreningar för olika grenar samt föreningar som arrangerar övrig motion.
Mer information om motionsmöjligheter i Karleby finns på Karleby stads webbplats.
Läs mer:
Motion.
Idrottstjänsterfinska _ svenska _ engelska
Motionsplatserfinska _ svenska
Gym för äldrefinska
Karlebynejdens institutfinska _ svenska
Att röra sig i naturen
Att röra sig i naturen är en traditionell och populär form av avkoppling för finländarna under alla årstider.
I Finland kan man med stöd av allemansrätten plocka bär och svamp i skogen och röra sig till fots, med cykel eller skidor vintertid.
Det är inte tillåtet att beträda folks gårdar utan lov.
För fiske krävs fiskelov, med undantag för mete och pilkning.
Även jakt fordrar jakttillstånd.
Allemansrätten ger inte rätt att skräpa ner i naturen, skada träd eller växter, störa eller skada fågelbon eller fågelungar, köra motorfordon utan markägarens tillstånd eller bygga ens tillfälliga byggen.
Mer information om motionsrutterna, rastplatser, möjligheter till fiske och båtliv samt exempelvis fågeltorn i Karleby finns på stadens webbplats.
Rutterna för camping, paddling, vandring, cykling och övriga rutter i Karleby finns i karttjänsten på nätet.
I karttjänsten visas även var största delen av motionsplatserna finns.
Du kan köpa friluftskartor över Karleby hos Karleby Turism: Salutorget 5, 67100 Karleby.
Läs mer: Att röra sig i naturen.
linkkiMiljöförvaltningen:
Allemansrättenfinska _ svenska _ engelska _ ryska
Motionskarta över Karlebyfinska _ svenska
Motionsrutter i Karlebyfinska _ svenska
Teater och film
Karleby är en teaterstad med långa anor, som erbjuder scenkonst på hög nivå framförd av både proffs och amatörer.
Karleby stadsteater finns i det stämningsfulla Vartiolinna (Torggatan 48).
Du kan läsa mer om amatörteatrarnas verksamhet på deras webbplats och i evenemangskalendern.
I Karleby finns biografen Bio Rex, vars två salar använder digital- och 3D-teknik.
Bio Rex program finns under länken här intill.
Läs mer: Teater och film.
Stadsteaternfinska
Biograffinska
Teater och danskonst i Karlebyfinska _ svenska _ engelska
Evenemangskalenderfinska
Museer
I hjärtat av staden, i det anrika Rooska gården, finns K.H.Renlunds museum.
Karleby stad grundade museet 1909 utgående från en testamentsgåva av affärsmannen Karl Herman Renlund (1850–1908) .
På museet finns Renlunds samling av finländsk konst från guldåldern och tillfälliga utställningar i en kulturhistorisk miljö.
Även i museikvarterens övriga byggnader finns utställningar om stadens kulturhistoria och utställningar med ITE-konst.
På K.H.Renlunds museums webbplats finns mer information om museets tjänster, utställningar samt aktuell verksamhet.
Utöver K.H.Renlunds museum lönar det sig att besöka det naturhistoriska museet Kieppi (Kieppi är stängt tills vidare på grund av brand) samt de många hembygdsmuseerna och övriga de historiska resmålen i regionen.
Exempelvis i Konst-Vionoja-centret presenteras konstnären Veikko Vionojas verk.
I Kelviå, ca 10 km norrut från Karleby, finns Toivonen djurpark och drängmuseum.
Mer information om dessa museer finns under länkarna här intill.
Läs mer: Museer.
Museer och traditionsarbetefinska _ svenska _ engelska
K.H. Renlunds museum - Mellersta Österbottens landskapsmuseumfinska _ svenska _ engelska
Kieppi, Karleby naturvetenskapliga museumfinska _ svenska _ engelska
linkkiToivonens djurpark och drängmuseum :
Toivonens djurpark och drängmuseum finska _ svenska _ engelska
Konst Vionojafinska
Hobbyer för barn och unga
Flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet.
Flera olika föreningar samt kommunala institut ger unga möjlighet att studera idrott och kultur samt bl.a. språk och hantverk.
Barn och unga kan delta i grundläggande undervisning i musik, dans, bildkonst och hantverk.
Dessutom erbjuder stadens ungdomstjänster en rockskola.
Stadens ungdomstjänster driver sju ungdomsgårdar runt om i Karleby.
De rusmedels- och rökfria ungdomslokalerna erbjuder handledd verksamhet för barn i årskurserna 3–6 och unga i åldern 13–17 år i olika delar av Karleby.
Information om hobbyverksamheter för barn och unga finns på stadens webbplats.
Rådgivningen vid Ungdomsgården Vinge ger aktuell information om bl.a. internationalisering, studier, arbetsliv, hälsa, hobbyverksamhet och boende.
Karlebynejdens institut erbjuder barn och unga olika former av hobbyverksamhet, exempelvis i konstämnen och musik.
Kontrollera vilka kurser som är aktuella i institutets webbtjänst.
Karleby evangelisk-lutherska församlingar erbjuder även hobbyverksamhet för barn och unga, såsom lekparksträffar, klubbar, musikverksamhet och läger.
Mer information om verksamheten finns på Karleby församlingssammanslutnings webbplats.
Ungdomsgården Vinge
67100 Karleby
Läs mer: Hobbyer för barn och unga.
Övrig undervisning i Karlebyfinska _ svenska
Ungdomstjänsterfinska _ svenska _ engelska
Karlebynejdens institutfinska _ svenska
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
Föreningar
Karleby har ett aktivt och mångsidigt föreningsliv för invånare i alla åldrar.
Läs mer: Föreningar.
Bibliotek
Motion
Att röra sig i naturen
Teater och film
Museer
Hobbyer för barn och unga
Föreningar
Karleby är en gammal sjöstad som erbjuder mångsidiga möjligheter för utfärder och friluftsliv.
Personer ntresserad av friluftsliv bör läsa mer om allemansrätten under rubriken ”Att röra sig i naturen” i denna tjänst.
Flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet.
Föreningar och organisationer samt hobbygrupper och kommunala institut erbjuder kurser i idrott och kultur samt bl.a. språk och hantverk.
I Snellman-salen och i stadens övriga kulturlokaler erbjuds kulturevenemang av varierande slag.
Årliga evenemang i Karleby är bland annat Veneziansk afton i slutet av sommaren, Kokkola Cup för fotbollsjuniorer, Stadsfestivalen Karleby sommarveckor, Lochteå kyrkomusikfest samt Vinterdans i Karleby och festivalen Karleby Vinterharmonika.
Mer information om fritidstjänsterna i Karleby finns på Karleby stads webbplats.
På stadens webbplats finns även en länk till Evenemangskalendern med daglig information om stadens kultur- och motionsevenemang.
Läs mer: Fritid.
Evenemangskalenderfinska
Kulturtjänsterfinska _ svenska _ engelska
Idrottstjänsterfinska _ svenska _ engelska
Bibliotek
Karleby stadsbibliotek finns i stadens centrum.
Närbiblioteken finns i Björkhagen, Kelviå, Lochteå samt Ullava kyrkby och Rahkonen.
Information om bibliotekets öppettider och tjänster finns på dess webbplats.
Biblioteket finns även på nätet.
Där kan kunderna bläddra i bibliotekets samlingar, reservera material, förnya sina lån, beställa fjärrlån och låna e-böcker under alla tider på dygnet.
Tack vare det effektiva biblioteksnätverket i Finland är nästan alla finländska biblioteks samlingar tillgängliga för bibliotekskunderna i Karleby.
Karleby stadsbibliotek/huvudbiblioteket
Storgatan 3, 67100 Karleby
Telefon: 040 806 5124, 040 806 5133
Läs mer: Bibliotek.
Bibliotekstjänsterfinska _ svenska _ engelska
Motion
I Karleby finns mångsidiga motionsmöjligheter året runt.
Staden anordnar ledda aktiviteter i Simcentret VesiVeijari och motionshallarna.
Dessutom finns det gym av flera olika slag.
Gym anpassade för äldre finns i Furuåsens aktivitetscenter och Kuusikumpu servicehus.
Staden underhåller cykelvägar, motionsrutter, joggingbanor, skidspår, badstränder, bollplaner och skridskobanor samt platser för närmotion.
I Karlebynejdens instituts nättjänst finns information om institutets mångsidiga motionsutbud.
I Karleby finns nära på hundra idrottsföreningar för olika grenar samt föreningar som arrangerar övrig motion.
Mer information om motionsmöjligheter i Karleby finns på Karleby stads webbplats.
Läs mer:
Motion.
Idrottstjänsterfinska _ svenska _ engelska
Motionsplatserfinska _ svenska
Gym för äldrefinska
Karlebynejdens institutfinska _ svenska
Att röra sig i naturen
Att röra sig i naturen är en traditionell och populär form av avkoppling för finländarna under alla årstider.
I Finland kan man med stöd av allemansrätten plocka bär och svamp i skogen och röra sig till fots, med cykel eller skidor vintertid.
Det är inte tillåtet att beträda folks gårdar utan lov.
För fiske krävs fiskelov, med undantag för mete och pilkning.
Även jakt fordrar jakttillstånd.
Allemansrätten ger inte rätt att skräpa ner i naturen, skada träd eller växter, störa eller skada fågelbon eller fågelungar, köra motorfordon utan markägarens tillstånd eller bygga ens tillfälliga byggen.
Mer information om motionsrutterna, rastplatser, möjligheter till fiske och båtliv samt exempelvis fågeltorn i Karleby finns på stadens webbplats.
Rutterna för camping, paddling, vandring, cykling och övriga rutter i Karleby finns i karttjänsten på nätet.
I karttjänsten visas även var största delen av motionsplatserna finns.
Du kan köpa friluftskartor över Karleby hos Karleby Turism: Salutorget 5, 67100 Karleby.
Läs mer: Att röra sig i naturen.
linkkiMiljöförvaltningen:
Allemansrättenfinska _ svenska _ engelska _ ryska
Motionskarta över Karlebyfinska _ svenska
Motionsrutter i Karlebyfinska _ svenska
Teater och film
Karleby är en teaterstad med långa anor, som erbjuder scenkonst på hög nivå framförd av både proffs och amatörer.
Karleby stadsteater finns i det stämningsfulla Vartiolinna (Torggatan 48).
Du kan läsa mer om amatörteatrarnas verksamhet på deras webbplats och i evenemangskalendern.
I Karleby finns biografen Bio Rex, vars två salar använder digital- och 3D-teknik.
Bio Rex program finns under länken här intill.
Läs mer: Teater och film.
Stadsteaternfinska
Biograffinska
Teater och danskonst i Karlebyfinska _ svenska _ engelska
Evenemangskalenderfinska
Museer
I hjärtat av staden, i det anrika Rooska gården, finns K.H.Renlunds museum.
Karleby stad grundade museet 1909 utgående från en testamentsgåva av affärsmannen Karl Herman Renlund (1850–1908) .
På museet finns Renlunds samling av finländsk konst från guldåldern och tillfälliga utställningar i en kulturhistorisk miljö.
Även i museikvarterens övriga byggnader finns utställningar om stadens kulturhistoria och utställningar med ITE-konst.
På K.H.Renlunds museums webbplats finns mer information om museets tjänster, utställningar samt aktuell verksamhet.
Utöver K.H.Renlunds museum lönar det sig att besöka det naturhistoriska museet Kieppi (Kieppi är stängt tills vidare på grund av brand) samt de många hembygdsmuseerna och övriga de historiska resmålen i regionen.
Exempelvis i Konst-Vionoja-centret presenteras konstnären Veikko Vionojas verk.
I Kelviå, ca 10 km norrut från Karleby, finns Toivonen djurpark och drängmuseum.
Mer information om dessa museer finns under länkarna här intill.
Läs mer: Museer.
Museer och traditionsarbetefinska _ svenska _ engelska
K.H. Renlunds museum - Mellersta Österbottens landskapsmuseumfinska _ svenska _ engelska
Kieppi, Karleby naturvetenskapliga museumfinska _ svenska _ engelska
linkkiToivonens djurpark och drängmuseum :
Toivonens djurpark och drängmuseum finska _ svenska _ engelska
Konst Vionojafinska
Hobbyer för barn och unga
Flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet.
Flera olika föreningar samt kommunala institut ger unga möjlighet att studera idrott och kultur samt bl.a. språk och hantverk.
Barn och unga kan delta i grundläggande undervisning i musik, dans, bildkonst och hantverk.
Dessutom erbjuder stadens ungdomstjänster en rockskola.
Stadens ungdomstjänster driver sju ungdomsgårdar runt om i Karleby.
De rusmedels- och rökfria ungdomslokalerna erbjuder handledd verksamhet för barn i årskurserna 3–6 och unga i åldern 13–17 år i olika delar av Karleby.
Information om hobbyverksamheter för barn och unga finns på stadens webbplats.
Rådgivningen vid Ungdomsgården Vinge ger aktuell information om bl.a. internationalisering, studier, arbetsliv, hälsa, hobbyverksamhet och boende.
Karlebynejdens institut erbjuder barn och unga olika former av hobbyverksamhet, exempelvis i konstämnen och musik.
Kontrollera vilka kurser som är aktuella i institutets webbtjänst.
Karleby evangelisk-lutherska församlingar erbjuder även hobbyverksamhet för barn och unga, såsom lekparksträffar, klubbar, musikverksamhet och läger.
Mer information om verksamheten finns på Karleby församlingssammanslutnings webbplats.
Ungdomsgården Vinge
67100 Karleby
Läs mer: Hobbyer för barn och unga.
Övrig undervisning i Karlebyfinska _ svenska
Ungdomstjänsterfinska _ svenska _ engelska
Karlebynejdens institutfinska _ svenska
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
Föreningar
Karleby har ett aktivt och mångsidigt föreningsliv för invånare i alla åldrar.
Läs mer: Föreningar.
Bibliotek
Motion
Att röra sig i naturen
Teater och film
Museer
Hobbyer för barn och unga
Föreningar
Karleby är en gammal sjöstad som erbjuder mångsidiga möjligheter för utfärder och friluftsliv.
Personer ntresserad av friluftsliv bör läsa mer om allemansrätten under rubriken ”Att röra sig i naturen” i denna tjänst.
Flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet.
Föreningar och organisationer samt hobbygrupper och kommunala institut erbjuder kurser i idrott och kultur samt bl.a. språk och hantverk.
I Snellman-salen och i stadens övriga kulturlokaler erbjuds kulturevenemang av varierande slag.
Årliga evenemang i Karleby är bland annat Veneziansk afton i slutet av sommaren, Kokkola Cup för fotbollsjuniorer, Stadsfestivalen Karleby sommarveckor, Lochteå kyrkomusikfest samt Vinterdans i Karleby och festivalen Karleby Vinterharmonika.
Mer information om fritidstjänsterna i Karleby finns på Karleby stads webbplats.
På stadens webbplats finns även en länk till Evenemangskalendern med daglig information om stadens kultur- och motionsevenemang.
Läs mer: Fritid.
Evenemangskalenderfinska
Kulturtjänsterfinska _ svenska _ engelska
Idrottstjänsterfinska _ svenska _ engelska
Bibliotek
Karleby stadsbibliotek finns i stadens centrum.
Närbiblioteken finns i Björkhagen, Kelviå, Lochteå samt Ullava kyrkby och Rahkonen.
Information om bibliotekets öppettider och tjänster finns på dess webbplats.
Biblioteket finns även på nätet.
Där kan kunderna bläddra i bibliotekets samlingar, reservera material, förnya sina lån, beställa fjärrlån och låna e-böcker under alla tider på dygnet.
Tack vare det effektiva biblioteksnätverket i Finland är nästan alla finländska biblioteks samlingar tillgängliga för bibliotekskunderna i Karleby.
Karleby stadsbibliotek/huvudbiblioteket
Storgatan 3, 67100 Karleby
Telefon: 040 806 5124, 040 806 5133
Läs mer: Bibliotek.
Bibliotekstjänsterfinska _ svenska _ engelska
Motion
I Karleby finns mångsidiga motionsmöjligheter året runt.
Staden anordnar ledda aktiviteter i Simcentret VesiVeijari och motionshallarna.
Dessutom finns det gym av flera olika slag.
Gym anpassade för äldre finns i Furuåsens aktivitetscenter och Kuusikumpu servicehus.
Staden underhåller cykelvägar, motionsrutter, joggingbanor, skidspår, badstränder, bollplaner och skridskobanor samt platser för närmotion.
I Karlebynejdens instituts nättjänst finns information om institutets mångsidiga motionsutbud.
I Karleby finns nära på hundra idrottsföreningar för olika grenar samt föreningar som arrangerar övrig motion.
Mer information om motionsmöjligheter i Karleby finns på Karleby stads webbplats.
Läs mer:
Motion.
Idrottstjänsterfinska _ svenska _ engelska
Motionsplatserfinska _ svenska
Gym för äldrefinska
Karlebynejdens institutfinska _ svenska
Att röra sig i naturen
Att röra sig i naturen är en traditionell och populär form av avkoppling för finländarna under alla årstider.
I Finland kan man med stöd av allemansrätten plocka bär och svamp i skogen och röra sig till fots, med cykel eller skidor vintertid.
Det är inte tillåtet att beträda folks gårdar utan lov.
För fiske krävs fiskelov, med undantag för mete och pilkning.
Även jakt fordrar jakttillstånd.
Allemansrätten ger inte rätt att skräpa ner i naturen, skada träd eller växter, störa eller skada fågelbon eller fågelungar, köra motorfordon utan markägarens tillstånd eller bygga ens tillfälliga byggen.
Mer information om motionsrutterna, rastplatser, möjligheter till fiske och båtliv samt exempelvis fågeltorn i Karleby finns på stadens webbplats.
Rutterna för camping, paddling, vandring, cykling och övriga rutter i Karleby finns i karttjänsten på nätet.
I karttjänsten visas även var största delen av motionsplatserna finns.
Du kan köpa friluftskartor över Karleby hos Karleby Turism: Salutorget 5, 67100 Karleby.
Läs mer: Att röra sig i naturen.
linkkiMiljöförvaltningen:
Allemansrättenfinska _ svenska _ engelska _ ryska
Motionskarta över Karlebyfinska _ svenska
Motionsrutter i Karlebyfinska _ svenska
Teater och film
Karleby är en teaterstad med långa anor, som erbjuder scenkonst på hög nivå framförd av både proffs och amatörer.
Karleby stadsteater finns i det stämningsfulla Vartiolinna (Torggatan 48).
Du kan läsa mer om amatörteatrarnas verksamhet på deras webbplats och i evenemangskalendern.
I Karleby finns biografen Bio Rex, vars två salar använder digital- och 3D-teknik.
Bio Rex program finns under länken här intill.
Läs mer: Teater och film.
Stadsteaternfinska
Biograffinska
Teater och danskonst i Karlebyfinska _ svenska _ engelska
Evenemangskalenderfinska
Museer
I hjärtat av staden, i det anrika Rooska gården, finns K.H.Renlunds museum.
Karleby stad grundade museet 1909 utgående från en testamentsgåva av affärsmannen Karl Herman Renlund (1850–1908) .
På museet finns Renlunds samling av finländsk konst från guldåldern och tillfälliga utställningar i en kulturhistorisk miljö.
Även i museikvarterens övriga byggnader finns utställningar om stadens kulturhistoria och utställningar med ITE-konst.
På K.H.Renlunds museums webbplats finns mer information om museets tjänster, utställningar samt aktuell verksamhet.
Utöver K.H.Renlunds museum lönar det sig att besöka det naturhistoriska museet Kieppi (Kieppi är stängt tills vidare på grund av brand) samt de många hembygdsmuseerna och övriga de historiska resmålen i regionen.
Exempelvis i Konst-Vionoja-centret presenteras konstnären Veikko Vionojas verk.
I Kelviå, ca 10 km norrut från Karleby, finns Toivonen djurpark och drängmuseum.
Mer information om dessa museer finns under länkarna här intill.
Läs mer: Museer.
Museer och traditionsarbetefinska _ svenska _ engelska
K.H. Renlunds museum - Mellersta Österbottens landskapsmuseumfinska _ svenska _ engelska
Kieppi, Karleby naturvetenskapliga museumfinska _ svenska _ engelska
linkkiToivonens djurpark och drängmuseum :
Toivonens djurpark och drängmuseum finska _ svenska _ engelska
Konst Vionojafinska
Hobbyer för barn och unga
Flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet.
Flera olika föreningar samt kommunala institut ger unga möjlighet att studera idrott och kultur samt bl.a. språk och hantverk.
Barn och unga kan delta i grundläggande undervisning i musik, dans, bildkonst och hantverk.
Dessutom erbjuder stadens ungdomstjänster en rockskola.
Stadens ungdomstjänster driver sju ungdomsgårdar runt om i Karleby.
De rusmedels- och rökfria ungdomslokalerna erbjuder handledd verksamhet för barn i årskurserna 3–6 och unga i åldern 13–17 år i olika delar av Karleby.
Information om hobbyverksamheter för barn och unga finns på stadens webbplats.
Rådgivningen vid Ungdomsgården Vinge ger aktuell information om bl.a. internationalisering, studier, arbetsliv, hälsa, hobbyverksamhet och boende.
Karlebynejdens institut erbjuder barn och unga olika former av hobbyverksamhet, exempelvis i konstämnen och musik.
Kontrollera vilka kurser som är aktuella i institutets webbtjänst.
Karleby evangelisk-lutherska församlingar erbjuder även hobbyverksamhet för barn och unga, såsom lekparksträffar, klubbar, musikverksamhet och läger.
Mer information om verksamheten finns på Karleby församlingssammanslutnings webbplats.
Ungdomsgården Vinge
67100 Karleby
Läs mer: Hobbyer för barn och unga.
Övrig undervisning i Karlebyfinska _ svenska
Ungdomstjänsterfinska _ svenska _ engelska
Karlebynejdens institutfinska _ svenska
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
Föreningar
Karleby har ett aktivt och mångsidigt föreningsliv för invånare i alla åldrar.
Läs mer: Föreningar.
Problem med uppehållstillstånd
Brott
Våld
Diskriminering och rasism
Behöver du en jurist?
Död
Problem i äktenskap eller parförhållande
Skilsmässa
Problem med den mentala hälsan
Missbruksproblem
I en krissituation kan du ringa nödcentralen på numret 112.
De slussar vid behov dig vidare till socialjouren.
Du ska endast ringa nödcentralen i brådskande nödsituationer, där liv, egendom eller miljön är i fara.
Problem med uppehållstillstånd
Om du har problem eller oklarheter med ditt uppehållstillstånd kan du kontakta Migrationsverket.
Migrationsverket
Korsholmsesplanaden 45
Vasa
Läs mer: Problem med uppehållstillstånd.
Brott
Om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112.
Ring inte nödnumret om det inte är fråga om en nödsituation.
Du kan göra en polisanmälan på nätet.
Mer information finns på Polisens webbplats.
Du kan även skriva ut anmälningsblanketten på nätet och lämna in den till polisstationen.
Karleby polisstation
Karlebygatan 74
67100 Karleby
Läs mer: Brott.
Tidsbokningfinska _ svenska _ engelska
Polisamälanfinska _ svenska _ engelska
Våld
Om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112.
Läs mer: Våld.
Diskriminering och rasism
Om du misstänker att du blivit utsatt för diskriminering då du sökt arbete eller på arbetsplatsen ska du först ta upp detta på din arbetsplats.
Om saken inte kan lösas på arbetsplatsen ska du kontakta arbetarskyddet vid Regionförvaltningsverket i Västra och Inre Finland.
Besöksadress:
Regionförvaltningsverket i Västra och Inre Finland
Wollfskavägen 35
65101 Vasa
Telefon: 0295 018 450
Om du utsätts för diskriminering kan du be om hjälp av Diskrimineringsombudsmannen.
Om du fallit offer för ett rasistiskt motiverat brott kan du göra en polisanmälan på nätet eller polisstationen.
Läs mer: Diskriminering och rasism.
linkkiRegionförvaltningsverket i Västra och Inre Finland:
Regionförvaltningsverket i Västra och Inre Finlandfinska _ svenska _ engelska
Hjälp och information för personer som drabbats av etnisk diskrimineringfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Behöver du en jurist?
Juridiska tjänster är avgiftsbelagda men om du har små eller medelstora inkomster, kan du få helt eller delvis avgiftsfri rättshjälp från statens rättshjälpsbyrå.
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
Besöksadress: Ämbetshuset, Torggatan 40, 67100 Karleby
Telefon: 029 566 1270
Information om enskilda jurister finns bland annat på Finlands Advokatförbunds webbplats.
Läs mer:
Behöver du en jurist?
linkkiFinlands advokatförbund:
Finlands advokatförbundfinska _ svenska _ engelska
Död
Den evangelisk-lutherska kyrkans församlingars begravningsplatser fungerar som allmänna begravningsplatser.
Där kan även avlidna som inte är medlemmar i kyrkan begravas.
De är alltså avsedda för alla invånare i staden.
Mer information finns på Karleby kyrkliga samfällighets webbplats.
Om en närstående plötsligt dör kan du söka krishjälp vid din egen hälsostation, eller utanför tjänstetid vid samjouren för Mellersta Österbottens centralsjukhus.
De evangelisk-lutherska församlingarna i Karlebynejden erbjuder även sorggrupper.
Även församlingarnas diakonimottagningar erbjuder samtalshjälp för sorgearbetet.
Läs mer: Död.
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Problem i äktenskap eller parförhållande
Vid problem i äktenskap eller parförhållande får du hjälp av Mellersta Österbottens familjerådgivningscentral som underhålls av Karleby kyrkliga samfällighets och Mellersta Österbottens social- och hälsovårdssamkommun Soites familjerådgivning.
Familjerågivningscentralen
Telefon: 050 3147 464.
Karleby familjerådgivning
67100 Karleby
tel. 044 730 7640
Läs mer: Problem i äktenskap eller parförhållande.
linkkiMellersta Österbottens Familjerådgivningscentral:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
Skilsmässa
Skilsmässa kan sökas av kvinnan, av mannen eller av båda makarna tillsammans.
Man ansöker om skilsmässa i tingsrätten.
Till att börja med görs en skriftlig skilsmässoansökan.
Österbottens tingsrätt Karleby kansli
Besöksadress: Karlebygatan 27, 67100 Karleby
Telefon: 029 56 49294
Läs mer: Skilsmässa.
Hälsovårdaren på barnrådgivningsbyrån ger råd i frågor som gäller små barns hälsa, tillväxt och utveckling.
Barnrådgivningsbyrån ger information om platser som erbjuder hjälp vid behov.
Vid problem hos unga i skolåldern hjälper exempelvis skolans hälsovårdare eller skolkuratorn.
Läs mer: Barns och ungas problem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Skolhälsovårdfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barnrådgivningarfinska _ svenska
Du kan ta upp problem med hälsovårdaren på skolan eller studieplatsen eller vuxna på ungdomsgården.
Mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats.
Föräldrar eller unga själva kan kontakta familjerådgivningen.
Där kan man tala om problem och få hjälp och stöd.
Mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats.
Familjerådgivningens telefonnummer: 044 730 7640.
Läs mer: Barns och ungas problem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Studerandehälsovårdfinska _ svenska
Ungdomsgårdar och -lokaler finska _ svenska
Problem med den mentala hälsan
Om du behöver hjälp och stöd för din mentala hälsa kan du boka en läkartid vid hälsostationen.
Läkaren bedömer situationen.
Vid behov skriver läkaren en remiss till psykiatrisk specialsjukvård.
Läs mer: Mental hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Mentalvårdstjänsterfinska _ svenska
Om du har ekonomiska problem kan du be om råd hos Mellersta Österbottens social- och hälsovårdssamkommun Soites enheter för socialarbete eller utkomststöd, tfn 040 806 5095 eller tjänstestyrningen, tfn 040 806 5093.
Om du har problem med skulder, kontakta rättshjälpsbyrån.
Du kan anlita vilken som helst rättshjälpsbyrå oberoende av din hemkommun.
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
Telefon: 029 566 1270
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Servicehandledningfinska _ svenska
Missbruksproblem
Om du har problem med alkohol, droger, läkemedel eller hasardspel kan du få vård och rehabilitering vid Porten, Mellersta Österbottens social- och hälsovårdssamkommun Soites center för missbruksproblem.
Du kan ta upp problemet med proffs inom hälsovården eller företagshälsovården, som kan slussa dig vidare i vårdsystemet, eller direkt kontakta Soites missbrukstjänster, tfn 040 8068 101.
För tillnyktrings- och avgiftningsvård debiteras en patientavgift liksom även för korttidsrehabilitering, öppen rehabilitering är gratis.
Även Karleby evangelisk-lutherska församlingssammanslutnings specialdiakoner erbjuder samtalshjälp vid missbruksproblem.
Kontaktuppgifter
Hälsovägen 4
67200 Karleby
Telefon: 040 806 8101
Läs mer: Missbruksproblem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Service för missbrukarefinska _ svenska
linkkiKarleby evangelisk-lutherska församlingssammansutning:
Karleby evangelisk-lutherska församlings arbete bland missbrukarefinska _ svenska
Problem med uppehållstillstånd
Brott
Våld
Diskriminering och rasism
Behöver du en jurist?
Död
Problem i äktenskap eller parförhållande
Skilsmässa
Problem med den mentala hälsan
Missbruksproblem
I en krissituation kan du ringa nödcentralen på numret 112.
De slussar vid behov dig vidare till socialjouren.
Du ska endast ringa nödcentralen i brådskande nödsituationer, där liv, egendom eller miljön är i fara.
Problem med uppehållstillstånd
Om du har problem eller oklarheter med ditt uppehållstillstånd kan du kontakta Migrationsverket.
Migrationsverket
Korsholmsesplanaden 45
Vasa
Läs mer: Problem med uppehållstillstånd.
Brott
Om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112.
Ring inte nödnumret om det inte är fråga om en nödsituation.
Du kan göra en polisanmälan på nätet.
Mer information finns på Polisens webbplats.
Du kan även skriva ut anmälningsblanketten på nätet och lämna in den till polisstationen.
Karleby polisstation
Karlebygatan 74
67100 Karleby
Läs mer: Brott.
Tidsbokningfinska _ svenska _ engelska
Polisamälanfinska _ svenska _ engelska
Våld
Om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112.
Läs mer: Våld.
Diskriminering och rasism
Om du misstänker att du blivit utsatt för diskriminering då du sökt arbete eller på arbetsplatsen ska du först ta upp detta på din arbetsplats.
Om saken inte kan lösas på arbetsplatsen ska du kontakta arbetarskyddet vid Regionförvaltningsverket i Västra och Inre Finland.
Besöksadress:
Regionförvaltningsverket i Västra och Inre Finland
Wollfskavägen 35
65101 Vasa
Telefon: 0295 018 450
Om du utsätts för diskriminering kan du be om hjälp av Diskrimineringsombudsmannen.
Om du fallit offer för ett rasistiskt motiverat brott kan du göra en polisanmälan på nätet eller polisstationen.
Läs mer: Diskriminering och rasism.
linkkiRegionförvaltningsverket i Västra och Inre Finland:
Regionförvaltningsverket i Västra och Inre Finlandfinska _ svenska _ engelska
Hjälp och information för personer som drabbats av etnisk diskrimineringfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Behöver du en jurist?
Juridiska tjänster är avgiftsbelagda men om du har små eller medelstora inkomster, kan du få helt eller delvis avgiftsfri rättshjälp från statens rättshjälpsbyrå.
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
Besöksadress: Ämbetshuset, Torggatan 40, 67100 Karleby
Telefon: 029 566 1270
Information om enskilda jurister finns bland annat på Finlands Advokatförbunds webbplats.
Läs mer:
Behöver du en jurist?
linkkiFinlands advokatförbund:
Finlands advokatförbundfinska _ svenska _ engelska
Död
Den evangelisk-lutherska kyrkans församlingars begravningsplatser fungerar som allmänna begravningsplatser.
Där kan även avlidna som inte är medlemmar i kyrkan begravas.
De är alltså avsedda för alla invånare i staden.
Mer information finns på Karleby kyrkliga samfällighets webbplats.
Om en närstående plötsligt dör kan du söka krishjälp vid din egen hälsostation, eller utanför tjänstetid vid samjouren för Mellersta Österbottens centralsjukhus.
De evangelisk-lutherska församlingarna i Karlebynejden erbjuder även sorggrupper.
Även församlingarnas diakonimottagningar erbjuder samtalshjälp för sorgearbetet.
Läs mer: Död.
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Problem i äktenskap eller parförhållande
Vid problem i äktenskap eller parförhållande får du hjälp av Mellersta Österbottens familjerådgivningscentral som underhålls av Karleby kyrkliga samfällighets och Mellersta Österbottens social- och hälsovårdssamkommun Soites familjerådgivning.
Familjerågivningscentralen
Telefon: 050 3147 464.
Karleby familjerådgivning
67100 Karleby
tel. 044 730 7640
Läs mer: Problem i äktenskap eller parförhållande.
linkkiMellersta Österbottens Familjerådgivningscentral:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
Skilsmässa
Skilsmässa kan sökas av kvinnan, av mannen eller av båda makarna tillsammans.
Man ansöker om skilsmässa i tingsrätten.
Till att börja med görs en skriftlig skilsmässoansökan.
Österbottens tingsrätt Karleby kansli
Besöksadress: Karlebygatan 27, 67100 Karleby
Telefon: 029 56 49294
Läs mer: Skilsmässa.
Hälsovårdaren på barnrådgivningsbyrån ger råd i frågor som gäller små barns hälsa, tillväxt och utveckling.
Barnrådgivningsbyrån ger information om platser som erbjuder hjälp vid behov.
Vid problem hos unga i skolåldern hjälper exempelvis skolans hälsovårdare eller skolkuratorn.
Läs mer: Barns och ungas problem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Skolhälsovårdfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barnrådgivningarfinska _ svenska
Du kan ta upp problem med hälsovårdaren på skolan eller studieplatsen eller vuxna på ungdomsgården.
Mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats.
Föräldrar eller unga själva kan kontakta familjerådgivningen.
Där kan man tala om problem och få hjälp och stöd.
Mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats.
Familjerådgivningens telefonnummer: 044 730 7640.
Läs mer: Barns och ungas problem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Studerandehälsovårdfinska _ svenska
Ungdomsgårdar och -lokaler finska _ svenska
Problem med den mentala hälsan
Om du behöver hjälp och stöd för din mentala hälsa kan du boka en läkartid vid hälsostationen.
Läkaren bedömer situationen.
Vid behov skriver läkaren en remiss till psykiatrisk specialsjukvård.
Läs mer: Mental hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Mentalvårdstjänsterfinska _ svenska
Om du har ekonomiska problem kan du be om råd hos Mellersta Österbottens social- och hälsovårdssamkommun Soites enheter för socialarbete eller utkomststöd, tfn 040 806 5095 eller tjänstestyrningen, tfn 040 806 5093.
Om du har problem med skulder, kontakta rättshjälpsbyrån.
Du kan anlita vilken som helst rättshjälpsbyrå oberoende av din hemkommun.
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
Telefon: 029 566 1270
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Servicehandledningfinska _ svenska
Missbruksproblem
Om du har problem med alkohol, droger, läkemedel eller hasardspel kan du få vård och rehabilitering vid Porten, Mellersta Österbottens social- och hälsovårdssamkommun Soites center för missbruksproblem.
Du kan ta upp problemet med proffs inom hälsovården eller företagshälsovården, som kan slussa dig vidare i vårdsystemet, eller direkt kontakta Soites missbrukstjänster, tfn 040 8068 101.
För tillnyktrings- och avgiftningsvård debiteras en patientavgift liksom även för korttidsrehabilitering, öppen rehabilitering är gratis.
Även Karleby evangelisk-lutherska församlingssammanslutnings specialdiakoner erbjuder samtalshjälp vid missbruksproblem.
Kontaktuppgifter
Hälsovägen 4
67200 Karleby
Telefon: 040 806 8101
Läs mer: Missbruksproblem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Service för missbrukarefinska _ svenska
linkkiKarleby evangelisk-lutherska församlingssammansutning:
Karleby evangelisk-lutherska församlings arbete bland missbrukarefinska _ svenska
Problem med uppehållstillstånd
Brott
Våld
Diskriminering och rasism
Behöver du en jurist?
Död
Problem i äktenskap eller parförhållande
Skilsmässa
Problem med den mentala hälsan
Missbruksproblem
I en krissituation kan du ringa nödcentralen på numret 112.
De slussar vid behov dig vidare till socialjouren.
Du ska endast ringa nödcentralen i brådskande nödsituationer, där liv, egendom eller miljön är i fara.
Problem med uppehållstillstånd
Om du har problem eller oklarheter med ditt uppehållstillstånd kan du kontakta Migrationsverket.
Migrationsverket
Korsholmsesplanaden 45
Vasa
Läs mer: Problem med uppehållstillstånd.
Brott
Om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112.
Ring inte nödnumret om det inte är fråga om en nödsituation.
Du kan göra en polisanmälan på nätet.
Mer information finns på Polisens webbplats.
Du kan även skriva ut anmälningsblanketten på nätet och lämna in den till polisstationen.
Karleby polisstation
Karlebygatan 74
67100 Karleby
Läs mer: Brott.
Tidsbokningfinska _ svenska _ engelska
Polisamälanfinska _ svenska _ engelska
Våld
Om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112.
Läs mer: Våld.
Diskriminering och rasism
Om du misstänker att du blivit utsatt för diskriminering då du sökt arbete eller på arbetsplatsen ska du först ta upp detta på din arbetsplats.
Om saken inte kan lösas på arbetsplatsen ska du kontakta arbetarskyddet vid Regionförvaltningsverket i Västra och Inre Finland.
Besöksadress:
Regionförvaltningsverket i Västra och Inre Finland
Wollfskavägen 35
65101 Vasa
Telefon: 0295 018 450
Om du utsätts för diskriminering kan du be om hjälp av Diskrimineringsombudsmannen.
Om du fallit offer för ett rasistiskt motiverat brott kan du göra en polisanmälan på nätet eller polisstationen.
Läs mer: Diskriminering och rasism.
linkkiRegionförvaltningsverket i Västra och Inre Finland:
Regionförvaltningsverket i Västra och Inre Finlandfinska _ svenska _ engelska
Hjälp och information för personer som drabbats av etnisk diskrimineringfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Behöver du en jurist?
Juridiska tjänster är avgiftsbelagda men om du har små eller medelstora inkomster, kan du få helt eller delvis avgiftsfri rättshjälp från statens rättshjälpsbyrå.
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
Besöksadress: Ämbetshuset, Torggatan 40, 67100 Karleby
Telefon: 029 566 1270
Information om enskilda jurister finns bland annat på Finlands Advokatförbunds webbplats.
Läs mer:
Behöver du en jurist?
linkkiFinlands advokatförbund:
Finlands advokatförbundfinska _ svenska _ engelska
Död
Den evangelisk-lutherska kyrkans församlingars begravningsplatser fungerar som allmänna begravningsplatser.
Där kan även avlidna som inte är medlemmar i kyrkan begravas.
De är alltså avsedda för alla invånare i staden.
Mer information finns på Karleby kyrkliga samfällighets webbplats.
Om en närstående plötsligt dör kan du söka krishjälp vid din egen hälsostation, eller utanför tjänstetid vid samjouren för Mellersta Österbottens centralsjukhus.
De evangelisk-lutherska församlingarna i Karlebynejden erbjuder även sorggrupper.
Även församlingarnas diakonimottagningar erbjuder samtalshjälp för sorgearbetet.
Läs mer: Död.
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Problem i äktenskap eller parförhållande
Vid problem i äktenskap eller parförhållande får du hjälp av Mellersta Österbottens familjerådgivningscentral som underhålls av Karleby kyrkliga samfällighets och Mellersta Österbottens social- och hälsovårdssamkommun Soites familjerådgivning.
Familjerågivningscentralen
Telefon: 050 3147 464.
Karleby familjerådgivning
67100 Karleby
tel. 044 730 7640
Läs mer: Problem i äktenskap eller parförhållande.
linkkiMellersta Österbottens Familjerådgivningscentral:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
Skilsmässa
Skilsmässa kan sökas av kvinnan, av mannen eller av båda makarna tillsammans.
Man ansöker om skilsmässa i tingsrätten.
Till att börja med görs en skriftlig skilsmässoansökan.
Österbottens tingsrätt Karleby kansli
Besöksadress: Karlebygatan 27, 67100 Karleby
Telefon: 029 56 49294
Läs mer: Skilsmässa.
Hälsovårdaren på barnrådgivningsbyrån ger råd i frågor som gäller små barns hälsa, tillväxt och utveckling.
Barnrådgivningsbyrån ger information om platser som erbjuder hjälp vid behov.
Vid problem hos unga i skolåldern hjälper exempelvis skolans hälsovårdare eller skolkuratorn.
Läs mer: Barns och ungas problem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Skolhälsovårdfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barnrådgivningarfinska _ svenska
Du kan ta upp problem med hälsovårdaren på skolan eller studieplatsen eller vuxna på ungdomsgården.
Mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats.
Föräldrar eller unga själva kan kontakta familjerådgivningen.
Där kan man tala om problem och få hjälp och stöd.
Mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats.
Familjerådgivningens telefonnummer: 044 730 7640.
Läs mer: Barns och ungas problem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Studerandehälsovårdfinska _ svenska
Ungdomsgårdar och -lokaler finska _ svenska
Problem med den mentala hälsan
Om du behöver hjälp och stöd för din mentala hälsa kan du boka en läkartid vid hälsostationen.
Läkaren bedömer situationen.
Vid behov skriver läkaren en remiss till psykiatrisk specialsjukvård.
Läs mer: Mental hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Mentalvårdstjänsterfinska _ svenska
Om du har ekonomiska problem kan du be om råd hos Mellersta Österbottens social- och hälsovårdssamkommun Soites enheter för socialarbete eller utkomststöd, tfn 040 806 5095 eller tjänstestyrningen, tfn 040 806 5093.
Om du har problem med skulder, kontakta rättshjälpsbyrån.
Du kan anlita vilken som helst rättshjälpsbyrå oberoende av din hemkommun.
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
Telefon: 029 566 1270
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Servicehandledningfinska _ svenska
Missbruksproblem
Om du har problem med alkohol, droger, läkemedel eller hasardspel kan du få vård och rehabilitering vid Porten, Mellersta Österbottens social- och hälsovårdssamkommun Soites center för missbruksproblem.
Du kan ta upp problemet med proffs inom hälsovården eller företagshälsovården, som kan slussa dig vidare i vårdsystemet, eller direkt kontakta Soites missbrukstjänster, tfn 040 8068 101.
För tillnyktrings- och avgiftningsvård debiteras en patientavgift liksom även för korttidsrehabilitering, öppen rehabilitering är gratis.
Även Karleby evangelisk-lutherska församlingssammanslutnings specialdiakoner erbjuder samtalshjälp vid missbruksproblem.
Kontaktuppgifter
Hälsovägen 4
67200 Karleby
Telefon: 040 806 8101
Läs mer: Missbruksproblem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Service för missbrukarefinska _ svenska
linkkiKarleby evangelisk-lutherska församlingssammansutning:
Karleby evangelisk-lutherska församlings arbete bland missbrukarefinska _ svenska
Äktenskap
Skilsmässa
Barn vid skilsmässa
När du väntar barn
Vård av barnet
Vård av barnet i hemmet
Äktenskap
Innan äktenskapet ingås ska du skriftligen be om prövning av äktenskapshinder.
Prövningen görs vid magistraten. Du kan lämna in ansökan om prövning vid vilken magistrat som helst.
Civilvigsel äger rum vid magistraten.
Magistraten i Västra Finland
Karleby enhet
Karlebygatan 27, PB 581
67701 Karleby
Telefon: 029 553 9451
Läs mer:
Äktenskap.
Skilsmässa
Skilsmässa kan sökas av kvinnan, av mannen eller av båda makarna tillsammans.
Man ansöker om skilsmässa i tingsrätten.
Till att börja med görs en skriftlig skilsmässoansökan.
Österbottens tingsrätt Karleby kansli
Besöksadress: Karlebygatan 27, 67100 Karleby
Telefon: 029 56 49294
Läs mer: Skilsmässa.
Barn vid skilsmässa
Om du har barn och går igenom en skilsmässa ska du ta kontakt med barnatillsyningsmannen.
Barnatillsyningsmannen bekräftar överenskommelsen om var barnen ska bo, vården av barnen, umgängesrätt och underhållsbidrag.
Barnatillsyningsmannen
67100 Karleby
Telefontid och tidsbokning
tel. 06 826 4111
Läs mer: Barn vid skilsmässa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barnatillsyningsmannenfinska _ svenska
När du väntar barn
Ta kontakt med rådgivningen då du märker att du är gravid.
På rådgivningen följer man med moderns, barnets och hela familjens välmående under graviditeten.
Du kan be om råd per telefon (06) 826 4477.
Läs mer:
När du väntar barn.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Mödrarådgivningfinska _ svenska
Vård av barnet
I Karleby finns stadens daghem, gruppfamiljedaghem, familjedagvårdare samt barnklubbar.
Dessutom finns det daghem som köptjänst (svenskspråkiga), ett privat daghem och privata familjedagvårdare i Karleby.
Du kan ansöka om plats inom småbarnspedagogiken för ditt barn elektroniskt via tjänsten suomi.fi eller med en blankett på stadens webbplats (ansökan om småbarnspedagogik).
Ansökan ska lämnas in fyra månader innan du behöver plats inom småbarnspedagogiken.
Det är möjligt att få en plats snabbare om den behövs för att du exempelvis erhållit arbete eller studieplats.
Ansökan kan returneras till platsen för småbarnspedagogik, kontorstjänster för småbarnspedagogik eller lämnas i brevlådan i den nedre aulan i Bildningscentralen.
Du kan ansöka om en plats i stadens barnklubbar med blanketten som finns på stadens webbplats.
Ansökan kan även skickas per post till följande adress:
Bildningscentralen
Tjänster för småbarnspedagogik
Strandgatan16
67100 Karleby
Läs mer:
Daghem och andra dagvårdsplatserfinska _ svenska
Gruppfamiljedaghemfinska _ svenska
Dagvårdsblanketterfinska _ svenska
Att ansöka om kommunal dagvårdfinska _ svenska
Vård av barnet i hemmet
Om familjens yngsta barn är yngre än tre år kan föräldern få hemvårdsstöd för vård av barnet i hemmet.
Om du har rätt till stödet kan du ansöka om stödet hos FPA.
Du kan fylla i ansökan på nätet eller skicka den per post till FPA.
Du kan även besöka FPA:s kontor.
Karleby stad betalar extra Karlebystöd för de familjer som tar hand om barn under tre år i hemmet.
Du kan ansöka om Karlebystödet om den ena av föräldrarna vårdar samtliga av familjens barn under skolåldern i hemmet.
Om din familj fyller villkoren, beviljas Karlebystödet i samband med beviljandet av vårdnadsbidraget.
Läs mer:
Stöd för vård av barn i hemmet.
Karlebystödfinska _ svenska
Information om FPA:s hemvårdsstödfinska _ svenska _ engelska
FPA kontaktuppgifterfinska _ svenska _ engelska
Äktenskap
Skilsmässa
Barn vid skilsmässa
När du väntar barn
Vård av barnet
Vård av barnet i hemmet
Äktenskap
Innan äktenskapet ingås ska du skriftligen be om prövning av äktenskapshinder.
Prövningen görs vid magistraten. Du kan lämna in ansökan om prövning vid vilken magistrat som helst.
Civilvigsel äger rum vid magistraten.
Magistraten i Västra Finland
Karleby enhet
Karlebygatan 27, PB 581
67701 Karleby
Telefon: 029 553 9451
Läs mer:
Äktenskap.
Skilsmässa
Skilsmässa kan sökas av kvinnan, av mannen eller av båda makarna tillsammans.
Man ansöker om skilsmässa i tingsrätten.
Till att börja med görs en skriftlig skilsmässoansökan.
Österbottens tingsrätt Karleby kansli
Besöksadress: Karlebygatan 27, 67100 Karleby
Telefon: 029 56 49294
Läs mer: Skilsmässa.
Barn vid skilsmässa
Om du har barn och går igenom en skilsmässa ska du ta kontakt med barnatillsyningsmannen.
Barnatillsyningsmannen bekräftar överenskommelsen om var barnen ska bo, vården av barnen, umgängesrätt och underhållsbidrag.
Barnatillsyningsmannen
67100 Karleby
Telefontid och tidsbokning
tel. 06 826 4111
Läs mer: Barn vid skilsmässa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barnatillsyningsmannenfinska _ svenska
När du väntar barn
Ta kontakt med rådgivningen då du märker att du är gravid.
På rådgivningen följer man med moderns, barnets och hela familjens välmående under graviditeten.
Du kan be om råd per telefon (06) 826 4477.
Läs mer:
När du väntar barn.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Mödrarådgivningfinska _ svenska
Vård av barnet
I Karleby finns stadens daghem, gruppfamiljedaghem, familjedagvårdare samt barnklubbar.
Dessutom finns det daghem som köptjänst (svenskspråkiga), ett privat daghem och privata familjedagvårdare i Karleby.
Du kan ansöka om plats inom småbarnspedagogiken för ditt barn elektroniskt via tjänsten suomi.fi eller med en blankett på stadens webbplats (ansökan om småbarnspedagogik).
Ansökan ska lämnas in fyra månader innan du behöver plats inom småbarnspedagogiken.
Det är möjligt att få en plats snabbare om den behövs för att du exempelvis erhållit arbete eller studieplats.
Ansökan kan returneras till platsen för småbarnspedagogik, kontorstjänster för småbarnspedagogik eller lämnas i brevlådan i den nedre aulan i Bildningscentralen.
Du kan ansöka om en plats i stadens barnklubbar med blanketten som finns på stadens webbplats.
Ansökan kan även skickas per post till följande adress:
Bildningscentralen
Tjänster för småbarnspedagogik
Strandgatan16
67100 Karleby
Läs mer:
Daghem och andra dagvårdsplatserfinska _ svenska
Gruppfamiljedaghemfinska _ svenska
Dagvårdsblanketterfinska _ svenska
Att ansöka om kommunal dagvårdfinska _ svenska
Vård av barnet i hemmet
Om familjens yngsta barn är yngre än tre år kan föräldern få hemvårdsstöd för vård av barnet i hemmet.
Om du har rätt till stödet kan du ansöka om stödet hos FPA.
Du kan fylla i ansökan på nätet eller skicka den per post till FPA.
Du kan även besöka FPA:s kontor.
Karleby stad betalar extra Karlebystöd för de familjer som tar hand om barn under tre år i hemmet.
Du kan ansöka om Karlebystödet om den ena av föräldrarna vårdar samtliga av familjens barn under skolåldern i hemmet.
Om din familj fyller villkoren, beviljas Karlebystödet i samband med beviljandet av vårdnadsbidraget.
Läs mer:
Stöd för vård av barn i hemmet.
Karlebystödfinska _ svenska
Information om FPA:s hemvårdsstödfinska _ svenska _ engelska
FPA kontaktuppgifterfinska _ svenska _ engelska
Äktenskap
Skilsmässa
Barn vid skilsmässa
När du väntar barn
Vård av barnet
Vård av barnet i hemmet
Äktenskap
Innan äktenskapet ingås ska du skriftligen be om prövning av äktenskapshinder.
Prövningen görs vid magistraten. Du kan lämna in ansökan om prövning vid vilken magistrat som helst.
Civilvigsel äger rum vid magistraten.
Magistraten i Västra Finland
Karleby enhet
Karlebygatan 27, PB 581
67701 Karleby
Telefon: 029 553 9451
Läs mer:
Äktenskap.
Skilsmässa
Skilsmässa kan sökas av kvinnan, av mannen eller av båda makarna tillsammans.
Man ansöker om skilsmässa i tingsrätten.
Till att börja med görs en skriftlig skilsmässoansökan.
Österbottens tingsrätt Karleby kansli
Besöksadress: Karlebygatan 27, 67100 Karleby
Telefon: 029 56 49294
Läs mer: Skilsmässa.
Barn vid skilsmässa
Om du har barn och går igenom en skilsmässa ska du ta kontakt med barnatillsyningsmannen.
Barnatillsyningsmannen bekräftar överenskommelsen om var barnen ska bo, vården av barnen, umgängesrätt och underhållsbidrag.
Barnatillsyningsmannen
67100 Karleby
Telefontid och tidsbokning
tel. 06 826 4111
Läs mer: Barn vid skilsmässa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barnatillsyningsmannenfinska _ svenska
När du väntar barn
Ta kontakt med rådgivningen då du märker att du är gravid.
På rådgivningen följer man med moderns, barnets och hela familjens välmående under graviditeten.
Du kan be om råd per telefon (06) 826 4477.
Läs mer: Graviditet och förlossning.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Mödrarådgivningfinska _ svenska
Vård av barnet
I Karleby finns stadens daghem, gruppfamiljedaghem, familjedagvårdare samt barnklubbar.
Dessutom finns det daghem som köptjänst (svenskspråkiga), ett privat daghem och privata familjedagvårdare i Karleby.
Du kan ansöka om plats inom småbarnspedagogiken för ditt barn elektroniskt via tjänsten suomi.fi eller med en blankett på stadens webbplats (ansökan om småbarnspedagogik).
Ansökan ska lämnas in fyra månader innan du behöver plats inom småbarnspedagogiken.
Det är möjligt att få en plats snabbare om den behövs för att du exempelvis erhållit arbete eller studieplats.
Ansökan kan returneras till platsen för småbarnspedagogik, kontorstjänster för småbarnspedagogik eller lämnas i brevlådan i den nedre aulan i Bildningscentralen.
Du kan ansöka om en plats i stadens barnklubbar med blanketten som finns på stadens webbplats.
Ansökan kan även skickas per post till följande adress:
Bildningscentralen
Tjänster för småbarnspedagogik
Strandgatan16
67100 Karleby
Läs mer:
Vård av barnet.
Daghem och andra dagvårdsplatserfinska _ svenska
Gruppfamiljedaghemfinska _ svenska
Dagvårdsblanketterfinska _ svenska
Att ansöka om kommunal dagvårdfinska _ svenska
Vård av barnet i hemmet
Om familjens yngsta barn är yngre än tre år kan föräldern få hemvårdsstöd för vård av barnet i hemmet.
Om du har rätt till stödet kan du ansöka om stödet hos FPA.
Du kan fylla i ansökan på nätet eller skicka den per post till FPA.
Du kan även besöka FPA:s kontor.
Karleby stad betalar extra Karlebystöd för de familjer som tar hand om barn under tre år i hemmet.
Du kan ansöka om Karlebystödet om den ena av föräldrarna vårdar samtliga av familjens barn under skolåldern i hemmet.
Om din familj fyller villkoren, beviljas Karlebystödet i samband med beviljandet av vårdnadsbidraget.
Läs mer:
Stöd för vård av barn i hemmet.
Karlebystödfinska _ svenska
Information om FPA:s hemvårdsstödfinska _ svenska _ engelska
FPA kontaktuppgifterfinska _ svenska _ engelska
Hälsovårdstjänster i Karleby
Äldre människors hälsa
Tandvård
Mental hälsa
Sexuell hälsa
När du väntar barn
Förlossning
Läkemedel
Handikappade personer
Ett handikappat barn
Hälsovårdstjänster i Karleby
I Karleby finns hälsostationer i olika delar av staden.
Varje hälsostation har ett eget telefonnummer för tidsbokning, som man kan ringa för att boka tid till sjukskötare eller läkare.
Kontaktuppgifter:
Karleby huvudhälsostation
Mariegatan 28
67200 Karleby
Telefon: (06) 8287 580
På Karleby huvudhälsostationen styrs patienterna till mottagningen på basis av hur akuta deras symptom är.
Klienten får en tid till akutvården, mottagningen eller Min Soite-mottagningen.
Samtal till huvudhälsostationen styrs till ett och samma telefonnummer, (06) 8287 310.
67800 Karleby
Telefon: (06) 8287 580
Mottagning /Kelviå
Ellfolkgatan 5
68300 Kelviå
Telefon: (06) 8287 701
Mottagning /Lochteå
Telefon: (06) 8287 750
Mottagning /Ullava
Ullavavägen 701
68370 Ullava
Telefon: (06) 8287 639
Om du kommer som flykting till Finland ska du komma överens om en hälsokontroll med Utlänningsbyrån.
Läs mer: Hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
Under kvällar och helger är hälsostationerna stängda.
Då hanteras plötsliga sjukdomar och olyckor vid jouren.
Jouren är avsedd för patienter vars sjukdom kräver brådskande bedömning och vård.
I livshotande situationer ska du ringa nödnumret 112.
Om du besöker jouren kvällstid eller under helger ska du först ringa jourens telefonrådgivning (06) 826 4500.
Samjourens adress:
Mellersta Österbottens centralsjukhus
Mariegatan 16–20 (l-flygeln, ingång B1)
67200 Karleby
Läs mer: Hälsovårdstjänster i Finland
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barns hälsa
Om ditt barn insjuknar ska du kontakta hälsostationen vid behov.
ådgivningarna erbjuder tjänster för gravida och barn under skolåldern.
Vid rådgivningarna utförs vaccinationer av barn och vuxna.
Du kan kontakta rådgivningen via den centraliserade telefontjänsten (06) 826 4477.
Genom regelbundna besök på barnrådgivningsbyrån följs barnets hälsa, tillväxt och utveckling upp.
På rådgivningen vårdas inte barn som insjuknar plötsligt, men du kan be om råd via den centraliserade telefontjänsten (06) 826 4477.
Skolhälsovårdaren har hand om skolelevers hälsa.
Mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats.
Läs mer: Barns hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barnrådgivningarfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Rådgivningarfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Skolhälsovårdfinska _ svenska
Äldre människors hälsa
Vid hälsopunkten Daalia ges vägledning och rådgivning för personer över 65 år om diet, motion och livsstil.
Vaccinering av personer över 65 år utförs vid seniorrådgivning.
Läs mer:
Äldre människors hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Seniorernas hälsopunkterfinska _ svenska
Tandvård
Om du behöver icke-brådskande tandvård ska du ringa munhälsans centraliserade tidsbokningen.
Centraliserad tidsbokning per telefon: (06) 8287 400
Huvudhälsostationens tandklinik
Mariegatan 28, 67200 Karleby
Björkhagens tandklinik
Storkisbackens tandklinik
Korpvägen 11, 67100 Karleby
Kelviå tandklinik
Ellfolkgatan 5, 68300, Kelviå
Lochteå tandklinik
Ullava tandklinik
Ullavavägen 701, 68370 Ullava
Vardagar kan tider till smärtjouren bokas enligt överenskommelse vid samtliga tandkliniker.
Brådskande tandvård/första hjälpen (kvälls-, vardags-, helg- och nattjour):
Vid smärtjouren får du första hjälpen vid plötslig tandvärk och tandolyckor.
Tandläkarjouren (kvälls-, vardags- och helgjour) ordnas vid polikliniken för tand- och munsjukdomar vid Mellersta Österbottens social- och hälsovårdssamkommun Soite, Mariegatan 16–20, 67200 Karleby (vån 1, del D), vardagkvällar kl. 16.00–21.00 samt veckoslut och helgdagar kl. 8.00–21.00.
Du kan i regel komma till jourmottagningen genom att först kontakta jouren via telefon.
För frågor gällande jouren ring tel. (06) 828 7450.
När du kommer till jourmottagningen ska du ta en kölapp, såvida du inte har en bokad tid.
Brådskande tandvård/första hjälpen (nattjour):
Allvarliga fall i samjour Uleåborgs universitetssjukhus (Oulun yliopistollinen sairaala OYS) kl. 21.00−8.00, tel. (08) 315 2655
Läs mer: Tandvård.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Munhälsovårdenfinska _ svenska
Mental hälsa
Vid problem med din mentala hälsa ska du i första hand kontakta din egen hälsostation eller företagshälsovårdens mottagning.
Vid brådskande problem, kontakta hälsovårdcentralens jour.
Läs mer: Mental hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
Sexuell hälsa
Om du känner att du behöver information om familjeplanering och prevention kan du kontakta din egen hälsostation.
Boka tid till hälsostationen om du behöver preventivmedel, överväger att göra en abort eller misstänker att du lider av en könssjukdom.
Du kan även boka en tid hos en allmänläkare för en gynekologisk eller urologisk undersökning.
I preventionsfrågor kan du kontakta den centraliserade telefontjänsten (06) 826 4477.
Läs mer:
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Preventivrådgivningfinska _ svenska
När du väntar barn
Ta kontakt med rådgivningen då du märker att du är gravid.
På rådgivningen följer man med moderns, barnets och hela familjens välmående under graviditeten.
Läs mer:
När du väntar barn.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Mödrarådgivningfinska _ svenska
Förlossning
Förlossningsavdelningen är öppen dygnet runt.
Om du önskar kan du ringa förlossningsavdelning då din förlossning satt igång eller om du vill fråga om råd.
Då du kommer till sjukhuset ska du använda centralsjukhusets huvudingång kl. 7–20 och övriga tider bör du använda den gemensamma jourens/poliklinikens dörr.
Kontaktuppgifter för förlossningsavdelningen:
Mariegatan 16–20,
67200 Karleby
Telefon: (06) 8264355.
Läs mer: Förlossning.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Förlossningarfinska _ svenska
Läkemedel
Du kan köpa läkemedel på apoteket.
Du kan besöka vilket apotek som helst.
Du kan även besöka apotek som inte finns i din egen kommun.
Läs mer: Läkemedel.
Handikappade personer
En handikappad person bosatt i Karleby har rätt att erhålla de tjänster han eller hon behöver på samma grunder som de övriga invånarna i kommunen.
Personen kan dock på grund av sitt handikapp eller sin sjukdom även behöva särskilda tjänster för handikappade för att klara vardagen.
För tjänsterna för handikappade i Karleby svarar Mellersta Österbottens social- och hälsovårdssamkommun Soite, där man kan ansöka om tjänster och stödfunktioner.
Tjänster av flera olika slag erbjuds även för personer med gravt handikapp.
Dessa tjänster inkluderar bland annat:
transporttjänster
ombyggnad och nödvändig utrustning för hemmet
maskiner och utrustning
personlig hjälp och dagverksamhet
stödboende
stöd för närståendevård av personer under 65 och arbetsverksamhet.
Dessutom är det möjligt att ansöka om specialboende, korttidsvård eller tillfällig vård samt handledning hos den öppna vården.
Mer information om tjänster för handikappade får du från Mellersta Österbottens social- och hälsovårdssamkommun Soites handikapptjänster per telefon: 040 804 2122.
Läs mer: Handikappade personer.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Tjänster för handikappadefinska _ svenska
Specialpedagogik i förskolanfinska _ svenska
Kontaktuppgifter för den grundläggande utbildningenfinska
Ett handikappat barn
Särskilt stöd erbjuds barn med handikapp inom småbarnspedagogiken och skolan.
Kontakta Karleby stads förskoleundervisning för information om specialsmåbarnspedagogiken.
Du kan be undervisningsväsendet om mer information om tjänster som skolan erbjuder.
Bildningscentralen
Strandgatan 16 (våning 5 och 6)
67100 Karleby
Telefon: 040 8065 149
Läs mer: Ett handikappat barn.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Tjänster för handikappadefinska _ svenska
Specialpedagogik i förskolanfinska _ svenska
Kontaktuppgifter för den grundläggande utbildningenfinska
Hälsovårdstjänster i Karleby
Äldre människors hälsa
Tandvård
Mental hälsa
Sexuell hälsa
När du väntar barn
Förlossning
Läkemedel
Handikappade personer
Ett handikappat barn
Hälsovårdstjänster i Karleby
I Karleby finns hälsostationer i olika delar av staden.
Varje hälsostation har ett eget telefonnummer för tidsbokning, som man kan ringa för att boka tid till sjukskötare eller läkare.
Kontaktuppgifter:
Karleby huvudhälsostation
Mariegatan 28
67200 Karleby
Telefon: (06) 8287 580
På Karleby huvudhälsostationen styrs patienterna till mottagningen på basis av hur akuta deras symptom är.
Klienten får en tid till akutvården, mottagningen eller Min Soite-mottagningen.
Samtal till huvudhälsostationen styrs till ett och samma telefonnummer, (06) 8287 310.
67800 Karleby
Telefon: (06) 8287 580
Mottagning /Kelviå
Ellfolkgatan 5
68300 Kelviå
Telefon: (06) 8287 701
Mottagning /Lochteå
Telefon: (06) 8287 750
Mottagning /Ullava
Ullavavägen 701
68370 Ullava
Telefon: (06) 8287 639
Om du kommer som flykting till Finland ska du komma överens om en hälsokontroll med Utlänningsbyrån.
Läs mer: Hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
Under kvällar och helger är hälsostationerna stängda.
Då hanteras plötsliga sjukdomar och olyckor vid jouren.
Jouren är avsedd för patienter vars sjukdom kräver brådskande bedömning och vård.
I livshotande situationer ska du ringa nödnumret 112.
Om du besöker jouren kvällstid eller under helger ska du först ringa jourens telefonrådgivning (06) 826 4500.
Samjourens adress:
Mellersta Österbottens centralsjukhus
Mariegatan 16–20 (l-flygeln, ingång B1)
67200 Karleby
Läs mer: Hälsovårdstjänster i Finland
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barns hälsa
Om ditt barn insjuknar ska du kontakta hälsostationen vid behov.
ådgivningarna erbjuder tjänster för gravida och barn under skolåldern.
Vid rådgivningarna utförs vaccinationer av barn och vuxna.
Du kan kontakta rådgivningen via den centraliserade telefontjänsten (06) 826 4477.
Genom regelbundna besök på barnrådgivningsbyrån följs barnets hälsa, tillväxt och utveckling upp.
På rådgivningen vårdas inte barn som insjuknar plötsligt, men du kan be om råd via den centraliserade telefontjänsten (06) 826 4477.
Skolhälsovårdaren har hand om skolelevers hälsa.
Mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats.
Läs mer: Barns hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barnrådgivningarfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Rådgivningarfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Skolhälsovårdfinska _ svenska
Äldre människors hälsa
Vid hälsopunkten Daalia ges vägledning och rådgivning för personer över 65 år om diet, motion och livsstil.
Vaccinering av personer över 65 år utförs vid seniorrådgivning.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Seniorernas hälsopunkterfinska _ svenska
Tandvård
Om du behöver icke-brådskande tandvård ska du ringa munhälsans centraliserade tidsbokningen.
Centraliserad tidsbokning per telefon: (06) 8287 400
Huvudhälsostationens tandklinik
Mariegatan 28, 67200 Karleby
Björkhagens tandklinik
Storkisbackens tandklinik
Korpvägen 11, 67100 Karleby
Kelviå tandklinik
Ellfolkgatan 5, 68300, Kelviå
Lochteå tandklinik
Ullava tandklinik
Ullavavägen 701, 68370 Ullava
Vardagar kan tider till smärtjouren bokas enligt överenskommelse vid samtliga tandkliniker.
Brådskande tandvård/första hjälpen (kvälls-, vardags-, helg- och nattjour):
Vid smärtjouren får du första hjälpen vid plötslig tandvärk och tandolyckor.
Tandläkarjouren (kvälls-, vardags- och helgjour) ordnas vid polikliniken för tand- och munsjukdomar vid Mellersta Österbottens social- och hälsovårdssamkommun Soite, Mariegatan 16–20, 67200 Karleby (vån 1, del D), vardagkvällar kl. 16.00–21.00 samt veckoslut och helgdagar kl. 8.00–21.00.
Du kan i regel komma till jourmottagningen genom att först kontakta jouren via telefon.
För frågor gällande jouren ring tel. (06) 828 7450.
När du kommer till jourmottagningen ska du ta en kölapp, såvida du inte har en bokad tid.
Brådskande tandvård/första hjälpen (nattjour):
Allvarliga fall i samjour Uleåborgs universitetssjukhus (Oulun yliopistollinen sairaala OYS) kl. 21.00−8.00, tel. (08) 315 2655
Läs mer: Tandvård.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Munhälsovårdenfinska _ svenska
Mental hälsa
Vid problem med din mentala hälsa ska du i första hand kontakta din egen hälsostation eller företagshälsovårdens mottagning.
Vid brådskande problem, kontakta hälsovårdcentralens jour.
Läs mer: Mental hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
Sexuell hälsa
Om du känner att du behöver information om familjeplanering och prevention kan du kontakta din egen hälsostation.
Boka tid till hälsostationen om du behöver preventivmedel, överväger att göra en abort eller misstänker att du lider av en könssjukdom.
Du kan även boka en tid hos en allmänläkare för en gynekologisk eller urologisk undersökning.
I preventionsfrågor kan du kontakta den centraliserade telefontjänsten (06) 826 4477.
Läs mer:
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Preventivrådgivningfinska _ svenska
När du väntar barn
Ta kontakt med rådgivningen då du märker att du är gravid.
På rådgivningen följer man med moderns, barnets och hela familjens välmående under graviditeten.
Läs mer:
När du väntar barn.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Mödrarådgivningfinska _ svenska
Förlossning
Förlossningsavdelningen är öppen dygnet runt.
Om du önskar kan du ringa förlossningsavdelning då din förlossning satt igång eller om du vill fråga om råd.
Då du kommer till sjukhuset ska du använda centralsjukhusets huvudingång kl. 7–20 och övriga tider bör du använda den gemensamma jourens/poliklinikens dörr.
Kontaktuppgifter för förlossningsavdelningen:
Mariegatan 16–20,
67200 Karleby
Telefon: (06) 8264355.
Läs mer: Förlossning.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Förlossningarfinska _ svenska
Läkemedel
Du kan köpa läkemedel på apoteket.
Du kan besöka vilket apotek som helst.
Du kan även besöka apotek som inte finns i din egen kommun.
Läs mer: Läkemedel.
Handikappade personer
En handikappad person bosatt i Karleby har rätt att erhålla de tjänster han eller hon behöver på samma grunder som de övriga invånarna i kommunen.
Personen kan dock på grund av sitt handikapp eller sin sjukdom även behöva särskilda tjänster för handikappade för att klara vardagen.
För tjänsterna för handikappade i Karleby svarar Mellersta Österbottens social- och hälsovårdssamkommun Soite, där man kan ansöka om tjänster och stödfunktioner.
Tjänster av flera olika slag erbjuds även för personer med gravt handikapp.
Dessa tjänster inkluderar bland annat:
transporttjänster
ombyggnad och nödvändig utrustning för hemmet
maskiner och utrustning
personlig hjälp och dagverksamhet
stödboende
stöd för närståendevård av personer under 65 och arbetsverksamhet.
Dessutom är det möjligt att ansöka om specialboende, korttidsvård eller tillfällig vård samt handledning hos den öppna vården.
Mer information om tjänster för handikappade får du från Mellersta Österbottens social- och hälsovårdssamkommun Soites handikapptjänster per telefon: 040 804 2122.
Läs mer: Handikappade personer.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Tjänster för handikappadefinska _ svenska
Specialpedagogik i förskolanfinska _ svenska
Kontaktuppgifter för den grundläggande utbildningenfinska
Ett handikappat barn
Särskilt stöd erbjuds barn med handikapp inom småbarnspedagogiken och skolan.
Kontakta Karleby stads förskoleundervisning för information om specialsmåbarnspedagogiken.
Du kan be undervisningsväsendet om mer information om tjänster som skolan erbjuder.
Bildningscentralen
Strandgatan 16 (våning 5 och 6)
67100 Karleby
Telefon: 040 8065 149
Läs mer: Ett handikappat barn.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Tjänster för handikappadefinska _ svenska
Specialpedagogik i förskolanfinska _ svenska
Kontaktuppgifter för den grundläggande utbildningenfinska
Hälsovårdstjänster i Karleby
Äldre människors hälsa
Tandvård
Mental hälsa
Sexuell hälsa
När du väntar barn
Förlossning
Läkemedel
Handikappade personer
Ett handikappat barn
Hälsovårdstjänster i Karleby
I Karleby finns hälsostationer i olika delar av staden.
Varje hälsostation har ett eget telefonnummer för tidsbokning, som man kan ringa för att boka tid till sjukskötare eller läkare.
Kontaktuppgifter:
Karleby huvudhälsostation
Mariegatan 28
67200 Karleby
Telefon: (06) 8287 580
På Karleby huvudhälsostationen styrs patienterna till mottagningen på basis av hur akuta deras symptom är.
Klienten får en tid till akutvården, mottagningen eller Min Soite-mottagningen.
Samtal till huvudhälsostationen styrs till ett och samma telefonnummer, (06) 8287 310.
67800 Karleby
Telefon: (06) 8287 580
Mottagning /Kelviå
Ellfolkgatan 5
68300 Kelviå
Telefon: (06) 8287 701
Mottagning /Lochteå
Telefon: (06) 8287 750
Mottagning /Ullava
Ullavavägen 701
68370 Ullava
Telefon: (06) 8287 639
Om du kommer som flykting till Finland ska du komma överens om en hälsokontroll med Utlänningsbyrån.
Läs mer: Hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
Under kvällar och helger är hälsostationerna stängda.
Då hanteras plötsliga sjukdomar och olyckor vid jouren.
Jouren är avsedd för patienter vars sjukdom kräver brådskande bedömning och vård.
I livshotande situationer ska du ringa nödnumret 112.
Om du besöker jouren kvällstid eller under helger ska du först ringa jourens telefonrådgivning (06) 826 4500.
Samjourens adress:
Mellersta Österbottens centralsjukhus
Mariegatan 16–20 (l-flygeln, ingång B1)
67200 Karleby
Läs mer: Hälsovårdstjänster i Finland
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barns hälsa
Om ditt barn insjuknar ska du kontakta hälsostationen vid behov.
ådgivningarna erbjuder tjänster för gravida och barn under skolåldern.
Vid rådgivningarna utförs vaccinationer av barn och vuxna.
Du kan kontakta rådgivningen via den centraliserade telefontjänsten (06) 826 4477.
Genom regelbundna besök på barnrådgivningsbyrån följs barnets hälsa, tillväxt och utveckling upp.
På rådgivningen vårdas inte barn som insjuknar plötsligt, men du kan be om råd via den centraliserade telefontjänsten (06) 826 4477.
Skolhälsovårdaren har hand om skolelevers hälsa.
Mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats.
Läs mer: Barns hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barnrådgivningarfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Rådgivningarfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Skolhälsovårdfinska _ svenska
Äldre människors hälsa
Vid hälsopunkten Daalia ges vägledning och rådgivning för personer över 65 år om diet, motion och livsstil.
Vaccinering av personer över 65 år utförs vid seniorrådgivning.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Seniorernas hälsopunkterfinska _ svenska
Tandvård
Om du behöver icke-brådskande tandvård ska du ringa munhälsans centraliserade tidsbokningen.
Centraliserad tidsbokning per telefon: (06) 8287 400
Huvudhälsostationens tandklinik
Mariegatan 28, 67200 Karleby
Björkhagens tandklinik
Storkisbackens tandklinik
Korpvägen 11, 67100 Karleby
Kelviå tandklinik
Ellfolkgatan 5, 68300, Kelviå
Lochteå tandklinik
Ullava tandklinik
Ullavavägen 701, 68370 Ullava
Vardagar kan tider till smärtjouren bokas enligt överenskommelse vid samtliga tandkliniker.
Brådskande tandvård/första hjälpen (kvälls-, vardags-, helg- och nattjour):
Vid smärtjouren får du första hjälpen vid plötslig tandvärk och tandolyckor.
Tandläkarjouren (kvälls-, vardags- och helgjour) ordnas vid polikliniken för tand- och munsjukdomar vid Mellersta Österbottens social- och hälsovårdssamkommun Soite, Mariegatan 16–20, 67200 Karleby (vån 1, del D), vardagkvällar kl. 16.00–21.00 samt veckoslut och helgdagar kl. 8.00–21.00.
Du kan i regel komma till jourmottagningen genom att först kontakta jouren via telefon.
För frågor gällande jouren ring tel. (06) 828 7450.
När du kommer till jourmottagningen ska du ta en kölapp, såvida du inte har en bokad tid.
Brådskande tandvård/första hjälpen (nattjour):
Allvarliga fall i samjour Uleåborgs universitetssjukhus (Oulun yliopistollinen sairaala OYS) kl. 21.00−8.00, tel. (08) 315 2655
Läs mer: Tandvård.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Munhälsovårdenfinska _ svenska
Mental hälsa
Vid problem med din mentala hälsa ska du i första hand kontakta din egen hälsostation eller företagshälsovårdens mottagning.
Vid brådskande problem, kontakta hälsovårdcentralens jour.
Läs mer: Mental hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
Sexuell hälsa
Om du känner att du behöver information om familjeplanering och prevention kan du kontakta din egen hälsostation.
Boka tid till hälsostationen om du behöver preventivmedel, överväger att göra en abort eller misstänker att du lider av en könssjukdom.
Du kan även boka en tid hos en allmänläkare för en gynekologisk eller urologisk undersökning.
I preventionsfrågor kan du kontakta den centraliserade telefontjänsten (06) 826 4477.
Läs mer:
Sexuell hälsa och prevention.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Preventivrådgivningfinska _ svenska
När du väntar barn
Ta kontakt med rådgivningen då du märker att du är gravid.
På rådgivningen följer man med moderns, barnets och hela familjens välmående under graviditeten.
Läs mer: Graviditet och förlossning.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Mödrarådgivningfinska _ svenska
Förlossning
Förlossningsavdelningen är öppen dygnet runt.
Om du önskar kan du ringa förlossningsavdelning då din förlossning satt igång eller om du vill fråga om råd.
Då du kommer till sjukhuset ska du använda centralsjukhusets huvudingång kl. 7–20 och övriga tider bör du använda den gemensamma jourens/poliklinikens dörr.
Kontaktuppgifter för förlossningsavdelningen:
Mariegatan 16–20,
67200 Karleby
Telefon: (06) 8264355.
Läs mer: Graviditet och förlossning.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Förlossningarfinska _ svenska
Läkemedel
Du kan köpa läkemedel på apoteket.
Du kan besöka vilket apotek som helst.
Du kan även besöka apotek som inte finns i din egen kommun.
Läs mer: Läkemedel.
Handikappade personer
En handikappad person bosatt i Karleby har rätt att erhålla de tjänster han eller hon behöver på samma grunder som de övriga invånarna i kommunen.
Personen kan dock på grund av sitt handikapp eller sin sjukdom även behöva särskilda tjänster för handikappade för att klara vardagen.
För tjänsterna för handikappade i Karleby svarar Mellersta Österbottens social- och hälsovårdssamkommun Soite, där man kan ansöka om tjänster och stödfunktioner.
Tjänster av flera olika slag erbjuds även för personer med gravt handikapp.
Dessa tjänster inkluderar bland annat:
transporttjänster
ombyggnad och nödvändig utrustning för hemmet
maskiner och utrustning
personlig hjälp och dagverksamhet
stödboende
stöd för närståendevård av personer under 65 och arbetsverksamhet.
Dessutom är det möjligt att ansöka om specialboende, korttidsvård eller tillfällig vård samt handledning hos den öppna vården.
Mer information om tjänster för handikappade får du från Mellersta Österbottens social- och hälsovårdssamkommun Soites handikapptjänster per telefon: 040 804 2122.
Läs mer: Handikappade personer.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Tjänster för handikappadefinska _ svenska
Specialpedagogik i förskolanfinska _ svenska
Kontaktuppgifter för den grundläggande utbildningenfinska
Ett handikappat barn
Särskilt stöd erbjuds barn med handikapp inom småbarnspedagogiken och skolan.
Kontakta Karleby stads förskoleundervisning för information om specialsmåbarnspedagogiken.
Du kan be undervisningsväsendet om mer information om tjänster som skolan erbjuder.
Bildningscentralen
Strandgatan 16 (våning 5 och 6)
67100 Karleby
Telefon: 040 8065 149
Läs mer: Ett handikappat barn.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Tjänster för handikappadefinska _ svenska
Specialpedagogik i förskolanfinska _ svenska
Kontaktuppgifter för den grundläggande utbildningenfinska
Småbarnspedagogik
Förskoleundervisning
Grundläggande utbildning
Undervisning i det egna modersmålet för invandrare
Yrkesutbildning
Gymnasium
Unga utan studieplats
Högskoleutbildning
Andra studiemöjligheter
Småbarnspedagogik
I Karleby finns stadens egna daghem, gruppfamiljedaghem, familjedagvårdare samt barnklubbar.
Dessutom finns det daghem som köptjänst (svenskspråkiga), ett privat daghem och privata familjedagvårdare i Karleby.
Du kan ansöka om plats inom småbarnspedagogiken för ditt barn elektroniskt via tjänsten Suomi.fi eller med en blankett på stadens webbplats (ansökan till småbarnspedagogiken).
Ansökan ska lämnas in fyra månader innan du behöver plats inom småbarnspedagogiken.
Det är möjligt att få en plats snabbare om den behövs för att du exempelvis erhållit arbete eller studieplats.
Ansökan kan returneras till platsen för småbarnspedagogik, kontorstjänster för småbarnspedagogik eller lämnas i brevlådan i den nedre aulan i Bildningscentralen.
Du kan ansöka om en plats i stadens barnklubbar med blanketten som finns på stadens webbplats.
Ansökan kan även skickas per post till följande adress:
Bildningscentralen
Tjänster för småbarnspedagogik
Strandgatan16
67100 Karleby
Läs mer:
Daghem och andra dagvårdsplatserfinska _ svenska
Gruppfamiljedaghemfinska _ svenska
Dagvårdsblanketterfinska _ svenska
Att ansöka om kommunal dagvårdfinska _ svenska
Förskoleundervisning
Karleby stad erbjuder gratis förskoleundervisning för alla 6 år fyllda barn.
Förskoleundervisningen ges av lärare med utbildning i pedagogik i minst 700 timmar om året, dvs. cirka fyra timmar om dagen, enligt skolans arbetstider.
Förskoleundervisningen är gratis.
Om barnet dessutom behöver avgiftsbelagd småbarnspedagogisk verksamhet arrangeras denna på samma ställe som förskoleundervisningen, dock med undantag för skiftesvård.
Anmälningar till förskoleundervisningen sker i januari–februari.
Detta meddelas i lokaltidningarna och på stadens webbplats.
Om du inte fått ett brev om förskoleplats eller ansöker om förskoleplats under annan tid på året, ta kontakt med kontorstjänster för småbarnspedagogik per telefon på numret 040 806 5089.
Läs mer: Förskoleundervisning.
Förskoleundervisningfinska _ svenska
Grundläggande utbildning
I Finland har alla barn som fyllt 7 år läroplikt, vilket innebär att de måste delta i den grundläggande utbildningen.
Läroplikten upphör i slutet av det läsår då barnet fyller 17.
Det är föräldrarna som har ansvaret för att barnet går i skolan.
Anmälan till grundskolan sker i början av året.
På stadens webbplats finns skolornas kontaktuppgifter och mer information om anmälan.
Om du har frågor om den grundläggande utbildningen kan du även kontakta stadens undervisningstjänster.
Varje barn och ung person har rätt att gå i skola.
Om barnet flyttar till Karleby under läsåret kan han eller hon genast börja i skolan.
Om barnet saknar tillräckliga färdigheter i finska eller svenska för att delta i undervisningen i klassen inleder han eller hon studierna i förberedande undervisning i en egen grupp eller i klassen enligt det egna studieprogrammet.
I Karleby finns grupper för den förberedande utbildningen i lågstadiet i Hollihaan koulu och Koivuhaan koulu och i högstadiet i Stenängens skola.
Övergången till den vanliga undervisningen sker steg för steg enligt elevens förutsättningar.
Undervisning i enlighet med lärokursen finska som andra språk och litteratur stödjer en helhetsmässig utveckling av språket.
Stöd för lärande arrangeras i mån av möjlighet på elevens eget modersmål i skolan.
Mer information om den förberedande undervisningen för invandrare får du av stadens undervisningstjänster.
Läs mer: Grundläggande utbildning.
Kontaktuppgifter för den grundläggande utbildningenfinska
Undervisning i det egna modersmålet för invandrare
Undervisning i elevens eget modersmål arrangeras i Karleby på flera olika språk, till exempel under läsåret 2017–2018 arrangerades undervisning på nio olika språk.
Undervisningsgruppen ska ha minst fyra elever.
Undervisningen sker vanligtvis i de skolor där det finns flest elever som talar språket i fråga.
Som elevens egen religion undervisas bland annat islam, buddhism och ortodox religion, beroende på antalet elever.
Information om undervisning i elevens eget modersmål och religion får du av koordinatoren för undervisningen för olika språk- och kulturgrupper:
Tfn 040 489 2129
Utbildning för invandrarefinska
Yrkesutbildning
Mellersta Österbottens yrkesinstitut erbjuder yrkesutbildning i Karleby, Kelviå, Kannus, Kaustby, Perho och Jakobstad.
Yrkesinstitutet anordnar även handledande utbildning för grundläggande yrkesutbildning, dvs. VALMA-utbildning samt förberedande utbildningar för vuxna invandrare vid Mellersta Österbottens folkhögskola i Kelviå.
Läs mer: Yrkesutbildning.
linkkiMellersta Österbottens utbildningskoncern:
Mellersta Österbottens utbildningskoncernfinska _ engelska
linkkiMellersta Österbottens utbildningskoncern:
Utbildning för invandrarefinska _ engelska
linkkiMellersta Österbottens folkhögskola:
Folkhögskolans invandrarlinjefinska
Gymnasium
I Karleby ges gymnasieutbildning för ungdomar vid Karleby finska gymnasium och Karleby svenska gymnasium, samt för vuxna vid Karleby vuxengymnasium.
Till gymnasieutbildning för ungdomar ansöker man under våren via gemensam ansökning för gymnasierna och man kan bli antagen om man i slutbetyget från grundskolan har tillräckligt högt snittbetyg i läsämnena.
Du kan ansöka till vuxenutbildningen direkt hos vuxengymnasiet året runt.
Karleby finska gymnasium erbjuder förberedande undervisning för gymnasiet även för invandrare.
Den förberedande undervisningen för gymnasiet är ett läsår och målet med den är att förbättra möjligheterna för elever med ett annat modersmål att klara av gymnasiestudierna.
Varje år fattas ett skilt beslut om undervisningens start.
För varje studerande utarbetas ett eget studieprogram.
Man ansöker till förberedande undervisning för gymnasiet under sommaren på webbsidan Opintopolku.fi.
Undervisningsspråket i vid Karleby finska gymnasium och Karleby vuxengymnasium är finska och svenska vid Karleby svenska gymnasium.
Vid Karleby finska gymnasium anordnas undervisning i finska som andraspråk för invandrare invandrare.
Målet är att invandrarna ska klara av gymnasiestudierna och efter gymnasiet kunna söka sig till fortsatta studier.
Mer information om gymnasieskolorna och den förberedande undervisningen för gymnasiet fås av stadens undervisningstjänster.
Kontaktuppgifterna för gymnasierna finns på stadens undervisningstjänsters webbplats.
Bildningscentralen
Strandgatan 16 (våning 5 och 6)
67100 Karleby
Telefon: 044 756 7673
Läs mer:
Gymnasium.
Gymnasie- och yrkesutbildningfinska _ svenska
Unga utan studieplats
Unga som saknar studieplats eller arbete kan få hjälp av det uppsökande ungdomsarbetet.
Det uppsökande ungdomsarbetet hjälper unga i åldern 15–28 år hitta rätt tjänster till stöd för utbildning, arbete och utkomst.
De anställda inom uppsökande ungdomsarbete hjälper med att klara upp den ungas livssituation, hantera praktiska ärenden, såsom besök hos olika myndigheter, och ger personlig handledning enligt den ungas önskemål.
Uppsökande ungdomsarbetefinska _ svenska
Högskoleutbildning
Vid Centria yrkeshögskola kan man avlägga högskoleexamen i teknik, företagsekonomi, social- och hälsovård.
Man kan även avlägga en examen inom musikpedagogik och samhällspedagogik.
Det är dessutom möjligt att studera vid den öppna yrkeshögskolan.
Vid Karleby universitetscenter Chydenius kan man avlägga såväl högre högskoleexamen som doktorsexamen.
Vid Chydenius anordnas även vuxenutbildning och vetenskaplig forskning bedrivs.
Läs mer: Högskoleutbildning.
Högskole- och universitetsutbildningfinska
linkkiCentria yrkeshögskola:
Centria yrkeshögskolafinska _ svenska _ engelska
Universitetscentret Chydeniusfinska _ svenska _ engelska
Andra studiemöjligheter
Karlebynejdens institut, som ägs och drivs av Karleby stad, är ett tvåspråkigt (finska och svenska) medborgarinstitut.
Institutet erbjuder undervisning i datateknik, musik, idrott och dans, konstämnen, hantverk, matlagning och första hjälpen.
Institutet erbjuder även undervisning i flera olika språk, bland annat finska, svenska, engelska, tyska, franska, ryska, spanska och italienska.
Undervisningsutbudet varierar från år till år, så det lönar sig att kontrollera aktuella kurser på institutets webbplats.
Invandrare ges rabatt på vissa kurser.
I kursuppgifterna anges om det är möjligt att få rabatt på kursen.
Kontrollera på institutets webbplats vilka kurser som är aktuella.
Vasavägen 7
67100 Karleby
Telefon: 040 8065 169, 040 8065 168
Vid Mellersta Österbottens sommaruniversitet kan du läsa kurser på universitetsnivå vid det öppna universitetet, delta i kompletterande yrkesutbildning samt läsa språk- och kulturkurser.
Under sommaren är det möjligt att repetera gymnasiestudier vid sommaruniversitetet.
Dessutom är det även möjligt att läsa normala gymnasiekurser vid sommaruniversitetets sommargymnasium.
Sommaruniversitets kurser är avgiftsbelagda för deltagarna.
Läs mer:
Studier som hobby, Arbetskraftsutbildning
Karlebynejdens institutfinska _ svenska
linkkiArbets- och näringsbyråns tjänster:
Offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiMellersta Österbottens sommaruniversitet:
Mellersta Österbottens sommaruniversitetfinska
Övrig undervisning i Karlebyfinska _ svenska
Småbarnspedagogik
Förskoleundervisning
Grundläggande utbildning
Undervisning i det egna modersmålet för invandrare
Yrkesutbildning
Gymnasium
Unga utan studieplats
Högskoleutbildning
Andra studiemöjligheter
Småbarnspedagogik
I Karleby finns stadens egna daghem, gruppfamiljedaghem, familjedagvårdare samt barnklubbar.
Dessutom finns det daghem som köptjänst (svenskspråkiga), ett privat daghem och privata familjedagvårdare i Karleby.
Du kan ansöka om plats inom småbarnspedagogiken för ditt barn elektroniskt via tjänsten Suomi.fi eller med en blankett på stadens webbplats (ansökan till småbarnspedagogiken).
Ansökan ska lämnas in fyra månader innan du behöver plats inom småbarnspedagogiken.
Det är möjligt att få en plats snabbare om den behövs för att du exempelvis erhållit arbete eller studieplats.
Ansökan kan returneras till platsen för småbarnspedagogik, kontorstjänster för småbarnspedagogik eller lämnas i brevlådan i den nedre aulan i Bildningscentralen.
Du kan ansöka om en plats i stadens barnklubbar med blanketten som finns på stadens webbplats.
Ansökan kan även skickas per post till följande adress:
Bildningscentralen
Tjänster för småbarnspedagogik
Strandgatan16
67100 Karleby
Läs mer:
Daghem och andra dagvårdsplatserfinska _ svenska
Gruppfamiljedaghemfinska _ svenska
Dagvårdsblanketterfinska _ svenska
Att ansöka om kommunal dagvårdfinska _ svenska
Förskoleundervisning
Karleby stad erbjuder gratis förskoleundervisning för alla 6 år fyllda barn.
Förskoleundervisningen ges av lärare med utbildning i pedagogik i minst 700 timmar om året, dvs. cirka fyra timmar om dagen, enligt skolans arbetstider.
Förskoleundervisningen är gratis.
Om barnet dessutom behöver avgiftsbelagd småbarnspedagogisk verksamhet arrangeras denna på samma ställe som förskoleundervisningen, dock med undantag för skiftesvård.
Anmälningar till förskoleundervisningen sker i januari–februari.
Detta meddelas i lokaltidningarna och på stadens webbplats.
Om du inte fått ett brev om förskoleplats eller ansöker om förskoleplats under annan tid på året, ta kontakt med kontorstjänster för småbarnspedagogik per telefon på numret 040 806 5089.
Läs mer: Förskoleundervisning.
Förskoleundervisningfinska _ svenska
Grundläggande utbildning
I Finland har alla barn som fyllt 7 år läroplikt, vilket innebär att de måste delta i den grundläggande utbildningen.
Läroplikten upphör i slutet av det läsår då barnet fyller 17.
Det är föräldrarna som har ansvaret för att barnet går i skolan.
Anmälan till grundskolan sker i början av året.
På stadens webbplats finns skolornas kontaktuppgifter och mer information om anmälan.
Om du har frågor om den grundläggande utbildningen kan du även kontakta stadens undervisningstjänster.
Varje barn och ung person har rätt att gå i skola.
Om barnet flyttar till Karleby under läsåret kan han eller hon genast börja i skolan.
Om barnet saknar tillräckliga färdigheter i finska eller svenska för att delta i undervisningen i klassen inleder han eller hon studierna i förberedande undervisning i en egen grupp eller i klassen enligt det egna studieprogrammet.
I Karleby finns grupper för den förberedande utbildningen i lågstadiet i Hollihaan koulu och Koivuhaan koulu och i högstadiet i Stenängens skola.
Övergången till den vanliga undervisningen sker steg för steg enligt elevens förutsättningar.
Undervisning i enlighet med lärokursen finska som andra språk och litteratur stödjer en helhetsmässig utveckling av språket.
Stöd för lärande arrangeras i mån av möjlighet på elevens eget modersmål i skolan.
Mer information om den förberedande undervisningen för invandrare får du av stadens undervisningstjänster.
Läs mer: Grundläggande utbildning.
Kontaktuppgifter för den grundläggande utbildningenfinska
Undervisning i det egna modersmålet för invandrare
Undervisning i elevens eget modersmål arrangeras i Karleby på flera olika språk, till exempel under läsåret 2017–2018 arrangerades undervisning på nio olika språk.
Undervisningsgruppen ska ha minst fyra elever.
Undervisningen sker vanligtvis i de skolor där det finns flest elever som talar språket i fråga.
Som elevens egen religion undervisas bland annat islam, buddhism och ortodox religion, beroende på antalet elever.
Information om undervisning i elevens eget modersmål och religion får du av koordinatoren för undervisningen för olika språk- och kulturgrupper:
Tfn 040 489 2129
Utbildning för invandrarefinska
Yrkesutbildning
Mellersta Österbottens yrkesinstitut erbjuder yrkesutbildning i Karleby, Kelviå, Kannus, Kaustby, Perho och Jakobstad.
Yrkesinstitutet anordnar även handledande utbildning för grundläggande yrkesutbildning, dvs. VALMA-utbildning samt förberedande utbildningar för vuxna invandrare vid Mellersta Österbottens folkhögskola i Kelviå.
Läs mer: Yrkesutbildning.
linkkiMellersta Österbottens utbildningskoncern:
Mellersta Österbottens utbildningskoncernfinska _ engelska
linkkiMellersta Österbottens utbildningskoncern:
Utbildning för invandrarefinska _ engelska
linkkiMellersta Österbottens folkhögskola:
Folkhögskolans invandrarlinjefinska
Gymnasium
I Karleby ges gymnasieutbildning för ungdomar vid Karleby finska gymnasium och Karleby svenska gymnasium, samt för vuxna vid Karleby vuxengymnasium.
Till gymnasieutbildning för ungdomar ansöker man under våren via gemensam ansökning för gymnasierna och man kan bli antagen om man i slutbetyget från grundskolan har tillräckligt högt snittbetyg i läsämnena.
Du kan ansöka till vuxenutbildningen direkt hos vuxengymnasiet året runt.
Karleby finska gymnasium erbjuder förberedande undervisning för gymnasiet även för invandrare.
Den förberedande undervisningen för gymnasiet är ett läsår och målet med den är att förbättra möjligheterna för elever med ett annat modersmål att klara av gymnasiestudierna.
Varje år fattas ett skilt beslut om undervisningens start.
För varje studerande utarbetas ett eget studieprogram.
Man ansöker till förberedande undervisning för gymnasiet under sommaren på webbsidan Opintopolku.fi.
Undervisningsspråket i vid Karleby finska gymnasium och Karleby vuxengymnasium är finska och svenska vid Karleby svenska gymnasium.
Vid Karleby finska gymnasium anordnas undervisning i finska som andraspråk för invandrare invandrare.
Målet är att invandrarna ska klara av gymnasiestudierna och efter gymnasiet kunna söka sig till fortsatta studier.
Mer information om gymnasieskolorna och den förberedande undervisningen för gymnasiet fås av stadens undervisningstjänster.
Kontaktuppgifterna för gymnasierna finns på stadens undervisningstjänsters webbplats.
Bildningscentralen
Strandgatan 16 (våning 5 och 6)
67100 Karleby
Telefon: 044 756 7673
Läs mer:
Gymnasium.
Gymnasie- och yrkesutbildningfinska _ svenska
Unga utan studieplats
Unga som saknar studieplats eller arbete kan få hjälp av det uppsökande ungdomsarbetet.
Det uppsökande ungdomsarbetet hjälper unga i åldern 15–28 år hitta rätt tjänster till stöd för utbildning, arbete och utkomst.
De anställda inom uppsökande ungdomsarbete hjälper med att klara upp den ungas livssituation, hantera praktiska ärenden, såsom besök hos olika myndigheter, och ger personlig handledning enligt den ungas önskemål.
Uppsökande ungdomsarbetefinska _ svenska
Högskoleutbildning
Vid Centria yrkeshögskola kan man avlägga högskoleexamen i teknik, företagsekonomi, social- och hälsovård.
Man kan även avlägga en examen inom musikpedagogik och samhällspedagogik.
Det är dessutom möjligt att studera vid den öppna yrkeshögskolan.
Vid Karleby universitetscenter Chydenius kan man avlägga såväl högre högskoleexamen som doktorsexamen.
Vid Chydenius anordnas även vuxenutbildning och vetenskaplig forskning bedrivs.
Läs mer: Högskoleutbildning.
Högskole- och universitetsutbildningfinska
linkkiCentria yrkeshögskola:
Centria yrkeshögskolafinska _ svenska _ engelska
Universitetscentret Chydeniusfinska _ svenska _ engelska
Andra studiemöjligheter
Karlebynejdens institut, som ägs och drivs av Karleby stad, är ett tvåspråkigt (finska och svenska) medborgarinstitut.
Institutet erbjuder undervisning i datateknik, musik, idrott och dans, konstämnen, hantverk, matlagning och första hjälpen.
Institutet erbjuder även undervisning i flera olika språk, bland annat finska, svenska, engelska, tyska, franska, ryska, spanska och italienska.
Undervisningsutbudet varierar från år till år, så det lönar sig att kontrollera aktuella kurser på institutets webbplats.
Invandrare ges rabatt på vissa kurser.
I kursuppgifterna anges om det är möjligt att få rabatt på kursen.
Kontrollera på institutets webbplats vilka kurser som är aktuella.
Vasavägen 7
67100 Karleby
Telefon: 040 8065 169, 040 8065 168
Vid Mellersta Österbottens sommaruniversitet kan du läsa kurser på universitetsnivå vid det öppna universitetet, delta i kompletterande yrkesutbildning samt läsa språk- och kulturkurser.
Under sommaren är det möjligt att repetera gymnasiestudier vid sommaruniversitetet.
Dessutom är det även möjligt att läsa normala gymnasiekurser vid sommaruniversitetets sommargymnasium.
Sommaruniversitets kurser är avgiftsbelagda för deltagarna.
Läs mer:
Studier som hobby, Arbetskraftsutbildning
Karlebynejdens institutfinska _ svenska
linkkiArbets- och näringsbyråns tjänster:
Offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiMellersta Österbottens sommaruniversitet:
Mellersta Österbottens sommaruniversitetfinska
Övrig undervisning i Karlebyfinska _ svenska
Småbarnspedagogik
Förskoleundervisning
Grundläggande utbildning
Undervisning i det egna modersmålet för invandrare
Yrkesutbildning
Gymnasium
Unga utan studieplats
Högskoleutbildning
Andra studiemöjligheter
Småbarnspedagogik
I Karleby finns stadens egna daghem, gruppfamiljedaghem, familjedagvårdare samt barnklubbar.
Dessutom finns det daghem som köptjänst (svenskspråkiga), ett privat daghem och privata familjedagvårdare i Karleby.
Du kan ansöka om plats inom småbarnspedagogiken för ditt barn elektroniskt via tjänsten Suomi.fi eller med en blankett på stadens webbplats (ansökan till småbarnspedagogiken).
Ansökan ska lämnas in fyra månader innan du behöver plats inom småbarnspedagogiken.
Det är möjligt att få en plats snabbare om den behövs för att du exempelvis erhållit arbete eller studieplats.
Ansökan kan returneras till platsen för småbarnspedagogik, kontorstjänster för småbarnspedagogik eller lämnas i brevlådan i den nedre aulan i Bildningscentralen.
Du kan ansöka om en plats i stadens barnklubbar med blanketten som finns på stadens webbplats.
Ansökan kan även skickas per post till följande adress:
Bildningscentralen
Tjänster för småbarnspedagogik
Strandgatan16
67100 Karleby
Läs mer:
Småbarnspedagogik.
Daghem och andra dagvårdsplatserfinska _ svenska
Gruppfamiljedaghemfinska _ svenska
Dagvårdsblanketterfinska _ svenska
Att ansöka om kommunal dagvårdfinska _ svenska
Förskoleundervisning
Karleby stad erbjuder gratis förskoleundervisning för alla 6 år fyllda barn.
Förskoleundervisningen ges av lärare med utbildning i pedagogik i minst 700 timmar om året, dvs. cirka fyra timmar om dagen, enligt skolans arbetstider.
Förskoleundervisningen är gratis.
Om barnet dessutom behöver avgiftsbelagd småbarnspedagogisk verksamhet arrangeras denna på samma ställe som förskoleundervisningen, dock med undantag för skiftesvård.
Anmälningar till förskoleundervisningen sker i januari–februari.
Detta meddelas i lokaltidningarna och på stadens webbplats.
Om du inte fått ett brev om förskoleplats eller ansöker om förskoleplats under annan tid på året, ta kontakt med kontorstjänster för småbarnspedagogik per telefon på numret 040 806 5089.
Läs mer: Förskoleundervisning.
Förskoleundervisningfinska _ svenska
Grundläggande utbildning
I Finland har alla barn som fyllt 7 år läroplikt, vilket innebär att de måste delta i den grundläggande utbildningen.
Läroplikten upphör i slutet av det läsår då barnet fyller 17.
Det är föräldrarna som har ansvaret för att barnet går i skolan.
Anmälan till grundskolan sker i början av året.
På stadens webbplats finns skolornas kontaktuppgifter och mer information om anmälan.
Om du har frågor om den grundläggande utbildningen kan du även kontakta stadens undervisningstjänster.
Varje barn och ung person har rätt att gå i skola.
Om barnet flyttar till Karleby under läsåret kan han eller hon genast börja i skolan.
Om barnet saknar tillräckliga färdigheter i finska eller svenska för att delta i undervisningen i klassen inleder han eller hon studierna i förberedande undervisning i en egen grupp eller i klassen enligt det egna studieprogrammet.
I Karleby finns grupper för den förberedande utbildningen i lågstadiet i Hollihaan koulu och Koivuhaan koulu och i högstadiet i Stenängens skola.
Övergången till den vanliga undervisningen sker steg för steg enligt elevens förutsättningar.
Undervisning i enlighet med lärokursen finska som andra språk och litteratur stödjer en helhetsmässig utveckling av språket.
Stöd för lärande arrangeras i mån av möjlighet på elevens eget modersmål i skolan.
Mer information om den förberedande undervisningen för invandrare får du av stadens undervisningstjänster.
Läs mer: Grundläggande utbildning.
Kontaktuppgifter för den grundläggande utbildningenfinska
Undervisning i det egna modersmålet för invandrare
Undervisning i elevens eget modersmål arrangeras i Karleby på flera olika språk, till exempel under läsåret 2017–2018 arrangerades undervisning på nio olika språk.
Undervisningsgruppen ska ha minst fyra elever.
Undervisningen sker vanligtvis i de skolor där det finns flest elever som talar språket i fråga.
Som elevens egen religion undervisas bland annat islam, buddhism och ortodox religion, beroende på antalet elever.
Information om undervisning i elevens eget modersmål och religion får du av koordinatoren för undervisningen för olika språk- och kulturgrupper:
Tfn 040 489 2129
Utbildning för invandrarefinska
Yrkesutbildning
Mellersta Österbottens yrkesinstitut erbjuder yrkesutbildning i Karleby, Kelviå, Kannus, Kaustby, Perho och Jakobstad.
Yrkesinstitutet anordnar även handledande utbildning för grundläggande yrkesutbildning, dvs. VALMA-utbildning samt förberedande utbildningar för vuxna invandrare vid Mellersta Österbottens folkhögskola i Kelviå.
Läs mer: Yrkesutbildning.
linkkiMellersta Österbottens utbildningskoncern:
Mellersta Österbottens utbildningskoncernfinska _ engelska
linkkiMellersta Österbottens utbildningskoncern:
Utbildning för invandrarefinska _ engelska
linkkiMellersta Österbottens folkhögskola:
Folkhögskolans invandrarlinjefinska
Gymnasium
I Karleby ges gymnasieutbildning för ungdomar vid Karleby finska gymnasium och Karleby svenska gymnasium, samt för vuxna vid Karleby vuxengymnasium.
Till gymnasieutbildning för ungdomar ansöker man under våren via gemensam ansökning för gymnasierna och man kan bli antagen om man i slutbetyget från grundskolan har tillräckligt högt snittbetyg i läsämnena.
Du kan ansöka till vuxenutbildningen direkt hos vuxengymnasiet året runt.
Karleby finska gymnasium erbjuder förberedande undervisning för gymnasiet även för invandrare.
Den förberedande undervisningen för gymnasiet är ett läsår och målet med den är att förbättra möjligheterna för elever med ett annat modersmål att klara av gymnasiestudierna.
Varje år fattas ett skilt beslut om undervisningens start.
För varje studerande utarbetas ett eget studieprogram.
Man ansöker till förberedande undervisning för gymnasiet under sommaren på webbsidan Opintopolku.fi.
Undervisningsspråket i vid Karleby finska gymnasium och Karleby vuxengymnasium är finska och svenska vid Karleby svenska gymnasium.
Vid Karleby finska gymnasium anordnas undervisning i finska som andraspråk för invandrare invandrare.
Målet är att invandrarna ska klara av gymnasiestudierna och efter gymnasiet kunna söka sig till fortsatta studier.
Mer information om gymnasieskolorna och den förberedande undervisningen för gymnasiet fås av stadens undervisningstjänster.
Kontaktuppgifterna för gymnasierna finns på stadens undervisningstjänsters webbplats.
Bildningscentralen
Strandgatan 16 (våning 5 och 6)
67100 Karleby
Telefon: 044 756 7673
Läs mer:
Gymnasium.
Gymnasie- och yrkesutbildningfinska _ svenska
Unga utan studieplats
Unga som saknar studieplats eller arbete kan få hjälp av det uppsökande ungdomsarbetet.
Det uppsökande ungdomsarbetet hjälper unga i åldern 15–28 år hitta rätt tjänster till stöd för utbildning, arbete och utkomst.
De anställda inom uppsökande ungdomsarbete hjälper med att klara upp den ungas livssituation, hantera praktiska ärenden, såsom besök hos olika myndigheter, och ger personlig handledning enligt den ungas önskemål.
Uppsökande ungdomsarbetefinska _ svenska
Högskoleutbildning
Vid Centria yrkeshögskola kan man avlägga högskoleexamen i teknik, företagsekonomi, social- och hälsovård.
Man kan även avlägga en examen inom musikpedagogik och samhällspedagogik.
Det är dessutom möjligt att studera vid den öppna yrkeshögskolan.
Vid Karleby universitetscenter Chydenius kan man avlägga såväl högre högskoleexamen som doktorsexamen.
Vid Chydenius anordnas även vuxenutbildning och vetenskaplig forskning bedrivs.
Läs mer:
Yrkeshögskolor, Universitet.
Högskole- och universitetsutbildningfinska
linkkiCentria yrkeshögskola:
Centria yrkeshögskolafinska _ svenska _ engelska
Universitetscentret Chydeniusfinska _ svenska _ engelska
Andra studiemöjligheter
Karlebynejdens institut, som ägs och drivs av Karleby stad, är ett tvåspråkigt (finska och svenska) medborgarinstitut.
Institutet erbjuder undervisning i datateknik, musik, idrott och dans, konstämnen, hantverk, matlagning och första hjälpen.
Institutet erbjuder även undervisning i flera olika språk, bland annat finska, svenska, engelska, tyska, franska, ryska, spanska och italienska.
Undervisningsutbudet varierar från år till år, så det lönar sig att kontrollera aktuella kurser på institutets webbplats.
Invandrare ges rabatt på vissa kurser.
I kursuppgifterna anges om det är möjligt att få rabatt på kursen.
Kontrollera på institutets webbplats vilka kurser som är aktuella.
Vasavägen 7
67100 Karleby
Telefon: 040 8065 169, 040 8065 168
Vid Mellersta Österbottens sommaruniversitet kan du läsa kurser på universitetsnivå vid det öppna universitetet, delta i kompletterande yrkesutbildning samt läsa språk- och kulturkurser.
Under sommaren är det möjligt att repetera gymnasiestudier vid sommaruniversitetet.
Dessutom är det även möjligt att läsa normala gymnasiekurser vid sommaruniversitetets sommargymnasium.
Sommaruniversitets kurser är avgiftsbelagda för deltagarna.
Läs mer:
Studier som hobby, Arbetskraftsutbildning
Karlebynejdens institutfinska _ svenska
linkkiArbets- och näringsbyråns tjänster:
Offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiMellersta Österbottens sommaruniversitet:
Mellersta Österbottens sommaruniversitetfinska
Övrig undervisning i Karlebyfinska _ svenska
Hyresbostad
Ägarbostad
Tillfälligt boende
Stöd- och serviceboende
Bostadslöshet
Avfallshantering för bostaden
Hyresbostad
Karleby stads blankett för ansökan om hyresbostad kan fyllas i och skickas in på nätet.
Bilagor till ansökningen ska tillhandahållas då bostad erbjuds, men kan även lämnas in tidigare.
Man kan även lämna in bostadsansökan på papper.
Ansökningsblanketterna kan hämtas från och lämnas in till Kokkolan Vuokra Asunnot Oy:s verksamhetsställen.
67800 Karleby
Telefon: 040 1817 400
Studiebostäder hyrs ut av Kiinteistöyhtiö Tankkari, som erbjuder möblerade kollektivbostäder samt familjebostäder i olika storlek.
En familjebostad är en omöblerad lägenhet som endast hyrs ut till personer i samma hushåll.
Såväl individer som sambor/gifta par kan ansöka om en hyresetta.
Bondegatan 2
67100 Karleby
Telefon: 040 193 6468
Läs mer:
Hyresbostad.
Hyresbostäderfinska _ svenska
Ansökan om Karleby stads hyresbostadfinska _ svenska _ engelska
Hyresbostäder enligt stadsdelfinska _ svenska
Studiebostäderfinska _ engelska
Privata hyresbostäderfinska _ svenska
Ägarbostad
De flesta finländarna bor i en ägarbostad, alltså i en bostad som de själva äger.
På lång sikt är det ofta förmånligare att köpa sin egen bostad än att hyra.
Bland annat hos bostadsförmedlingen, på internet och i lokala tidningar finns annonser om bostäder som är till salu.
Läs mer:
Ägarbostad.
Tillfälligt boende
I Karlebynejden erbjuds olika inkvarteringsalternativ.
Kontaktuppgifterna finns under länkarna nedan.
Läs mer:
Tillfälligt boende.
Övernattningsalternativ i Karlebyfinska _ svenska _ engelska
Om du saknar boende på grund av kris eller olycka ska du kontakta Kokkolan Vuokra Asunnot Oy eller bostadsbyrån.
Om din bostad har skadats, till exempel till följd av brand eller vattenskada, kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
Kontakta ditt försäkringsbolag direkt när skadan har inträffat.
Om en familjemedlem är våldsam eller hotar med våld, ta kontakt med Karleby mödra- och skyddshem.
Du kan ringa skyddshemmet under alla tider på dygnet.
Du behöver inte uppge ditt namn då du ringer.
Karleby mödra- och skyddshem
Telefon: 044 336 0056
Hyresbostäderfinska _ svenska
Karleby mödra- och skyddshemfinska
Stöd- och serviceboende
Äldre människor erbjuds boendeservice anordnad av Mellersta Österbottens social- och hälsovårdssamkommun Soite samt privata servicebostäder.
Serviceboende för äldre är avsett för personer över 65 år som behöver vård och omsorg dygnet runt.
Serviceboende är lämpat för personer som inte längre klarar sig på egen hand med tjänster som tillhandahålls i hemmet.
Mer information om boendeservice anordnad av Mellersta Österbottens social- och hälsovårdssamkommun Soite får du av bland annat samkommunens servicestyrcentral, tfn 040 806 5093.
För handikappade och personer som återhämtar sig från mentala problem erbjuds bostäder som beaktar invånarnas särskilda behov.
Hemvårdens stödtjänster erbjuds personer som har svårigheter med att klara vardagen utan hjälp, såsom äldre och handikappade personer.
Tjänster av detta slag är bland annat måltidstjänst och transporttjänst.
Målet med hemvården är att erbjuda trygg vård och omsorg samt främja invånarnas ork, handlingskraft och företagsamhet.
Läs mer:
Stöd- och serviceboende.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Servicehandledningscentretfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Seniorernas tjänster, hemvårdfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Seniorernas tjänster, serviceboendet och anstaltsvårdenfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Boendetjänster för utvecklingsstörda och handikappadefinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Socialrådgivningfinska _ svenska
Bostadslöshet
Om du blir bostadslös bör du kontakta Kokkolan Vuokra Asunnot Oy eller bostadsbyrån.
Hyresbostäderfinska _ svenska
Avfallshantering för bostaden
Med bioavfall avses bl.a.:
matrester
skämda och torra livsmedel
skal från frukt och grönsaker
Separat insamlat bioavfall packas i en papperspåse, en påse vikt av en dagstidning eller en plastkasse. Kassen eller påsen får vara högst 30l stor.
En full sopsäck ska tillslutas noggrant.
Med energiavfall avses bl.a.:
bakplåtspapper, hushållspapper och våtservetter
kläder (inte skor, regnställ eller läderplagg)
små plastleksaker och bruksföremål i plast såsom disk- och tandborstar.
Separat insamlat energiavfall ska packas i plastkasse eller papperspåsar.
Kassen eller påsen får vara högst 30 l stor.
Påsen tillsluts noga.
Avfall som inte får läggas i det egna husets sopbehållare kan föras till återvinningsstationer.
Kontrollera på förhand vilken typ av avfall stationen tar emot.
Mer information om avfallshanteringen i Karlebynejden finns på Karleby stads och på Ab Ekorosk Oy:s (kommunalt avfallshanteringsbolag) webbplats.
Läs mer: Avfallshantering och återvinning.
Avfallshantering för bostaden finska _ svenska
Ett kommunalt avfallshanteringsbolagfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ vietnamesiska _ polska _ kroatiska
Hyresbostad
Köpa bostad
Tillfälligt boende
Stöd- och serviceboende
Bostadslöshet
Avfallshantering för bostaden
Hyresbostad
Karleby stads blankett för ansökan om hyresbostad kan fyllas i och skickas in på nätet.
Bilagor till ansökningen ska tillhandahållas då bostad erbjuds, men kan även lämnas in tidigare.
Man kan även lämna in bostadsansökan på papper.
Ansökningsblanketterna kan hämtas från och lämnas in till Kokkolan Vuokra Asunnot Oy:s verksamhetsställen.
67800 Karleby
Telefon: 040 1817 400
Studiebostäder hyrs ut av Kiinteistöyhtiö Tankkari, som erbjuder möblerade kollektivbostäder samt familjebostäder i olika storlek.
En familjebostad är en omöblerad lägenhet som endast hyrs ut till personer i samma hushåll.
Såväl individer som sambor/gifta par kan ansöka om en hyresetta.
Bondegatan 2
67100 Karleby
Telefon: 040 193 6468
Läs mer: Hyresbostad.
Hyresbostäderfinska _ svenska
Ansökan om Karleby stads hyresbostadfinska _ svenska _ engelska
Hyresbostäder enligt stadsdelfinska _ svenska
Studiebostäderfinska _ engelska
Privata hyresbostäderfinska _ svenska
Köpa bostad
De flesta finländarna bor i en ägarbostad, alltså i en bostad som de själva äger.
På lång sikt är det ofta förmånligare att köpa sin egen bostad än att hyra.
Bland annat hos bostadsförmedlingen, på internet och i lokala tidningar finns annonser om bostäder som är till salu.
Läs mer: Köpa bostad.
Tillfälligt boende
I Karlebynejden erbjuds olika inkvarteringsalternativ.
Kontaktuppgifterna finns under länkarna nedan.
Läs mer:
Tillfälligt boende.
Övernattningsalternativ i Karlebyfinska _ svenska _ engelska
Om du saknar boende på grund av kris eller olycka ska du kontakta Kokkolan Vuokra Asunnot Oy eller bostadsbyrån.
Om din bostad har skadats, till exempel till följd av brand eller vattenskada, kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
Kontakta ditt försäkringsbolag direkt när skadan har inträffat.
Om en familjemedlem är våldsam eller hotar med våld, ta kontakt med Karleby mödra- och skyddshem.
Du kan ringa skyddshemmet under alla tider på dygnet.
Du behöver inte uppge ditt namn då du ringer.
Karleby mödra- och skyddshem
Telefon: 044 336 0056
Läs mer: Boende.
Hyresbostäderfinska _ svenska
Karleby mödra- och skyddshemfinska
Stöd- och serviceboende
Äldre människor erbjuds boendeservice anordnad av Mellersta Österbottens social- och hälsovårdssamkommun Soite samt privata servicebostäder.
Serviceboende för äldre är avsett för personer över 65 år som behöver vård och omsorg dygnet runt.
Serviceboende är lämpat för personer som inte längre klarar sig på egen hand med tjänster som tillhandahålls i hemmet.
Mer information om boendeservice anordnad av Mellersta Österbottens social- och hälsovårdssamkommun Soite får du av bland annat samkommunens servicestyrcentral, tfn 040 806 5093.
För handikappade och personer som återhämtar sig från mentala problem erbjuds bostäder som beaktar invånarnas särskilda behov.
Hemvårdens stödtjänster erbjuds personer som har svårigheter med att klara vardagen utan hjälp, såsom äldre och handikappade personer.
Tjänster av detta slag är bland annat måltidstjänst och transporttjänst.
Målet med hemvården är att erbjuda trygg vård och omsorg samt främja invånarnas ork, handlingskraft och företagsamhet.
Läs mer:
Stöd- och serviceboende.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Servicehandledningscentretfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Seniorernas tjänster, hemvårdfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Seniorernas tjänster, serviceboendet och anstaltsvårdenfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Boendetjänster för utvecklingsstörda och handikappadefinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Socialrådgivningfinska _ svenska
Bostadslöshet
Om du blir bostadslös bör du kontakta Kokkolan Vuokra Asunnot Oy eller bostadsbyrån.
Läs mer: Bostadslöshet.
Hyresbostäderfinska _ svenska
Avfallshantering för bostaden
Med bioavfall avses bl.a.:
matrester
skämda och torra livsmedel
skal från frukt och grönsaker
Separat insamlat bioavfall packas i en papperspåse, en påse vikt av en dagstidning eller en plastkasse. Kassen eller påsen får vara högst 30l stor.
En full sopsäck ska tillslutas noggrant.
Med energiavfall avses bl.a.:
bakplåtspapper, hushållspapper och våtservetter
kläder (inte skor, regnställ eller läderplagg)
små plastleksaker och bruksföremål i plast såsom disk- och tandborstar.
Separat insamlat energiavfall ska packas i plastkasse eller papperspåsar.
Kassen eller påsen får vara högst 30 l stor.
Påsen tillsluts noga.
Avfall som inte får läggas i det egna husets sopbehållare kan föras till återvinningsstationer.
Kontrollera på förhand vilken typ av avfall stationen tar emot.
Mer information om avfallshanteringen i Karlebynejden finns på Karleby stads och på Ab Ekorosk Oy:s (kommunalt avfallshanteringsbolag) webbplats.
Läs mer: Avfallshantering och återvinning.
Avfallshantering för bostaden finska _ svenska
Ett kommunalt avfallshanteringsbolagfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ vietnamesiska _ polska _ kroatiska
Hyresbostad
Köpa bostad
Tillfälligt boende
Stöd- och serviceboende
Bostadslöshet
Avfallshantering för bostaden
Hyresbostad
Karleby stads blankett för ansökan om hyresbostad kan fyllas i och skickas in på nätet.
Bilagor till ansökningen ska tillhandahållas då bostad erbjuds, men kan även lämnas in tidigare.
Man kan även lämna in bostadsansökan på papper.
Ansökningsblanketterna kan hämtas från och lämnas in till Kokkolan Vuokra Asunnot Oy:s verksamhetsställen.
67800 Karleby
Telefon: 040 1817 400
Studiebostäder hyrs ut av Kiinteistöyhtiö Tankkari, som erbjuder möblerade kollektivbostäder samt familjebostäder i olika storlek.
En familjebostad är en omöblerad lägenhet som endast hyrs ut till personer i samma hushåll.
Såväl individer som sambor/gifta par kan ansöka om en hyresetta.
Bondegatan 2
67100 Karleby
Telefon: 040 193 6468
Läs mer: Hyresbostad.
Hyresbostäderfinska _ svenska
Ansökan om Karleby stads hyresbostadfinska _ svenska _ engelska
Hyresbostäder enligt stadsdelfinska _ svenska
Studiebostäderfinska _ engelska
Privata hyresbostäderfinska _ svenska
Köpa bostad
De flesta finländarna bor i en ägarbostad, alltså i en bostad som de själva äger.
På lång sikt är det ofta förmånligare att köpa sin egen bostad än att hyra.
Bland annat hos bostadsförmedlingen, på internet och i lokala tidningar finns annonser om bostäder som är till salu.
Läs mer: Köpa bostad.
Tillfälligt boende
I Karlebynejden erbjuds olika inkvarteringsalternativ.
Kontaktuppgifterna finns under länkarna nedan.
Läs mer:
Tillfälligt boende.
Övernattningsalternativ i Karlebyfinska _ svenska _ engelska
Om du saknar boende på grund av kris eller olycka ska du kontakta Kokkolan Vuokra Asunnot Oy eller bostadsbyrån.
Om din bostad har skadats, till exempel till följd av brand eller vattenskada, kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
Kontakta ditt försäkringsbolag direkt när skadan har inträffat.
Om en familjemedlem är våldsam eller hotar med våld, ta kontakt med Karleby mödra- och skyddshem.
Du kan ringa skyddshemmet under alla tider på dygnet.
Du behöver inte uppge ditt namn då du ringer.
Karleby mödra- och skyddshem
Telefon: 044 336 0056
Läs mer: Boende.
Hyresbostäderfinska _ svenska
Karleby mödra- och skyddshemfinska
Stöd- och serviceboende
Äldre människor erbjuds boendeservice anordnad av Mellersta Österbottens social- och hälsovårdssamkommun Soite samt privata servicebostäder.
Serviceboende för äldre är avsett för personer över 65 år som behöver vård och omsorg dygnet runt.
Serviceboende är lämpat för personer som inte längre klarar sig på egen hand med tjänster som tillhandahålls i hemmet.
Mer information om boendeservice anordnad av Mellersta Österbottens social- och hälsovårdssamkommun Soite får du av bland annat samkommunens servicestyrcentral, tfn 040 806 5093.
För handikappade och personer som återhämtar sig från mentala problem erbjuds bostäder som beaktar invånarnas särskilda behov.
Hemvårdens stödtjänster erbjuds personer som har svårigheter med att klara vardagen utan hjälp, såsom äldre och handikappade personer.
Tjänster av detta slag är bland annat måltidstjänst och transporttjänst.
Målet med hemvården är att erbjuda trygg vård och omsorg samt främja invånarnas ork, handlingskraft och företagsamhet.
Läs mer:
Stöd- och serviceboende.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Servicehandledningscentretfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Seniorernas tjänster, hemvårdfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Seniorernas tjänster, serviceboendet och anstaltsvårdenfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Boendetjänster för utvecklingsstörda och handikappadefinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Socialrådgivningfinska _ svenska
Bostadslöshet
Om du blir bostadslös bör du kontakta Kokkolan Vuokra Asunnot Oy eller bostadsbyrån.
Läs mer: Bostadslöshet.
Hyresbostäderfinska _ svenska
Avfallshantering för bostaden
Med bioavfall avses bl.a.:
matrester
skämda och torra livsmedel
skal från frukt och grönsaker
Separat insamlat bioavfall packas i en papperspåse, en påse vikt av en dagstidning eller en plastkasse. Kassen eller påsen får vara högst 30l stor.
En full sopsäck ska tillslutas noggrant.
Med energiavfall avses bl.a.:
bakplåtspapper, hushållspapper och våtservetter
kläder (inte skor, regnställ eller läderplagg)
små plastleksaker och bruksföremål i plast såsom disk- och tandborstar.
Separat insamlat energiavfall ska packas i plastkasse eller papperspåsar.
Kassen eller påsen får vara högst 30 l stor.
Påsen tillsluts noga.
Avfall som inte får läggas i det egna husets sopbehållare kan föras till återvinningsstationer.
Kontrollera på förhand vilken typ av avfall stationen tar emot.
Mer information om avfallshanteringen i Karlebynejden finns på Karleby stads och på Ab Ekorosk Oy:s (kommunalt avfallshanteringsbolag) webbplats.
Läs mer: Avfallshantering och återvinning.
Avfallshantering för bostaden finska _ svenska
Ett kommunalt avfallshanteringsbolagfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ vietnamesiska _ polska _ kroatiska
Möjligheter att studera finska eller svenska
Karlebynejdens institut erbjuder undervisning i finska och svenska från grundnivå.
Mellersta Österbottens utbildningskoncern erbjuder kurser i finska vid Mellersta Österbottens folkhögskola i Kelviå inom utbildningen i läs- och skrivfärdigheter och den förberedande utbildningen för vuxna invandrare. Det går också att studera finska inom utbildningen som handleder för yrkesutbildning (VALMA) vid Mellersta Österbottens Vuxeninstitut.
Vuxenutbildningen anordnar även förberedande utbildning för vuxna invandrare vid Mellersta Österbottens folkhögskola i Kelviå.
Vid Kronoby folkhögskola kan du studera finska och svenska på grund- och påbyggnadsnivå.
Om du är berättigad till integrationsstöd ska du kontakta TE-byrån innan du ansöker.
Du kan be om information om undervisning i finska och svenska för invandrare hos utlänningsbyrån.
Läs mer: Finska och svenska språket
Karlebynejdens institutfinska _ svenska
linkkiMellersta Österbottens utbildningskoncern:
Utbildning för invandrarefinska _ engelska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Utlänningsbyrånfinska _ svenska
linkkiKronoby folkhögskola:
Kronoby folkhögskolafinska _ svenska _ engelska
Möjligheter att studera finska eller svenska
Karlebynejdens institut erbjuder undervisning i finska och svenska från grundnivå.
Mellersta Österbottens utbildningskoncern erbjuder kurser i finska vid Mellersta Österbottens folkhögskola i Kelviå inom utbildningen i läs- och skrivfärdigheter och den förberedande utbildningen för vuxna invandrare. Det går också att studera finska inom utbildningen som handleder för yrkesutbildning (VALMA) vid Mellersta Österbottens Vuxeninstitut.
Vuxenutbildningen anordnar även förberedande utbildning för vuxna invandrare vid Mellersta Österbottens folkhögskola i Kelviå.
Vid Kronoby folkhögskola kan du studera finska och svenska på grund- och påbyggnadsnivå.
Om du är berättigad till integrationsstöd ska du kontakta TE-byrån innan du ansöker.
Du kan be om information om undervisning i finska och svenska för invandrare hos utlänningsbyrån.
Läs mer: Finska och svenska språket
Karlebynejdens institutfinska _ svenska
linkkiMellersta Österbottens utbildningskoncern:
Utbildning för invandrarefinska _ engelska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Utlänningsbyrånfinska _ svenska
linkkiKronoby folkhögskola:
Kronoby folkhögskolafinska _ svenska _ engelska
Möjligheter att studera finska eller svenska
Karlebynejdens institut erbjuder undervisning i finska och svenska från grundnivå.
Mellersta Österbottens utbildningskoncern erbjuder kurser i finska vid Mellersta Österbottens folkhögskola i Kelviå inom utbildningen i läs- och skrivfärdigheter och den förberedande utbildningen för vuxna invandrare. Det går också att studera finska inom utbildningen som handleder för yrkesutbildning (VALMA) vid Mellersta Österbottens Vuxeninstitut.
Vuxenutbildningen anordnar även förberedande utbildning för vuxna invandrare vid Mellersta Österbottens folkhögskola i Kelviå.
Vid Kronoby folkhögskola kan du studera finska och svenska på grund- och påbyggnadsnivå.
Om du är berättigad till integrationsstöd ska du kontakta TE-byrån innan du ansöker.
Du kan be om information om undervisning i finska och svenska för invandrare hos utlänningsbyrån.
Läs mer: Finska och svenska språket
Karlebynejdens institutfinska _ svenska
linkkiMellersta Österbottens utbildningskoncern:
Utbildning för invandrarefinska _ engelska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Utlänningsbyrånfinska _ svenska
linkkiKronoby folkhögskola:
Kronoby folkhögskolafinska _ svenska _ engelska
Var hittar jag jobb?
Att grunda ett företag
Beskattning
Om du blir arbetslös
Var hittar jag jobb?
Du kan söka arbetsplatser på internet och i tidningar.
På internet hittar du jobbsajter när du skriver ”avoimet työpaikat” (lediga jobb) i sökmotorns textfält.
På många jobbsajter kan du spara din jobbansökan och meritförteckning (CV) så att arbetsgivaren kan läsa dem.
Vid Österbottens TE-byrå (arbets- och näringsbyrå) får du hjälp med att hitta en arbetsplats.
Du behöver inte alltid boka tid för att besöka TE-byrån.
I Mina e-tjänster på nätet kan du bl.a. ändra dina uppgifter som arbetssökande och kontrollera giltighetstiden för jobbsökningen och utlåtandet om arbetslöshetsförsäkring.
Om du behöver boka en tid till TE-byrån ska du kontakta TE-byrån direkt per telefon eller boka en tid på plats.
Var även direkt i kontakt med TE-byrån om du önskar ändra en tidsbokning.
Du kan ringa TE-telefonservice då du behöver information om TE-byråns tjänster eller vägledning i tjänsterna på nätet.
Telefonnumret till TE-telefonservice är 0295 025 500 på finska, 0295 025 510 på svenska, 0295 020 713 på engelska och 0295 020 715 på ryska.
TE-byrån i Österbotten betjänar i Karleby, Kaustby, Jakobstad, Närpes, Kristinestad och Vasa.
Du kan fritt välja vilken TE-byrå du besöker.
Adressen för TE-byrån i Karleby är
67100 Karleby.
På TE-byråns jobbsajt finns tusentals arbetsplatser runt om i Finland.
Du hittar lediga arbetsplatser i din kommun genom att skriva kommunens namn i sökfältet ”Region”.
Läs mer:
Var hittar jag jobb?
linkkiArbets- och näringsbyråns tjänster:
Offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiArbets- och näringsbyråns tjänster:
Österbottens TE-byråfinska _ svenska
linkkiArbets- och näringsbyråns tjänster:
TE-telefonservicefinska _ svenska _ engelska _ ryska
linkkiArbets- och näringsbyråns tjänster:
Arbets- och näringsbyråns arbetsplatssajtfinska _ svenska
Att grunda ett företag
KOSEK (Karlebynejdens Utveckling Ab) erbjuder tjänster som nyttar företaget under hela dess livscykel, från och med att starta företagsverksamhet.
KOSEKs experter hjälper bland annat med att utarbeta en affärsverksamhetsplan och att ansöka startpeng.
Tjänsterna är avgiftsfria.
Verksamheten av Mellersta Österbottens Nyföretagarcentral FIRMAXI fortsätter som en del av KOSEKs tjänster.
Du kan besöka Karlebynejdens Utveckling Ab om du behöver information om att grunda ett företag.
Detta kan exempelvis inkludera
företagsfinansiering
rekrytering av anställda
samarbetsnätverk
verksamhetslokaler
Läs mer:
Att grunda ett företag.
linkkiNyföretagarcentralen Firmaxi:
Nyföretagarcentralen Firmaxifinska
Karlebynejdens Utveckling Abfinska _ svenska _ engelska
Beskattning
Om du behöver ett skattekort eller skattenummer kan du besöka Västra Finlands skattebyrå.
Skattebyråns kontaktuppgifter:
PB 1002, 67101 Karleby
Besöksadress: Karlebygatan 27, Karleby
Skatteförvaltningens riksomfattande telefontjänst: 029 497 050
Läs mer: Beskattning.
Om du blir arbetslös
Medborgare i EU- och EES-länderna kan anmäla sig som arbetslösa på nätet i TE-byråns ”Mina e-tjänster”.
Du kan besöka TE-byrån om du inte kan anmäla dig som arbetssökande på nätet eller om du är medborgare i något annat land.
Du kan ringa till riksomfattande servicenummer om du behöver hjälp med att använda e-tjänsterna eller mer information om TE-byråns tjänster.
Det riksomfattande servicenumret är 0295 025 500 på finska, 0295 025 510 på svenska, 0295 020 713 på engelska och 0295 020 715 på ryska.
TE-byrån i Österbotten betjänar i Karleby, Kaustby, Jakobstad, Närpes, Kristinestad och Vasa.
Du kan fritt välja vilken TE-byrå du besöker.
TE-byråns adress i Karleby
Läs mer: Arbetslöshetsförsäkring.
linkkiArbets- och näringsbyråns tjänster:
Offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiArbets- och näringsbyråns tjänster:
Österbottens TE-byråfinska _ svenska
linkkiArbets- och näringsbyråns tjänster:
TE-telefonservicefinska _ svenska _ engelska _ ryska
Fennovoima bygger kärnkraftverksenheten Hanhikivi 1 i Pyhäjoki.
Kärnkraftverket levereras av RAOS Project Oy, ett bolag som ingår i den ryska Rosatom-koncernen.
Enligt den överenskomna tidtabellen kommer kärnkraftverket att producera el år 2024.
Planeringen och konstruktionen av kärnkraftverket är ett omfattande projekt som tar cirka 10 år att slutföra.
Under tiden kärnkraftverket uppförs kommer som mest upp till 3 000–4 000 personer att arbeta på området.
Arbetsgivaren arrangerar logi för merparten av arbetstagarna, och man strävar efter att ordna inkvartering så nära bygget som möjligt.
I kärnkraftverkets omedelbara närhet byggs ett inkvarteringsområde för 1 000 personer.
I Pyhäjoki och det omgivande området har man förberett sig på kärnkraftverksprojektet redan i flera års tid.
Information om området har sammanställts bl.a. i Hanhikivi-guiden som publicerats på finska, engelska, svenska och ryska.
Elektroniska versioner av guiden finns på storprojektets webbplats.
Den tryckta guiden finns i företagsservicecentralerna i kommunerna på området.
Som en del av förberedelserna för kärnkraftverksprojektet finns information samlad om tjänsterna på området på dessa lokala InfoFinland-sidor.
Mer information om Fennovoimas kärnkraftverksprojekt i Pyhäjoki:
Fennovoima Oyfinska _ engelska
linkkiBrahestadsregionens företagstjänster:
Information om storprojekt som förverkligas i regionen och förberedelserna för dessafinska _ engelska _ ryska
Karlebynejdens Utveckling Abfinska _ svenska _ engelska
linkkiPyhäjoki kommun:
Pyhäjoki kommunfinska _ svenska _ engelska
Information om verksamhetsmiljön för kärnkraftverksprojektetfinska _ svenska _ engelska _ ryska
Var hittar jag jobb?
Att grunda ett företag
Beskattning
Om du blir arbetslös
Var hittar jag jobb?
Du kan söka arbetsplatser på internet och i tidningar.
På internet hittar du jobbsajter när du skriver ”avoimet työpaikat” (lediga jobb) i sökmotorns textfält.
På många jobbsajter kan du spara din jobbansökan och meritförteckning (CV) så att arbetsgivaren kan läsa dem.
Vid Österbottens TE-byrå (arbets- och näringsbyrå) får du hjälp med att hitta en arbetsplats.
Du behöver inte alltid boka tid för att besöka TE-byrån.
I Mina e-tjänster på nätet kan du bl.a. ändra dina uppgifter som arbetssökande och kontrollera giltighetstiden för jobbsökningen och utlåtandet om arbetslöshetsförsäkring.
Om du behöver boka en tid till TE-byrån ska du kontakta TE-byrån direkt per telefon eller boka en tid på plats.
Var även direkt i kontakt med TE-byrån om du önskar ändra en tidsbokning.
Du kan ringa TE-telefonservice då du behöver information om TE-byråns tjänster eller vägledning i tjänsterna på nätet.
Telefonnumret till TE-telefonservice är 0295 025 500 på finska, 0295 025 510 på svenska, 0295 020 713 på engelska och 0295 020 715 på ryska.
TE-byrån i Österbotten betjänar i Karleby, Kaustby, Jakobstad, Närpes, Kristinestad och Vasa.
Du kan fritt välja vilken TE-byrå du besöker.
Adressen för TE-byrån i Karleby är
67100 Karleby.
På TE-byråns jobbsajt finns tusentals arbetsplatser runt om i Finland.
Du hittar lediga arbetsplatser i din kommun genom att skriva kommunens namn i sökfältet ”Region”.
Läs mer:
Var hittar jag jobb?
linkkiArbets- och näringsbyråns tjänster:
Offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiArbets- och näringsbyråns tjänster:
Österbottens TE-byråfinska _ svenska
linkkiArbets- och näringsbyråns tjänster:
TE-telefonservicefinska _ svenska _ engelska _ ryska
linkkiArbets- och näringsbyråns tjänster:
Arbets- och näringsbyråns arbetsplatssajtfinska _ svenska
Att grunda ett företag
KOSEK (Karlebynejdens Utveckling Ab) erbjuder tjänster som nyttar företaget under hela dess livscykel, från och med att starta företagsverksamhet.
KOSEKs experter hjälper bland annat med att utarbeta en affärsverksamhetsplan och att ansöka startpeng.
Tjänsterna är avgiftsfria.
Verksamheten av Mellersta Österbottens Nyföretagarcentral FIRMAXI fortsätter som en del av KOSEKs tjänster.
Du kan besöka Karlebynejdens Utveckling Ab om du behöver information om att grunda ett företag.
Detta kan exempelvis inkludera
företagsfinansiering
rekrytering av anställda
samarbetsnätverk
verksamhetslokaler
Läs mer:
Att grunda ett företag.
linkkiNyföretagarcentralen Firmaxi:
Nyföretagarcentralen Firmaxifinska
Karlebynejdens Utveckling Abfinska _ svenska _ engelska
Beskattning
Om du behöver ett skattekort eller skattenummer kan du besöka Västra Finlands skattebyrå.
Skattebyråns kontaktuppgifter:
PB 1002, 67101 Karleby
Besöksadress: Karlebygatan 27, Karleby
Skatteförvaltningens riksomfattande telefontjänst: 029 497 050
Läs mer: Beskattning.
Om du blir arbetslös
Medborgare i EU- och EES-länderna kan anmäla sig som arbetslösa på nätet i TE-byråns ”Mina e-tjänster”.
Du kan besöka TE-byrån om du inte kan anmäla dig som arbetssökande på nätet eller om du är medborgare i något annat land.
Du kan ringa till riksomfattande servicenummer om du behöver hjälp med att använda e-tjänsterna eller mer information om TE-byråns tjänster.
Det riksomfattande servicenumret är 0295 025 500 på finska, 0295 025 510 på svenska, 0295 020 713 på engelska och 0295 020 715 på ryska.
TE-byrån i Österbotten betjänar i Karleby, Kaustby, Jakobstad, Närpes, Kristinestad och Vasa.
Du kan fritt välja vilken TE-byrå du besöker.
TE-byråns adress i Karleby
Läs mer: Arbetslöshetsförsäkring.
linkkiArbets- och näringsbyråns tjänster:
Offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiArbets- och näringsbyråns tjänster:
Österbottens TE-byråfinska _ svenska
linkkiArbets- och näringsbyråns tjänster:
TE-telefonservicefinska _ svenska _ engelska _ ryska
Fennovoima bygger kärnkraftverksenheten Hanhikivi 1 i Pyhäjoki.
Kärnkraftverket levereras av RAOS Project Oy, ett bolag som ingår i den ryska Rosatom-koncernen.
Enligt den överenskomna tidtabellen kommer kärnkraftverket att producera el år 2024.
Planeringen och konstruktionen av kärnkraftverket är ett omfattande projekt som tar cirka 10 år att slutföra.
Under tiden kärnkraftverket uppförs kommer som mest upp till 3 000–4 000 personer att arbeta på området.
Arbetsgivaren arrangerar logi för merparten av arbetstagarna, och man strävar efter att ordna inkvartering så nära bygget som möjligt.
I kärnkraftverkets omedelbara närhet byggs ett inkvarteringsområde för 1 000 personer.
I Pyhäjoki och det omgivande området har man förberett sig på kärnkraftverksprojektet redan i flera års tid.
Information om området har sammanställts bl.a. i Hanhikivi-guiden som publicerats på finska, engelska, svenska och ryska.
Elektroniska versioner av guiden finns på storprojektets webbplats.
Den tryckta guiden finns i företagsservicecentralerna i kommunerna på området.
Som en del av förberedelserna för kärnkraftverksprojektet finns information samlad om tjänsterna på området på dessa lokala InfoFinland-sidor.
Mer information om Fennovoimas kärnkraftverksprojekt i Pyhäjoki:
Fennovoima Oyfinska _ engelska
linkkiBrahestadsregionens företagstjänster:
Information om storprojekt som förverkligas i regionen och förberedelserna för dessafinska _ engelska _ ryska
Karlebynejdens Utveckling Abfinska _ svenska _ engelska
linkkiPyhäjoki kommun:
Pyhäjoki kommunfinska _ svenska _ engelska
Information om verksamhetsmiljön för kärnkraftverksprojektetfinska _ svenska _ engelska _ ryska
Var hittar jag jobb?
Att grunda ett företag
Beskattning
Om du blir arbetslös
Var hittar jag jobb?
Du kan söka arbetsplatser på internet och i tidningar.
På internet hittar du jobbsajter när du skriver ”avoimet työpaikat” (lediga jobb) i sökmotorns textfält.
På många jobbsajter kan du spara din jobbansökan och meritförteckning (CV) så att arbetsgivaren kan läsa dem.
Vid Österbottens TE-byrå (arbets- och näringsbyrå) får du hjälp med att hitta en arbetsplats.
Du behöver inte alltid boka tid för att besöka TE-byrån.
I Mina e-tjänster på nätet kan du bl.a. ändra dina uppgifter som arbetssökande och kontrollera giltighetstiden för jobbsökningen och utlåtandet om arbetslöshetsförsäkring.
Om du behöver boka en tid till TE-byrån ska du kontakta TE-byrån direkt per telefon eller boka en tid på plats.
Var även direkt i kontakt med TE-byrån om du önskar ändra en tidsbokning.
Du kan ringa TE-telefonservice då du behöver information om TE-byråns tjänster eller vägledning i tjänsterna på nätet.
Telefonnumret till TE-telefonservice är 0295 025 500 på finska, 0295 025 510 på svenska, 0295 020 713 på engelska och 0295 020 715 på ryska.
TE-byrån i Österbotten betjänar i Karleby, Kaustby, Jakobstad, Närpes, Kristinestad och Vasa.
Du kan fritt välja vilken TE-byrå du besöker.
Adressen för TE-byrån i Karleby är
67100 Karleby.
På TE-byråns jobbsajt finns tusentals arbetsplatser runt om i Finland.
Du hittar lediga arbetsplatser i din kommun genom att skriva kommunens namn i sökfältet ”Region”.
Läs mer:
Var hittar jag jobb?
linkkiArbets- och näringsbyråns tjänster:
Offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiArbets- och näringsbyråns tjänster:
Österbottens TE-byråfinska _ svenska
linkkiArbets- och näringsbyråns tjänster:
TE-telefonservicefinska _ svenska _ engelska _ ryska
linkkiArbets- och näringsbyråns tjänster:
Arbets- och näringsbyråns arbetsplatssajtfinska _ svenska
Att grunda ett företag
KOSEK (Karlebynejdens Utveckling Ab) erbjuder tjänster som nyttar företaget under hela dess livscykel, från och med att starta företagsverksamhet.
KOSEKs experter hjälper bland annat med att utarbeta en affärsverksamhetsplan och att ansöka startpeng.
Tjänsterna är avgiftsfria.
Verksamheten av Mellersta Österbottens Nyföretagarcentral FIRMAXI fortsätter som en del av KOSEKs tjänster.
Du kan besöka Karlebynejdens Utveckling Ab om du behöver information om att grunda ett företag.
Detta kan exempelvis inkludera
företagsfinansiering
rekrytering av anställda
samarbetsnätverk
verksamhetslokaler
Läs mer:
Att grunda ett företag.
linkkiNyföretagarcentralen Firmaxi:
Nyföretagarcentralen Firmaxifinska
Karlebynejdens Utveckling Abfinska _ svenska _ engelska
Beskattning
Om du behöver ett skattekort eller skattenummer kan du besöka Västra Finlands skattebyrå.
Skattebyråns kontaktuppgifter:
PB 1002, 67101 Karleby
Besöksadress: Karlebygatan 27, Karleby
Skatteförvaltningens riksomfattande telefontjänst: 029 497 050
Läs mer: Beskattning.
Om du blir arbetslös
Medborgare i EU- och EES-länderna kan anmäla sig som arbetslösa på nätet i TE-byråns ”Mina e-tjänster”.
Du kan besöka TE-byrån om du inte kan anmäla dig som arbetssökande på nätet eller om du är medborgare i något annat land.
Du kan ringa till riksomfattande servicenummer om du behöver hjälp med att använda e-tjänsterna eller mer information om TE-byråns tjänster.
Det riksomfattande servicenumret är 0295 025 500 på finska, 0295 025 510 på svenska, 0295 020 713 på engelska och 0295 020 715 på ryska.
TE-byrån i Österbotten betjänar i Karleby, Kaustby, Jakobstad, Närpes, Kristinestad och Vasa.
Du kan fritt välja vilken TE-byrå du besöker.
TE-byråns adress i Karleby
Läs mer: Arbetslöshetsförsäkring.
linkkiArbets- och näringsbyråns tjänster:
Offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiArbets- och näringsbyråns tjänster:
Österbottens TE-byråfinska _ svenska
linkkiArbets- och näringsbyråns tjänster:
TE-telefonservicefinska _ svenska _ engelska _ ryska
Fennovoima bygger kärnkraftverksenheten Hanhikivi 1 i Pyhäjoki.
Kärnkraftverket levereras av RAOS Project Oy, ett bolag som ingår i den ryska Rosatom-koncernen.
Enligt den överenskomna tidtabellen kommer kärnkraftverket att producera el år 2024.
Planeringen och konstruktionen av kärnkraftverket är ett omfattande projekt som tar cirka 10 år att slutföra.
Under tiden kärnkraftverket uppförs kommer som mest upp till 3 000–4 000 personer att arbeta på området.
Arbetsgivaren arrangerar logi för merparten av arbetstagarna, och man strävar efter att ordna inkvartering så nära bygget som möjligt.
I kärnkraftverkets omedelbara närhet byggs ett inkvarteringsområde för 1 000 personer.
I Pyhäjoki och det omgivande området har man förberett sig på kärnkraftverksprojektet redan i flera års tid.
Information om området har sammanställts bl.a. i Hanhikivi-guiden som publicerats på finska, engelska, svenska och ryska.
Elektroniska versioner av guiden finns på storprojektets webbplats.
Den tryckta guiden finns i företagsservicecentralerna i kommunerna på området.
Som en del av förberedelserna för kärnkraftverksprojektet finns information samlad om tjänsterna på området på dessa lokala InfoFinland-sidor.
Mer information om Fennovoimas kärnkraftverksprojekt i Pyhäjoki:
Fennovoima Oyfinska _ engelska
linkkiBrahestadsregionens företagstjänster:
Information om storprojekt som förverkligas i regionen och förberedelserna för dessafinska _ engelska _ ryska
Karlebynejdens Utveckling Abfinska _ svenska _ engelska
linkkiPyhäjoki kommun:
Pyhäjoki kommunfinska _ svenska _ engelska
Information om verksamhetsmiljön för kärnkraftverksprojektetfinska _ svenska _ engelska _ ryska
Rådgivning och integration för invandrare
Inledande kartläggning och integrationsplan
Behöver du en tolk?
Rådgivning och integration för invandrare
Då du flyttar till Finland kan du använda dig av TE-byråns (arbets- och näringsbyrån) tjänster som hjälper dig att göra dig hemmastadd i Finland och hitta en arbetsplats.
Tjänster särskilt avsedda för invandrare är:
handledning och rådgivning för invandrare
inledande kartläggning
integrationsutbildning
Österbottens TE-byrå
67100 Karleby
Telefonväxel: 0295 025 500
Karleby evangelisk-lutherska församlingssammanslutnings invandrararbete stöder invandrares integrering i det finländska samhället.
linkkiArbets- och näringsbyråns tjänster:
Offentliga arbets- och näringstjänsterfinska _ svenska
linkkiArbets- och näringsministeriet:
Guiden Välkommen till Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
linkkiKarleby evangelisk-lutherska församlingssammansutning:
Karleby evangelisk-lutherska församlings invandrararbetefinska _ svenska _ engelska _ ryska
Inledande kartläggning och integrationsplan
En inledande kartläggning och integrationsplan utarbetas för dig i arbets- och näringsbyrån. Om du kommit till
Finland som flykting utarbetas en inledande kartläggning och integrationsplan för dig vid utlänningsbyrån.
Du kan fråga mer om kartläggningen och integrationsplanen vid utlänningsbyrån eller TE-byrån.
Utlänningsbyrån
Vasavägen 6 C
67100 Karleby
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Utlänningsbyrånfinska _ svenska
Behöver du en tolk?
Om du måste sköta ärenden med finländska myndigheter, men inte kan finska eller svenska och det inte heller finns något annat språk som både du och myndigheten talar, kan du i vissa fall ha rätt till tolkning.
Myndigheten beställer tolken om du på förhand uppgett att du behöver en tolk.
I detta fall är det gratis för dig att använda dig av tolk.
Du kan använda tolken när du själv önskar om du betalar kostnaderna och beställer tolken själv.
Läs mer:
Behöver du en tolk?
Rådgivning och integration för invandrare
Inledande kartläggning och integrationsplan
Behöver du en tolk?
Rådgivning och integration för invandrare
Då du flyttar till Finland kan du använda dig av TE-byråns (arbets- och näringsbyrån) tjänster som hjälper dig att göra dig hemmastadd i Finland och hitta en arbetsplats.
Tjänster särskilt avsedda för invandrare är:
handledning och rådgivning för invandrare
inledande kartläggning
integrationsutbildning
Österbottens TE-byrå
67100 Karleby
Telefonväxel: 0295 025 500
Karleby evangelisk-lutherska församlingssammanslutnings invandrararbete stöder invandrares integrering i det finländska samhället.
linkkiArbets- och näringsbyråns tjänster:
Offentliga arbets- och näringstjänsterfinska _ svenska
linkkiArbets- och näringsministeriet:
Guiden Välkommen till Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
linkkiKarleby evangelisk-lutherska församlingssammansutning:
Karleby evangelisk-lutherska församlings invandrararbetefinska _ svenska _ engelska _ ryska
Inledande kartläggning och integrationsplan
En inledande kartläggning och integrationsplan utarbetas för dig i arbets- och näringsbyrån. Om du kommit till
Finland som flykting utarbetas en inledande kartläggning och integrationsplan för dig vid utlänningsbyrån.
Du kan fråga mer om kartläggningen och integrationsplanen vid utlänningsbyrån eller TE-byrån.
Utlänningsbyrån
Vasavägen 6 C
67100 Karleby
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Utlänningsbyrånfinska _ svenska
Behöver du en tolk?
Om du måste sköta ärenden med finländska myndigheter, men inte kan finska eller svenska och det inte heller finns något annat språk som både du och myndigheten talar, kan du i vissa fall ha rätt till tolkning.
Myndigheten beställer tolken om du på förhand uppgett att du behöver en tolk.
I detta fall är det gratis för dig att använda dig av tolk.
Du kan använda tolken när du själv önskar om du betalar kostnaderna och beställer tolken själv.
Läs mer:
Behöver du en tolk?
Rådgivning och integration för invandrare
Inledande kartläggning och integrationsplan
Behöver du en tolk?
Rådgivning och integration för invandrare
Då du flyttar till Finland kan du använda dig av TE-byråns (arbets- och näringsbyrån) tjänster som hjälper dig att göra dig hemmastadd i Finland och hitta en arbetsplats.
Tjänster särskilt avsedda för invandrare är:
handledning och rådgivning för invandrare
inledande kartläggning
integrationsutbildning
Österbottens TE-byrå
67100 Karleby
Telefonväxel: 0295 025 500
Karleby evangelisk-lutherska församlingssammanslutnings invandrararbete stöder invandrares integrering i det finländska samhället.
linkkiArbets- och näringsbyråns tjänster:
Offentliga arbets- och näringstjänsterfinska _ svenska
linkkiArbets- och näringsministeriet:
Guiden Välkommen till Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
linkkiKarleby evangelisk-lutherska församlingssammansutning:
Karleby evangelisk-lutherska församlings invandrararbetefinska _ svenska _ engelska _ ryska
Inledande kartläggning och integrationsplan
En inledande kartläggning och integrationsplan utarbetas för dig i arbets- och näringsbyrån. Om du kommit till
Finland som flykting utarbetas en inledande kartläggning och integrationsplan för dig vid utlänningsbyrån.
Du kan fråga mer om kartläggningen och integrationsplanen vid utlänningsbyrån eller TE-byrån.
Utlänningsbyrån
Vasavägen 6 C
67100 Karleby
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Utlänningsbyrånfinska _ svenska
Behöver du en tolk?
Om du måste sköta ärenden med finländska myndigheter, men inte kan finska eller svenska och det inte heller finns något annat språk som både du och myndigheten talar, kan du i vissa fall ha rätt till tolkning.
Myndigheten beställer tolken om du på förhand uppgett att du behöver en tolk.
I detta fall är det gratis för dig att använda dig av tolk.
Du kan använda tolken när du själv önskar om du betalar kostnaderna och beställer tolken själv.
Läs mer:
Behöver du en tolk?
Registrering som invånare
Om du vill flytta till Finland behöver du vanligtvis ett uppehållstillstånd.
Uppehållstillståndsärenden hanteras av Finlands beskickningar i utlandet och Migrationsverket.
Läs mer: Flytta till Finland.
Då du flyttar till Karleby (Kokkola) ska du registrera dig som invånare i kommunen.
Du kan personligen registrera dig på Karleby enheten för Magistraten i Västra Finland:
Magistraten i Västra Finland
Karleby enhet
Karlebygatan 27
67701 Karleby
Telefon: 029 553 9451
När du går till magistraten ska du ta med dig
uppehållstillstånd och uppehållskort (om du behöver ett uppehållstillstånd i Finland)
registreringsintyget över uppehållsrätt för EU-medborgare (om du är EU-medborgare)
äktenskapsbevis
födelseattester för dina barn
Observera att officiella handlingar som tagits med från utlandet ska vara legaliserade och i original samt översatta till finska, svenska eller engelska.
Mer information om legalisering av handlingar får du hos magistraten eller hos ditt lands beskickning i Finland.
Läs mer:
Registrering som invånare.
Magistratens kontaktuppgifterfinska _ svenska _ engelska
Fortsatt uppehållstillstånd
Du ska ansöka om fortsatt uppehållstillstånd innan ditt tidigare uppehållstillstånd går ut.
Du ansöker om tillståndet vid Migrationsverkets servicesställen.
Du kan endast ansöka om fortsatt uppehållstillstånd i Finland.
Migrationsverket
Korsholmsesplanaden 45
Vasa
Läs mer: Fortsatt uppehållstillstånd.
Registrering som invånare
Om du vill flytta till Finland behöver du vanligtvis ett uppehållstillstånd.
Uppehållstillståndsärenden hanteras av Finlands beskickningar i utlandet och Migrationsverket.
Läs mer: Flytta till Finland.
Då du flyttar till Karleby (Kokkola) ska du registrera dig som invånare i kommunen.
Du kan personligen registrera dig på Karleby enheten för Magistraten i Västra Finland:
Magistraten i Västra Finland
Karleby enhet
Karlebygatan 27
67701 Karleby
Telefon: 029 553 9451
När du går till magistraten ska du ta med dig
uppehållstillstånd och uppehållskort (om du behöver ett uppehållstillstånd i Finland)
registreringsintyget över uppehållsrätt för EU-medborgare (om du är EU-medborgare)
äktenskapsbevis
födelseattester för dina barn
Observera att officiella handlingar som tagits med från utlandet ska vara legaliserade och i original samt översatta till finska, svenska eller engelska.
Mer information om legalisering av handlingar får du hos magistraten eller hos ditt lands beskickning i Finland.
Läs mer:
Registrering som invånare.
Magistratens kontaktuppgifterfinska _ svenska _ engelska
Fortsatt uppehållstillstånd
Du ska ansöka om fortsatt uppehållstillstånd innan ditt tidigare uppehållstillstånd går ut.
Du ansöker om tillståndet vid Migrationsverkets servicesställen.
Du kan endast ansöka om fortsatt uppehållstillstånd i Finland.
Migrationsverket
Korsholmsesplanaden 45
Vasa
Läs mer: Fortsatt uppehållstillstånd.
Registrering som invånare
Om du vill flytta till Finland behöver du vanligtvis ett uppehållstillstånd.
Uppehållstillståndsärenden hanteras av Finlands beskickningar i utlandet och Migrationsverket.
Läs mer: Flytta till Finland.
Då du flyttar till Karleby (Kokkola) ska du registrera dig som invånare i kommunen.
Du kan personligen registrera dig på Karleby enheten för Magistraten i Västra Finland:
Magistraten i Västra Finland
Karleby enhet
Karlebygatan 27
67701 Karleby
Telefon: 029 553 9451
När du går till magistraten ska du ta med dig
uppehållstillstånd och uppehållskort (om du behöver ett uppehållstillstånd i Finland)
registreringsintyget över uppehållsrätt för EU-medborgare (om du är EU-medborgare)
äktenskapsbevis
födelseattester för dina barn
Observera att officiella handlingar som tagits med från utlandet ska vara legaliserade och i original samt översatta till finska, svenska eller engelska.
Mer information om legalisering av handlingar får du hos magistraten eller hos ditt lands beskickning i Finland.
Läs mer:
Registrering som invånare.
Magistratens kontaktuppgifterfinska _ svenska _ engelska
Fortsatt uppehållstillstånd
Du ska ansöka om fortsatt uppehållstillstånd innan ditt tidigare uppehållstillstånd går ut.
Du ansöker om tillståndet vid Migrationsverkets servicesställen.
Du kan endast ansöka om fortsatt uppehållstillstånd i Finland.
Migrationsverket
Korsholmsesplanaden 45
Vasa
Läs mer: Fortsatt uppehållstillstånd.
InfoFinland finansieras av Samarbetskommunerna och staten.
Åren 2017–2020 var statens finansiärer arbets- och näringsministeriet, undervisnings- och kulturministeriet, miljöministeriet, FPA och Skatteförvaltningen.
InfoFinland utvecklas i samarbete med finansiärerna.
Den som planerar att flytta till Finland med hjälp av Infobanken hittar lätt information om att leva, bo, arbeta och studera i Finland på många olika språk.
Staten
Arbets- och näringsministeriet
Arbets- och näringsministeriet svarar för beredningen av ärenden i anslutning till integrationen av invandrare i Finland.
Kompetenscentret för integration av invandrare stöder arbete som främjar integrationen av invandrare lokalt, regionalt och riksomfattande.
linkkiArbets- och näringsministeriet :
Integration av invandrarefinska _ svenska _ engelska
Undervisnings- och kulturministeriet
Undervisnings- och kulturministeriet svarar för utvecklingen av och det internationella samarbetet inom utbildnings-, vetenskaps-, kultur-, motions- och ungdomspolitiken.
linkkiUndervisnings- och kulturministeriet:
Webbsidorfinska _ svenska _ engelska
Miljöministeriet
linkkiMiljöministeriet:
Webbsidorfinska _ svenska _ engelska
FPA
FPA sköter grundtryggheten i olika skeden av livet för dem som bor i Finland.
FPA:s kunder är alla personer som bor i Finland och utomlands och som omfattas av socialskyddet i Finland.
FPA och Skatteförvaltningen erbjuder information till utländska anställda på servicestället In To Finland i Helsingfors.
Flyttning till eller från Finlandfinska _ svenska _ engelska
Skatteförvaltningen
linkkiSkatteförvaltningen:
Webbsidorfinska _ svenska _ engelska
Kommunerna
Helsingfors stad
Publicerar och administrerar InfoFinland.
Kommuner som är med i samarbetsavtalet
InfoFinlands samarbetsavtal
InfoFinlands finansiärer har ingått ett samarbetsavtal med vilket man överenskommit om principerna för genomförandet och finansieringen av nättjänsten InfoFinland (tidigare Infobanken) för åren 2017–2020.
Samarbetet möjliggör riksomfattande webbinformation för invandrare och personer som planerar att flytta till Finland och för myndigheter inom invandrarsektorn på ett sätt som också stöder behovet av information i kommunerna.
Det är lätt att på ett pålitligt sätt hitta väsentlig information om integration av invandrare och om att bo i Finland på ett ställe, www.infofinland.fi.
Avtalsparterna driver och utvecklar tjänsten tillsammans.
De vill dessutom stärka InfoFinlands riksomfattande ställning, så att det är möjligt för nya kommuner och andra organisationer att ansluta sig till tjänsten också i fortsättningen.
Kommunernas finansieringsandelar fastställs utgående från antalet invånare.
Genomförandet av avtalet följs upp av en styrgrupp.
Nya aktörer är välkomna att utveckla den flerspråkiga informationen till invandrare och ansluta sig till InfoFinlands samarbetsavtal.
Närmare information om hur man ansluter sig till avtalet ger InfoFinlands chefredaktör Eija Kyllönen-Saarnio, eija.kyllonen-saarnio(snabel-a)hel.fi, tfn 050 363 3285.
InfoFinland finansieras av Samarbetskommunerna och staten.
Åren 2017–2020 var statens finansiärer arbets- och näringsministeriet, undervisnings- och kulturministeriet, miljöministeriet, FPA och Skatteförvaltningen.
InfoFinland utvecklas i samarbete med finansiärerna.
Den som planerar att flytta till Finland med hjälp av Infobanken hittar lätt information om att leva, bo, arbeta och studera i Finland på många olika språk.
Staten
Arbets- och näringsministeriet
Arbets- och näringsministeriet svarar för beredningen av ärenden i anslutning till integrationen av invandrare i Finland.
Kompetenscentret för integration av invandrare stöder arbete som främjar integrationen av invandrare lokalt, regionalt och riksomfattande.
linkkiArbets- och näringsministeriet :
Integration av invandrarefinska _ svenska _ engelska
Undervisnings- och kulturministeriet
Undervisnings- och kulturministeriet svarar för utvecklingen av och det internationella samarbetet inom utbildnings-, vetenskaps-, kultur-, motions- och ungdomspolitiken.
linkkiUndervisnings- och kulturministeriet:
Webbsidorfinska _ svenska _ engelska
Miljöministeriet
linkkiMiljöministeriet:
Webbsidorfinska _ svenska _ engelska
FPA
FPA sköter grundtryggheten i olika skeden av livet för dem som bor i Finland.
FPA:s kunder är alla personer som bor i Finland och utomlands och som omfattas av socialskyddet i Finland.
FPA och Skatteförvaltningen erbjuder information till utländska anställda på servicestället In To Finland i Helsingfors.
Flyttning till eller från Finlandfinska _ svenska _ engelska
Skatteförvaltningen
linkkiSkatteförvaltningen:
Webbsidorfinska _ svenska _ engelska
Kommunerna
Helsingfors stad
Publicerar och administrerar InfoFinland.
Kommuner som är med i samarbetsavtalet
InfoFinlands samarbetsavtal
InfoFinlands finansiärer har ingått ett samarbetsavtal med vilket man överenskommit om principerna för genomförandet och finansieringen av nättjänsten InfoFinland (tidigare Infobanken) för åren 2017–2020.
Samarbetet möjliggör riksomfattande webbinformation för invandrare och personer som planerar att flytta till Finland och för myndigheter inom invandrarsektorn på ett sätt som också stöder behovet av information i kommunerna.
Det är lätt att på ett pålitligt sätt hitta väsentlig information om integration av invandrare och om att bo i Finland på ett ställe, www.infofinland.fi.
Avtalsparterna driver och utvecklar tjänsten tillsammans.
De vill dessutom stärka InfoFinlands riksomfattande ställning, så att det är möjligt för nya kommuner och andra organisationer att ansluta sig till tjänsten också i fortsättningen.
Kommunernas finansieringsandelar fastställs utgående från antalet invånare.
Genomförandet av avtalet följs upp av en styrgrupp.
Nya aktörer är välkomna att utveckla den flerspråkiga informationen till invandrare och ansluta sig till InfoFinlands samarbetsavtal.
Närmare information om hur man ansluter sig till avtalet ger InfoFinlands chefredaktör Eija Kyllönen-Saarnio, eija.kyllonen-saarnio(snabel-a)hel.fi, tfn 050 363 3285.
InfoFinland finansieras av Samarbetskommunerna och staten.
Åren 2017–2020 var statens finansiärer arbets- och näringsministeriet, undervisnings- och kulturministeriet, miljöministeriet, FPA och Skatteförvaltningen.
InfoFinland utvecklas i samarbete med finansiärerna.
Den som planerar att flytta till Finland med hjälp av Infobanken hittar lätt information om att leva, bo, arbeta och studera i Finland på många olika språk.
Staten
Arbets- och näringsministeriet
Arbets- och näringsministeriet svarar för beredningen av ärenden i anslutning till integrationen av invandrare i Finland.
Kompetenscentret för integration av invandrare stöder arbete som främjar integrationen av invandrare lokalt, regionalt och riksomfattande.
linkkiArbets- och näringsministeriet :
Integration av invandrarefinska _ svenska _ engelska
Undervisnings- och kulturministeriet
Undervisnings- och kulturministeriet svarar för utvecklingen av och det internationella samarbetet inom utbildnings-, vetenskaps-, kultur-, motions- och ungdomspolitiken.
linkkiUndervisnings- och kulturministeriet:
Webbsidorfinska _ svenska _ engelska
Miljöministeriet
linkkiMiljöministeriet:
Webbsidorfinska _ svenska _ engelska
FPA
FPA sköter grundtryggheten i olika skeden av livet för dem som bor i Finland.
FPA:s kunder är alla personer som bor i Finland och utomlands och som omfattas av socialskyddet i Finland.
FPA och Skatteförvaltningen erbjuder information till utländska anställda på servicestället In To Finland i Helsingfors.
Flyttning till eller från Finlandfinska _ svenska _ engelska
Skatteförvaltningen
linkkiSkatteförvaltningen:
Webbsidorfinska _ svenska _ engelska
Kommunerna
Helsingfors stad
Publicerar och administrerar InfoFinland.
Kommuner som är med i samarbetsavtalet
InfoFinlands samarbetsavtal
InfoFinlands finansiärer har ingått ett samarbetsavtal med vilket man överenskommit om principerna för genomförandet och finansieringen av nättjänsten InfoFinland (tidigare Infobanken) för åren 2017–2020.
Samarbetet möjliggör riksomfattande webbinformation för invandrare och personer som planerar att flytta till Finland och för myndigheter inom invandrarsektorn på ett sätt som också stöder behovet av information i kommunerna.
Det är lätt att på ett pålitligt sätt hitta väsentlig information om integration av invandrare och om att bo i Finland på ett ställe, www.infofinland.fi.
Avtalsparterna driver och utvecklar tjänsten tillsammans.
De vill dessutom stärka InfoFinlands riksomfattande ställning, så att det är möjligt för nya kommuner och andra organisationer att ansluta sig till tjänsten också i fortsättningen.
Kommunernas finansieringsandelar fastställs utgående från antalet invånare.
Genomförandet av avtalet följs upp av en styrgrupp.
Nya aktörer är välkomna att utveckla den flerspråkiga informationen till invandrare och ansluta sig till InfoFinlands samarbetsavtal.
Närmare information om hur man ansluter sig till avtalet ger InfoFinlands chefredaktör Eija Kyllönen-Saarnio, eija.kyllonen-saarnio(snabel-a)hel.fi, tfn 050 363 3285.
Alla texter som publicerats på InfoFinlands webbplats på alla språk är fritt tillgängliga i enlighet med licensen Creative Commons Erkännande 4.0.
Du har tillstånd att:
Dela – kopiera och vidaredistribuera materialet oavsett medium eller format
Bearbeta – remixa, transformera, och bygga vidare på materialet för alla ändamål, även kommersiellt.
På följande villkor:
Erkännande (BY) – Du måste nämna källan InfoFinland.fi.
Ange en länk till webbplatsen InfoFinland.fi och nämn licensen CC BY 4.0.
Ange om bearbetningar är gjorda.
Du behöver göra så i enlighet med god sed, och inte på ett sätt som ger en bild av att InfoFinland stödjer dig eller ditt användande.
Inga ytterligare begränsningar – Du får inte tillämpa lagliga begränsningar eller teknologiska metoder som juridiskt begränsar andra från att gör något som licensen tillåter.
Erkännande 4.0 Internationellfinska _ svenska _ engelska _ ryska _ franska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ japanska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ grekiska
_ tjeckiska
Öppet programmeringsgränssnitt (API)
Vi erbjuder allt textinnehåll i InfoFinland via ett öppet programmeringsgränssnitt (API).
Med hjälp av gränssnittet kan du visa InfoFinlands innehåll på andra webbplatser eller skapa olika applikationer.
Information om gränssnittetfinska _ engelska
Öppet programmeringsgränssnittfinska
Alla texter som publicerats på InfoFinlands webbplats på alla språk är fritt tillgängliga i enlighet med licensen Creative Commons Erkännande 4.0.
Du har tillstånd att:
Dela – kopiera och vidaredistribuera materialet oavsett medium eller format
Bearbeta – remixa, transformera, och bygga vidare på materialet för alla ändamål, även kommersiellt.
På följande villkor:
Erkännande (BY) – Du måste nämna källan InfoFinland.fi.
Ange en länk till webbplatsen InfoFinland.fi och nämn licensen CC BY 4.0.
Ange om bearbetningar är gjorda.
Du behöver göra så i enlighet med god sed, och inte på ett sätt som ger en bild av att InfoFinland stödjer dig eller ditt användande.
Inga ytterligare begränsningar – Du får inte tillämpa lagliga begränsningar eller teknologiska metoder som juridiskt begränsar andra från att gör något som licensen tillåter.
Erkännande 4.0 Internationellfinska _ svenska _ engelska _ ryska _ franska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ japanska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ grekiska
_ tjeckiska
Öppet programmeringsgränssnitt (API)
Vi erbjuder allt textinnehåll i InfoFinland via ett öppet programmeringsgränssnitt (API).
Med hjälp av gränssnittet kan du visa InfoFinlands innehåll på andra webbplatser eller skapa olika applikationer.
Information om gränssnittetfinska _ engelska
Öppet programmeringsgränssnittfinska
Användning av InfoFinland-texterna på andra ställen
Texterna ur webbtjänsten InfoFinland.fi används i följande tjänster:
linkkiArbets- och näringsministeriet:
Guiden Välkommen till Finland(pdf, 3,40 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
Alla texter som publicerats på InfoFinlands webbplats på alla språk är fritt tillgängliga i enlighet med licensen Creative Commons Erkännande 4.0.
Du har tillstånd att:
Dela – kopiera och vidaredistribuera materialet oavsett medium eller format
Bearbeta – remixa, transformera, och bygga vidare på materialet för alla ändamål, även kommersiellt.
På följande villkor:
Erkännande (BY) – Du måste nämna källan InfoFinland.fi.
Ange en länk till webbplatsen InfoFinland.fi och nämn licensen CC BY 4.0.
Ange om bearbetningar är gjorda.
Du behöver göra så i enlighet med god sed, och inte på ett sätt som ger en bild av att InfoFinland stödjer dig eller ditt användande.
Inga ytterligare begränsningar – Du får inte tillämpa lagliga begränsningar eller teknologiska metoder som juridiskt begränsar andra från att gör något som licensen tillåter.
Erkännande 4.0 Internationellfinska _ svenska _ engelska _ ryska _ franska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ japanska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ grekiska
_ tjeckiska
Öppet programmeringsgränssnitt (API)
Vi erbjuder allt textinnehåll i InfoFinland via ett öppet programmeringsgränssnitt (API).
Med hjälp av gränssnittet kan du visa InfoFinlands innehåll på andra webbplatser eller skapa olika applikationer.
Information om gränssnittetfinska _ engelska
Öppet programmeringsgränssnittfinska
Användning av InfoFinland-texterna på andra ställen
Texterna ur webbtjänsten InfoFinland.fi används i följande tjänster:
linkkiArbets- och näringsministeriet:
Guiden Välkommen till Finland(pdf, 3,40 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
Medlemskommunerna har själv hand om översättningen av de övriga kommunsidorna.
Översättningsanvisning:
Översättningsanvisningen är på finska.
Översättningsanvisning:
Översättningsanvisningen är på finska.
Översättningsanvisning:
Översättningsanvisningen är på finska.
Trafik
Beslutsfattande och påverkan
Religion
Grundläggande information
Historia
Trafik
Huvudstadsregionen har goda kollektivtrafikförbindelser.
I Grankulla finns en järnvägsstation och i staden finns många busslinjer.
Du kan söka information om rutterna i tjänsten Reseplaneraren.
Tjänsten ger dig förslag på olika kollektivtrafikförbindelser från ett ställe till ett annat.
Reseplanerarefinska _ svenska _ engelska _ ryska
Inom kollektivtrafiken kan du betala med kontanter eller resekort.
I närtågen måste du köpa biljetten i förväg.
Du kan köpa resekortet på Grankulla stadshus.
Du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat.
Stadshuset
Grankullavägen 10
Mån–fre kl. 8.00–15.00; tis, ons, tors även kl. 17.00–19.30
Den närmaste flygstationen är Helsingfors–Vanda flygplats.
Flygplatsenfinska _ svenska _ engelska _ ryska _ kinesiska
Läs mer:
Trafiken i Finland.
Beslutsfattande och påverkan
I Grankulla beslutas ärenden av stadsfullmäktige.
I stadsfullmäktige sitter 35 ledamöter som representerar olika politiska grupper.
Fullmäktige väljs var fjärde år genom kommunalval.
På Grankulla stads webbplats kan du skicka respons till förvaltningen.
Du kan också lämna initiativ och ställa frågor samt kommentera ärenden på finska och på svenska.
Även engelskspråkiga frågor besvaras.
Delta och påverkafinska _ svenska
Religion
Många religiösa samfund är verksamma i Esbo och Helsingfors.
I tjänsten Uskonnot Suomessa kan du söka information enligt det religiösa samfundet och orten.
Religiösa samfundfinska _ engelska
linkkiHelsingfors ortodoxa församling:
Ortodoxa församlingenfinska _ ryska
I Grankulla finns en evangelisk-luthersk kyrka med två församlingar, en finskspråkig och en svenskspråkig.
Församlingarfinska _ svenska
Läs mer: Kulturer och religioner i Finland.
Grundläggande information
Grankulla är en av de fyra kommunerna i huvudstadsregionen.
Den ligger mitt i Esbo, 15 kilometer västerut från Helsingfors.
Grankulla har cirka 9 600 invånare, varav 60 procent har finska, 36 procent svenska och 4 procent ett annat språk som modersmål.
Grankullas areal är 6,0 km2.
Information om stadenfinska _ svenska _ engelska
Historia
År 1906 grundades ett aktiebolag i Grankulla som sålde villatomter till invånarna i huvudstadsregionen.
Området hade en direkt förbindelse till Helsingfors.
År 1920 blev villasamhället en köping.
Till en början var största delen av invånarna svenskspråkiga.
År 1972 fick köpingen stadsrättigheter.
Nätmuseetfinska _ svenska
Trafik
Beslutsfattande och påverkan
Religion
Grundläggande information
Historia
Trafik
Huvudstadsregionen har goda kollektivtrafikförbindelser.
I Grankulla finns en järnvägsstation och i staden finns många busslinjer.
Du kan söka information om rutterna i tjänsten Reseplaneraren.
Tjänsten ger dig förslag på olika kollektivtrafikförbindelser från ett ställe till ett annat.
Reseplanerarefinska _ svenska _ engelska _ ryska
Inom kollektivtrafiken kan du betala med kontanter eller resekort.
I närtågen måste du köpa biljetten i förväg.
Du kan köpa resekortet på Grankulla stadshus.
Du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat.
Stadshuset
Grankullavägen 10
Mån–fre kl. 8.00–15.00; tis, ons, tors även kl. 17.00–19.30
Den närmaste flygstationen är Helsingfors–Vanda flygplats.
Flygplatsenfinska _ svenska _ engelska _ ryska _ kinesiska
Läs mer:
Trafiken i Finland.
Beslutsfattande och påverkan
I Grankulla beslutas ärenden av stadsfullmäktige.
I stadsfullmäktige sitter 35 ledamöter som representerar olika politiska grupper.
Fullmäktige väljs var fjärde år genom kommunalval.
På Grankulla stads webbplats kan du skicka respons till förvaltningen.
Du kan också lämna initiativ och ställa frågor samt kommentera ärenden på finska och på svenska.
Även engelskspråkiga frågor besvaras.
Delta och påverkafinska _ svenska
Religion
Många religiösa samfund är verksamma i Esbo och Helsingfors.
I tjänsten Uskonnot Suomessa kan du söka information enligt det religiösa samfundet och orten.
Religiösa samfundfinska _ engelska
linkkiHelsingfors ortodoxa församling:
Ortodoxa församlingenfinska _ ryska
I Grankulla finns en evangelisk-luthersk kyrka med två församlingar, en finskspråkig och en svenskspråkig.
Församlingarfinska _ svenska
Läs mer: Kulturer och religioner i Finland.
Grundläggande information
Grankulla är en av de fyra kommunerna i huvudstadsregionen.
Den ligger mitt i Esbo, 15 kilometer västerut från Helsingfors.
Grankulla har cirka 9 600 invånare, varav 60 procent har finska, 36 procent svenska och 4 procent ett annat språk som modersmål.
Grankullas areal är 6,0 km2.
Information om stadenfinska _ svenska _ engelska
Historia
År 1906 grundades ett aktiebolag i Grankulla som sålde villatomter till invånarna i huvudstadsregionen.
Området hade en direkt förbindelse till Helsingfors.
År 1920 blev villasamhället en köping.
Till en början var största delen av invånarna svenskspråkiga.
År 1972 fick köpingen stadsrättigheter.
Nätmuseetfinska _ svenska
Trafik
Beslutsfattande och påverkan
Religion
Grundläggande information
Historia
Trafik
Huvudstadsregionen har goda kollektivtrafikförbindelser.
I Grankulla finns en järnvägsstation och i staden finns många busslinjer.
Du kan söka information om rutterna i tjänsten Reseplaneraren.
Tjänsten ger dig förslag på olika kollektivtrafikförbindelser från ett ställe till ett annat.
Reseplanerarefinska _ svenska _ engelska
Inom kollektivtrafiken kan du betala med kontanter eller resekort.
I närtågen måste du köpa biljetten i förväg.
Du kan köpa resekortet på Grankulla stadshus.
Du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat.
Stadshuset
Grankullavägen 10
Mån–fre kl. 8.00–15.00; tis, ons, tors även kl. 17.00–19.30
Den närmaste flygstationen är Helsingfors–Vanda flygplats.
Flygplatsenfinska _ svenska _ engelska _ ryska _ kinesiska
Läs mer:
Trafiken i Finland.
Beslutsfattande och påverkan
I Grankulla beslutas ärenden av stadsfullmäktige.
I stadsfullmäktige sitter 35 ledamöter som representerar olika politiska grupper.
Fullmäktige väljs var fjärde år genom kommunalval.
På Grankulla stads webbplats kan du skicka respons till förvaltningen.
Du kan också lämna initiativ och ställa frågor samt kommentera ärenden på finska och på svenska.
Även engelskspråkiga frågor besvaras.
Delta och påverkafinska _ svenska
Religion
Många religiösa samfund är verksamma i Esbo och Helsingfors.
I tjänsten Uskonnot Suomessa kan du söka information enligt det religiösa samfundet och orten.
Religiösa samfundfinska _ engelska
linkkiHelsingfors ortodoxa församling:
Ortodoxa församlingenfinska _ ryska
I Grankulla finns en evangelisk-luthersk kyrka med två församlingar, en finskspråkig och en svenskspråkig.
Församlingarfinska _ svenska
Läs mer: Kulturer och religioner i Finland.
Grundläggande information
Grankulla är en av de fyra kommunerna i huvudstadsregionen.
Den ligger mitt i Esbo, 15 kilometer västerut från Helsingfors.
Grankulla har cirka 9 600 invånare, varav 60 procent har finska, 36 procent svenska och 4 procent ett annat språk som modersmål.
Grankullas areal är 6,0 km2.
Information om stadenfinska _ svenska _ engelska
Historia
År 1906 grundades ett aktiebolag i Grankulla som sålde villatomter till invånarna i huvudstadsregionen.
Området hade en direkt förbindelse till Helsingfors.
År 1920 blev villasamhället en köping.
Till en början var största delen av invånarna svenskspråkiga.
År 1972 fick köpingen stadsrättigheter.
Nätmuseetfinska _ svenska
Evenemang
Bibliotek
Fritidsverksamhet för barn och unga
Föreningar
Evenemang
Evenemang i Grankullafinska _ svenska _ engelska
Vid medborgarinstitutet kan man till exempel skapa konst, göra handarbeten, laga mat, dansa eller motionera.
Man kan även studera språk.
Medborgarinstitutetfinska _ svenska _ engelska
Vid musikinstitutet kan man musicera.
Information om Musikinstitutetfinska _ svenska
Grankulla stad ordnar mångsidig kulturverksamhet.
Kulturtjänsterfinska _ svenska _ engelska
I staden finns också många idrottsmöjligheter.
Idrottstjänsterfinska _ svenska _ engelska
Det finns en biograf i Grankulla.
linkkiBio Grani:
Biograffinska
Läs mer: Fritid.
Bibliotek
På Grankulla stadsbibliotek kan du låna böcker, tidningar, musik, filmer, spel och mycket annat.
I biblioteket kan du också använda dator.
Stadsbiblioteketfinska _ svenska _ engelska
Huvudstadsregionens gemensamma bibliotekstjänstfinska _ svenska _ engelska _ somaliska _ persiska _ arabiska
Läs mer: Bibliotek
Flerspråkiga biblioteket
Flerspråkiga biblioteket ligger i Böle i Helsingfors
Här finns böcker, musik, tidningar och tidskrifter samt ljudböcker på flera olika språk.
Du kan åka till Böle eller beställa material till ditt eget närbibliotek.
linkkiHelsingfors stadsbibliotek:
Flerspråkiga biblioteketfinska _ svenska _ engelska
Hobbyer för barn och unga
Barn och ungdomar kan studera musik vid Grankulla musikinstitut och bildkonst vid Grankulla konstskola.
I Grankulla kan man också motionera på många olika sätt.
På Grankulla ungdomsgård ordnas många olika slags verksamheter.
Ungdomsgårdenfinska _ svenska _ engelska
Läs mer: Hobbyer för barn och unga
Föreningar
I Grankulla finns många olika föreningar, till exempel kulturföreningar och idrottsklubbar.
Föreningarfinska _ svenska
Läs mer: Föreningar.
Läs mer: Fritid i Esbo
Evenemang
Bibliotek
Fritidsverksamhet för barn och unga
Föreningar
Evenemang
Evenemang i Grankullafinska _ svenska _ engelska
Vid medborgarinstitutet kan man till exempel skapa konst, göra handarbeten, laga mat, dansa eller motionera.
Man kan även studera språk.
Medborgarinstitutetfinska _ svenska _ engelska
Vid musikinstitutet kan man musicera.
Information om Musikinstitutetfinska _ svenska
Grankulla stad ordnar mångsidig kulturverksamhet.
Kulturtjänsterfinska _ svenska _ engelska
I staden finns också många idrottsmöjligheter.
Idrottstjänsterfinska _ svenska _ engelska
Det finns en biograf i Grankulla.
linkkiBio Grani:
Biograffinska
Läs mer: Fritid.
Bibliotek
På Grankulla stadsbibliotek kan du låna böcker, tidningar, musik, filmer, spel och mycket annat.
I biblioteket kan du också använda dator.
Stadsbiblioteketfinska _ svenska _ engelska
Huvudstadsregionens gemensamma bibliotekstjänstfinska _ svenska _ engelska _ somaliska _ persiska _ arabiska
Läs mer: Bibliotek
Flerspråkiga biblioteket
Flerspråkiga biblioteket ligger i Böle i Helsingfors
Här finns böcker, musik, tidningar och tidskrifter samt ljudböcker på flera olika språk.
Du kan åka till Böle eller beställa material till ditt eget närbibliotek.
linkkiHelsingfors stadsbibliotek:
Flerspråkiga biblioteketfinska _ svenska _ engelska
Hobbyer för barn och unga
Barn och ungdomar kan studera musik vid Grankulla musikinstitut och bildkonst vid Grankulla konstskola.
I Grankulla kan man också motionera på många olika sätt.
På Grankulla ungdomsgård ordnas många olika slags verksamheter.
Ungdomsgårdenfinska _ svenska _ engelska
Läs mer: Hobbyer för barn och unga
Föreningar
I Grankulla finns många olika föreningar, till exempel kulturföreningar och idrottsklubbar.
Föreningarfinska _ svenska
Läs mer: Föreningar.
Läs mer: Fritid i Esbo
Evenemang
Bibliotek
Fritidsverksamhet för barn och unga
Föreningar
Evenemang
Evenemang i Grankullafinska _ svenska _ engelska
Vid medborgarinstitutet kan man till exempel skapa konst, göra handarbeten, laga mat, dansa eller motionera.
Man kan även studera språk.
Medborgarinstitutetfinska _ svenska _ engelska
Vid musikinstitutet kan man musicera.
Information om Musikinstitutetfinska _ svenska
Grankulla stad ordnar mångsidig kulturverksamhet.
Kulturtjänsterfinska _ svenska _ engelska
I staden finns också många idrottsmöjligheter.
Idrottstjänsterfinska _ svenska _ engelska
Det finns en biograf i Grankulla.
linkkiBio Grani:
Biograffinska
Läs mer: Fritid.
Bibliotek
På Grankulla stadsbibliotek kan du låna böcker, tidningar, musik, filmer, spel och mycket annat.
I biblioteket kan du också använda dator.
Stadsbiblioteketfinska _ svenska _ engelska
Huvudstadsregionens gemensamma bibliotekstjänstfinska _ svenska _ engelska _ somaliska _ persiska _ arabiska
Läs mer: Bibliotek
Flerspråkiga biblioteket
Flerspråkiga biblioteket ligger i Böle i Helsingfors
Här finns böcker, musik, tidningar och tidskrifter samt ljudböcker på flera olika språk.
Du kan åka till Böle eller beställa material till ditt eget närbibliotek.
linkkiHelsingfors stadsbibliotek:
Flerspråkiga biblioteketfinska _ svenska _ engelska
Hobbyer för barn och unga
Barn och ungdomar kan studera musik vid Grankulla musikinstitut och bildkonst vid Grankulla konstskola.
I Grankulla kan man också motionera på många olika sätt.
På Grankulla ungdomsgård ordnas många olika slags verksamheter.
Ungdomsgårdenfinska _ svenska _ engelska
Läs mer: Hobbyer för barn och unga
Föreningar
I Grankulla finns många olika föreningar, till exempel kulturföreningar och idrottsklubbar.
Föreningarfinska _ svenska
Läs mer: Föreningar.
Läs mer: Fritid i Esbo
Social- och krisjouren
Problem med uppehållstillstånd
Brott
Våld
Problem i äktenskap och parförhållande
Behöver du juristhjälp? Barns och ungas problem
Död
Ring nödnumret 112 om det är fråga om en nödsituation.
Via nödnumret kan du tillkalla polis, ambulans eller brandkår.
Ring inte nödnumret om det inte är en nödsituation.
Social- och krisjouren
Social- och krisjouren vid Jorv sjukhus i Esbo hjälper dygnet runt om du eller din familj behöver hjälp i en akut krissituation, till exempel vid våld, problem med barnen eller psykiska problem.
I krissituationer kan du ringa eller åka till jouren.
Esbo social- och krisjour
Jorv sjukhus, Åbovägen 150, Esbo
Tfn (09) 816 42439
Vardagar kl. 15–08, fre–sön och helgdagar dygnet runt
linkkiEsbo stad:
Social- och krisjourenfinska _ svenska _ engelska
linkkiFöreningen för mental hälsa i Finland:
Krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Problem med uppehållstillstånd
Om du har problem med eller det råder oklarheter kring uppehållstillståndet kan du ta kontakt med Migrationsverket, Flyktingrådgivningen eller Helsingfors stads Helsinki-info.
Läs mer: Problem med uppehållstillstånd
Information om uppehållstillståndfinska _ svenska _ engelska
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Helsingfors-infofinska _ svenska _ engelska
Brott
Om du blir utsatt för ett brott, gör en brottsanmälan hos polisen.
Du kan göra brottsanmälan på internet.
Du kan även fylla i en blankett och lämna den till Esbo huvudpolisstation.
Esbo huvudpolisstation
Knektbrovägen 4
Läs mer: Brott
Kontaktuppgifterfinska _ svenska _ engelska
Elektronisk polisanmälanfinska _ svenska _ engelska
Behöver du en jurist?
Västra Nylands rättshjälpsbyrå betjänar invånarna i Grankulla.
Västra Nylands rättshjälpsbyrå
Östanvindsvägen 1 A
Tfn 029 56 61820.
linkkiVästra Nylands rättshjälpsbyrå:
Läs mer:
Behöver du en jurist?
Våld
Om du behöver brådskande hjälp av polisen i nödsituationer, ring nödnumret 112.
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kontakta ett skyddshem.
Tfn (09) 4777 180 (24h)
Hjälp till offer för familjevåldfinska
Föreningen Monika-Naiset Liitto har en jourtelefon för invandrarkvinnor som blivit utsatta för våld.
Tfn 0800 05058
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Invandrarmän som har problem med våld kan få hjälp via tjänsten Miehen linja.
Tfn (09) 276 62899
Hjälp för invandrarmänfinska _ engelska
Läs mer: Våld
Problem i äktenskap och parförhållande
Vid problem i äktenskap och parförhållande kan du få hjälp vid familjerådgivningen.
Familjerådgivningen betjänar invånarna i Grankulla.
Familjerådgivningen
Tfn (09) 5056 297
Familjerådgivningfinska _ svenska
Problem i äktenskap och parförhållande
Barns och ungas problem
Vid problem som gäller barn under skolåldern, kontakta barnrådgivningen.
Barnrådgivningen
Tfn (09) 5056 357 eller (09) 5056 358
Rådgivningsbyråerfinska _ svenska _ engelska
Vid problem som gäller barn i skolåldern hjälper till exempel skolans hälsovårdare.
Skolhälsovårdenfinska _ svenska
Om du behöver råd i frågor kring barns psykiska tillväxt och utveckling, kan du boka en tid hos familjerådgivningen.
Familjerådgivningfinska _ svenska
Du kan prata om dina problem med skolans eller läroanstaltens hälsovårdare eller de vuxna vid ungdomsgården.
Den unga själv eller föräldrarna kan också kontakta familjerådgivningen.
En ung som inte är trygg i sitt eget hem kan kontakta Finlands Röda Kors De ungas skyddshus.
Skyddshuset finns i Stensvik.
De ungas skyddshus
Tfn (09) 8195 5360
linkkiFinlands Röda Kors:
De ungas skyddshusfinska
Läs mer: Barns och ungas problem
Död
Om en nära anhörig till dig avlider oväntat, kan du få stöd av Grankullas grupp för krisbearbetning, tfn 050 344 6652.
Grankulla stad har en egen begravningsplats i Kasabergsområdet.
Den är avsedd för stadens invånare.
Läs mer: Död
Social- och krisjouren
Problem med uppehållstillstånd
Brott
Våld
Problem i äktenskap och parförhållande
Behöver du juristhjälp? Barns och ungas problem
Död
Ring nödnumret 112 om det är fråga om en nödsituation.
Via nödnumret kan du tillkalla polis, ambulans eller brandkår.
Ring inte nödnumret om det inte är en nödsituation.
Social- och krisjouren
Social- och krisjouren vid Jorv sjukhus i Esbo hjälper dygnet runt om du eller din familj behöver hjälp i en akut krissituation, till exempel vid våld, problem med barnen eller psykiska problem.
I krissituationer kan du ringa eller åka till jouren.
Esbo social- och krisjour
Jorv sjukhus, Åbovägen 150, Esbo
Tfn (09) 816 42439
Vardagar kl. 15–08, fre–sön och helgdagar dygnet runt
linkkiEsbo stad:
Social- och krisjourenfinska _ svenska _ engelska
linkkiFöreningen för mental hälsa i Finland:
Krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Problem med uppehållstillstånd
Om du har problem med eller det råder oklarheter kring uppehållstillståndet kan du ta kontakt med Migrationsverket, Flyktingrådgivningen eller Helsingfors stads Helsinki-info.
Läs mer: Problem med uppehållstillstånd
Information om uppehållstillståndfinska _ svenska _ engelska
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Helsingfors-infofinska _ svenska _ engelska
Brott
Om du blir utsatt för ett brott, gör en brottsanmälan hos polisen.
Du kan göra brottsanmälan på internet.
Du kan även fylla i en blankett och lämna den till Esbo huvudpolisstation.
Esbo huvudpolisstation
Knektbrovägen 4
Läs mer: Brott
Kontaktuppgifterfinska _ svenska _ engelska
Elektronisk polisanmälanfinska _ svenska _ engelska
Behöver du en jurist?
Västra Nylands rättshjälpsbyrå betjänar invånarna i Grankulla.
Västra Nylands rättshjälpsbyrå
Östanvindsvägen 1 A
Tfn 029 56 61820.
linkkiVästra Nylands rättshjälpsbyrå:
Läs mer:
Behöver du en jurist?
Våld
Om du behöver brådskande hjälp av polisen i nödsituationer, ring nödnumret 112.
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kontakta ett skyddshem.
Tfn (09) 4777 180 (24h)
Hjälp till offer för familjevåldfinska
Föreningen Monika-Naiset Liitto har en jourtelefon för invandrarkvinnor som blivit utsatta för våld.
Tfn 0800 05058
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Invandrarmän som har problem med våld kan få hjälp via tjänsten Miehen linja.
Tfn (09) 276 62899
Hjälp för invandrarmänfinska _ engelska
Läs mer: Våld
Problem i äktenskap och parförhållande
Vid problem i äktenskap och parförhållande kan du få hjälp vid familjerådgivningen.
Familjerådgivningen betjänar invånarna i Grankulla.
Familjerådgivningen
Tfn (09) 5056 297
Familjerådgivningfinska _ svenska
Problem i äktenskap och parförhållande
Barns och ungas problem
Vid problem som gäller barn under skolåldern, kontakta barnrådgivningen.
Barnrådgivningen
Tfn (09) 5056 357 eller (09) 5056 358
Rådgivningsbyråerfinska _ svenska _ engelska
Vid problem som gäller barn i skolåldern hjälper till exempel skolans hälsovårdare.
Skolhälsovårdenfinska _ svenska
Om du behöver råd i frågor kring barns psykiska tillväxt och utveckling, kan du boka en tid hos familjerådgivningen.
Familjerådgivningfinska _ svenska
Du kan prata om dina problem med skolans eller läroanstaltens hälsovårdare eller de vuxna vid ungdomsgården.
Den unga själv eller föräldrarna kan också kontakta familjerådgivningen.
En ung som inte är trygg i sitt eget hem kan kontakta Finlands Röda Kors De ungas skyddshus.
Skyddshuset finns i Stensvik.
De ungas skyddshus
Tfn (09) 8195 5360
linkkiFinlands Röda Kors:
De ungas skyddshusfinska
Läs mer: Barns och ungas problem
Död
Om en nära anhörig till dig avlider oväntat, kan du få stöd av Grankullas grupp för krisbearbetning, tfn 050 344 6652.
Grankulla stad har en egen begravningsplats i Kasabergsområdet.
Den är avsedd för stadens invånare.
Läs mer: Död
Social- och krisjouren
Problem med uppehållstillstånd
Brott
Våld
Problem i äktenskap och parförhållande
Behöver du juristhjälp? Barns och ungas problem
Död
Ring nödnumret 112 om det är fråga om en nödsituation.
Via nödnumret kan du tillkalla polis, ambulans eller brandkår.
Ring inte nödnumret om det inte är en nödsituation.
Social- och krisjouren
Social- och krisjouren vid Jorv sjukhus i Esbo hjälper dygnet runt om du eller din familj behöver hjälp i en akut krissituation, till exempel vid våld, problem med barnen eller psykiska problem.
I krissituationer kan du ringa eller åka till jouren.
Esbo social- och krisjour
Jorv sjukhus, Åbovägen 150, Esbo
Tfn (09) 816 42439
Vardagar kl. 15–08, fre–sön och helgdagar dygnet runt
linkkiEsbo stad:
Social- och krisjourenfinska _ svenska _ engelska
linkkiFöreningen för mental hälsa i Finland:
Krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Problem med uppehållstillstånd
Om du har problem med eller det råder oklarheter kring uppehållstillståndet kan du ta kontakt med Migrationsverket, Flyktingrådgivningen eller Helsingfors stads Helsinki-info.
Läs mer: Problem med uppehållstillstånd
Information om uppehållstillståndfinska _ svenska _ engelska
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Helsingfors-infofinska _ svenska _ engelska
Brott
Om du blir utsatt för ett brott, gör en brottsanmälan hos polisen.
Du kan göra brottsanmälan på internet.
Du kan även fylla i en blankett och lämna den till Esbo huvudpolisstation.
Esbo huvudpolisstation
Knektbrovägen 4
Läs mer: Brott
Kontaktuppgifterfinska _ svenska _ engelska
Elektronisk polisanmälanfinska _ svenska _ engelska
Behöver du en jurist?
Västra Nylands rättshjälpsbyrå betjänar invånarna i Grankulla.
Västra Nylands rättshjälpsbyrå
Östanvindsvägen 1 A
Tfn 029 56 61820.
linkkiVästra Nylands rättshjälpsbyrå:
Läs mer:
Behöver du en jurist?
Våld
Om du behöver brådskande hjälp av polisen i nödsituationer, ring nödnumret 112.
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kontakta ett skyddshem.
Tfn (09) 4777 180 (24h)
Hjälp till offer för familjevåldfinska
Föreningen Monika-Naiset Liitto har en jourtelefon för invandrarkvinnor som blivit utsatta för våld.
Tfn 0800 05058
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Invandrarmän som har problem med våld kan få hjälp via tjänsten Miehen linja.
Tfn (09) 276 62899
Hjälp för invandrarmänfinska _ engelska
Läs mer: Våld
Problem i äktenskap och parförhållande
Vid problem i äktenskap och parförhållande kan du få hjälp vid familjerådgivningen.
Familjerådgivningen betjänar invånarna i Grankulla.
Familjerådgivningen
Tfn (09) 5056 297
Familjerådgivningfinska _ svenska
Problem i äktenskap och parförhållande
Barns och ungas problem
Vid problem som gäller barn under skolåldern, kontakta barnrådgivningen.
Barnrådgivningen
Tfn (09) 5056 357 eller (09) 5056 358
Rådgivningsbyråerfinska _ svenska _ engelska
Vid problem som gäller barn i skolåldern hjälper till exempel skolans hälsovårdare.
Skolhälsovårdenfinska _ svenska
Om du behöver råd i frågor kring barns psykiska tillväxt och utveckling, kan du boka en tid hos familjerådgivningen.
Familjerådgivningfinska _ svenska
Du kan prata om dina problem med skolans eller läroanstaltens hälsovårdare eller de vuxna vid ungdomsgården.
Den unga själv eller föräldrarna kan också kontakta familjerådgivningen.
En ung som inte är trygg i sitt eget hem kan kontakta Finlands Röda Kors De ungas skyddshus.
Skyddshuset finns i Stensvik.
De ungas skyddshus
Tfn (09) 8195 5360
linkkiFinlands Röda Kors:
De ungas skyddshusfinska
Läs mer: Barns och ungas problem
Död
Om en nära anhörig till dig avlider oväntat, kan du få stöd av Grankullas grupp för krisbearbetning, tfn 050 344 6652.
Grankulla stad har en egen begravningsplats i Kasabergsområdet.
Den är avsedd för stadens invånare.
Läs mer: Död
Äktenskap
Skilsmässa
Barn vid skilsmässa
Vård av barnet
Äktenskap
Före äktenskapet ska du skriftligt begära prövning av hinder mot äktenskap.
Hindersprövningen görs i magistraten.
Läs mer: Prövning av hinder mot äktenskap, Äktenskap
Kontaktuppgifter till magistratfinska _ svenska _ engelska
Skilsmässa
Kvinnan eller mannen kan lämna in skilsmässoansökan i Västra Nylands tingsrätts kansli.
Du kan också söka skilsmässa ensam, utan din makes eller makas samtycke.
Du kan skicka in ansökan till tingsrättens kansli per post, fax eller via e-post.
Västra Nylands tingsrätt
Tfn 029 5645 000
Läs mer: Skilsmässa
linkkiVästra Nylands tingsrätt:
Kontaktuppgifterfinska _ svenska
Barn vid skilsmässa
Om du har barn och ska skilja dig, ta kontakt med barnatillsyningsmannen.
Socialväsendet bekräftar ett avtal om barnens boende, vårdnad, umgängesrätt och underhållsbidrag.
Läs mer: Barn vid skilsmässa
Vårdnad om barn och umgängesrättfinska _ svenska
Vård av barnet
På InfoFinlands sida Utbildning i Grankulla finns information om dagvård för barn.
Vård av barnet i hemmet
Om du sköter ditt barn hemma kan du delta i Grankulla stads öppna familjeverksamhet. Där kan du träffa andra barnfamiljer.
Läs mer: Stöd för vård av barn i hemmet
Öppen familjeverksamhetfinska _ svenska
Stöd för hemvård av barnfinska _ svenska
Äktenskap
Skilsmässa
Barn vid skilsmässa
Vård av barnet
Äktenskap
Före äktenskapet ska du skriftligt begära prövning av hinder mot äktenskap.
Hindersprövningen görs i magistraten.
Läs mer: Prövning av hinder mot äktenskap, Äktenskap
Kontaktuppgifter till magistratfinska _ svenska _ engelska
Skilsmässa
Kvinnan eller mannen kan lämna in skilsmässoansökan i Västra Nylands tingsrätts kansli.
Du kan också söka skilsmässa ensam, utan din makes eller makas samtycke.
Du kan skicka in ansökan till tingsrättens kansli per post, fax eller via e-post.
Västra Nylands tingsrätt
Tfn 029 5645 000
Läs mer: Skilsmässa
linkkiVästra Nylands tingsrätt:
Kontaktuppgifterfinska _ svenska
Barn vid skilsmässa
Om du har barn och ska skilja dig, ta kontakt med barnatillsyningsmannen.
Socialväsendet bekräftar ett avtal om barnens boende, vårdnad, umgängesrätt och underhållsbidrag.
Läs mer: Barn vid skilsmässa
Vårdnad om barn och umgängesrättfinska _ svenska
Vård av barnet
På InfoFinlands sida Utbildning i Grankulla finns information om dagvård för barn.
Vård av barnet i hemmet
Om du sköter ditt barn hemma kan du delta i Grankulla stads öppna familjeverksamhet. Där kan du träffa andra barnfamiljer.
Läs mer: Stöd för vård av barn i hemmet
Öppen familjeverksamhetfinska _ svenska
Stöd för hemvård av barnfinska _ svenska
Äktenskap
Skilsmässa
Barn vid skilsmässa
Vård av barnet
Äktenskap
Före äktenskapet ska du skriftligt begära prövning av hinder mot äktenskap.
Hindersprövningen görs i magistraten.
Läs mer: Prövning av hinder mot äktenskap, Äktenskap
Kontaktuppgifter till magistratfinska _ svenska _ engelska
Skilsmässa
Kvinnan eller mannen kan lämna in skilsmässoansökan i Västra Nylands tingsrätts kansli.
Du kan också söka skilsmässa ensam, utan din makes eller makas samtycke.
Du kan skicka in ansökan till tingsrättens kansli per post, fax eller via e-post.
Västra Nylands tingsrätt
Tfn 029 5645 000
Läs mer: Skilsmässa
linkkiVästra Nylands tingsrätt:
Kontaktuppgifterfinska _ svenska
Barn vid skilsmässa
Om du har barn och ska skilja dig, ta kontakt med barnatillsyningsmannen.
Socialväsendet bekräftar ett avtal om barnens boende, vårdnad, umgängesrätt och underhållsbidrag.
Läs mer: Barn vid skilsmässa
Vårdnad om barn och umgängesrättfinska _ svenska
Vård av barnet
På InfoFinlands sida Utbildning i Grankulla finns information om dagvård för barn.
Vård av barnet i hemmet
Om du sköter ditt barn hemma kan du delta i Grankulla stads öppna familjeverksamhet. Där kan du träffa andra barnfamiljer.
Läs mer: Stöd för vård av barn i hemmet
Öppen familjeverksamhetfinska _ svenska
Stöd för hemvård av barnfinska _ svenska
Hälsovårdstjänsterna i Grankulla
Barns hälsa
Äldre människors hälsa
Tandvård
Mental hälsa
Sexualhälsa
När du väntar barn
Handikappade personer
Ring nödnumret 112 om det är fråga om en brådskande nödsituation.
Ring nödnumret till exempel vid en allvarlig olycka eller när någon drabbas av en sjukdomsattack.
Ring inte nödnumret om det inte är en nödsituation.
Om du har din hemkommun i Grankulla, kan du utnyttja de offentliga hälso- och sjukvårdstjänsterna.
Offentliga hälso- och sjukvårdstjänster tillhandahålls till exempel vid hälsostationer, tandkliniker, rådgivningsbyråer och sjukhus.
Om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna, kan du söka dig till en privat läkarstation.
På en privat läkarstation måste du betala samtliga kostnader själv.
Läs mer: Hälsa
Hälsovårdstjänsterna i Grankulla
I Grankulla tillhandahålls offentliga hälso- och sjukvårdstjänster på hälsostationen.
På hälsostationen finns läkarens, sjukskötarens och hälsovårdarens mottagningar.
Hälsostationen har öppet vardagar kl. 8.00–16.00.
Om du behöver vård under samma dag ska du kontakta hälsostationen direkt på morgonen när hälsostationen öppnar.
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
Tfn (09) 8789 1300
Hälsostationenfinska _ svenska _ engelska
Privata hälsotjänster
Information om privata hälsotjänster hittar du på sidorna Hälsa i Esbo och Hälsa i Helsingfors.
Läkemedel
Du kan köpa läkemedel på apoteket.
Adressen till apoteket i Grankulla är Kyrkovägen 15, Grankulla.
Läs mer: Läkemedel.
Apotekfinska _ svenska
linkkiApotekareförbundet:
Hälsovård för papperslösa
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärvård.
Tfn 044 977 4547
Kontaktuppgifterfinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Läs mer: Hälsovårdstjänster i Finland
Kvällstid och under veckoslut har hälsostationen stängt.
Då vårdas akuta sjukdomar och olycksfall på jourmottagningen.
Den närmaste jourmottagningen finns vid Jorv sjukhus i Esbo.
Ring den kostnadsfria Jourhjälpen på tfn 116 117 innan du kommer till jourmottagningen.
Jouren vid Jorv sjukhus
Åbovägen 150
Tfn (09) 4711
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Jourfinska _ svenska _ engelska
Läs mer: Hälsovårdstjänster i Finland
Barns hälsa
I hälso- och sjukvården av barn under skolåldern får man hjälp av rådgivningens hälsovårdare och läkare.
Dem kan du fråga om råd och få stöd i föräldraskapet och fostran av barn.
På rådgivningsbyrån följs barnets hälsa och tillväxt.
Rådgivningsbyråerfinska _ svenska _ engelska
När barnet blir sjukt ska du vid behov kontakta Grankulla hälsostation.
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
Tfn (09) 8789 1300
Hälsostationenfinska _ svenska _ engelska
Skolhälsovårdaren tar hand om skolbarns hälsa.
Skolhälsovårdenfinska _ svenska
Under kvällar och veckoslut finns jourmottagningen för barn under 16 år vid Jorv sjukhus i Esbo och på Barnkliniken i Helsingfors.
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Jourmottagning för barnfinska _ svenska _ engelska
Läs mer: Barns hälsa
Äldre människors hälsa
Om du är över 65 år kan du kontakta seniorrådgivningen vid Grankulla hälsostation.
Seniorrådgivningenfinska _ svenska
Serviceguide för seniorer(pdf, 1,8 MB)finska _ svenska
Tandvård
Tidsbeställningen till tandkliniken vid Grankulla hälsostation mån–fre:
Tfn (09) 505 6379
Jourmottagningen vid Haartmanska sjukhuset har öppet vardagar kl. 14–21 och lör–sön kl. 8–21.
Tfn (09) 310 49999
Mun- och tandhälsovårdenfinska _ svenska
Privat tandvård
I Grankulla finns också privata tandläkare.
Om om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna, kan du gå till en privat tandläkare.
Privat tandvård är dyrare än offentlig tandvård.
Privat tandläkarefinska _ svenska
Läs mer: Tandvård
Mental hälsa
Om du behöver psykisk hjälp och psykiskt stöd kan du kontakta hälsostationen.
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
Tfn (09) 5056 600
Mental hälsafinska _ svenska
Esbo social- och krisjour vid Jorv sjukhus betjänar personer som bor i Grankulla.
I krissituationer kan du ringa eller åka till jouren.
Esbo social- och krisjour
Jorv sjukhus, Åbovägen 150, Esbo
Tfn (09) 816 42439
Vardagar kl. 15–08, fre–sön och helgdagar dygnet runt
Kristjänsterfinska _ svenska
Läs mer: Mental hälsa
Sexualhälsa
Vid mödra- och preventivrådgivningen får du hjälp med graviditetsprevention och familjeplanering.
Könssjukdomar behandlas på hälsostationen och på polikliniken för könssjukdomar i Helsingfors. .
Hälsostationenfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Polikliniken för könssjukdomarfinska _ svenska _ engelska
När du väntar barn
Vid mödrarådgivningen följs moderns, fostrets och hela familjens hälsotillstånd under graviditeten.
Kontakta rådgivningsbyrån när du upptäcker att du är gravid.
Tidsbokning vardagar kl. 12–13
Tfn (09) 8789 1344
Rådgivningsbyråerfinska _ svenska _ engelska
Det närmaste förlossningssjukhuset är Jorv sjukhus i Esbo.
Om du vill kan du även föda barnet på något annat sjukhus inom Helsingfors och Nylands sjukvårdsdistrikt (HNS).
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Val av förlossningssjukhusfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Läs mer: Förlossning
Handikappade personer
Grankulla stad erbjuder olika tjänster för handikappade, till exempel hjälpmedel och dagverksamhet.
Du kan fråga om tjänsterna för handikappade hos socialarbetaren för ditt område.
Tjänster inom handikappvårdenfinska _ svenska
Läs mer: Handikappade personer
Hälsovårdstjänsterna i Grankulla
Barns hälsa
Äldre människors hälsa
Tandvård
Mental hälsa
Sexualhälsa
När du väntar barn
Handikappade personer
Ring nödnumret 112 om det är fråga om en brådskande nödsituation.
Ring nödnumret till exempel vid en allvarlig olycka eller när någon drabbas av en sjukdomsattack.
Ring inte nödnumret om det inte är en nödsituation.
Om du har din hemkommun i Grankulla, kan du utnyttja de offentliga hälso- och sjukvårdstjänsterna.
Offentliga hälso- och sjukvårdstjänster tillhandahålls till exempel vid hälsostationer, tandkliniker, rådgivningsbyråer och sjukhus.
Om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna, kan du söka dig till en privat läkarstation.
På en privat läkarstation måste du betala samtliga kostnader själv.
Läs mer: Hälsa
Hälsovårdstjänsterna i Grankulla
I Grankulla tillhandahålls offentliga hälso- och sjukvårdstjänster på hälsostationen.
På hälsostationen finns läkarens, sjukskötarens och hälsovårdarens mottagningar.
Hälsostationen har öppet vardagar kl. 8.00–16.00.
Om du behöver vård under samma dag ska du kontakta hälsostationen direkt på morgonen när hälsostationen öppnar.
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
Tfn (09) 8789 1300
Hälsostationenfinska _ svenska _ engelska
Privata hälsotjänster
Information om privata hälsotjänster hittar du på sidorna Hälsa i Esbo och Hälsa i Helsingfors.
Läkemedel
Du kan köpa läkemedel på apoteket.
Adressen till apoteket i Grankulla är Kyrkovägen 15, Grankulla.
Läs mer: Läkemedel.
Apotekfinska _ svenska
linkkiApotekareförbundet:
Hälsovård för papperslösa
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärvård.
Tfn 044 977 4547
Kontaktuppgifterfinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Läs mer: Hälsovårdstjänster i Finland
Kvällstid och under veckoslut har hälsostationen stängt.
Då vårdas akuta sjukdomar och olycksfall på jourmottagningen.
Den närmaste jourmottagningen finns vid Jorv sjukhus i Esbo.
Ring den kostnadsfria Jourhjälpen på tfn 116 117 innan du kommer till jourmottagningen.
Jouren vid Jorv sjukhus
Åbovägen 150
Tfn (09) 4711
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Jourfinska _ svenska _ engelska
Läs mer: Hälsovårdstjänster i Finland
Barns hälsa
I hälso- och sjukvården av barn under skolåldern får man hjälp av rådgivningens hälsovårdare och läkare.
Dem kan du fråga om råd och få stöd i föräldraskapet och fostran av barn.
På rådgivningsbyrån följs barnets hälsa och tillväxt.
Rådgivningsbyråerfinska _ svenska _ engelska
När barnet blir sjukt ska du vid behov kontakta Grankulla hälsostation.
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
Tfn (09) 8789 1300
Hälsostationenfinska _ svenska _ engelska
Skolhälsovårdaren tar hand om skolbarns hälsa.
Skolhälsovårdenfinska _ svenska
Under kvällar och veckoslut finns jourmottagningen för barn under 16 år vid Jorv sjukhus i Esbo och på Barnkliniken i Helsingfors.
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Jourmottagning för barnfinska _ svenska _ engelska
Läs mer: Barns hälsa
Äldre människors hälsa
Om du är över 65 år kan du kontakta seniorrådgivningen vid Grankulla hälsostation.
Information om tjänster för äldrefinska _ svenska
Serviceguide för seniorer(pdf, 1,8 MB)finska _ svenska
Äldre människor
Tandvård
Tidsbeställningen till tandkliniken vid Grankulla hälsostation mån–fre:
Tfn (09) 505 6379
Jourmottagningen vid Haartmanska sjukhuset har öppet vardagar kl. 14–21 och lör–sön kl. 8–21.
Tfn (09) 310 49999
Mun- och tandhälsovårdenfinska _ svenska
Privat tandvård
I Grankulla finns också privata tandläkare.
Om om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna, kan du gå till en privat tandläkare.
Privat tandvård är dyrare än offentlig tandvård.
Privat tandläkarefinska _ svenska
Läs mer: Tandvård
Mental hälsa
Om du behöver psykisk hjälp och psykiskt stöd kan du kontakta hälsostationen.
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
Tfn (09) 5056 600
Mental hälsafinska _ svenska
Esbo social- och krisjour vid Jorv sjukhus betjänar personer som bor i Grankulla.
I krissituationer kan du ringa eller åka till jouren.
Esbo social- och krisjour
Jorv sjukhus, Åbovägen 150, Esbo
Tfn (09) 816 42439
Vardagar kl. 15–08, fre–sön och helgdagar dygnet runt
Kristjänsterfinska _ svenska
Läs mer: Mental hälsa
Sexualhälsa
Vid mödra- och preventivrådgivningen får du hjälp med graviditetsprevention och familjeplanering.
Könssjukdomar behandlas på hälsostationen och på polikliniken för könssjukdomar i Helsingfors. .
Hälsostationenfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Polikliniken för könssjukdomarfinska _ svenska _ engelska
När du väntar barn
Vid mödrarådgivningen följs moderns, fostrets och hela familjens hälsotillstånd under graviditeten.
Kontakta rådgivningsbyrån när du upptäcker att du är gravid.
Tidsbokning vardagar kl. 12–13
Tfn (09) 8789 1344
Rådgivningsbyråerfinska _ svenska _ engelska
Det närmaste förlossningssjukhuset är Jorv sjukhus i Esbo.
Om du vill kan du även föda barnet på något annat sjukhus inom Helsingfors och Nylands sjukvårdsdistrikt (HNS).
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Val av förlossningssjukhusfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Läs mer: Förlossning
Handikappade personer
Grankulla stad erbjuder olika tjänster för handikappade, till exempel hjälpmedel och dagverksamhet.
Du kan fråga om tjänsterna för handikappade hos socialarbetaren för ditt område.
Tjänster inom handikappvårdenfinska _ svenska
Läs mer: Handikappade personer
Hälsovårdstjänsterna i Grankulla
Barns hälsa
Äldre människors hälsa
Tandvård
Mental hälsa
Sexualhälsa
När du väntar barn
Handikappade personer
Ring nödnumret 112 om det är fråga om en brådskande nödsituation.
Ring nödnumret till exempel vid en allvarlig olycka eller när någon drabbas av en sjukdomsattack.
Ring inte nödnumret om det inte är en nödsituation.
Om du har din hemkommun i Grankulla, kan du utnyttja de offentliga hälso- och sjukvårdstjänsterna.
Offentliga hälso- och sjukvårdstjänster tillhandahålls till exempel vid hälsostationer, tandkliniker, rådgivningsbyråer och sjukhus.
Om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna, kan du söka dig till en privat läkarstation.
På en privat läkarstation måste du betala samtliga kostnader själv.
Läs mer: Hälsa
Hälsovårdstjänsterna i Grankulla
I Grankulla tillhandahålls offentliga hälso- och sjukvårdstjänster på hälsostationen.
På hälsostationen finns läkarens, sjukskötarens och hälsovårdarens mottagningar.
Hälsostationen har öppet vardagar kl. 8.00–16.00.
Om du behöver vård under samma dag ska du kontakta hälsostationen direkt på morgonen när hälsostationen öppnar.
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
Tfn (09) 8789 1300
Hälsostationenfinska _ svenska
Privata hälsotjänster
Information om privata hälsotjänster hittar du på sidorna Hälsa i Esbo och Hälsa i Helsingfors.
Läkemedel
Du kan köpa läkemedel på apoteket.
Adressen till apoteket i Grankulla är Kyrkovägen 15, Grankulla.
Läs mer: Läkemedel.
Apotekfinska _ svenska
linkkiApotekareförbundet:
Hälsovård för papperslösa
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärvård.
Tfn 044 977 4547
Kontaktuppgifterfinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Läs mer: Hälsovårdstjänster i Finland
Kvällstid och under veckoslut har hälsostationen stängt.
Då vårdas akuta sjukdomar och olycksfall på jourmottagningen.
Den närmaste jourmottagningen finns vid Jorv sjukhus i Esbo.
Ring den kostnadsfria Jourhjälpen på tfn 116 117 innan du kommer till jourmottagningen.
Jouren vid Jorv sjukhus
Åbovägen 150
Tfn (09) 4711
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Jourfinska _ svenska _ engelska
Läs mer: Hälsovårdstjänster i Finland
Barns hälsa
I hälso- och sjukvården av barn under skolåldern får man hjälp av rådgivningens hälsovårdare och läkare.
Dem kan du fråga om råd och få stöd i föräldraskapet och fostran av barn.
På rådgivningsbyrån följs barnets hälsa och tillväxt.
Rådgivningsbyråerfinska _ svenska _ engelska
När barnet blir sjukt ska du vid behov kontakta Grankulla hälsostation.
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
Tfn (09) 8789 1300
Hälsostationenfinska _ svenska
Skolhälsovårdaren tar hand om skolbarns hälsa.
Skolhälsovårdenfinska _ svenska
Under kvällar och veckoslut finns jourmottagningen för barn under 16 år vid Jorv sjukhus i Esbo och på Barnkliniken i Helsingfors.
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Jourmottagning för barnfinska _ svenska _ engelska
Läs mer: Barns hälsa
Äldre människors hälsa
Om du är över 65 år kan du kontakta seniorrådgivningen vid Grankulla hälsostation.
Information om tjänster för äldrefinska _ svenska
Äldre människor
Tandvård
Tidsbeställningen till tandkliniken vid Grankulla hälsostation mån–fre:
Tfn (09) 505 6379
Jourmottagningen vid Haartmanska sjukhuset har öppet vardagar kl. 14–21 och lör–sön kl. 8–21.
Tfn (09) 310 49999
Mun- och tandhälsovårdenfinska _ svenska
Privat tandvård
I Grankulla finns också privata tandläkare.
Om om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna, kan du gå till en privat tandläkare.
Privat tandvård är dyrare än offentlig tandvård.
Privat tandläkarefinska _ svenska
Läs mer: Tandvård
Mental hälsa
Om du behöver psykisk hjälp och psykiskt stöd kan du kontakta hälsostationen.
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
Tfn (09) 5056 600
Mental hälsafinska _ svenska
Esbo social- och krisjour vid Jorv sjukhus betjänar personer som bor i Grankulla.
I krissituationer kan du ringa eller åka till jouren.
Esbo social- och krisjour
Jorv sjukhus, Åbovägen 150, Esbo
Tfn (09) 816 42439
Vardagar kl. 15–08, fre–sön och helgdagar dygnet runt
Kristjänsterfinska _ svenska
Läs mer: Mental hälsa
Sexualhälsa
Vid mödra- och preventivrådgivningen får du hjälp med graviditetsprevention och familjeplanering.
Könssjukdomar behandlas på hälsostationen och på polikliniken för könssjukdomar i Helsingfors. .
Hälsostationenfinska _ svenska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Polikliniken för könssjukdomarfinska _ svenska _ engelska
När du väntar barn
Vid mödrarådgivningen följs moderns, fostrets och hela familjens hälsotillstånd under graviditeten.
Kontakta rådgivningsbyrån när du upptäcker att du är gravid.
Tidsbokning vardagar kl. 12–13
Tfn (09) 8789 1344
Rådgivningsbyråerfinska _ svenska _ engelska
Det närmaste förlossningssjukhuset är Jorv sjukhus i Esbo.
Om du vill kan du även föda barnet på något annat sjukhus inom Helsingfors och Nylands sjukvårdsdistrikt (HNS).
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Val av förlossningssjukhusfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Läs mer: Förlossning
Handikappade personer
Grankulla stad erbjuder olika tjänster för handikappade, till exempel hjälpmedel och dagverksamhet.
Du kan fråga om tjänsterna för handikappade hos socialarbetaren för ditt område.
Tjänster inom handikappvårdenfinska _ svenska
Läs mer: Handikappade personer
Dagvård
Förskoleundervisning
Grundläggande utbildning
Yrkesutbildning
Gymnasium
Högskoleutbildning
Andra studiemöjligheter
Dagvård
I Grankulla finns stadens egna daghem, privata daghem och privata familjedagvårdare.
Dagvård fås på finska och på svenska.
I Grankulla finns också ett engelskspråkigt daghem.
Ansök om dagvårdsplats för ditt barn minst fyra månader innan barnet ska börja i dagvården.
Om du ansöker om dagvårdplats för första gången ska du använda den elektroniska ansökan.
Du kan också hämta ansökningsblanketten på daghemmet eller vid informationen i stadshuset.
Lämna in ansökan till daghemmet eller stadshuset.
Familjer som bor i Grankulla kan också söka dagvårdsplats till sitt barn i Esbo, Helsingfors eller Vanda.
Du ska ändå lämna in din ansökan i Grankulla.
Mer information finns på tjänsten HelsingforsRegionen.fi.
Läs mer: Dagvård
Dagvård och förskoleundervisningfinska _ svenska _ engelska
Ansökan om dagvårdsplatsfinska _ svenska
Engelsk-finskspråkigt daghemfinska _ engelska
Dagvårdens samanvändningsområdefinska _ svenska _ engelska
Förskoleundervisning
I Grankulla anordnas förskoleundervisningen i daghemmen.
Förskoleundervisningen börjar i augusti och ansökningstiden är i januari.
Läs mer: Förskoleundervisning
Information om förskoleundervisningenfinska _ svenska _ engelska
Grundläggande utbildning
I Grankulla finns både en finsk- och en svenskspråkig grundskola. Anmälan till grundskolan ska ske i början av året.
Om du har frågor om den grundläggande utbildningen kan du kontakta skolbyrån.
Skolbyrån
Grankulla stadshus
Grankullavägen 10
02700 Grankulla
Tfn (09) 50 561 (växel)
Grundläggande utbildning
Grundläggande utbildning och gymnasiumfinska _ svenska _ engelska
Internationella skolor i huvudstadsregionenfinska
linkkiExpatFinland.fi:
Internationella skolor i huvudstadsregionenengelska
Yrkesutbildning
De närmaste yrkesläroanstalterna finns i Esbo och Helsingfors.
Läs mer: Yrkesutbildning
Yrkesutbildningfinska _ engelska
Yrkesinriktad utbildningfinska
Gymnasium
I Grankulla finns två gymnasier, ett finskspråkigt och ett svenskspråkigt.
I Esbo finns ett vuxengymnasium där vuxna kan avlägga gymnasiet och studentexamen.
Läs mer: Gymnasium
Grundläggande utbildning och gymnasiumfinska _ svenska _ engelska
linkkiEsbo stad:
Vuxengymnasietfinska
Högskoleutbildning
I anslutning till folkhögskolan Työväen Akatemia i Grankulla finns en enhet för Humanistiska Yrkeshögskolan, där du kan avlägga yrkeshögskoleexamen för kulturproducenter.
Vid yrkeshögskolorna och universiteten i Esbo och Helsingfors kan du studera inom många områden.
Mer information om högskolorna i Esbo och Helsingfors hittar du på städernas webbplatser.
Läs mer: Högskoleutbildning
linkkiHumanistiska yrkeshögskolan:
Information om Humanistiska yrkeshögskolanfinska _ engelska
linkkiEsbo stad:
Högskolorfinska _ engelska
Högskolorfinska
Andra studiemöjligheter
Vid Grankulla medborgarinstitut kan du studera till exempel språk, handarbete och matlagning eller delta i ledd motion.
Medborgarinstitutetfinska _ svenska _ engelska
Vid Grankulla konstskola kan barn och unga studera bildkonst och vid Grankulla musikinstitut kan barn och vuxna studera musik.
Information om Konstskolanfinska _ svenska
Information om Musikinstitutetfinska _ svenska
I Grankulla ligger Finska Bibelinstitutet.
Vid institutet kan du avlägga enskilda kurser eller studera på någon av institutets studielinjer.
Studierna på studielinjerna pågår i 1–2 år.
Vid bibelinstitutet finns även en studielinje som är särskilt avsedd för invandrare.
Kristliga folkhögskolanfinska _ engelska
Folkhögskolan Työväen Akatemia tillhandahåller undervisning inom många akademiska discipliner samt träning för dem som vill läsa på universitet.
Information om Työväen Akatemiafinska _ engelska
Läs mer: Andra studiemöjligheter
Dagvård
Förskoleundervisning
Grundläggande utbildning
Yrkesutbildning
Gymnasium
Högskoleutbildning
Andra studiemöjligheter
Dagvård
I Grankulla finns stadens egna daghem, privata daghem och privata familjedagvårdare.
Dagvård fås på finska och på svenska.
I Grankulla finns också ett engelskspråkigt daghem.
Ansök om dagvårdsplats för ditt barn minst fyra månader innan barnet ska börja i dagvården.
Om du ansöker om dagvårdplats för första gången ska du använda den elektroniska ansökan.
Du kan också hämta ansökningsblanketten på daghemmet eller vid informationen i stadshuset.
Lämna in ansökan till daghemmet eller stadshuset.
Familjer som bor i Grankulla kan också söka dagvårdsplats till sitt barn i Esbo, Helsingfors eller Vanda.
Du ska ändå lämna in din ansökan i Grankulla.
Mer information finns på tjänsten HelsingforsRegionen.fi.
Läs mer: Dagvård
Dagvård och förskoleundervisningfinska _ svenska _ engelska
Ansökan om dagvårdsplatsfinska _ svenska
Engelsk-finskspråkigt daghemfinska _ engelska
Dagvårdens samanvändningsområdefinska _ svenska _ engelska
Förskoleundervisning
I Grankulla anordnas förskoleundervisningen i daghemmen.
Förskoleundervisningen börjar i augusti och ansökningstiden är i januari.
Läs mer: Förskoleundervisning
Information om förskoleundervisningenfinska _ svenska _ engelska
Grundläggande utbildning
I Grankulla finns både en finsk- och en svenskspråkig grundskola. Anmälan till grundskolan ska ske i början av året.
Om du har frågor om den grundläggande utbildningen kan du kontakta skolbyrån.
Skolbyrån
Grankulla stadshus
Grankullavägen 10
02700 Grankulla
Tfn (09) 50 561 (växel)
Grundläggande utbildning
Grundläggande utbildning och gymnasiumfinska _ svenska _ engelska
Internationella skolor i huvudstadsregionenfinska
linkkiExpatFinland.fi:
Internationella skolor i huvudstadsregionenengelska
Yrkesutbildning
De närmaste yrkesläroanstalterna finns i Esbo och Helsingfors.
Läs mer: Yrkesutbildning
Yrkesutbildningfinska _ engelska
Yrkesinriktad utbildningfinska
Gymnasium
I Grankulla finns två gymnasier, ett finskspråkigt och ett svenskspråkigt.
I Esbo finns ett vuxengymnasium där vuxna kan avlägga gymnasiet och studentexamen.
Läs mer: Gymnasium
Grundläggande utbildning och gymnasiumfinska _ svenska _ engelska
linkkiEsbo stad:
Vuxengymnasietfinska
Högskoleutbildning
I anslutning till folkhögskolan Työväen Akatemia i Grankulla finns en enhet för Humanistiska Yrkeshögskolan, där du kan avlägga yrkeshögskoleexamen för kulturproducenter.
Vid yrkeshögskolorna och universiteten i Esbo och Helsingfors kan du studera inom många områden.
Mer information om högskolorna i Esbo och Helsingfors hittar du på städernas webbplatser.
Läs mer: Högskoleutbildning
linkkiHumanistiska yrkeshögskolan:
Information om Humanistiska yrkeshögskolanfinska _ engelska
linkkiEsbo stad:
Högskolorfinska _ engelska
Högskolorfinska
Andra studiemöjligheter
Vid Grankulla medborgarinstitut kan du studera till exempel språk, handarbete och matlagning eller delta i ledd motion.
Medborgarinstitutetfinska _ svenska _ engelska
Vid Grankulla konstskola kan barn och unga studera bildkonst och vid Grankulla musikinstitut kan barn och vuxna studera musik.
Information om Konstskolanfinska _ svenska
Information om Musikinstitutetfinska _ svenska
I Grankulla ligger Finska Bibelinstitutet.
Vid institutet kan du avlägga enskilda kurser eller studera på någon av institutets studielinjer.
Studierna på studielinjerna pågår i 1–2 år.
Vid bibelinstitutet finns även en studielinje som är särskilt avsedd för invandrare.
Kristliga folkhögskolanfinska _ engelska
Folkhögskolan Työväen Akatemia tillhandahåller undervisning inom många akademiska discipliner samt träning för dem som vill läsa på universitet.
Information om Työväen Akatemiafinska _ engelska
Läs mer: Andra studiemöjligheter
Dagvård
Förskoleundervisning
Grundläggande utbildning
Yrkesutbildning
Gymnasium
Högskoleutbildning
Andra studiemöjligheter
Dagvård
I Grankulla finns stadens egna daghem, privata daghem och privata familjedagvårdare.
Dagvård fås på finska och på svenska.
I Grankulla finns också ett engelskspråkigt daghem.
Ansök om dagvårdsplats för ditt barn minst fyra månader innan barnet ska börja i dagvården.
Om du ansöker om dagvårdplats för första gången ska du använda den elektroniska ansökan.
Du kan också hämta ansökningsblanketten på daghemmet eller vid informationen i stadshuset.
Lämna in ansökan till daghemmet eller stadshuset.
Familjer som bor i Grankulla kan också söka dagvårdsplats till sitt barn i Esbo, Helsingfors eller Vanda.
Du ska ändå lämna in din ansökan i Grankulla.
Mer information finns på tjänsten HelsingforsRegionen.fi.
Läs mer: Dagvård
Dagvård och förskoleundervisningfinska _ svenska _ engelska
Ansökan om dagvårdsplatsfinska _ svenska
Engelsk-finskspråkigt daghemfinska _ engelska
Dagvårdens samanvändningsområdefinska _ svenska _ engelska
Förskoleundervisning
I Grankulla anordnas förskoleundervisningen i daghemmen.
Förskoleundervisningen börjar i augusti och ansökningstiden är i januari.
Läs mer: Förskoleundervisning
Information om förskoleundervisningenfinska _ svenska _ engelska
Grundläggande utbildning
I Grankulla finns både en finsk- och en svenskspråkig grundskola. Anmälan till grundskolan ska ske i början av året.
Om du har frågor om den grundläggande utbildningen kan du kontakta skolbyrån.
Skolbyrån
Grankulla stadshus
Grankullavägen 10
02700 Grankulla
Tfn (09) 50 561 (växel)
Grundläggande utbildning
Grundläggande utbildning och gymnasiumfinska _ svenska _ engelska
Internationella skolor i huvudstadsregionenfinska
linkkiExpatFinland.fi:
Internationella skolor i huvudstadsregionenengelska
Yrkesutbildning
De närmaste yrkesläroanstalterna finns i Esbo och Helsingfors.
Läs mer: Yrkesutbildning
Yrkesutbildningfinska _ engelska
Yrkesinriktad utbildningfinska
Gymnasium
I Grankulla finns två gymnasier, ett finskspråkigt och ett svenskspråkigt.
I Esbo finns ett vuxengymnasium där vuxna kan avlägga gymnasiet och studentexamen.
Läs mer: Gymnasium
Grundläggande utbildning och gymnasiumfinska _ svenska _ engelska
linkkiEsbo stad:
Vuxengymnasietfinska
Högskoleutbildning
I anslutning till folkhögskolan Työväen Akatemia i Grankulla finns en enhet för Humanistiska Yrkeshögskolan, där du kan avlägga yrkeshögskoleexamen för kulturproducenter.
Vid yrkeshögskolorna och universiteten i Esbo och Helsingfors kan du studera inom många områden.
Mer information om högskolorna i Esbo och Helsingfors hittar du på städernas webbplatser.
Läs mer: Högskoleutbildning
linkkiHumanistiska yrkeshögskolan:
Information om Humanistiska yrkeshögskolanfinska _ engelska
linkkiEsbo stad:
Högskolorfinska _ engelska
Högskolorfinska
Andra studiemöjligheter
Vid Grankulla medborgarinstitut kan du studera till exempel språk, handarbete och matlagning eller delta i ledd motion.
Medborgarinstitutetfinska _ svenska _ engelska
Vid Grankulla konstskola kan barn och unga studera bildkonst och vid Grankulla musikinstitut kan barn och vuxna studera musik.
Information om Konstskolanfinska _ svenska
Information om Musikinstitutetfinska _ svenska
I Grankulla ligger Finska Bibelinstitutet.
Vid institutet kan du avlägga enskilda kurser eller studera på någon av institutets studielinjer.
Studierna på studielinjerna pågår i 1–2 år.
Vid bibelinstitutet finns även en studielinje som är särskilt avsedd för invandrare.
Kristliga folkhögskolanfinska _ engelska
Folkhögskolan Työväen Akatemia tillhandahåller undervisning inom många akademiska discipliner samt träning för dem som vill läsa på universitet.
Information om Työväen Akatemiafinska _ engelska
Läs mer: Andra studiemöjligheter
Hyresbostad
Ägarbostad
Stöd- och serviceboende
Avfallshantering i bostaden
Hyresbostad
Hyresbostäderna är dyra i huvudstadsregionen.
Stadens hyresbostäder är förmånligare än bostäder som hyrs ut av företag och privatpersoner.
Privata hyresbostäder
Du hittar bostäder som hyrs ut av företag och privatpersoner via bostadssidor på internet.
Sökning av hyresbostäderfinska
Sökning av hyresbostäderfinska _ engelska
Stadens hyresbostäder
Om du vill söka en av stadens hyresbostäder ska du fylla i en ansökningsblankett för hyresbostäder.
Blanketten får du antingen vid informationen på Grankulla stadshus, på socialbyrån eller på Grankulla stads webbplats.
På stadens webbplats hittar du också anvisningar om hur du söker hyresbostad.
Skicka din ansökan till adressen:
PB 52
02701 Grankulla
Stadens hyresbostäderfinska _ svenska _ engelska
Om du är studerande kan du få en hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS.
linkkiHOAS:
Hyresbostäder för studerandefinska _ svenska _ engelska
Läs mer: Hyresbostad
Ägarbostad
På internet finns många annonser om bostäder som är till salu.
Bostäderna i Grankulla är tämligen dyra.
Information om köp av bostad hittar du på InfoFinlands sida Ägarbostad.
Om du blir bostadslös på grund av en kris eller en olycka, ska du kontakta socialbyrån.
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta ett skyddshem.
Steniusvägen 20
Du kan ringa skyddshemmet dygnet runt, telefonnumret är 09 4777 180.
Du behöver inte uppge ditt namn när du ringer.
Om du är ung och har problem hemma, kan du kontakta Finlands Röda Kors De ungas skyddshus.
Det närmaste skyddshuset finns i Esbo.
De ungas skyddshus
Tfn 09 819 55360
Hjälp till offer för familjevåldfinska
linkkiFörbundet för mödra- och skyddshem:
Information om skyddshem och mödrahemfinska
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Stöd- och serviceboende
Personer som har svårt att klara av de dagliga sysslorna utan hjälp, till exempel äldre eller personer med funktionsnedsättning, kan få ta del av hemvårdens stödtjänster.
En person som inte kan bo på egen hand kan bo på en anstalt.
På Grankulla socialbyrå kan du fråga mer om hemvårdens stödtjänster och boende på anstalt.
Grankulla socialbyrå
Köpcentret Grani
Grankullavägen 7 02700 Grankulla
Tfn 09 505 61
Läs mer: Stöd- och serviceboende
Information om hemvårdens stödtjänsterfinska _ svenska
Information om boende på anstaltfinska _ svenska
Avfallshantering och återvinning
På InfoFinlands sida Avfallshantering och återvinning hittar du information om sopsortering.
linkkiHelsingforsregionens miljötjänster:
Sopsorteringsanvisningarfinska _ svenska _ engelska
Avfallsinsamlingsstationerfinska
Hyresbostad
Ägarbostad
Stöd- och serviceboende
Avfallshantering i bostaden
Hyresbostad
Hyresbostäderna är dyra i huvudstadsregionen.
Stadens hyresbostäder är förmånligare än bostäder som hyrs ut av företag och privatpersoner.
Privata hyresbostäder
Du hittar bostäder som hyrs ut av företag och privatpersoner via bostadssidor på internet.
Sökning av hyresbostäderfinska
Sökning av hyresbostäderfinska _ engelska
Stadens hyresbostäder
Om du vill söka en av stadens hyresbostäder ska du fylla i en ansökningsblankett för hyresbostäder.
Blanketten får du antingen vid informationen på Grankulla stadshus, på socialbyrån eller på Grankulla stads webbplats.
På stadens webbplats hittar du också anvisningar om hur du söker hyresbostad.
Skicka din ansökan till adressen:
PB 52
02701 Grankulla
Stadens hyresbostäderfinska _ svenska _ engelska
Om du är studerande kan du få en hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS.
linkkiHOAS:
Hyresbostäder för studerandefinska _ svenska _ engelska
Läs mer: Hyresbostad
Ägarbostad
På internet finns många annonser om bostäder som är till salu.
Bostäderna i Grankulla är tämligen dyra.
Information om köp av bostad hittar du på InfoFinlands sida Ägarbostad.
Om du blir bostadslös på grund av en kris eller en olycka, ska du kontakta socialbyrån.
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta ett skyddshem.
Steniusvägen 20
Du kan ringa skyddshemmet dygnet runt, telefonnumret är 09 4777 180.
Du behöver inte uppge ditt namn när du ringer.
Om du är ung och har problem hemma, kan du kontakta Finlands Röda Kors De ungas skyddshus.
Det närmaste skyddshuset finns i Esbo.
De ungas skyddshus
Tfn 09 819 55360
Hjälp till offer för familjevåldfinska
linkkiFörbundet för mödra- och skyddshem:
Information om skyddshem och mödrahemfinska
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Stöd- och serviceboende
Personer som har svårt att klara av de dagliga sysslorna utan hjälp, till exempel äldre eller personer med funktionsnedsättning, kan få ta del av hemvårdens stödtjänster.
En person som inte kan bo på egen hand kan bo på en anstalt.
På Grankulla socialbyrå kan du fråga mer om hemvårdens stödtjänster och boende på anstalt.
Grankulla socialbyrå
Köpcentret Grani
Grankullavägen 7 02700 Grankulla
Tfn 09 505 61
Läs mer: Stöd- och serviceboende
Information om hemvårdens stödtjänsterfinska _ svenska
Information om boende på anstaltfinska _ svenska
Avfallshantering och återvinning
På InfoFinlands sida Avfallshantering och återvinning hittar du information om sopsortering.
linkkiHelsingforsregionens miljötjänster:
Sopsorteringsanvisningarfinska _ svenska _ engelska
Avfallsinsamlingsstationerfinska
Hyresbostad
Ägarbostad
Stöd- och serviceboende
Avfallshantering i bostaden
Hyresbostad
Hyresbostäderna är dyra i huvudstadsregionen.
Stadens hyresbostäder är förmånligare än bostäder som hyrs ut av företag och privatpersoner.
Privata hyresbostäder
Du hittar bostäder som hyrs ut av företag och privatpersoner via bostadssidor på internet.
Sökning av hyresbostäderfinska
Sökning av hyresbostäderfinska _ engelska
Stadens hyresbostäder
Om du vill söka en av stadens hyresbostäder ska du fylla i en ansökningsblankett för hyresbostäder.
Blanketten får du antingen vid informationen på Grankulla stadshus, på socialbyrån eller på Grankulla stads webbplats.
På stadens webbplats hittar du också anvisningar om hur du söker hyresbostad.
Skicka din ansökan till adressen:
PB 52
02701 Grankulla
Stadens hyresbostäderfinska _ svenska _ engelska
Om du är studerande kan du få en hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS.
linkkiHOAS:
Hyresbostäder för studerandefinska _ svenska _ engelska
Läs mer: Hyresbostad
Ägarbostad
På internet finns många annonser om bostäder som är till salu.
Bostäderna i Grankulla är tämligen dyra.
Information om köp av bostad hittar du på InfoFinlands sida Ägarbostad.
Om du blir bostadslös på grund av en kris eller en olycka, ska du kontakta socialbyrån.
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta ett skyddshem.
Steniusvägen 20
Du kan ringa skyddshemmet dygnet runt, telefonnumret är 09 4777 180.
Du behöver inte uppge ditt namn när du ringer.
Om du är ung och har problem hemma, kan du kontakta Finlands Röda Kors De ungas skyddshus.
Det närmaste skyddshuset finns i Esbo.
De ungas skyddshus
Tfn 09 819 55360
Hjälp till offer för familjevåldfinska
linkkiFörbundet för mödra- och skyddshem:
Information om skyddshem och mödrahemfinska
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Stöd- och serviceboende
Personer som har svårt att klara av de dagliga sysslorna utan hjälp, till exempel äldre eller personer med funktionsnedsättning, kan få ta del av hemvårdens stödtjänster.
En person som inte kan bo på egen hand kan bo på en anstalt.
På Grankulla socialbyrå kan du fråga mer om hemvårdens stödtjänster och boende på anstalt.
Grankulla socialbyrå
Köpcentret Grani
Grankullavägen 7 02700 Grankulla
Tfn 09 505 61
Läs mer: Stöd- och serviceboende
Information om hemvårdens stödtjänsterfinska _ svenska
Information om boende på anstaltfinska _ svenska
Avfallshantering och återvinning
På InfoFinlands sida Avfallshantering och återvinning hittar du information om sopsortering.
linkkiHelsingforsregionens miljötjänster:
Sopsorteringsanvisningarfinska _ svenska _ engelska
Avfallsinsamlingsstationerfinska
Språkkurser
Med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors, Vanda, Esbo eller Grankulla.
I tjänsten finns också information om kurser i svenska.
Kurser i finska och svenska språketfinska _ engelska _ ryska
I Grankulla ordnas kurser i finska och svenska av Grankulla medborgarinstitut.
Du kan anmäla dig till medborgarinstitutets kurser per telefon eller via internet.
Medborgarinstitutetfinska _ svenska _ engelska
Läs mer: Studier i finska och svenska
Svenska språket i Finland.
Diskutera på finska
Information om bibliotekens språkkaféer och andra finska samtalsgrupper hittar du på InfoFinlands sidor Finska och svenska språket i Esbo och Finska och svenska språket i Helsingfors.
Allmän språkexamen
Du kan avlägga allmän språkexamen i finska eller svenska till exempel i Esbo och Helsingfors.
På Utbildningsstyrelsens webbplats finns en sökmotor med vilken du kan kontrollera var och när du kan avlägga examen.
Läs mer: Officiellt intyg på språkkunskaper.
linkkiUtbildningsstyrelsen:
Allmänna språkexaminafinska _ svenska _ engelska
Språkkurser
Med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors, Vanda, Esbo eller Grankulla.
I tjänsten finns också information om kurser i svenska.
Kurser i finska och svenska språketfinska _ engelska _ ryska
I Grankulla ordnas kurser i finska och svenska av Grankulla medborgarinstitut.
Du kan anmäla dig till medborgarinstitutets kurser per telefon eller via internet.
Medborgarinstitutetfinska _ svenska _ engelska
Läs mer: Studier i finska och svenska
Svenska språket i Finland.
Diskutera på finska
Information om bibliotekens språkkaféer och andra finska samtalsgrupper hittar du på InfoFinlands sidor Finska och svenska språket i Esbo och Finska och svenska språket i Helsingfors.
Allmän språkexamen
Du kan avlägga allmän språkexamen i finska eller svenska till exempel i Esbo och Helsingfors.
På Utbildningsstyrelsens webbplats finns en sökmotor med vilken du kan kontrollera var och när du kan avlägga examen.
Läs mer: Officiellt intyg på språkkunskaper.
linkkiUtbildningsstyrelsen:
Allmänna språkexaminafinska _ svenska _ engelska
Språkkurser
Med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors, Vanda, Esbo eller Grankulla.
I tjänsten finns också information om kurser i svenska.
Kurser i finska och svenska språketfinska _ engelska _ ryska
I Grankulla ordnas kurser i finska och svenska av Grankulla medborgarinstitut.
Du kan anmäla dig till medborgarinstitutets kurser per telefon eller via internet.
Medborgarinstitutetfinska _ svenska _ engelska
Läs mer: Studier i finska och svenska
Svenska språket i Finland.
Diskutera på finska
Information om bibliotekens språkkaféer och andra finska samtalsgrupper hittar du på InfoFinlands sidor Finska och svenska språket i Esbo och Finska och svenska språket i Helsingfors.
Allmän språkexamen
Du kan avlägga allmän språkexamen i finska eller svenska till exempel i Esbo och Helsingfors.
På Utbildningsstyrelsens webbplats finns en sökmotor med vilken du kan kontrollera var och när du kan avlägga examen.
Läs mer: Officiellt intyg på språkkunskaper.
linkkiUtbildningsstyrelsen:
Allmänna språkexaminafinska _ svenska _ engelska
Var hittar jag jobb?
Att grunda ett företag
Beskattning
Var hittar jag jobb?
Nylands arbets- och näringsbyrå hjälper invånare i Grankulla att söka jobb.
Den närmaste byrån finns i Esbo.
Nylands arbets- och näringsbyrå, Esbo
Läs mer: Arbete och entreprenörskap i Esbo
Information om arbets- och näringsbyråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös.
Information om jobbsökning i Finland hittar du på InfoFinlands sida Var hittar jag jobb?
Seure erbjuder kortvariga jobb vid Helsingfors, Vanda, Esbo och Grankulla städer.
Jobben finns till exempel på skolor, daghem och sjukhus.
Arbetsplatser i kommunernafinska _ svenska
Lediga jobbfinska _ svenska _ engelska
Arbetslöshetsersättning
Information om att ansöka om arbetslöshetsersättning hittar du på InfoFinlands sida Arbetslöshetsförsäkring.
Att grunda ett företag
På InfoFinlands sida Att grunda ett företag hittar du information om hur man grundar ett företag i Finland.
Bekanta dig med de lokala tjänsterna på sidorna Arbete och entreprenörskap i Esbo och Arbete och entreprenörskap i Helsingfors.
Om du är företagare kan du bli medlem i företagarnas intressebevakningsorganisation Grankulla företagare rf som erbjuder sina medlemmar utbildning, nätverk och rådgivning.
Information för företagarefinska
Beskattning
Huvudstadsregionens skattebyrå ligger på Alexandersgatan 9 i Gloet i Helsingfors.
linkkiSkatteförvaltningen:
Kontaktuppgifter till skattebyråerfinska _ svenska _ engelska
Du kan även besöka servicestället In To Finland i Kampen i Helsingfors för att fråga om beskattningen.
Servicestället betjänar invandrare som kommer till Finland för att arbeta i ärenden som berör beskattning och social trygghet.
Albertsgatan 25
Lär mer Beskattning
Var hittar jag jobb?
Att grunda ett företag
Beskattning
Var hittar jag jobb?
Nylands arbets- och näringsbyrå hjälper invånare i Grankulla att söka jobb.
Den närmaste byrån finns i Esbo.
Nylands arbets- och näringsbyrå, Esbo
Läs mer: Arbete och entreprenörskap i Esbo
Information om arbets- och näringsbyråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös.
Information om jobbsökning i Finland hittar du på InfoFinlands sida Var hittar jag jobb?
Seure erbjuder kortvariga jobb vid Helsingfors, Vanda, Esbo och Grankulla städer.
Jobben finns till exempel på skolor, daghem och sjukhus.
Arbetsplatser i kommunernafinska _ svenska
Lediga jobbfinska _ svenska _ engelska
Arbetslöshetsersättning
Information om att ansöka om arbetslöshetsersättning hittar du på InfoFinlands sida Arbetslöshetsförsäkring.
Att grunda ett företag
På InfoFinlands sida Att grunda ett företag hittar du information om hur man grundar ett företag i Finland.
Bekanta dig med de lokala tjänsterna på sidorna Arbete och entreprenörskap i Esbo och Arbete och entreprenörskap i Helsingfors.
Om du är företagare kan du bli medlem i företagarnas intressebevakningsorganisation Grankulla företagare rf som erbjuder sina medlemmar utbildning, nätverk och rådgivning.
Information för företagarefinska
Beskattning
Huvudstadsregionens skattebyrå ligger på Alexandersgatan 9 i Gloet i Helsingfors.
linkkiSkatteförvaltningen:
Kontaktuppgifter till skattebyråerfinska _ svenska _ engelska
Invandrare kan även sköta ärenden vid servicestället International House Helsinki.
På servicestället hjälper FPA:s och Skatteförvaltningens experter invandrare som kommer till Finland för att arbeta i frågor som rör beskattning och social trygghet.
Lär mer Beskattning
Var hittar jag jobb?
Att grunda ett företag
Beskattning
Var hittar jag jobb?
Nylands arbets- och näringsbyrå hjälper invånare i Grankulla att söka jobb.
Den närmaste byrån finns i Esbo.
Nylands arbets- och näringsbyrå, Esbo
Läs mer: Arbete och entreprenörskap i Esbo
Information om arbets- och näringsbyråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös.
Information om jobbsökning i Finland hittar du på InfoFinlands sida Var hittar jag jobb?
Seure erbjuder kortvariga jobb vid Helsingfors, Vanda, Esbo och Grankulla städer.
Jobben finns till exempel på skolor, daghem och sjukhus.
Arbetsplatser i kommunernafinska _ svenska _ engelska
Lediga jobbfinska _ svenska _ engelska
Arbetslöshetsersättning
Information om att ansöka om arbetslöshetsersättning hittar du på InfoFinlands sida Arbetslöshetsförsäkring.
Att grunda ett företag
På InfoFinlands sida Att grunda ett företag hittar du information om hur man grundar ett företag i Finland.
Bekanta dig med de lokala tjänsterna på sidorna Arbete och entreprenörskap i Esbo och Arbete och entreprenörskap i Helsingfors.
Om du är företagare kan du bli medlem i företagarnas intressebevakningsorganisation Grankulla företagare rf som erbjuder sina medlemmar utbildning, nätverk och rådgivning.
Information för företagarefinska
Beskattning
Huvudstadsregionens skattebyrå ligger på Alexandersgatan 9 i Gloet i Helsingfors.
linkkiSkatteförvaltningen:
Kontaktuppgifter till skattebyråerfinska _ svenska _ engelska
Invandrare kan även sköta ärenden vid servicestället International House Helsinki.
På servicestället hjälper FPA:s och Skatteförvaltningens experter invandrare som kommer till Finland för att arbeta i frågor som rör beskattning och social trygghet.
IHH – serviceställe för dig som flyttar till Finland engelska
Lär mer Beskattning
Rådgivning för och integration av invandrare
Inledande kartläggning och integrationsplan
Behöver du en tolk?
Rådgivning för och integration av invandrare
Om du har frågor om tjänsterna vid Grankulla stad kan du kontakta stadens rådgivningstjänst via e-post på adressen neuvontapalvelu(at)kauniainen.fi.
Du kan skriva på finska, svenska eller engelska.
Helsingfors stads rådgivning för invandrare, Helsingfors-info, betjänar alla invandrare i huvudstadsregionen.
Helsingfors-infofinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
IHH – serviceställe för dig som flyttar till Finland engelska
Inledande kartläggning och integrationsplan
Tillsammans med en anställd vid arbets- och näringsbyrån (TE-byrån) gör du en inledande kartläggning och en integrationsplan i samband med att du registrerar dig som arbetssökande.
linkkiArbets- och näringsministeriet:
Arbets- och näringsbyråerna i Nylandfinska _ svenska
Om du inte är kund hos arbets- och näringsbyrån görs den inledande kartläggningen och integrationsplanen på socialbyrån.
Kontaktuppgifter till socialbyrån:
Köpcentret Grani
Grankullavägen 7
02700 Grankulla
Tfn (09) 50 561
Socialbyrånfinska _ svenska
Behöver du en tolk?
Om du inte kan finska eller svenska kan du anlita en tolk när du sköter ärenden med myndigheter.
Du kan anlita en tolk när som helst om du bokar tolken och betalar kostnaderna själv.
I vissa fall får du en tolk via myndigheten.
Då är tolkningen avgiftsfri för dig.
Läs mer: Behöver du en tolk?
linkkiFinlands översättar- och tolkförbund:
Sök tolk eller översättarefinska _ svenska _ engelska
Rådgivning för och integration av invandrare
Inledande kartläggning och integrationsplan
Behöver du en tolk?
Rådgivning för och integration av invandrare
Om du har frågor om tjänsterna vid Grankulla stad kan du kontakta stadens rådgivningstjänst via e-post på adressen neuvontapalvelu(at)kauniainen.fi.
Du kan skriva på finska, svenska eller engelska.
Helsingfors stads rådgivning för invandrare, Helsingfors-info, betjänar alla invandrare i huvudstadsregionen.
Helsingfors-infofinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
IHH – serviceställe för dig som flyttar till Finland engelska
Inledande kartläggning och integrationsplan
Tillsammans med en anställd vid arbets- och näringsbyrån (TE-byrån) gör du en inledande kartläggning och en integrationsplan i samband med att du registrerar dig som arbetssökande.
linkkiArbets- och näringsministeriet:
Arbets- och näringsbyråerna i Nylandfinska _ svenska
Om du inte är kund hos arbets- och näringsbyrån görs den inledande kartläggningen och integrationsplanen på socialbyrån.
Kontaktuppgifter till socialbyrån:
Köpcentret Grani
Grankullavägen 7
02700 Grankulla
Tfn (09) 50 561
Socialbyrånfinska _ svenska
Behöver du en tolk?
Om du inte kan finska eller svenska kan du anlita en tolk när du sköter ärenden med myndigheter.
Du kan anlita en tolk när som helst om du bokar tolken och betalar kostnaderna själv.
I vissa fall får du en tolk via myndigheten.
Då är tolkningen avgiftsfri för dig.
Läs mer: Behöver du en tolk?
linkkiFinlands översättar- och tolkförbund:
Sök tolk eller översättarefinska _ svenska _ engelska
Rådgivning för och integration av invandrare
Inledande kartläggning och integrationsplan
Behöver du en tolk?
Rådgivning för och integration av invandrare
Om du har frågor om tjänsterna vid Grankulla stad kan du kontakta stadens rådgivningstjänst via e-post på adressen neuvontapalvelu(at)kauniainen.fi.
Du kan skriva på finska, svenska eller engelska.
Helsingfors stads rådgivning för invandrare, Helsingfors-info, betjänar alla invandrare i huvudstadsregionen.
Helsingfors-infofinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
IHH – serviceställe för dig som flyttar till Finland engelska
Inledande kartläggning och integrationsplan
Tillsammans med en anställd vid arbets- och näringsbyrån (TE-byrån) gör du en inledande kartläggning och en integrationsplan i samband med att du registrerar dig som arbetssökande.
linkkiArbets- och näringsministeriet:
Arbets- och näringsbyråerna i Nylandfinska _ svenska
Om du inte är kund hos arbets- och näringsbyrån görs den inledande kartläggningen och integrationsplanen på socialbyrån.
Kontaktuppgifter till socialbyrån:
Köpcentret Grani
Grankullavägen 7
02700 Grankulla
Tfn (09) 50 561
Socialbyrånfinska _ svenska
Behöver du en tolk?
Om du inte kan finska eller svenska kan du anlita en tolk när du sköter ärenden med myndigheter.
Du kan anlita en tolk när som helst om du bokar tolken och betalar kostnaderna själv.
I vissa fall får du en tolk via myndigheten.
Då är tolkningen avgiftsfri för dig.
Läs mer: Behöver du en tolk?
linkkiFinlands översättar- och tolkförbund:
Sök tolk eller översättarefinska _ svenska _ engelska
Tillståndsärenden
På Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU-medborgarens uppehållsrätt.
Boka en tid i förväg.
Adress:
Göksgränd 3A
Elektronisk tidsbokningfinska _ svenska _ engelska
Du kan också ansöka om många slags uppehållstillstånd och EU-registrering på internet i tjänsten Enter Finland.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Läs mer: Flytta till Finland.
Registrering som invånare
Om du flyttar ditt stadigvarande boende till Grankulla, ska du registrera dig som invånare i kommunen.
Du kan registrera dig vid Helsingfors enhet vid magistraten i Nyland.
Helsingfors enhet
Albertsgatan 25
Tfn 029 55 39391
När du går till magistraten ska du ta med dig
legitimation (till exempel pass)
uppehållstillstånd och uppehållskort (om du behöver uppehållstillstånd i Finland)
registreringsintyget över uppehållsrätten (om du är EU-medborgare)
äktenskapsintyg
dina barns födelseattester.
Observera att utländska handlingar ska vara legaliserade samt översatta till finska eller svenska.
Läs mer: Registrering som invånare
Hemkommun i Finland
Registrering av utlänningarfinska _ svenska _ engelska
IHH – serviceställe för dig som flyttar till Finland engelska
Tillståndsärenden
På Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU-medborgarens uppehållsrätt.
Boka en tid i förväg.
Adress:
Göksgränd 3A
Elektronisk tidsbokningfinska _ svenska _ engelska
Du kan också ansöka om många slags uppehållstillstånd och EU-registrering på internet i tjänsten Enter Finland.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Läs mer: Flytta till Finland.
Registrering som invånare
Om du flyttar ditt stadigvarande boende till Grankulla, ska du registrera dig som invånare i kommunen.
Du kan registrera dig vid Helsingfors enhet vid magistraten i Nyland.
Helsingfors enhet
Tfn 029 55 39391
När du går till magistraten ska du ta med dig
legitimation (till exempel pass)
uppehållstillstånd och uppehållskort (om du behöver uppehållstillstånd i Finland)
registreringsintyget över uppehållsrätten (om du är EU-medborgare)
äktenskapsintyg
dina barns födelseattester.
Observera att utländska handlingar ska vara legaliserade samt översatta till finska eller svenska.
Läs mer: Registrering som invånare
Hemkommun i Finland
Registrering av utlänningarfinska _ svenska _ engelska
IHH – serviceställe för dig som flyttar till Finland engelska
Tillståndsärenden
På Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU-medborgarens uppehållsrätt.
Boka en tid i förväg.
Adress:
Göksgränd 3A
Elektronisk tidsbokningfinska _ svenska _ engelska
Du kan också ansöka om många slags uppehållstillstånd och EU-registrering på internet i tjänsten Enter Finland.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Läs mer: Flytta till Finland.
Registrering som invånare
Om du flyttar ditt stadigvarande boende till Grankulla, ska du registrera dig som invånare i kommunen.
Du kan registrera dig vid Helsingfors enhet vid magistraten i Nyland.
Helsingfors enhet
Tfn 029 55 39391
När du går till magistraten ska du ta med dig
legitimation (till exempel pass)
uppehållstillstånd och uppehållskort (om du behöver uppehållstillstånd i Finland)
registreringsintyget över uppehållsrätten (om du är EU-medborgare)
äktenskapsintyg
dina barns födelseattester.
Observera att utländska handlingar ska vara legaliserade samt översatta till finska eller svenska.
Läs mer: Registrering som invånare
Hemkommun i Finland
Registrering av utlänningarfinska _ svenska _ engelska
IHH – serviceställe för dig som flyttar till Finland engelska
Trafik
Beslutsfattande och påverkan
Religion
Grundläggande information
Historia
Trafik
Kollektivtrafiken
Vanda och hela huvudstadsregionen har goda kollektivtrafikförbindelser.
Längs stambanan och Mårtensdals bana finns flera tågstationer.
I staden finns flera busslinjer.
Vanda tillhör samkommunen Helsingforsregionens trafik (HRT) (Helsingin seudun liikenne -kuntayhtymä (HSL)), som ordnar kollektivtrafiken i huvudstadsregionen.
Mer information hittar du på HRT:s webbplats.
Du kan söka information om rutterna i Reseplaneraren (Reittiopas).
Tjänsten ger dig förslag på olika kollektivtrafikförbindelser från ett ställe till ett annat.
I kollektivtrafiken kan du betala med kontanter eller resekort.
I närtågen måste du köpa biljetten i förväg.
Du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat.
Reseplanerarefinska _ svenska _ engelska _ ryska
Resekort
Med ett resekort (matkakortti) reser du förmånligare än med kontanter.
Resekortet gäller i lokaltrafikens bussar, närtågen, metron, spårvagnarna och Sveaborgsfärjorna.
Det finns två slags resekort.
Det är det billigaste sättet att resa.
Ett innehavarkort (haltijakohtainen kortti) kan användas av flera personer.
Innan du skaffar dig ett personligt kort ska du registrera dig som invånare i någon av kommunerna inom HRT-området.
Du kan köpa resekort vid HRT:s försäljningsställen (myyntipiste) eller serviceställen (palvelupiste).
De finns runtom i huvudstadsregionen.
Personligt resekort kan du köpa vid serviceställena.
Ta med dig identitetsbevis om du ska köpa personligt resekort.
Om du har finska nätbankskoder kan du även köpa personligt resekort på HRT:s webbplats.
Du kan resa med resekortet när du laddar kortet med period (kausi) eller värde (arvo).
En period betyder tid: till exempel en månad.
Värde betyder pengar.
Om du använder kollektivtrafiken ofta tjänar du på att ladda kortet med period.
Du kan ladda resekortet på vilket serviceställe för resekort (matkakortin latauspiste) som helst.
Du hittar mer information på HRT:s webbplats.
Ansökan om försäljningsplatserfinska _ svenska _ engelska
Information och råd till resenärerfinska _ svenska _ engelska
Biljetter och priserfinska _ svenska _ engelska
Att gå och cykla
Om du vill gå eller cykla i Vanda kan du söka en lämplig rutt i reseplaneraren för cykling och gång.
En cykelkarta i pappersformat för Vanda kan du hämta i Vandainfo.
Cykelkartorna är kostnadsfria.
linkkiVanda stad:
Vandainfofinska _ svenska _ engelska
Bil och flyg
Helsingfors-Vanda internationella flygplats ligger i Vanda.
Flygplatsen har goda trafikförbindelser till exempel med bil, buss och tåg.
Du kan parkera bilen på många järnvägsstationer och fortsätta färden med kollektivtrafiken.
Tidtabellerna för bussar och tåg hittar du enkelt i reseplaneraren.
Läs mer: Trafik.
Flygplatsenfinska _ svenska _ engelska _ ryska _ kinesiska
Beslutsfattande och påverkan
I Vanda beslutas ärenden av stadsfullmäktige (kaupunginvaltuusto).
I stadsfullmäktige sitter 67 ledamöter som representerar olika politiska grupper.
Fullmäktige väljs var fjärde år genom kommunalval (kunnallisvaalit).
Invånarna i Vanda kan påverka beslutsfattandet och beredning av ärenden på många olika sätt.
På Vandakanalen kan du följa fullmäktiges sammanträden och få mer information om beslutsfattandet.
I Vanda finns en delegation för mångkulturella frågor (monikulttuurisuusasiain neuvottelukunta) som lägger fram propositioner i ärenden som rör invandrare.
Läs mer på Vanda stads webbplats.
I Vanda finns många politiska föreningar, invandrarföreningar och andra föreningar via vilka du också kan påverka beslutsfattandet.
Mer information om föreningarna hittar du på sidan Vantaalla.info.
linkkiVanda stad:
Beslutsfattandefinska _ svenska _ engelska
linkkiVanda stad:
Delta och påverkafinska
Stadsfullmäktiges sammanträden på Internetfinska
linkkiVanda stad:
Delegationen för mångkulturella frågorfinska
Religion
Många religiösa samfund är verksamma i Vanda och Helsingfors.
Via tjänsten Uskonnot Suomessa kan du söka information efter det religiösa samfundet och orten.
Den evangelisk-lutherska kyrkan har sex finskspråkiga församlingar och en svenskspråkig församling i Vanda.
Läs mer på Vanda kyrkliga samfällighets webbplats.
I Dickursby finns en ortodox kyrka.
Mer information om verksamheten vid den ortodoxa kyrkan i Vanda hittar du på Helsingfors ortodoxa församlings webbplats.
Läs mer: Kulturer och religioner i Finland.
linkkiVanda kyrkliga samfällighet:
Evangelisk-lutherska församlingarfinska
linkkiHelsingfors ortodoxa församling:
Ortodoxa församlingenfinska _ ryska
Religiösa samfundfinska _ engelska
Grundläggande information
Vanda är en av de fyra kommunerna i huvudstadsregionen.
Den ligger intill Esbo och Helsingfors.
Vanda centrum ligger i Dickursby.
Därtill finns det andra stora tätorter i Vanda, till exempel Korso, Björkby-Havukoski, Myrbacka, Mårtensdal, Håkansböle, Västerkulla och Backas.
Vanda har drygt 205 000 invånare.
Av dem är cirka 2,8 procent svenskspråkiga och 11 procent har något annat modersmål än finska eller svenska.
Arealen är cirka 240 km2, varav cirka 2 km2 består av vatten.
linkkiVanda stad:
Grundläggande informationfinska _ svenska _ engelska
Historia
Vanda område har varit bebott länge.
Man har hittat upp till 7 000 år gamla lämningar efter bosättning.
Nuvarande Vanda har uppstått på ett område som förr var Helsingfors socken.
Helsingfors sockens historia sträcker sig ända till 1300-talet.
Helsingfors socken blev först Helsingfors landskommun, sedan Vanda köping år 1972 och till slut Vanda stad år 1974.
Läget som granne till huvudstaden Helsingfors har varit viktigt för Vanda.
Viktiga vägar, såsom vägen från Åbo via Helsingfors till Viborg och senare järnvägen norrut från Helsingfors, har gått genom Vanda.
Längs med vägarna och järnvägen har det utvecklats industrier och bostadsområden.
Vanda är än idag en viktig trafikknutpunkt.
Till exempel ligger Helsingfors-Vanda flygplats i Vanda.
linkkiVanda stad:
Information om Vandafinska
linkkiVanda stad:
Stadsmuseetfinska _ svenska _ engelska
Trafik
Beslutsfattande och påverkan
Religion
Grundläggande information
Historia
Trafik
Kollektivtrafiken
Vanda och hela huvudstadsregionen har goda kollektivtrafikförbindelser.
Längs stambanan och Mårtensdals bana finns flera tågstationer.
I staden finns flera busslinjer.
Vanda tillhör samkommunen Helsingforsregionens trafik (HRT) (Helsingin seudun liikenne -kuntayhtymä (HSL)), som ordnar kollektivtrafiken i huvudstadsregionen.
Mer information hittar du på HRT:s webbplats.
Du kan söka information om rutterna i Reseplaneraren (Reittiopas).
Tjänsten ger dig förslag på olika kollektivtrafikförbindelser från ett ställe till ett annat.
I kollektivtrafiken kan du betala med kontanter eller resekort.
I närtågen måste du köpa biljetten i förväg.
Du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat.
Reseplanerarefinska _ svenska _ engelska _ ryska
Resekort
Med ett resekort (matkakortti) reser du förmånligare än med kontanter.
Resekortet gäller i lokaltrafikens bussar, närtågen, metron, spårvagnarna och Sveaborgsfärjorna.
Det finns två slags resekort.
Det är det billigaste sättet att resa.
Ett innehavarkort (haltijakohtainen kortti) kan användas av flera personer.
Innan du skaffar dig ett personligt kort ska du registrera dig som invånare i någon av kommunerna inom HRT-området.
Du kan köpa resekort vid HRT:s försäljningsställen (myyntipiste) eller serviceställen (palvelupiste).
De finns runtom i huvudstadsregionen.
Personligt resekort kan du köpa vid serviceställena.
Ta med dig identitetsbevis om du ska köpa personligt resekort.
Om du har finska nätbankskoder kan du även köpa personligt resekort på HRT:s webbplats.
Du kan resa med resekortet när du laddar kortet med period (kausi) eller värde (arvo).
En period betyder tid: till exempel en månad.
Värde betyder pengar.
Om du använder kollektivtrafiken ofta tjänar du på att ladda kortet med period.
Du kan ladda resekortet på vilket serviceställe för resekort (matkakortin latauspiste) som helst.
Du hittar mer information på HRT:s webbplats.
Ansökan om försäljningsplatserfinska _ svenska _ engelska
Information och råd till resenärerfinska _ svenska _ engelska
Biljetter och priserfinska _ svenska _ engelska
Att gå och cykla
Om du vill gå eller cykla i Vanda kan du söka en lämplig rutt i reseplaneraren för cykling och gång.
En cykelkarta i pappersformat för Vanda kan du hämta i Vandainfo.
Cykelkartorna är kostnadsfria.
linkkiVanda stad:
Vandainfofinska _ svenska _ engelska
Bil och flyg
Helsingfors-Vanda internationella flygplats ligger i Vanda.
Flygplatsen har goda trafikförbindelser till exempel med bil, buss och tåg.
Du kan parkera bilen på många järnvägsstationer och fortsätta färden med kollektivtrafiken.
Tidtabellerna för bussar och tåg hittar du enkelt i reseplaneraren.
Läs mer: Trafik.
Flygplatsenfinska _ svenska _ engelska _ ryska _ kinesiska
Beslutsfattande och påverkan
I Vanda beslutas ärenden av stadsfullmäktige (kaupunginvaltuusto).
I stadsfullmäktige sitter 67 ledamöter som representerar olika politiska grupper.
Fullmäktige väljs var fjärde år genom kommunalval (kunnallisvaalit).
Invånarna i Vanda kan påverka beslutsfattandet och beredning av ärenden på många olika sätt.
På Vandakanalen kan du följa fullmäktiges sammanträden och få mer information om beslutsfattandet.
I Vanda finns en delegation för mångkulturella frågor (monikulttuurisuusasiain neuvottelukunta) som lägger fram propositioner i ärenden som rör invandrare.
Läs mer på Vanda stads webbplats.
I Vanda finns många politiska föreningar, invandrarföreningar och andra föreningar via vilka du också kan påverka beslutsfattandet.
Mer information om föreningarna hittar du på sidan Vantaalla.info.
linkkiVanda stad:
Beslutsfattandefinska _ svenska _ engelska
linkkiVanda stad:
Delta och påverkafinska
Stadsfullmäktiges sammanträden på Internetfinska
linkkiVanda stad:
Delegationen för mångkulturella frågorfinska
Religion
Många religiösa samfund är verksamma i Vanda och Helsingfors.
Via tjänsten Uskonnot Suomessa kan du söka information efter det religiösa samfundet och orten.
Den evangelisk-lutherska kyrkan har sex finskspråkiga församlingar och en svenskspråkig församling i Vanda.
Läs mer på Vanda kyrkliga samfällighets webbplats.
I Dickursby finns en ortodox kyrka.
Mer information om verksamheten vid den ortodoxa kyrkan i Vanda hittar du på Helsingfors ortodoxa församlings webbplats.
Läs mer: Kulturer och religioner i Finland.
linkkiVanda kyrkliga samfällighet:
Evangelisk-lutherska församlingarfinska
linkkiHelsingfors ortodoxa församling:
Ortodoxa församlingenfinska _ ryska
Religiösa samfundfinska _ engelska
Grundläggande information
Vanda är en av de fyra kommunerna i huvudstadsregionen.
Den ligger intill Esbo och Helsingfors.
Vanda centrum ligger i Dickursby.
Därtill finns det andra stora tätorter i Vanda, till exempel Korso, Björkby-Havukoski, Myrbacka, Mårtensdal, Håkansböle, Västerkulla och Backas.
Vanda har drygt 205 000 invånare.
Av dem är cirka 2,8 procent svenskspråkiga och 11 procent har något annat modersmål än finska eller svenska.
Arealen är cirka 240 km2, varav cirka 2 km2 består av vatten.
linkkiVanda stad:
Grundläggande informationfinska _ svenska _ engelska
Historia
Vanda område har varit bebott länge.
Man har hittat upp till 7 000 år gamla lämningar efter bosättning.
Nuvarande Vanda har uppstått på ett område som förr var Helsingfors socken.
Helsingfors sockens historia sträcker sig ända till 1300-talet.
Helsingfors socken blev först Helsingfors landskommun, sedan Vanda köping år 1972 och till slut Vanda stad år 1974.
Läget som granne till huvudstaden Helsingfors har varit viktigt för Vanda.
Viktiga vägar, såsom vägen från Åbo via Helsingfors till Viborg och senare järnvägen norrut från Helsingfors, har gått genom Vanda.
Längs med vägarna och järnvägen har det utvecklats industrier och bostadsområden.
Vanda är än idag en viktig trafikknutpunkt.
Till exempel ligger Helsingfors-Vanda flygplats i Vanda.
linkkiVanda stad:
Information om Vandafinska
linkkiVanda stad:
Stadsmuseetfinska _ svenska _ engelska
Trafik
Beslutsfattande och påverkan
Religion
Grundläggande information
Historia
Trafik
Kollektivtrafiken
Vanda och hela huvudstadsregionen har goda kollektivtrafikförbindelser.
Längs stambanan och Mårtensdals bana finns flera tågstationer.
I staden finns flera busslinjer.
Vanda tillhör samkommunen Helsingforsregionens trafik (HRT) (Helsingin seudun liikenne -kuntayhtymä (HSL)), som ordnar kollektivtrafiken i huvudstadsregionen.
Mer information hittar du på HRT:s webbplats.
Du kan söka information om rutterna i Reseplaneraren (Reittiopas).
Tjänsten ger dig förslag på olika kollektivtrafikförbindelser från ett ställe till ett annat.
I kollektivtrafiken kan du betala med kontanter eller resekort.
I närtågen måste du köpa biljetten i förväg.
Du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat.
Reseplanerarefinska _ svenska _ engelska
Resekort
Med ett resekort (matkakortti) reser du förmånligare än med kontanter.
Resekortet gäller i lokaltrafikens bussar, närtågen, metron, spårvagnarna och Sveaborgsfärjorna.
Det finns två slags resekort.
Det är det billigaste sättet att resa.
Ett innehavarkort (haltijakohtainen kortti) kan användas av flera personer.
Innan du skaffar dig ett personligt kort ska du registrera dig som invånare i någon av kommunerna inom HRT-området.
Du kan köpa resekort vid HRT:s försäljningsställen (myyntipiste) eller serviceställen (palvelupiste).
De finns runtom i huvudstadsregionen.
Personligt resekort kan du köpa vid serviceställena.
Ta med dig identitetsbevis om du ska köpa personligt resekort.
Om du har finska nätbankskoder kan du även köpa personligt resekort på HRT:s webbplats.
Du kan resa med resekortet när du laddar kortet med period (kausi) eller värde (arvo).
En period betyder tid: till exempel en månad.
Värde betyder pengar.
Om du använder kollektivtrafiken ofta tjänar du på att ladda kortet med period.
Du kan ladda resekortet på vilket serviceställe för resekort (matkakortin latauspiste) som helst.
Du hittar mer information på HRT:s webbplats.
Ansökan om försäljningsplatserfinska _ svenska _ engelska
Information och råd till resenärerfinska _ svenska _ engelska
Biljetter och priserfinska _ svenska _ engelska
Att gå och cykla
Om du vill gå eller cykla i Vanda kan du söka en lämplig rutt i reseplaneraren för cykling och gång.
En cykelkarta i pappersformat för Vanda kan du hämta i Vandainfo.
Cykelkartorna är kostnadsfria.
linkkiVanda stad:
Vandainfofinska _ svenska _ engelska
Bil och flyg
Helsingfors-Vanda internationella flygplats ligger i Vanda.
Flygplatsen har goda trafikförbindelser till exempel med bil, buss och tåg.
Du kan parkera bilen på många järnvägsstationer och fortsätta färden med kollektivtrafiken.
Tidtabellerna för bussar och tåg hittar du enkelt i reseplaneraren.
Läs mer: Trafik.
Flygplatsenfinska _ svenska _ engelska _ ryska _ kinesiska
Beslutsfattande och påverkan
I Vanda beslutas ärenden av stadsfullmäktige (kaupunginvaltuusto).
I stadsfullmäktige sitter 67 ledamöter som representerar olika politiska grupper.
Fullmäktige väljs var fjärde år genom kommunalval (kunnallisvaalit).
Invånarna i Vanda kan påverka beslutsfattandet och beredning av ärenden på många olika sätt.
På Vandakanalen kan du följa fullmäktiges sammanträden och få mer information om beslutsfattandet.
I Vanda finns en delegation för mångkulturella frågor (monikulttuurisuusasiain neuvottelukunta) som lägger fram propositioner i ärenden som rör invandrare.
Läs mer på Vanda stads webbplats.
I Vanda finns många politiska föreningar, invandrarföreningar och andra föreningar via vilka du också kan påverka beslutsfattandet.
Mer information om föreningarna hittar du på sidan Vantaalla.info.
linkkiVanda stad:
Beslutsfattandefinska _ svenska _ engelska
linkkiVanda stad:
Delta och påverkafinska
Stadsfullmäktiges sammanträden på Internetfinska
linkkiVanda stad:
Delegationen för mångkulturella frågorfinska
Religion
Många religiösa samfund är verksamma i Vanda och Helsingfors.
Via tjänsten Uskonnot Suomessa kan du söka information efter det religiösa samfundet och orten.
Den evangelisk-lutherska kyrkan har sex finskspråkiga församlingar och en svenskspråkig församling i Vanda.
Läs mer på Vanda kyrkliga samfällighets webbplats.
I Dickursby finns en ortodox kyrka.
Mer information om verksamheten vid den ortodoxa kyrkan i Vanda hittar du på Helsingfors ortodoxa församlings webbplats.
Läs mer: Kulturer och religioner i Finland.
linkkiVanda kyrkliga samfällighet:
Evangelisk-lutherska församlingarfinska
linkkiHelsingfors ortodoxa församling:
Ortodoxa församlingenfinska _ ryska
Religiösa samfundfinska _ engelska
Grundläggande information
Vanda är en av de fyra kommunerna i huvudstadsregionen.
Den ligger intill Esbo och Helsingfors.
Vanda centrum ligger i Dickursby.
Därtill finns det andra stora tätorter i Vanda, till exempel Korso, Björkby-Havukoski, Myrbacka, Mårtensdal, Håkansböle, Västerkulla och Backas.
Vanda har drygt 205 000 invånare.
Av dem är cirka 2,8 procent svenskspråkiga och 11 procent har något annat modersmål än finska eller svenska.
Arealen är cirka 240 km2, varav cirka 2 km2 består av vatten.
linkkiVanda stad:
Grundläggande informationfinska _ svenska _ engelska
Historia
Vanda område har varit bebott länge.
Man har hittat upp till 7 000 år gamla lämningar efter bosättning.
Nuvarande Vanda har uppstått på ett område som förr var Helsingfors socken.
Helsingfors sockens historia sträcker sig ända till 1300-talet.
Helsingfors socken blev först Helsingfors landskommun, sedan Vanda köping år 1972 och till slut Vanda stad år 1974.
Läget som granne till huvudstaden Helsingfors har varit viktigt för Vanda.
Viktiga vägar, såsom vägen från Åbo via Helsingfors till Viborg och senare järnvägen norrut från Helsingfors, har gått genom Vanda.
Längs med vägarna och järnvägen har det utvecklats industrier och bostadsområden.
Vanda är än idag en viktig trafikknutpunkt.
Till exempel ligger Helsingfors-Vanda flygplats i Vanda.
linkkiVanda stad:
Information om Vandafinska
linkkiVanda stad:
Stadsmuseetfinska _ svenska _ engelska
Bibliotek
Motion
Att röra sig i naturen
Teater och film
Museer
Fritidsverksamhet för barn och unga
Fritidsverksamhet för seniorer
Föreningar
Vid Vanda vuxenutbildningsinstitut (Vantaan Aikuisopisto) kan man till exempel skapa konst, handarbeten, laga mat eller dansa.
Man kan även studera språk.
I Vanda finns två kulturhus: konserthuset Martinus och allaktivitetscentret Myrbackahuset.
Dessutom ordnar allaktivitetscentret LUMO många evenemang.
Kulturhuset för barn och unga Fernissan, Konsthuset Pessi och Konsthuset Totem ordnar kulturevenemang för barn.
Läs mer: Fritid.
linkkiVanda vuxenutbildningsinstitut:
Studiehandbokfinska
linkkiVanda stad:
Kulturevenemangfinska _ svenska _ engelska
Konserterfinska _ svenska _ engelska
Evenemangfinska _ engelska
linkkiKulturhuset för barn och unga Fernissan:
Kulturevenemang för barnfinska
Kulturevenemang för barnfinska
Kulturevenemang för barnfinska _ svenska
linkkiVanda stad:
Evenemang och festivalerfinska _ engelska
Bibliotek
I Vanda finns 10 bibliotek (kirjasto) och två bokbussar (kirjastoauto).
På biblioteket kan du låna böcker, tidningar, musik, filmer, spel och mycket annat.
Böcker och annat material finns på flera olika språk.
På biblioteket kan du också använda dator.
På vissa bibliotek ordnas även språkcaféer i det finska språket för invandrare.
Biblioteken i Vanda är med i huvudstadsregionens bibliotekstjänst HelMet.
Du kan alltså använda samma bibliotekskort på stadsbiblioteken i Vanda, Esbo, Grankulla och Helsingfors.
I Helsingfors huvudbibliotek i Böle finns Flerspråkigt bibliotek.
Där hittar man böcker på över 60 olika språk.
Om du har ett Helmet-lånekort, kan du också låna böcker i Flerspråkiga biblioteket.
Läs mer: Bibliotek
linkkiVanda stad:
Information om bibliotekenfinska _ svenska _ engelska
linkkiHelsingfors stadsbibliotek:
Flerspråkiga biblioteketfinska _ svenska _ engelska
Motion
I Vanda finns fem kommunala simhallar.
Simhallen i Korso har ett eget simpass för invandrarkvinnor och -flickor.
I Vanda finns flera idrottshallar, idrottsplaner och andra idrottsplatser för olika idrottsgrenar.
På motionsslingorna kan man springa på somrarna och åka skidor på vintrarna.
Läs mer: Motion.
linkkiVanda stad:
Simhallarnas kontaktuppgifterfinska _ svenska _ engelska
linkkiVanda stad:
Simpass för invandrarkvinnorfinska _ engelska
linkkiVanda stad:
Idrottsklubbarfinska
Att röra sig i naturen
I Vanda finns många motionsslingor och naturstigar.
Du kan även röra dig i naturen i Petikkos rekreationsområde.
Du kan fiska på Vanda stads fiskeområden i Vanda å, Kervo å och på Finska viken.
Läs mer: Att röra sig i naturen.
linkkiVanda stad:
Rekreations- och campingområdenfinska _ svenska
linkkiVanda stad:
Idrottsplatser och friluftsområdenfinska _ svenska
Friluftsområdenfinska
linkkiVanda stad:
Fiske och båtlivfinska
Teater och film
I Vanda finns flera yrkes- och amatörteatrar.
I Vanda finns fyra biografer.
Mer information om filmerna hittar du på biografernas webbplatser.
Därtill ordnar Vanda stad filmvisningar.
Läs mer: Teater och film.
linkkiVanda stad:
Film, dans och teaterfinska _ engelska
Museer
I Vanda finns flera museer.
På Vanda konstmuseum ordnas växlande utställningar med inhemsk och utländsk modern konst.
Om de övriga museerna hittar du information på Vanda stads webbplats.
Läs mer: Museer.
linkkiVanda stad:
Museerfinska _ engelska
linkkiVanda stad:
Stadsmuseetfinska _ svenska _ engelska
linkkiVanda stad:
Konstmuseetfinska _ svenska _ engelska
Fritidsverksamhet för barn och unga
I Vanda finns flera läroanstalter som ger grundundervisning i konst speciellt för barn och unga.
Olika konstarter är musik, bildkonst, dans, teater, cirkuskonst, ordkonst, handarbete och arkitektur.
Stadens ungdomsgårdar är öppna för alla ungdomar i åldrarna 10–17 år.
Projektet Sport för alla (Sporttia kaikille-hanke) ordnar idrottsklubbar, turneringar och läger för barn och ungdomar med invandrarbakgrund.
Också föreningar och idrottsklubbar ordnar mycket verksamhet för ungdomar.
Mer information hittar du på Vanda stads webbplats.
Läs mer: Fritidsverksamhet för barn och unga.
linkkiVanda stad:
Information om hobbymöjligheter för ungdomarfinska
linkkiVanda stad:
Kultur för barn och ungafinska _ svenska _ engelska
linkkiVanda stad:
Information om konstundervisningfinska _ engelska
Ungdomsgårdarfinska
Motionsmöjligheterfinska
Hobbysökningfinska
linkkiVanda stad:
Delta och påverkafinska _ svenska
Fritidsverksamhet för seniorer
Om du har fyllt 70 år och Vanda är din hemkommun kan du kostnadsfritt använda Vanda stads simhallar och gym. Du kommer gratis in till idrottsanläggningarna om du har ett Sportkort (Sporttikortti).
Du kan avhämta Sportkortet kostnadsfritt vid Vanda-informationspunkterna.
Ta med dig identitetsbevis och ett foto när du ansöker om kortet.
På Seniorrådgivningen (seniorineuvonta) får du information om hobbyer och tjänster för seniorer som olika organisationer, företag och staden erbjuder.
Seniorrådgivningen
Tfn: (09) 8392 4202
Motionsmöjligheterfinska _ svenska
Föreningar
I Vanda finns många olika föreningar, till exempel kulturföreningar och idrottsklubbar.
Mer information hittar du på Vanda stads webbplats.
Läs mer: Föreningar.
linkkiVanda stad:
Kulturföreningarfinska
linkkiVanda stad:
Idrottsklubbarfinska
Bibliotek
Motion
Att röra sig i naturen
Teater och film
Museer
Fritidsverksamhet för barn och unga
Fritidsverksamhet för seniorer
Föreningar
Vid Vanda vuxenutbildningsinstitut (Vantaan Aikuisopisto) kan man till exempel skapa konst, handarbeten, laga mat eller dansa.
Man kan även studera språk.
I Vanda finns två kulturhus: konserthuset Martinus och allaktivitetscentret Myrbackahuset.
Dessutom ordnar allaktivitetscentret LUMO många evenemang.
Kulturhuset för barn och unga Fernissan, Konsthuset Pessi och Konsthuset Totem ordnar kulturevenemang för barn.
Läs mer: Fritid.
linkkiVanda vuxenutbildningsinstitut:
Studiehandbokfinska
linkkiVanda stad:
Kulturevenemangfinska _ svenska _ engelska
Konserterfinska _ svenska _ engelska
Evenemangfinska _ engelska
linkkiKulturhuset för barn och unga Fernissan:
Kulturevenemang för barnfinska
Kulturevenemang för barnfinska
Kulturevenemang för barnfinska _ svenska
linkkiVanda stad:
Evenemang och festivalerfinska _ engelska
Bibliotek
I Vanda finns 10 bibliotek (kirjasto) och två bokbussar (kirjastoauto).
På biblioteket kan du låna böcker, tidningar, musik, filmer, spel och mycket annat.
Böcker och annat material finns på flera olika språk.
På biblioteket kan du också använda dator.
På vissa bibliotek ordnas även språkcaféer i det finska språket för invandrare.
Biblioteken i Vanda är med i huvudstadsregionens bibliotekstjänst HelMet.
Du kan alltså använda samma bibliotekskort på stadsbiblioteken i Vanda, Esbo, Grankulla och Helsingfors.
I Helsingfors huvudbibliotek i Böle finns Flerspråkigt bibliotek.
Där hittar man böcker på över 60 olika språk.
Om du har ett Helmet-lånekort, kan du också låna böcker i Flerspråkiga biblioteket.
Läs mer: Bibliotek
linkkiVanda stad:
Information om bibliotekenfinska _ svenska _ engelska
linkkiHelsingfors stadsbibliotek:
Flerspråkiga biblioteketfinska _ svenska _ engelska
Motion
I Vanda finns fem kommunala simhallar.
Simhallen i Korso har ett eget simpass för invandrarkvinnor och -flickor.
I Vanda finns flera idrottshallar, idrottsplaner och andra idrottsplatser för olika idrottsgrenar.
På motionsslingorna kan man springa på somrarna och åka skidor på vintrarna.
Läs mer: Motion.
linkkiVanda stad:
Simhallarnas kontaktuppgifterfinska _ svenska _ engelska
linkkiVanda stad:
Simpass för invandrarkvinnorfinska _ engelska
linkkiVanda stad:
Idrottsklubbarfinska
Att röra sig i naturen
I Vanda finns många motionsslingor och naturstigar.
Du kan även röra dig i naturen i Petikkos rekreationsområde.
Du kan fiska på Vanda stads fiskeområden i Vanda å, Kervo å och på Finska viken.
Läs mer: Att röra sig i naturen.
linkkiVanda stad:
Rekreations- och campingområdenfinska _ svenska
linkkiVanda stad:
Idrottsplatser och friluftsområdenfinska _ svenska
Friluftsområdenfinska
linkkiVanda stad:
Fiske och båtlivfinska
Teater och film
I Vanda finns flera yrkes- och amatörteatrar.
I Vanda finns fyra biografer.
Mer information om filmerna hittar du på biografernas webbplatser.
Därtill ordnar Vanda stad filmvisningar.
Läs mer: Teater och film.
linkkiVanda stad:
Film, dans och teaterfinska _ engelska
Museer
I Vanda finns flera museer.
På Vanda konstmuseum ordnas växlande utställningar med inhemsk och utländsk modern konst.
Om de övriga museerna hittar du information på Vanda stads webbplats.
Läs mer: Museer.
linkkiVanda stad:
Museerfinska _ engelska
linkkiVanda stad:
Stadsmuseetfinska _ svenska _ engelska
linkkiVanda stad:
Konstmuseetfinska _ svenska _ engelska
Fritidsverksamhet för barn och unga
I Vanda finns flera läroanstalter som ger grundundervisning i konst speciellt för barn och unga.
Olika konstarter är musik, bildkonst, dans, teater, cirkuskonst, ordkonst, handarbete och arkitektur.
Stadens ungdomsgårdar är öppna för alla ungdomar i åldrarna 10–17 år.
Projektet Sport för alla (Sporttia kaikille-hanke) ordnar idrottsklubbar, turneringar och läger för barn och ungdomar med invandrarbakgrund.
Också föreningar och idrottsklubbar ordnar mycket verksamhet för ungdomar.
Mer information hittar du på Vanda stads webbplats.
Läs mer: Fritidsverksamhet för barn och unga.
linkkiVanda stad:
Information om hobbymöjligheter för ungdomarfinska
linkkiVanda stad:
Kultur för barn och ungafinska _ svenska _ engelska
linkkiVanda stad:
Information om konstundervisningfinska _ engelska
Ungdomsgårdarfinska
Motionsmöjligheterfinska
Hobbysökningfinska
linkkiVanda stad:
Delta och påverkafinska _ svenska
Fritidsverksamhet för seniorer
Om du har fyllt 70 år och Vanda är din hemkommun kan du kostnadsfritt använda Vanda stads simhallar och gym. Du kommer gratis in till idrottsanläggningarna om du har ett Sportkort (Sporttikortti).
Du kan avhämta Sportkortet kostnadsfritt vid Vanda-informationspunkterna.
Ta med dig identitetsbevis och ett foto när du ansöker om kortet.
På Seniorrådgivningen (seniorineuvonta) får du information om hobbyer och tjänster för seniorer som olika organisationer, företag och staden erbjuder.
Seniorrådgivningen
Tfn: (09) 8392 4202
Motionsmöjligheterfinska _ svenska
Föreningar
I Vanda finns många olika föreningar, till exempel kulturföreningar och idrottsklubbar.
Mer information hittar du på Vanda stads webbplats.
Läs mer: Föreningar.
linkkiVanda stad:
Kulturföreningarfinska
linkkiVanda stad:
Idrottsklubbarfinska
Bibliotek
Motion
Att röra sig i naturen
Teater och film
Museer
Fritidsverksamhet för barn och unga
Fritidsverksamhet för seniorer
Föreningar
Vid Vanda vuxenutbildningsinstitut (Vantaan Aikuisopisto) kan man till exempel skapa konst, handarbeten, laga mat eller dansa.
Man kan även studera språk.
I Vanda finns två kulturhus: konserthuset Martinus och allaktivitetscentret Myrbackahuset.
Dessutom ordnar allaktivitetscentret LUMO många evenemang.
Kulturhuset för barn och unga Fernissan, Konsthuset Pessi och Konsthuset Totem ordnar kulturevenemang för barn.
Läs mer: Fritid.
linkkiVanda vuxenutbildningsinstitut:
Studiehandbokfinska
linkkiVanda stad:
Kulturevenemangfinska _ svenska _ engelska
Konserterfinska _ svenska _ engelska
Evenemangfinska _ engelska
linkkiKulturhuset för barn och unga Fernissan:
Kulturevenemang för barnfinska
Kulturevenemang för barnfinska
Kulturevenemang för barnfinska _ svenska
linkkiVanda stad:
Evenemang och festivalerfinska _ engelska
Bibliotek
I Vanda finns 10 bibliotek (kirjasto) och två bokbussar (kirjastoauto).
På biblioteket kan du låna böcker, tidningar, musik, filmer, spel och mycket annat.
Böcker och annat material finns på flera olika språk.
På biblioteket kan du också använda dator.
På vissa bibliotek ordnas även språkcaféer i det finska språket för invandrare.
Biblioteken i Vanda är med i huvudstadsregionens bibliotekstjänst HelMet.
Du kan alltså använda samma bibliotekskort på stadsbiblioteken i Vanda, Esbo, Grankulla och Helsingfors.
I Helsingfors huvudbibliotek i Böle finns Flerspråkigt bibliotek.
Där hittar man böcker på över 60 olika språk.
Om du har ett Helmet-lånekort, kan du också låna böcker i Flerspråkiga biblioteket.
Läs mer: Bibliotek
linkkiVanda stad:
Information om bibliotekenfinska _ svenska _ engelska
linkkiHelsingfors stadsbibliotek:
Flerspråkiga biblioteketfinska _ svenska _ engelska
Motion
I Vanda finns fem kommunala simhallar.
Simhallen i Korso har ett eget simpass för invandrarkvinnor och -flickor.
I Vanda finns flera idrottshallar, idrottsplaner och andra idrottsplatser för olika idrottsgrenar.
På motionsslingorna kan man springa på somrarna och åka skidor på vintrarna.
Läs mer: Motion.
linkkiVanda stad:
Simhallarnas kontaktuppgifterfinska _ svenska _ engelska
linkkiVanda stad:
Simpass för invandrarkvinnorfinska _ engelska
linkkiVanda stad:
Idrottsklubbarfinska
Att röra sig i naturen
I Vanda finns många motionsslingor och naturstigar.
Du kan även röra dig i naturen i Petikkos rekreationsområde.
Du kan fiska på Vanda stads fiskeområden i Vanda å, Kervo å och på Finska viken.
Läs mer: Att röra sig i naturen.
linkkiVanda stad:
Rekreations- och campingområdenfinska _ svenska
linkkiVanda stad:
Idrottsplatser och friluftsområdenfinska _ svenska
Friluftsområdenfinska
linkkiVanda stad:
Fiske och båtlivfinska
Teater och film
I Vanda finns flera yrkes- och amatörteatrar.
I Vanda finns fyra biografer.
Mer information om filmerna hittar du på biografernas webbplatser.
Därtill ordnar Vanda stad filmvisningar.
Läs mer: Teater och film.
linkkiVanda stad:
Film, dans och teaterfinska _ engelska
Museer
I Vanda finns flera museer.
På Vanda konstmuseum ordnas växlande utställningar med inhemsk och utländsk modern konst.
Om de övriga museerna hittar du information på Vanda stads webbplats.
Läs mer: Museer.
linkkiVanda stad:
Museerfinska _ engelska
linkkiVanda stad:
Stadsmuseetfinska _ svenska _ engelska
linkkiVanda stad:
Konstmuseetfinska _ svenska _ engelska
Fritidsverksamhet för barn och unga
I Vanda finns flera läroanstalter som ger grundundervisning i konst speciellt för barn och unga.
Olika konstarter är musik, bildkonst, dans, teater, cirkuskonst, ordkonst, handarbete och arkitektur.
Stadens ungdomsgårdar är öppna för alla ungdomar i åldrarna 10–17 år.
Projektet Sport för alla (Sporttia kaikille-hanke) ordnar idrottsklubbar, turneringar och läger för barn och ungdomar med invandrarbakgrund.
Också föreningar och idrottsklubbar ordnar mycket verksamhet för ungdomar.
Mer information hittar du på Vanda stads webbplats.
Läs mer: Fritidsverksamhet för barn och unga.
linkkiVanda stad:
Information om hobbymöjligheter för ungdomarfinska
linkkiVanda stad:
Kultur för barn och ungafinska _ svenska _ engelska
linkkiVanda stad:
Information om konstundervisningfinska _ engelska
Ungdomsgårdarfinska
Motionsmöjligheterfinska
Hobbysökningfinska
linkkiVanda stad:
Delta och påverkafinska _ svenska
Fritidsverksamhet för seniorer
Om du har fyllt 70 år och Vanda är din hemkommun kan du kostnadsfritt använda Vanda stads simhallar och gym. Du kommer gratis in till idrottsanläggningarna om du har ett Sportkort (Sporttikortti).
Du kan avhämta Sportkortet kostnadsfritt vid Vanda-informationspunkterna.
Ta med dig identitetsbevis och ett foto när du ansöker om kortet.
På Seniorrådgivningen (seniorineuvonta) får du information om hobbyer och tjänster för seniorer som olika organisationer, företag och staden erbjuder.
Seniorrådgivningen
Tfn: (09) 8392 4202
Motionsmöjligheterfinska _ svenska
Föreningar
I Vanda finns många olika föreningar, till exempel kulturföreningar och idrottsklubbar.
Mer information hittar du på Vanda stads webbplats.
Läs mer: Föreningar.
linkkiVanda stad:
Kulturföreningarfinska
linkkiVanda stad:
Idrottsklubbarfinska
Problem med uppehållstillståndet
Brott
Behöver du en jurist?
Våld
Missbruksproblem och spelberoende
Dödsfall
Om du behöver brådskande hjälp av polisen, brandkåren eller ambulansen, ring nödnumret 112.
Du får ringa nödnumret endast i brådskande nödfall där liv, hälsa, egendom eller miljö är i fara.
Om du drabbas av en akut krissituation, såsom att en närstående avlider eller på grund av familjevåld, kan du kontakta social- och krisjouren (sosiaali- ja kriisipäivystys).
Du kan också söka hjälp för en familjemedlem eller en vän.
Social- och krisjouren har öppet dygnet runt varje dag.
Social- och krisjouren
Tfn (09) 8392 4005
linkkiNödcentralsverket:
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
linkkiVanda stad:
Social- och krisjourenfinska _ svenska _ engelska
Problem med uppehållstillståndet
Om du har problem eller oklarheter med uppehållstillståndet, kontakta Migrationsverket.
Du kan även fråga om råd på rådgivningstjänsterna för invandrare.
Information om tjänsterna finns på sidan Som invandrare i Vanda.
Migrationsverkets närmaste tjänsteställe finns i Helsingfors:
Göksgränd 3A
Läs mer: Problem med uppehållstillståndet
Olika tillståndfinska _ svenska _ engelska
Hälsovård för papperslösa
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärhälsovård.
Tjänsterna vid Global Clinic är avgiftsfria för kunderna.
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter.
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
Telefonnumret till Global Clinic i Helsingfors är 044 977 4547.
Samtalet besvaras av en sjukskötare eller en läkare.
E-postadressen är globalclinic.finland(at)gmail.com.
Läs mer: Problem med uppehållstillstånd
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Brott
Brottsanmälan (rikosilmoitus) kan göras per telefon eller personligen på polisstationen.
Du kan också göra brottsanmälan på internet om brottet i fråga är ringa och du inte behöver omedelbar hjälp av polisen.
Konvaljvägen 21
Tfn 0295 430291
Läs mer: Brott.
Kontaktuppgifterfinska _ svenska
Elektronisk polisanmälanfinska _ svenska _ engelska
Behöver du en jurist?
Östra Nylands rättshjälpsbyrå (Itä-Uudenmaan oikeusaputoimisto) betjänar invånarna i Vanda.
Pyrolavägen 37
Tfn 029 5660 160
Du kan också söka information om privata jurister på till exempel Finlands Juristförbunds (Suomen Asianajajaliitto) webbplats.
Läs mer: Behöver du en jurist?
linkkiÖstra Nylands rättshjälpsbyrå:
Information om rättshjälpfinska _ svenska _ engelska
linkkiFinlands Advokatförbund:
Advokaterfinska _ svenska _ engelska
Våld
I nödsituationer ringer du nödnumret 112.
I krissituationer får man även hjälp vid Vanda stads social- och krisjour (sosiaali- ja kriisipäivystys), som har öppet dygnet runt.
Social- och krisjouren
Tfn (09) 8392 4005
linkkiNödcentralsverket:
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
Skyddshem
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta ett skyddshem (turvakoti).
Skyddshemmen har jourmottagning dygnet runt.
Skyddshemmet Mona (turvakoti Mona) är ett skyddshem avsett för invandrarkvinnor och deras barn.
Tfn 045 639 6274
linkkiTurvakoti Mona:
Skyddshemfinska
Du kan även gå till Vanda skyddshem (Vantaan turvakoti) eller huvudstadsregionens skyddshem (pääkaupunkiseudun turvakoti).
Puh. (09) 8392 0071
Skyddshemfinska _ engelska
Steniusvägen 20
Tfn (09) 4777 180
Hjälp till offer för familjevåldfinska
Hjälp för invandrarkvinnor
Föreningen Monika-Naiset liitto (Monika-Naiset Liitto) ger råd och stöd till invandrarkvinnor.
Föreningen har ett resurscenter (voimavarakeskus) i Vanda där man får stöd och råd.
Tfn (09) 839 35013
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Hjälp för män
Män som har utövat våld mot sina familjemedlemmar eller har själva blivit offer för våld i hemmet, kan få hjälp från Jussi-arbetet i Vanda (Vantaan Jussi-työ).
Hjälp för män att sluta med våldsamt beteendefinska
Miehen linja (Miehen linja) hjälper invandrarmän som har problem med våld.
Tfn (09) 276 62899
Hjälp för män för att sluta med våldsamt beteendefinska _ engelska
Hjälp för unga
Finlands Röda Kors De ungas skyddshus (Suomen Punaisen Ristin Nuorten turvatalo) ger stöd och hjälp i krissituationer för 12–19-åringar.
Skyddshuset har öppet kl. 17–10, telefonjouren betjänar dygnet runt.
Sjukhusgatan 3 (Räckhals gård)
Tfn (09) 871 4043
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Läs mer: Våld
Problem i äktenskap eller parförhållande
Par med barn under 13 år kan vid problem i äktenskap och parförhållande få hjälp vid familjerådgivningen (perheneuvola).
Kontaktuppgifterna hittar du på Vanda stads webbplats.
Familjerådgivningens tjänster är konfidentiella och avgiftsfria.
Vid akuta krissituationer inom familjen kan du kontakta social- och krisjouren (sosiaali- ja kriisipäivystys), som har öppet dygnet runt varje dag.
Social- och krisjouren
Tfn (09) 8392 4005
Vid problem i parförhållandet och familjen får man även hjälp av familjerådgivningen vid Vanda församlingar (Vantaan seurakunnan perheneuvonta).
Läs mer: Problem i äktenskap och parförhållande
linkkiVanda stad:
Familjerådgivningarfinska _ svenska
linkkiVanda kyrkliga samfällighet:
Familjerådgivningfinska _ engelska
Barnrådgivningsbyråerna (lastenneuvola) och familjerådgivningsbyråerna (perheneuvola) ger råd i frågor som rör barns hälsa, uppväxt och utveckling.
Vid problem hos barn i skolåldern får man hjälp hos skolhälsovårdarna (kouluterveydenhoitaja), skolkuratorerna (koulukuraattori) och socialhandledarna (sosiaaliohjaaja).
Mer information hittar du på Vanda stads webbplats.
Läs mer: Barns och ungas problem
linkkiVanda stad:
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad:
Familjerådgivningarfinska _ svenska
linkkiVanda stad:
Information om tjänster för barn, ungdomar och familjerfinska _ svenska _ engelska
I skolan får de unga hjälp av skol- och studenthälsovårdarna (koulu- ja opiskeluterveydenhoitajat), skolkuratorerna (koulukuraattorit) och skolpsykologerna (koulupsykologit).
linkkiVanda stad:
Information om skolhälsovårdenfinska _ svenska _ engelska
linkkiVanda stad:
Skolkuratorerfinska _ svenska
linkkiVanda stad:
Skolpsykologerfinska _ svenska
Nuppi
13–21-åriga barn och ungdomar samt deras familjer kan få hjälp hos ungdomscentralen (nuortenkeskus).
På Nuppi kan du till exempel få hjälp med mentala problem och missbruksproblem.
Hjälp för ungafinska _ svenska _ engelska
Om du är under 30 år, kan du få råd och handledning via tjänsten Navigatorn.
Personalen vid Navigatorn hjälper dig om du inte har något arbete eller en studieplats.
Du kan även be om råd gällande andra saker, till exempel boende och ekonomi.
De ungas skyddshus
Finlands Röda Kors De ungas skyddshus (Suomen Punaisen Ristin Nuorten turvatalo) ger stöd och hjälp i krissituationer för 12–19-åringar.
Skyddshuset har öppet kl. 17–10, telefonjouren betjänar dygnet runt.
Sjukhusgatan 3
Tfn (09) 871 4043
Läs mer: Barns och ungas problem
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Vägledning och stöd för ungafinska _ svenska
Socialrådgivningen (sosiaalineuvonta) ger information om utkomststöd (toimeentulotuki) och andra bidrag om du har ekonomiska problem.
Tfn (09) 83 911.
linkkiVanda stad:
Socialrådgivningenfinska _ svenska _ engelska
Utkomststöd
Utkomststödet (toimeentulotuki) är avsett som en sista utväg då du inte har några andra inkomster eller medel, eller om dina inkomster är mycket låga.
Utkomststöd kan du få om du inte lyckas få tillräckliga inkomster genom eget arbete, andras omsorg eller på något annat sätt.
Du kan be om råd gällande ansökan om utkomststöd via den centraliserade telefontjänsten tfn (09) 8392 1119.
linkkiVanda stad:
Information om utkomststödfinska _ svenska _ engelska
Ekonomi- och skuldrådgivning
Om du inte kan betala dina räkningar eller skulder då de förfaller, ska du kontakta skuldrådgivningen (velkaneuvonta).
Tfn (09) 8392 2120.
linkkiVanda ekonomi- och skuldrådgivning:
Ekonomi- och skuldrådgivningfinska _ svenska _ engelska
Social kreditgivning
Om du har låga inkomster och är medellös samt har svårt att få lån, kan du ansöka om lån via den sociala kreditgivningen (sosiaalinen luototus).
Telefonnumret till kundrådgivningen och tidsbokningen är (09) 8392 0173.
linkkiVanda stad:
Information om social kreditgivningfinska _ svenska _ engelska
Missbruksproblem och spelberoende
Itä-Vantaan A-klinikka
Konvaljvägen 20 C vån.
tfn (09) 8392 3415
Länsi-Vantaan A-klinikka
tfn (09) 8393 5534
H-klinikka
Eldstadsvägen 7 B, vån.
Tfn (09) 839 21064
H-kliniken har också verksamhetsställen på Dickursby och Myrbacka hälsostationer.
Om du har spelproblem kan du söka hjälp vid Spelkliniken (Peliklinikka), som finns i centrala Helsingfors.
Peliklinikka
tfn 040 152 3918.
Ungdomscentralen Nuppi (nuortenkeskus Nuppi) hjälper ungdomar med missbruksproblem, Internetberoende eller spelberoende.
Nuppi ger också stöd till ungdomar som oroar sig för rusmedelsbruket hos någon närstående person.
Läs mer: Missbruksproblem.
linkkiVanda stad:
Hjälp med missbruksproblemfinska _ svenska _ engelska
linkkiVanda stad:
Information om vård av drogproblemfinska _ svenska _ engelska
Hjälp med penningspelproblemfinska
Hjälp för ungafinska _ svenska _ engelska
Dödsfall
I Vanda finns fyra begravningsplatser som tillhör de evangelisk-lutherska församlingarna.
I Furumo i Vanda finns dessutom Vandas och Helsingfors gemensamma begravningsplats för avlidna personer som inte har varit medlemmar i något religionssamfund.
Information om begravning får du på Vanda församlingars gravkontor (Vantaan seurakuntien hautaustoimisto) och vid privata begravningsbyråer (hautaustoimisto).
Vanda församlingars gravkontor
Prästgårdsgränden 5
Tfn (09) 8306 220
Om din närstående avlider plötsligt, kan du få hjälp med att återhämta dig från den chockartade upplevelsen och stöd i att klara dig efter förlusten av Vandas social- och krisjour (sosiaali- ja kriisipäivystys).
Jouren har öppet varje dag dygnet runt.
Social- och krisjouren
Tfn (09) 8392 4005
Läs mer: Död
linkkiVanda kyrkliga samfällighet:
Begravningsplatserfinska
linkkiHelsingfors kyrkliga samfällighet:
Konfessionslös begravningsplatsfinska
linkkiFinlands Begravningbyråers Förbund:
Begravningsbyråerfinska _ svenska _ engelska
När en närstående har avliditfinska _ svenska _ engelska
linkkiVanda stad:
Social- och krisjourenfinska _ svenska _ engelska
Problem med uppehållstillståndet
Brott
Behöver du en jurist?
Våld
Missbruksproblem och spelberoende
Dödsfall
Om du behöver brådskande hjälp av polisen, brandkåren eller ambulansen, ring nödnumret 112.
Du får ringa nödnumret endast i brådskande nödfall där liv, hälsa, egendom eller miljö är i fara.
Om du drabbas av en akut krissituation, såsom att en närstående avlider eller på grund av familjevåld, kan du kontakta social- och krisjouren (sosiaali- ja kriisipäivystys).
Du kan också söka hjälp för en familjemedlem eller en vän.
Social- och krisjouren har öppet dygnet runt varje dag.
Social- och krisjouren
Tfn (09) 8392 4005
linkkiNödcentralsverket:
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
linkkiVanda stad:
Social- och krisjourenfinska _ svenska _ engelska
Problem med uppehållstillståndet
Om du har problem eller oklarheter med uppehållstillståndet, kontakta Migrationsverket.
Du kan även fråga om råd på rådgivningstjänsterna för invandrare.
Information om tjänsterna finns på sidan Som invandrare i Vanda.
Migrationsverkets närmaste tjänsteställe finns i Helsingfors:
Göksgränd 3A
Läs mer: Problem med uppehållstillståndet
Olika tillståndfinska _ svenska _ engelska
Hälsovård för papperslösa
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärhälsovård.
Tjänsterna vid Global Clinic är avgiftsfria för kunderna.
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter.
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
Telefonnumret till Global Clinic i Helsingfors är 044 977 4547.
Samtalet besvaras av en sjukskötare eller en läkare.
E-postadressen är globalclinic.finland(at)gmail.com.
Läs mer: Problem med uppehållstillstånd
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Brott
Brottsanmälan (rikosilmoitus) kan göras per telefon eller personligen på polisstationen.
Du kan också göra brottsanmälan på internet om brottet i fråga är ringa och du inte behöver omedelbar hjälp av polisen.
Konvaljvägen 21
Tfn 0295 430291
Läs mer: Brott.
Kontaktuppgifterfinska _ svenska
Elektronisk polisanmälanfinska _ svenska _ engelska
Behöver du en jurist?
Östra Nylands rättshjälpsbyrå (Itä-Uudenmaan oikeusaputoimisto) betjänar invånarna i Vanda.
Pyrolavägen 37
Tfn 029 5660 160
Du kan också söka information om privata jurister på till exempel Finlands Juristförbunds (Suomen Asianajajaliitto) webbplats.
Läs mer: Behöver du en jurist?
linkkiÖstra Nylands rättshjälpsbyrå:
Information om rättshjälpfinska _ svenska _ engelska
linkkiFinlands Advokatförbund:
Advokaterfinska _ svenska _ engelska
Våld
I nödsituationer ringer du nödnumret 112.
I krissituationer får man även hjälp vid Vanda stads social- och krisjour (sosiaali- ja kriisipäivystys), som har öppet dygnet runt.
Social- och krisjouren
Tfn (09) 8392 4005
linkkiNödcentralsverket:
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
Skyddshem
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta ett skyddshem (turvakoti).
Skyddshemmen har jourmottagning dygnet runt.
Skyddshemmet Mona (turvakoti Mona) är ett skyddshem avsett för invandrarkvinnor och deras barn.
Tfn 045 639 6274
linkkiTurvakoti Mona:
Skyddshemfinska
Du kan även gå till Vanda skyddshem (Vantaan turvakoti) eller huvudstadsregionens skyddshem (pääkaupunkiseudun turvakoti).
Puh. (09) 8392 0071
Skyddshemfinska _ engelska
Steniusvägen 20
Tfn (09) 4777 180
Hjälp till offer för familjevåldfinska
Hjälp för invandrarkvinnor
Föreningen Monika-Naiset liitto (Monika-Naiset Liitto) ger råd och stöd till invandrarkvinnor.
Föreningen har ett resurscenter (voimavarakeskus) i Vanda där man får stöd och råd.
Tfn (09) 839 35013
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Hjälp för män
Män som har utövat våld mot sina familjemedlemmar eller har själva blivit offer för våld i hemmet, kan få hjälp från Jussi-arbetet i Vanda (Vantaan Jussi-työ).
Hjälp för män att sluta med våldsamt beteendefinska
Miehen linja (Miehen linja) hjälper invandrarmän som har problem med våld.
Tfn (09) 276 62899
Hjälp för män för att sluta med våldsamt beteendefinska _ engelska
Hjälp för unga
Finlands Röda Kors De ungas skyddshus (Suomen Punaisen Ristin Nuorten turvatalo) ger stöd och hjälp i krissituationer för 12–19-åringar.
Skyddshuset har öppet kl. 17–10, telefonjouren betjänar dygnet runt.
Sjukhusgatan 3 (Räckhals gård)
Tfn (09) 871 4043
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Läs mer: Våld
Problem i äktenskap eller parförhållande
Par med barn under 13 år kan vid problem i äktenskap och parförhållande få hjälp vid familjerådgivningen (perheneuvola).
Kontaktuppgifterna hittar du på Vanda stads webbplats.
Familjerådgivningens tjänster är konfidentiella och avgiftsfria.
Vid akuta krissituationer inom familjen kan du kontakta social- och krisjouren (sosiaali- ja kriisipäivystys), som har öppet dygnet runt varje dag.
Social- och krisjouren
Tfn (09) 8392 4005
Vid problem i parförhållandet och familjen får man även hjälp av familjerådgivningen vid Vanda församlingar (Vantaan seurakunnan perheneuvonta).
Läs mer: Problem i äktenskap och parförhållande
linkkiVanda stad:
Familjerådgivningarfinska _ svenska
linkkiVanda kyrkliga samfällighet:
Familjerådgivningfinska _ engelska
Barnrådgivningsbyråerna (lastenneuvola) och familjerådgivningsbyråerna (perheneuvola) ger råd i frågor som rör barns hälsa, uppväxt och utveckling.
Vid problem hos barn i skolåldern får man hjälp hos skolhälsovårdarna (kouluterveydenhoitaja), skolkuratorerna (koulukuraattori) och socialhandledarna (sosiaaliohjaaja).
Mer information hittar du på Vanda stads webbplats.
Läs mer: Barns och ungas problem
linkkiVanda stad:
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad:
Familjerådgivningarfinska _ svenska
linkkiVanda stad:
Information om tjänster för barn, ungdomar och familjerfinska _ svenska _ engelska
I skolan får de unga hjälp av skol- och studenthälsovårdarna (koulu- ja opiskeluterveydenhoitajat), skolkuratorerna (koulukuraattorit) och skolpsykologerna (koulupsykologit).
linkkiVanda stad:
Information om skolhälsovårdenfinska _ svenska _ engelska
linkkiVanda stad:
Skolkuratorerfinska _ svenska
linkkiVanda stad:
Skolpsykologerfinska _ svenska
Nuppi
13–21-åriga barn och ungdomar samt deras familjer kan få hjälp hos ungdomscentralen (nuortenkeskus).
På Nuppi kan du till exempel få hjälp med mentala problem och missbruksproblem.
Hjälp för ungafinska _ svenska _ engelska
Om du är under 30 år, kan du få råd och handledning via tjänsten Navigatorn.
Personalen vid Navigatorn hjälper dig om du inte har något arbete eller en studieplats.
Du kan även be om råd gällande andra saker, till exempel boende och ekonomi.
De ungas skyddshus
Finlands Röda Kors De ungas skyddshus (Suomen Punaisen Ristin Nuorten turvatalo) ger stöd och hjälp i krissituationer för 12–19-åringar.
Skyddshuset har öppet kl. 17–10, telefonjouren betjänar dygnet runt.
Sjukhusgatan 3
Tfn (09) 871 4043
Läs mer: Barns och ungas problem
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Vägledning och stöd för ungafinska _ svenska
Socialrådgivningen (sosiaalineuvonta) ger information om utkomststöd (toimeentulotuki) och andra bidrag om du har ekonomiska problem.
Tfn (09) 83 911.
linkkiVanda stad:
Socialrådgivningenfinska _ svenska _ engelska
Utkomststöd
Utkomststödet (toimeentulotuki) är avsett som en sista utväg då du inte har några andra inkomster eller medel, eller om dina inkomster är mycket låga.
Utkomststöd kan du få om du inte lyckas få tillräckliga inkomster genom eget arbete, andras omsorg eller på något annat sätt.
Du kan be om råd gällande ansökan om utkomststöd via den centraliserade telefontjänsten tfn (09) 8392 1119.
linkkiVanda stad:
Information om utkomststödfinska _ svenska _ engelska
Ekonomi- och skuldrådgivning
Om du inte kan betala dina räkningar eller skulder då de förfaller, ska du kontakta skuldrådgivningen (velkaneuvonta).
Tfn (09) 8392 2120.
linkkiVanda ekonomi- och skuldrådgivning:
Ekonomi- och skuldrådgivningfinska _ svenska _ engelska
Social kreditgivning
Om du har låga inkomster och är medellös samt har svårt att få lån, kan du ansöka om lån via den sociala kreditgivningen (sosiaalinen luototus).
Telefonnumret till kundrådgivningen och tidsbokningen är (09) 8392 0173.
linkkiVanda stad:
Information om social kreditgivningfinska _ svenska _ engelska
Missbruksproblem och spelberoende
Itä-Vantaan A-klinikka
Konvaljvägen 20 C vån.
tfn (09) 8392 3415
Länsi-Vantaan A-klinikka
tfn (09) 8393 5534
H-klinikka
Eldstadsvägen 7 B, vån.
Tfn (09) 839 21064
H-kliniken har också verksamhetsställen på Dickursby och Myrbacka hälsostationer.
Om du har spelproblem kan du söka hjälp vid Spelkliniken (Peliklinikka), som finns i centrala Helsingfors.
Peliklinikka
tfn 040 152 3918.
Ungdomscentralen Nuppi (nuortenkeskus Nuppi) hjälper ungdomar med missbruksproblem, Internetberoende eller spelberoende.
Nuppi ger också stöd till ungdomar som oroar sig för rusmedelsbruket hos någon närstående person.
Läs mer: Missbruksproblem.
linkkiVanda stad:
Hjälp med missbruksproblemfinska _ svenska _ engelska
linkkiVanda stad:
Information om vård av drogproblemfinska _ svenska _ engelska
Hjälp med penningspelproblemfinska
Hjälp för ungafinska _ svenska _ engelska
Dödsfall
I Vanda finns fyra begravningsplatser som tillhör de evangelisk-lutherska församlingarna.
I Furumo i Vanda finns dessutom Vandas och Helsingfors gemensamma begravningsplats för avlidna personer som inte har varit medlemmar i något religionssamfund.
Information om begravning får du på Vanda församlingars gravkontor (Vantaan seurakuntien hautaustoimisto) och vid privata begravningsbyråer (hautaustoimisto).
Vanda församlingars gravkontor
Prästgårdsgränden 5
Tfn (09) 8306 220
Om din närstående avlider plötsligt, kan du få hjälp med att återhämta dig från den chockartade upplevelsen och stöd i att klara dig efter förlusten av Vandas social- och krisjour (sosiaali- ja kriisipäivystys).
Jouren har öppet varje dag dygnet runt.
Social- och krisjouren
Tfn (09) 8392 4005
Läs mer: Död
linkkiVanda kyrkliga samfällighet:
Begravningsplatserfinska
linkkiHelsingfors kyrkliga samfällighet:
Konfessionslös begravningsplatsfinska
linkkiFinlands Begravningbyråers Förbund:
Begravningsbyråerfinska
När en närstående har avliditfinska _ svenska _ engelska
linkkiVanda stad:
Social- och krisjourenfinska _ svenska _ engelska
Problem med uppehållstillståndet
Brott
Behöver du en jurist?
Våld
Missbruksproblem och spelberoende
Dödsfall
Om du behöver brådskande hjälp av polisen, brandkåren eller ambulansen, ring nödnumret 112.
Du får ringa nödnumret endast i brådskande nödfall där liv, hälsa, egendom eller miljö är i fara.
Om du drabbas av en akut krissituation, såsom att en närstående avlider eller på grund av familjevåld, kan du kontakta social- och krisjouren (sosiaali- ja kriisipäivystys).
Du kan också söka hjälp för en familjemedlem eller en vän.
Social- och krisjouren har öppet dygnet runt varje dag.
Social- och krisjouren
Tfn (09) 8392 4005
linkkiNödcentralsverket:
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
linkkiVanda stad:
Social- och krisjourenfinska _ svenska _ engelska
Problem med uppehållstillståndet
Om du har problem eller oklarheter med uppehållstillståndet, kontakta Migrationsverket.
Du kan även fråga om råd på rådgivningstjänsterna för invandrare.
Information om tjänsterna finns på sidan Som invandrare i Vanda.
Migrationsverkets närmaste tjänsteställe finns i Helsingfors:
Göksgränd 3A
Läs mer: Problem med uppehållstillståndet
Olika tillståndfinska _ svenska _ engelska
Hälsovård för papperslösa
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärhälsovård.
Tjänsterna vid Global Clinic är avgiftsfria för kunderna.
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter.
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
Telefonnumret till Global Clinic i Helsingfors är 044 977 4547.
Samtalet besvaras av en sjukskötare eller en läkare.
E-postadressen är globalclinic.finland(at)gmail.com.
Läs mer: Problem med uppehållstillstånd
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Brott
Brottsanmälan (rikosilmoitus) kan göras per telefon eller personligen på polisstationen.
Du kan också göra brottsanmälan på internet om brottet i fråga är ringa och du inte behöver omedelbar hjälp av polisen.
Konvaljvägen 21
Tfn 0295 430291
Läs mer: Brott.
Kontaktuppgifterfinska _ svenska
Elektronisk polisanmälanfinska _ svenska _ engelska
Behöver du en jurist?
Östra Nylands rättshjälpsbyrå (Itä-Uudenmaan oikeusaputoimisto) betjänar invånarna i Vanda.
Pyrolavägen 37
Tfn 029 5660 160
Du kan också söka information om privata jurister på till exempel Finlands Juristförbunds (Suomen Asianajajaliitto) webbplats.
Läs mer: Behöver du en jurist?
linkkiÖstra Nylands rättshjälpsbyrå:
Information om rättshjälpfinska _ svenska _ engelska
linkkiFinlands Advokatförbund:
Advokaterfinska _ svenska _ engelska
Våld
I nödsituationer ringer du nödnumret 112.
I krissituationer får man även hjälp vid Vanda stads social- och krisjour (sosiaali- ja kriisipäivystys), som har öppet dygnet runt.
Social- och krisjouren
Tfn (09) 8392 4005
linkkiNödcentralsverket:
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
Skyddshem
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta ett skyddshem (turvakoti).
Skyddshemmen har jourmottagning dygnet runt.
Skyddshemmet Mona (turvakoti Mona) är ett skyddshem avsett för invandrarkvinnor och deras barn.
Tfn 045 639 6274
linkkiTurvakoti Mona:
Skyddshemfinska
Du kan även gå till Vanda skyddshem (Vantaan turvakoti) eller huvudstadsregionens skyddshem (pääkaupunkiseudun turvakoti).
Puh. (09) 8392 0071
Skyddshemfinska _ engelska
Steniusvägen 20
Tfn (09) 4777 180
Hjälp till offer för familjevåldfinska
Hjälp för invandrarkvinnor
Föreningen Monika-Naiset liitto (Monika-Naiset Liitto) ger råd och stöd till invandrarkvinnor.
Föreningen har ett resurscenter (voimavarakeskus) i Vanda där man får stöd och råd.
Tfn (09) 839 35013
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Hjälp för män
Män som har utövat våld mot sina familjemedlemmar eller har själva blivit offer för våld i hemmet, kan få hjälp från Jussi-arbetet i Vanda (Vantaan Jussi-työ).
Hjälp för män att sluta med våldsamt beteendefinska
Miehen linja (Miehen linja) hjälper invandrarmän som har problem med våld.
Tfn (09) 276 62899
Hjälp för män för att sluta med våldsamt beteendefinska _ engelska
Hjälp för unga
Finlands Röda Kors De ungas skyddshus (Suomen Punaisen Ristin Nuorten turvatalo) ger stöd och hjälp i krissituationer för 12–19-åringar.
Skyddshuset har öppet kl. 17–10, telefonjouren betjänar dygnet runt.
Sjukhusgatan 3 (Räckhals gård)
Tfn (09) 871 4043
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Läs mer: Våld
Problem i äktenskap eller parförhållande
Par med barn under 13 år kan vid problem i äktenskap och parförhållande få hjälp vid familjerådgivningen (perheneuvola).
Kontaktuppgifterna hittar du på Vanda stads webbplats.
Familjerådgivningens tjänster är konfidentiella och avgiftsfria.
Vid akuta krissituationer inom familjen kan du kontakta social- och krisjouren (sosiaali- ja kriisipäivystys), som har öppet dygnet runt varje dag.
Social- och krisjouren
Tfn (09) 8392 4005
Vid problem i parförhållandet och familjen får man även hjälp av familjerådgivningen vid Vanda församlingar (Vantaan seurakunnan perheneuvonta).
Läs mer: Problem i äktenskap och parförhållande
linkkiVanda stad:
Familjerådgivningarfinska _ svenska
linkkiVanda kyrkliga samfällighet:
Familjerådgivningfinska _ engelska
Barnrådgivningsbyråerna (lastenneuvola) och familjerådgivningsbyråerna (perheneuvola) ger råd i frågor som rör barns hälsa, uppväxt och utveckling.
Vid problem hos barn i skolåldern får man hjälp hos skolhälsovårdarna (kouluterveydenhoitaja), skolkuratorerna (koulukuraattori) och socialhandledarna (sosiaaliohjaaja).
Mer information hittar du på Vanda stads webbplats.
Läs mer: Barns och ungas problem
linkkiVanda stad:
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad:
Familjerådgivningarfinska _ svenska
linkkiVanda stad:
Information om tjänster för barn, ungdomar och familjerfinska _ svenska _ engelska
I skolan får de unga hjälp av skol- och studenthälsovårdarna (koulu- ja opiskeluterveydenhoitajat), skolkuratorerna (koulukuraattorit) och skolpsykologerna (koulupsykologit).
linkkiVanda stad:
Information om skolhälsovårdenfinska _ svenska _ engelska
linkkiVanda stad:
Skolkuratorerfinska _ svenska
linkkiVanda stad:
Skolpsykologerfinska _ svenska
Nuppi
13–21-åriga barn och ungdomar samt deras familjer kan få hjälp hos ungdomscentralen (nuortenkeskus).
På Nuppi kan du till exempel få hjälp med mentala problem och missbruksproblem.
Hjälp för ungafinska _ svenska _ engelska
Om du är under 30 år, kan du få råd och handledning via tjänsten Navigatorn.
Personalen vid Navigatorn hjälper dig om du inte har något arbete eller en studieplats.
Du kan även be om råd gällande andra saker, till exempel boende och ekonomi.
De ungas skyddshus
Finlands Röda Kors De ungas skyddshus (Suomen Punaisen Ristin Nuorten turvatalo) ger stöd och hjälp i krissituationer för 12–19-åringar.
Skyddshuset har öppet kl. 17–10, telefonjouren betjänar dygnet runt.
Sjukhusgatan 3
Tfn (09) 871 4043
Läs mer: Barns och ungas problem
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Vägledning och stöd för ungafinska _ svenska
Socialrådgivningen (sosiaalineuvonta) ger information om utkomststöd (toimeentulotuki) och andra bidrag om du har ekonomiska problem.
Tfn (09) 83 911.
linkkiVanda stad:
Socialrådgivningenfinska _ svenska _ engelska
Utkomststöd
Utkomststödet (toimeentulotuki) är avsett som en sista utväg då du inte har några andra inkomster eller medel, eller om dina inkomster är mycket låga.
Utkomststöd kan du få om du inte lyckas få tillräckliga inkomster genom eget arbete, andras omsorg eller på något annat sätt.
Du kan be om råd gällande ansökan om utkomststöd via den centraliserade telefontjänsten tfn (09) 8392 1119.
linkkiVanda stad:
Information om utkomststödfinska _ svenska _ engelska
Ekonomi- och skuldrådgivning
Om du inte kan betala dina räkningar eller skulder då de förfaller, ska du kontakta skuldrådgivningen (velkaneuvonta).
Tfn 029 566 0175.
linkkiVanda ekonomi- och skuldrådgivning:
Ekonomi- och skuldrådgivningfinska _ svenska _ engelska
Social kreditgivning
Om du har låga inkomster och är medellös samt har svårt att få lån, kan du ansöka om lån via den sociala kreditgivningen (sosiaalinen luototus).
Telefonnumret till kundrådgivningen och tidsbokningen är (09) 8392 0173.
linkkiVanda stad:
Information om social kreditgivningfinska _ svenska _ engelska
Missbruksproblem och spelberoende
Itä-Vantaan A-klinikka
Konvaljvägen 20 C vån.
tfn (09) 8392 3415
Länsi-Vantaan A-klinikka
tfn (09) 8393 5534
H-klinikka
Eldstadsvägen 7 B, vån.
Tfn (09) 839 21064
H-kliniken har också verksamhetsställen på Dickursby och Myrbacka hälsostationer.
Om du har spelproblem kan du söka hjälp vid Spelkliniken (Peliklinikka), som finns i centrala Helsingfors.
Peliklinikka
tfn 040 152 3918.
Ungdomscentralen Nuppi (nuortenkeskus Nuppi) hjälper ungdomar med missbruksproblem, Internetberoende eller spelberoende.
Nuppi ger också stöd till ungdomar som oroar sig för rusmedelsbruket hos någon närstående person.
Läs mer: Missbruksproblem.
linkkiVanda stad:
Hjälp med missbruksproblemfinska _ svenska _ engelska
linkkiVanda stad:
Information om vård av drogproblemfinska _ svenska _ engelska
Hjälp med penningspelproblemfinska
Hjälp för ungafinska _ svenska _ engelska
Dödsfall
I Vanda finns fyra begravningsplatser som tillhör de evangelisk-lutherska församlingarna.
I Furumo i Vanda finns dessutom Vandas och Helsingfors gemensamma begravningsplats för avlidna personer som inte har varit medlemmar i något religionssamfund.
Information om begravning får du på Vanda församlingars gravkontor (Vantaan seurakuntien hautaustoimisto) och vid privata begravningsbyråer (hautaustoimisto).
Vanda församlingars gravkontor
Prästgårdsgränden 5
Tfn (09) 8306 220
Om din närstående avlider plötsligt, kan du få hjälp med att återhämta dig från den chockartade upplevelsen och stöd i att klara dig efter förlusten av Vandas social- och krisjour (sosiaali- ja kriisipäivystys).
Jouren har öppet varje dag dygnet runt.
Social- och krisjouren
Tfn (09) 8392 4005
Läs mer: Död
linkkiVanda kyrkliga samfällighet:
Begravningsplatserfinska
linkkiHelsingfors kyrkliga samfällighet:
Konfessionslös begravningsplatsfinska
linkkiFinlands Begravningbyråers Förbund:
Begravningsbyråerfinska
När en närstående har avliditfinska _ svenska _ engelska
linkkiVanda stad:
Social- och krisjourenfinska _ svenska _ engelska
Äktenskap
Skilsmässa
Barnets födelse
Vård av barn
Problem i familjen
Äktenskap
Före äktenskapet ska du skriftligt begära hindersprövning (avioliiton esteiden tutkiminen).
Hindersprövningen görs på magistraten (maistraatti).
Du kan begära hindersprövning på vilken magistrat som helst.
Mer information hittar du på magistratens webbplats.
Också borgerliga vigslar förrättas på magistraten.
Konvaljvägen 15, PB 112
01301 Vanda
Läs mer: Äktenskap.
Anhållan om prövning av hinder mot äktenskapfinska _ svenska
Ingående av äktenskapfinska _ svenska _ engelska
linkkiVanda församlingar:
Information om kyrklig vigselfinska _ svenska _ engelska
linkkiHelsingfors ortodoxa församling:
Information om ortodox vigselfinska _ ryska
Skilsmässa
Kvinnan eller mannen kan lämna in skilsmässoansökan i Vanda tingsrätts kansli.
Makarna kan ansöka om skilsmässa tillsammans eller också kan den ena maken göra det ensam.
Ansökan kan lämnas till tingsrättens kansli eller skickas dit per post, fax eller via e-post.
Tfn 029 56 45200
Läs mer: Skilsmässa.
linkkiVanda stad:
Information om skilsmässafinska _ engelska
Att ansöka om skilsmässafinska _ svenska _ engelska
Om du har barn och ska skilja dig tar du kontakt med barnatillsyningsmannen (lastenvalvoja) vid Vanda stad.
Socialväsendet bekräftar ett avtal om barnens boende, vårdnad, umgängesrätt och underhållsbidrag.
Barnatillsyningsmännen ger även råd till föräldrar som ska skiljas.
Kontaktuppgifterna till barnatillsyningsmannen hittar du på Vanda stads webbplats.
Läs mer:
Barn vid skilsmässa.
linkkiVanda stad:
Kontaktuppgifter till barnatillsyningsmännenfinska _ svenska _ engelska
Barnets födelse
Uppgifterna om barnets födelse skickas från sjukhuset till befolkningsdataregistret i Finland.
Du ska meddela barnets namn, modersmål och andra erforderliga uppgifter till magistraten (Maistraatti) med en separat blankett som skickas hem till dig.
Du kan läsa mer om registrering av barnets födelse, faderskapserkännande och vårdnaden om barnet på InfoFinlands sida: När ett barn föds i Finland.
Vård av barn
Dagvård
På InfoFinlands sida Utbildning i Vanda hittar du information om dagvård för barn i Vanda.
Hemvårdsstöd
Om du tar hand om ett under treårigt barn, kan du få hemvårdsstöd (kotihoidon tuki).
Du ansöker om hemvårdsstödet hos FPA.
Vanda stad betalar dessutom ett kommuntillägg till hemvårdsstödet för barn till de familjer som vårdar ett under 1 ½-årigt barn i hemmet.
Du behöver inte ansöka separat om stödet, utan FPA betalar ut Vandatillägget (Vantaa-lisä) med hemvårdsstödet.
Information om hemvårdsstödfinska _ svenska _ engelska
linkkiVanda stad:
Information om hemvårdsstödets kommuntilläggfinska _ svenska _ engelska
Öppna daghem och invånarparker
Öppna daghem (avoin päiväkoti) är avsedda för barn under skolåldern och de föräldrar och vårdare som tar hand om dem.
Invånarparker (asukaspuistot) är avsedda för barn i alla åldrar och deras föräldrar eller vårdare.
Små barn kan delta i verksamheten tillsammans med sin förälder eller vårdare.
Verksamheten i öppna daghem och invånarparker är kostnadsfri och du behöver inte anmäla dig på förhand.
I verksamheten ingår lek och ledda aktiviteter, till exempel musik, motion och utflykter.
linkkiVanda stad:
Parker för invånare och öppna daghemfinska _ svenska _ engelska
Klubbar
Vanda stad ordnar även klubbar (kerho) för 2,5–5-åriga barn som vårdas i hemmet.
Klubbarna är avgiftsfria.
I klubben lär sig barnet tala finska, fungera i en grupp och där kan barnet träffa andra barn.
Till klubben ansöker du om plats med samma ansökan om småbarnsfostran (varhaiskasvatushakemus), med vilken du även ansöker om dagvårdsplats.
linkkiVanda stad:
Klubbverksamhetfinska _ svenska _ engelska
Barnpassningsservice för barn
Om du vårdar ditt barn i hemmet och behöver tillfälligt en vårdplats för barnet, till exempel när du ska sköta ärenden, kan du kontakta barnpassningsservicen (hoitoapupalvelu).
Barnpassningen är avgiftsbelagd.
linkkiVanda stad:
Barnpassningsservice för barnfinska _ engelska
Tillfällig barnpassning
Om du behöver tillfällig barnpassning i hemmet, kan du kontakta Mannerheims Barnskyddsförbund eller Väestöliitto.
Den tillfälliga barnpassningshjälpen är avgiftsbelagd.
Läs mer: Vård av barnet
linkkiMannerheims barnskyddsförbund:
Barnvaktshjälpfinska _ engelska
linkkiVanda stad:
Hjälp i hemmet för barnfamiljer(pdf, 500 kb)finska _ engelska
Problem i familjen
Om du misstänker att ditt barn eller din ungdom behöver barnskyddets (lastensuojelu) hjälp, ska du kontakta en socialarbetare.
Tfn växeln 09 83 911
mån–fre kl. 8.15–16.00
Kvällar och helger
Social- och krisjouren
tfn 09 8392 4005
linkkiVanda stad:
Barnskyddsanmälanfinska _ engelska
På InfoFinlands sida Problematiska situationer i Vanda hittar du information om var någonstans i Vanda det finns hjälp att få till barns och ungas problem.
Information om barns och ungas problem finns även på InfoFinlands sidor Barns och ungas problem och Barnskydd.
På InfoFinlands sida Problem i äktenskap och parförhållande finns information om var man kan få hjälp med problem i parförhållanden.
Äktenskap
Skilsmässa
Barnets födelse
Vård av barn
Problem i familjen
Äldre människor
Äktenskap
Före äktenskapet ska du skriftligt begära hindersprövning (avioliiton esteiden tutkiminen).
Hindersprövningen görs på magistraten (maistraatti).
Du kan begära hindersprövning på vilken magistrat som helst.
Mer information hittar du på magistratens webbplats.
Också borgerliga vigslar förrättas på magistraten.
Konvaljvägen 15, PB 112
01301 Vanda
Läs mer: Äktenskap.
Anhållan om prövning av hinder mot äktenskapfinska _ svenska
Ingående av äktenskapfinska _ svenska _ engelska
linkkiVanda församlingar:
Information om kyrklig vigselfinska _ svenska _ engelska
linkkiHelsingfors ortodoxa församling:
Information om ortodox vigselfinska _ ryska
Skilsmässa
Kvinnan eller mannen kan lämna in skilsmässoansökan i Vanda tingsrätts kansli.
Makarna kan ansöka om skilsmässa tillsammans eller också kan den ena maken göra det ensam.
Ansökan kan lämnas till tingsrättens kansli eller skickas dit per post, fax eller via e-post.
Tfn 029 56 45200
Läs mer: Skilsmässa.
linkkiVanda stad:
Information om skilsmässafinska _ engelska
Att ansöka om skilsmässafinska _ svenska _ engelska
Om du har barn och ska skilja dig tar du kontakt med barnatillsyningsmannen (lastenvalvoja) vid Vanda stad.
Socialväsendet bekräftar ett avtal om barnens boende, vårdnad, umgängesrätt och underhållsbidrag.
Barnatillsyningsmännen ger även råd till föräldrar som ska skiljas.
Kontaktuppgifterna till barnatillsyningsmannen hittar du på Vanda stads webbplats.
Läs mer:
Barn vid skilsmässa.
linkkiVanda stad:
Kontaktuppgifter till barnatillsyningsmännenfinska _ svenska _ engelska
Barnets födelse
Uppgifterna om barnets födelse skickas från sjukhuset till befolkningsdataregistret i Finland.
Du ska meddela barnets namn, modersmål och andra erforderliga uppgifter till magistraten (Maistraatti) med en separat blankett som skickas hem till dig.
Du kan läsa mer om registrering av barnets födelse, faderskapserkännande och vårdnaden om barnet på InfoFinlands sida: När ett barn föds i Finland.
Vård av barn
Dagvård
På InfoFinlands sida Utbildning i Vanda hittar du information om dagvård för barn i Vanda.
Hemvårdsstöd
Om du tar hand om ett under treårigt barn, kan du få hemvårdsstöd (kotihoidon tuki).
Du ansöker om hemvårdsstödet hos FPA.
Vanda stad betalar dessutom ett kommuntillägg till hemvårdsstödet för barn till de familjer som vårdar ett under 1 ½-årigt barn i hemmet.
Du behöver inte ansöka separat om stödet, utan FPA betalar ut Vandatillägget (Vantaa-lisä) med hemvårdsstödet.
Information om hemvårdsstödfinska _ svenska _ engelska
linkkiVanda stad:
Information om hemvårdsstödets kommuntilläggfinska _ svenska _ engelska
Öppna daghem och invånarparker
Öppna daghem (avoin päiväkoti) är avsedda för barn under skolåldern och de föräldrar och vårdare som tar hand om dem.
Invånarparker (asukaspuistot) är avsedda för barn i alla åldrar och deras föräldrar eller vårdare.
Små barn kan delta i verksamheten tillsammans med sin förälder eller vårdare.
Verksamheten i öppna daghem och invånarparker är kostnadsfri och du behöver inte anmäla dig på förhand.
I verksamheten ingår lek och ledda aktiviteter, till exempel musik, motion och utflykter.
linkkiVanda stad:
Parker för invånare och öppna daghemfinska _ svenska _ engelska
Klubbar
Vanda stad ordnar även klubbar (kerho) för 2,5–5-åriga barn som vårdas i hemmet.
Klubbarna är avgiftsfria.
I klubben lär sig barnet tala finska, fungera i en grupp och där kan barnet träffa andra barn.
Till klubben ansöker du om plats med samma ansökan om småbarnsfostran (varhaiskasvatushakemus), med vilken du även ansöker om dagvårdsplats.
linkkiVanda stad:
Klubbverksamhetfinska _ svenska _ engelska
Barnpassningsservice för barn
Om du vårdar ditt barn i hemmet och behöver tillfälligt en vårdplats för barnet, till exempel när du ska sköta ärenden, kan du kontakta barnpassningsservicen (hoitoapupalvelu).
Barnpassningen är avgiftsbelagd.
linkkiVanda stad:
Barnpassningsservice för barnfinska _ engelska
Tillfällig barnpassning
Om du behöver tillfällig barnpassning i hemmet, kan du kontakta Mannerheims Barnskyddsförbund eller Väestöliitto.
Den tillfälliga barnpassningshjälpen är avgiftsbelagd.
Läs mer: Vård av barnet
linkkiMannerheims barnskyddsförbund:
Barnvaktshjälpfinska _ engelska
linkkiVanda stad:
Hjälp i hemmet för barnfamiljer(pdf, 500 kb)finska _ engelska
Problem i familjen
Om du misstänker att ditt barn eller din ungdom behöver barnskyddets (lastensuojelu) hjälp, ska du kontakta en socialarbetare.
Tfn växeln 09 83 911
mån–fre kl. 8.15–16.00
Kvällar och helger
Social- och krisjouren
tfn 09 8392 4005
linkkiVanda stad:
Barnskyddsanmälanfinska _ engelska
På InfoFinlands sida Problematiska situationer i Vanda hittar du information om var någonstans i Vanda det finns hjälp att få till barns och ungas problem.
Information om barns och ungas problem finns även på InfoFinlands sidor Barns och ungas problem och Barnskydd.
På InfoFinlands sida Problem i äktenskap och parförhållande finns information om var man kan få hjälp med problem i parförhållanden.
Äldre människor
I Vanda finns tjänster som är särskilt avsedda för äldre.
Du får information om dem vid seniorrådgivningen.
Seniorrådgivningen Tfn: 09 8392 4202
När du tar hand om en anhörig i hemmet
När en familjemedlem behöver kontinuerlig hjälp och vården är både bindande och krävande, finns det möjlighet att få stöd för närståendevård av kommunen.
Seniorrådgivningen bedömer behovet av anhörigvård för en äldre person.
Läs mer: Äldre människor.
linkkiVanda stad:
Seniorrådgivningenfinska _ svenska _ engelska
Äktenskap
Skilsmässa
Barnets födelse
Vård av barn
Problem i familjen
Äldre människor
Äktenskap
Före äktenskapet ska du skriftligt begära hindersprövning (avioliiton esteiden tutkiminen).
Hindersprövningen görs på magistraten (maistraatti).
Du kan begära hindersprövning på vilken magistrat som helst.
Mer information hittar du på magistratens webbplats.
Också borgerliga vigslar förrättas på magistraten.
Konvaljvägen 15, PB 112
01301 Vanda
Läs mer: Äktenskap.
Anhållan om prövning av hinder mot äktenskapfinska _ svenska _ engelska
Ingående av äktenskapfinska _ svenska _ engelska
linkkiVanda församlingar:
Information om kyrklig vigselfinska _ svenska _ engelska
linkkiHelsingfors ortodoxa församling:
Information om ortodox vigselfinska _ ryska
Skilsmässa
Kvinnan eller mannen kan lämna in skilsmässoansökan i Vanda tingsrätts kansli.
Makarna kan ansöka om skilsmässa tillsammans eller också kan den ena maken göra det ensam.
Ansökan kan lämnas till tingsrättens kansli eller skickas dit per post, fax eller via e-post.
Tfn 029 56 45200
Läs mer: Skilsmässa.
linkkiVanda stad:
Information om skilsmässafinska _ engelska
Att ansöka om skilsmässafinska _ svenska _ engelska
Om du har barn och ska skilja dig tar du kontakt med barnatillsyningsmannen (lastenvalvoja) vid Vanda stad.
Socialväsendet bekräftar ett avtal om barnens boende, vårdnad, umgängesrätt och underhållsbidrag.
Barnatillsyningsmännen ger även råd till föräldrar som ska skiljas.
Kontaktuppgifterna till barnatillsyningsmannen hittar du på Vanda stads webbplats.
Läs mer:
Barn vid skilsmässa.
linkkiVanda stad:
Kontaktuppgifter till barnatillsyningsmännenfinska _ svenska _ engelska
Barnets födelse
Uppgifterna om barnets födelse skickas från sjukhuset till befolkningsdataregistret i Finland.
Du ska meddela barnets namn, modersmål och andra erforderliga uppgifter till magistraten (Maistraatti) med en separat blankett som skickas hem till dig.
Du kan läsa mer om registrering av barnets födelse, faderskapserkännande och vårdnaden om barnet på InfoFinlands sida: När ett barn föds i Finland.
Vård av barn
Dagvård
På InfoFinlands sida Utbildning i Vanda hittar du information om dagvård för barn i Vanda.
Hemvårdsstöd
Om du tar hand om ett under treårigt barn, kan du få hemvårdsstöd (kotihoidon tuki).
Du ansöker om hemvårdsstödet hos FPA.
Vanda stad betalar dessutom ett kommuntillägg till hemvårdsstödet för barn till de familjer som vårdar ett under 1 ½-årigt barn i hemmet.
Du behöver inte ansöka separat om stödet, utan FPA betalar ut Vandatillägget (Vantaa-lisä) med hemvårdsstödet.
Information om hemvårdsstödfinska _ svenska _ engelska
linkkiVanda stad:
Information om hemvårdsstödets kommuntilläggfinska _ svenska _ engelska
Öppna daghem och invånarparker
Öppna daghem (avoin päiväkoti) är avsedda för barn under skolåldern och de föräldrar och vårdare som tar hand om dem.
Invånarparker (asukaspuistot) är avsedda för barn i alla åldrar och deras föräldrar eller vårdare.
Små barn kan delta i verksamheten tillsammans med sin förälder eller vårdare.
Verksamheten i öppna daghem och invånarparker är kostnadsfri och du behöver inte anmäla dig på förhand.
I verksamheten ingår lek och ledda aktiviteter, till exempel musik, motion och utflykter.
linkkiVanda stad:
Parker för invånare och öppna daghemfinska _ svenska _ engelska
Klubbar
Vanda stad ordnar även klubbar (kerho) för 2,5–5-åriga barn som vårdas i hemmet.
Klubbarna är avgiftsfria.
I klubben lär sig barnet tala finska, fungera i en grupp och där kan barnet träffa andra barn.
Till klubben ansöker du om plats med samma ansökan om småbarnsfostran (varhaiskasvatushakemus), med vilken du även ansöker om dagvårdsplats.
linkkiVanda stad:
Klubbverksamhetfinska _ svenska _ engelska
Barnpassningsservice för barn
Om du vårdar ditt barn i hemmet och behöver tillfälligt en vårdplats för barnet, till exempel när du ska sköta ärenden, kan du kontakta barnpassningsservicen (hoitoapupalvelu).
Barnpassningen är avgiftsbelagd.
linkkiVanda stad:
Barnpassningsservice för barnfinska _ engelska
Tillfällig barnpassning
Om du behöver tillfällig barnpassning i hemmet, kan du kontakta Mannerheims Barnskyddsförbund eller Väestöliitto.
Den tillfälliga barnpassningshjälpen är avgiftsbelagd.
Läs mer: Vård av barnet
linkkiMannerheims barnskyddsförbund:
Barnvaktshjälpfinska _ engelska
linkkiVanda stad:
Hjälp i hemmet för barnfamiljer(pdf, 500 kb)finska _ engelska
Problem i familjen
Om du misstänker att ditt barn eller din ungdom behöver barnskyddets (lastensuojelu) hjälp, ska du kontakta en socialarbetare.
Tfn växeln 09 83 911
mån–fre kl. 8.15–16.00
Kvällar och helger
Social- och krisjouren
tfn 09 8392 4005
linkkiVanda stad:
Barnskyddsanmälanfinska _ engelska
På InfoFinlands sida Problematiska situationer i Vanda hittar du information om var någonstans i Vanda det finns hjälp att få till barns och ungas problem.
Information om barns och ungas problem finns även på InfoFinlands sidor Barns och ungas problem och Barnskydd.
På InfoFinlands sida Problem i äktenskap och parförhållande finns information om var man kan få hjälp med problem i parförhållanden.
Äldre människor
I Vanda finns tjänster som är särskilt avsedda för äldre.
Du får information om dem vid seniorrådgivningen.
Seniorrådgivningen Tfn: 09 8392 4202
När du tar hand om en anhörig i hemmet
När en familjemedlem behöver kontinuerlig hjälp och vården är både bindande och krävande, finns det möjlighet att få stöd för närståendevård av kommunen.
Seniorrådgivningen bedömer behovet av anhörigvård för en äldre person.
Läs mer: Äldre människor.
linkkiVanda stad:
Seniorrådgivningenfinska _ svenska _ engelska
Hälsotjänster i Vanda
Privata hälsotjänster
Barns hälsa
Äldre människors hälsa
Tandvård
Mental hälsa
Sexuell hälsa
När du väntar barn
Handikappade
Hälsotjänsterna i Vanda
Om du behöver information om hälsotjänsterna, kan du ringa hälsorådgivningstelefonen: Tfn (09) 839 10023, mån-fre kl. 8–16.
Via tjänsten kan du också fråga om anvisningar för vård av sjukdomar.
Du kan tala finska, svenska eller engelska.
Läs mer: Hälsa.
linkkiVanda stad:
Information om hälsorådgivningfinska _ svenska _ engelska
Offentliga hälsovårdstjänster
Om du har din hemkommun i Vanda, kan du utnyttja de offentliga hälsovårdstjänsterna.
Offentliga hälsovårdstjänster tillhandahålls till exempel vid hälsostationer, tandkliniker, rådgivningsbyråer och sjukhus.
Om du insjuknar plötsligt eller om du råkar ut för en olycka, får du akut sjukvård även om din hemkommun inte är Vanda.
I Vanda finns sju hälsostationer (terveysasema) som tillhandahåller offentliga hälsovårdstjänster.
Hälsostationerna har öppet vardagar kl. 8.00–16.00.
Hälsostationerna når du genom att ringa till respektive hälsostations eget telefonnummer eller hälsorådgivningens telefonnummer (09) 839 10023 och väljer din hälsostation med hjälpa av knappsatsen.
Om du behöver akut vård samma dag, ska du ringa hälsostationen direkt då den öppnar.
Hälsostationernas adresser:
Håkansböle hälsostation, Galoppbrinken 4
Korso hälsostation, Fjällrävsstigen 6
Västerkulla hälsostation, Kägelgränden 1
Myrbacka hälsostation, Jönsasvägen 4
Dickursby hälsostation, Konvaljvägen 11
Närmare information hittar du på hälsostationernas egna webbplatser.
linkkiVanda stad:
Hälsostationernafinska _ svenska _ engelska
Privata hälsotjänster
I Vanda finns flera läkarstationer som erbjuder privata hälsovårdstjänster.
Du kan gå till en privat läkarstation även om du inte har rätt att använda den offentliga hälsovårdens tjänster i Finland.
På en privat läkarstation måste du betala samtliga kostnader själv.
I vissa fall ersätter Kela en liten del av kostnaderna för privat sjukvård.
Privat läkarstationfinska _ svenska _ engelska
Privat läkarstationfinska _ svenska _ engelska _ ryska
Privat läkarstationfinska _ svenska _ engelska
linkkiAava:
Privat läkarstationfinska _ svenska _ engelska
Läkemedel
Information om köp av läkemedel hittar du på InfoFinlands sida Läkemedel.
linkkiApotekareförbundet:
Apotekens kontaktuppgifterfinska
Hälsovård för papperslösa
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärhälsovård.
Tjänsterna vid Global Clinic är avgiftsfria för kunderna.
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter.
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
Telefonnumret till Helsingfors Global Clinicin är 044 948 1698.
En sjuksköterska eller läkare svarar i telefonen.
Läs mer: Hälsovårdstjänster i Finland.
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
På kvällar, helger och storhelger är hälsostationerna stängda.
Då vårdas akuta sjukfall och olycksfall på jourmottagningen (päivystys).
Jourmottagningen är öppen alla dagar dygnet runt
I Vanda finns jourmottagningen på Pejas sjukhus (Peijaksen sairaala).
Adress:
Sjukhusgatan 1
Tfn 116 117
Om du blir akut sjuk, kan du även besöka någon annan jourmottagning i huvudstadsregionen.
Mer information om jourmottagningarna hittar du på Vanda stads webbplats om hälsovårdstjänster.
I nödsituationer ringer du det allmänna nödnumret 112.
Läs mer: Hälsovårdstjänster i Finland.
linkkiVanda stad:
Jourmottagningarfinska _ svenska _ engelska
Barns hälsa
I hälsovården av barn under skolåldern får man hjälp av rådgivningsbyråerna (neuvola).
Där kan du fråga om råd och få stöd i föräldraskapet och fostran av barn.
På rådgivningsbyrån följs barnets hälsa, tillväxt och utveckling upp och där ges även vaccinationerna.
Kontaktuppgifterna till rådgivningsbyråerna hittar du på Vanda webbplats.
Via rådgivningsbyråernas telefontjänst kan du boka tid på rådgivningsbyrån och fråga hälsovårdaren om råd beträffande graviditet och barns hälsa.
Numret till telefontjänsten är (09) 8392 5900.
Den är öppen mån-tors kl. 8–15 och fre kl. 8–13.
Skolhälsovården har hand om skolbarns hälsa.
Mer information hittar du på Vanda stads webbplats.
Om ett barn blir akut sjukt, ska du ta kontakt med hälsostationen eller jourmottagningen.
I nödsituationer ringer du det allmänna nödnumret 112.
Läs mer: Barns hälsa.
linkkiVanda stad:
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad:
Tidsbokning och rådgivningfinska _ svenska _ engelska
linkkiVanda stad:
Information om skolhälsovårdenfinska _ svenska _ engelska
linkkiVanda stad:
Hälsostationernafinska _ svenska _ engelska
linkkiVanda stad:
Jourmottagningarfinska _ svenska _ engelska
Äldre människors hälsa
Äldre människor använder samma hälsovårdstjänster som alla andra.
Dessutom finns det i Vanda särskilda tjänster för äldre som du får information om via seniorrådgivningen (seniorineuvonta).
Tfn: (09) 8392 4202
Mer information om tjänsterna för äldre hittar du på Vanda stads webbplats.
Läs mer: Äldre människors hälsa och Äldre människor.
linkkiVanda stad:
Seniorrådgivningenfinska _ svenska _ engelska
linkkiVanda stad:
Information om tjänster för äldrefinska _ svenska _ engelska
linkkiVanda stad:
Serviceguide för seniorer(pdf, 1 MB)finska
När du tar hand om en anhörig i hemmet
När en familjemedlem behöver kontinuerlig hjälp och vården är både bindande och krävande, finns det möjlighet att få stöd för närståendevård av kommunen.
Behovet av närståendevård bedöms inom seniorrådgivningen.
Tfn: (09) 8392 4202
Behovet av närståendevård för personer under 65 år bedöms inom handikapprådgivningen.
Tfn: (09) 8392 4682
linkkiVanda stad:
Stöd för närståendevårdfinska _ svenska
Tandvård
Offentlig tandvård
Tidsbokningsnumret till Vanda tandvård (hammashoito) är (09) 8393 5300.
Tidsbokningen kan du ringa:
Mån-tors 7.30–15
Fredagar och storhelgsaftnar 7.30–14.
Om ditt ärende inte är brådskande, ring efter kl. 10.00.
Om tjänsten är hårt belastad, kan du lämna ett meddelande om att bli uppringd vid ett senare tillfälle.
Om du behöver akut tandvård på en vardag, ska du ringa tidsbokningen så fort den öppnar.
linkkiVanda stad:
Information om tandvårdenfinska _ svenska _ engelska
linkkiVanda stad:
Tandklinikerfinska _ svenska
Tandvårdens jourmottagning
Under kvällar och veckoslut finns tandvårdsjouren (hammashoidon päivystys) vid Haartmanska sjukhuset i Helsingfors.
Tfn (09) 310 49999.
Tandvårdens nattjour (hammashoidon yöpäivystys) finns på Tölö sjukhus olycksfallsstation.
Tölö sjukhus olycksfallsstation, Oral och käkkirurgisk jourmottagning
Tfn 040 621 5699
Tandvårdens jourmottagning kvällar och veckoslutfinska _ svenska _ engelska
Barns tandvård
Om tandvården för barn under skolåldern får du information på barnrådgivningen (lastenneuvola) och vid tandklinikerna (hammashoitola).
Barn under 17 år kallas till tandkliniken för undersökning med cirka två års mellanrum.
linkkiVanda stad:
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad:
Information om tandvården för skolbarnfinska
Privata tandvårdstjänster
I Vanda finns också privata tandläkare.
Om du inte har rätt att använda de offentliga hälsovårdstjänsterna, kan du söka dig till en privat tandläkare.
Hos en privat tandläkare måste du betala samtliga kostnader själv.
I vissa fall ersätter Kela en liten del av kostnaderna för privat tandvård.
Läs mer: Tandvård.
Sök tandläkarefinska
Mental hälsa
Om du behöver psykisk hjälp eller stöd, ska du kontakta din hälsostation (terveysasema).
På hälsostationen behandlas de vanligaste psykiska problemen.
Från hälsostationen kan du remitteras vidare exempelvis till depressionsskötare.
Om hälsostationen inte har öppet och situationen är akut, ska du kontakta samjouren vid Pejas sjukhus (Peijaksen sairaalan yhteispäivystys).
Sjukhusgatan 1
Tfn (09) 4716 7060
Om du behöver omedelbar krishjälp, kan du också ta kontakt med social- och krisjouren.
Den har öppet dygnet runt.
Social- och krisjouren
Tfn (09) 8392 4005
Läs mer: Mental hälsa.
linkkiVanda stad:
Information om mentalvårdstjänsternafinska _ svenska _ engelska
linkkiVanda stad:
Hälsostationernafinska _ svenska _ engelska
linkkiVanda stad:
Jourmottagningarfinska _ svenska _ engelska
linkkiVanda stad:
Social- och krisjourenfinska _ svenska _ engelska
Sexuell hälsa
Om du vill har information om graviditetsprevention, abort, sexuell hälsa och könssjukdomar, kan du kontakta preventivmedels- och familjeplaneringsrådgivningen (ehkäisy- ja perhesuunnitteluneuvola).
Preventivmedels- och familjeplaneringsrådgivningarna betjänar kvinnor och män i alla åldrar.
Du måste beställa tid vid rådgivningarna.
Besöken är avgiftsfria för kunderna.
Information om kontaktuppgifter finns på Vanda stads webbplats.
Boka en tid hos preventivmedelsrådgivningens läkare eller hälsovårdare om du behöver preventivmedel (raskauden ehkäisy) eller om du överväger abort (abortti).
Boka en tid hos hälsostationens allmänläkare om du till exempel har problem med blödningar eller smärtor i underlivet.
Vid hälsostationerna vårdas även könssjukdomar (sukupuolitauti).
Vandabor kan även besöka polikliniken för könssjukdomar i Helsingfors.
linkkiVanda stad:
Rådgivningarna för familjeplaneringfinska _ svenska.
linkkiVanda stad:
Hälsostationernafinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Polikliniken för könssjukdomarfinska _ svenska _ engelska
När du väntar barn
Vid mödrarådgivningen (äitiysneuvola) följs moderns, fostrets och hela familjens hälsotillstånd under graviditeten.
Kontakta rådgivningsbyrån (neuvola) när du upptäcker att du är gravid.
Rådgivningarnas telefontjänst
mån-tors kl. 8–15 och fre kl. 8–13
Via rådgivningsbyråernas telefontjänst kan du boka tid på rådgivningsbyrån och fråga hälsovårdaren om råd beträffande graviditet och förlossning.
Mer information om graviditet och förlossning hittar du på Vanda stads mödra- och barnrådgivning på Internet (Nettineuvola).
Läs mer: När du väntar barn.
linkkiVanda stad:
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad:
Rådgivningarna för familjeplaneringfinska _ svenska
linkkiVanda stad:
Förlossningen
Läs mer: Förlossning.
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Förlossningfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Handikappade
Du kan få tjänster för handikappade (vammaispalvelut) om du eller en närstående till dig har en invaliditet eller en sjukdom som orsakar långvariga, betydande svårigheter att klara sig hemma och i livet utanför hemmet.
Tjänster för handikappade är till exempel personlig assistans, serviceboende, färdtjänst och ombyggnadsarbeten i bostaden.
Ta kontakt med handikapprådgivningen som utreder ditt behov av stöd, handledning och tjänster utifrån din situation.
Mån.-fre. kl. 9–15
Tfn: (09) 8392 4682
Läs mer: Handikappade personer.
linkkiVanda stad:
Information om handikapptjänsternafinska _ svenska _ engelska
Hälsotjänster i Vanda
Barns hälsa
Tandvård
Mental hälsa
Sexuell hälsa och prevention
Graviditet och förlossning
Handikappade
Hälsotjänsterna i Vanda
Det allmänna nödnumret är 112.
Ring nödnumret endast om det handlar om ett nödfall, till exempel en akut sjukdomsattack.
Om din hemkommun är Vanda kan du använda kommunens offentliga hälsovårdstjänster.
Offentliga hälsovårdstjänster tillhandahålls till exempel vid hälsostationer, tandkliniker, rådgivningsbyråer och sjukhus.
Om du insjuknar akut eller råkar ut för en olycka får du akut sjukvård även om din hemkommun inte är Vanda.
Om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna, kan du boka tid på en privat läkarstation.
Läs mer: Hälsovårdstjänster i Finland.
Offentliga hälsovårdstjänster
Telefonnumret till den gemensamma telefontjänsten för hälsostationerna i Vanda är 09 839 50 000.
Du kan ringa detta nummer om du behöver rådgivning i behandlingen av en sjukdom eller vill boka eller avboka en läkartid.
Tjänsten har öppet måndag till fredag kl. 8–16.
I Vanda finns sju hälsostationer som tillhandahåller offentliga hälsovårdstjänster.
På hälsostationerna finns läkarens, sjukskötarens och hälsovårdarens mottagningar.
Om du insjuknar akut kan du gå direkt till vilken som helst hälsostation.
Det är bäst att gå till hälsostationen direkt på morgonen.
Hälsostationerna har öppet vardagar kl. 8.00–16.00.
linkkiVanda stad:
Information om hälsorådgivningfinska _ svenska _ engelska
linkkiVanda stad:
Hälsostationernafinska _ svenska _ engelska
Privata hälsotjänster
I Vanda finns flera läkarstationer som erbjuder privata hälsovårdstjänster.
Du kan gå till en privat läkarstation även om du inte har rätt att använda den offentliga hälsovårdens tjänster i Finland.
På en privat läkarstation måste du betala samtliga kostnader själv.
I vissa fall ersätter Kela en liten del av kostnaderna för privat sjukvård.
Läs mer: Hälsovårdstjänster i Finland.
Privat läkarstationfinska _ svenska _ engelska
Privat läkarstationfinska _ svenska _ engelska _ ryska
Privat läkarstationfinska _ svenska _ engelska
linkkiAava:
Privat läkarstationfinska _ svenska _ engelska
Läkemedel
Information om köp av läkemedel hittar du på InfoFinlands sida Läkemedel.
linkkiApotekareförbundet:
Apotekens kontaktuppgifterfinska
Hälsovård för papperslösa
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärhälsovård.
Tjänsterna vid Global Clinic är avgiftsfria för kunderna.
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter.
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
Telefonnumret till Helsingfors Global Clinicin är 044 948 1698.
En sjuksköterska eller läkare svarar i telefonen.
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
På kvällar, helger och storhelger är hälsostationerna stängda.
Om du insjuknar akut eller råkar ut för en olycka och inte kan vänta tills hälsostationen öppnar, kontakta jourmottagningen.
I Vanda finns jourmottagningen på Pejas sjukhus (Peijaksen sairaala).
Adress:
Sjukhusgatan 1
Tfn 116 117
Om du blir akut sjuk, kan du även besöka någon annan jourmottagning i huvudstadsregionen.
Mer information om jourmottagningarna hittar du på Vanda stads webbplats om hälsovårdstjänster.
linkkiVanda stad:
Jourmottagningarfinska _ svenska _ engelska
Barns hälsa
I hälsovården av barn under skolåldern får man hjälp av rådgivningsbyråerna (neuvola).
Telefonnumret till rådgivningsbyråerna i Vanda är 09 8392 5900.
Du kan boka en tid på rådgivningen eller fråga om råd om du har frågor kring barnets hälsa.
Skolhälsovården har hand om skolbarns hälsa.
Mer information hittar du på Vanda stads webbplats.
Om ett barn insjuknar akut, ska du kontakta hälsostationen.
Hälsostationerna har öppet måndag till fredag kl. 8–16.
När hälsostationen har stängt ska du kontakta jourmottagningen vid Barnsjukhuset.
Jourmottagningen tar endast hand om barn med brådskande hjälpbehov.
Telefonnumret till jourmottagningen är 116 117.
Adress:
Barnsjukhuset
Stenbäcksgatan 9
Du kan även ta barnet till en privat läkarstation.
I Vanda finns många privata läkarstationer som även tar hand om barn.
Läs mer: Barns hälsa.
linkkiVanda stad:
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad:
Tidsbokning och rådgivningfinska _ svenska _ engelska
linkkiVanda stad:
Information om skolhälsovårdenfinska _ svenska _ engelska
linkkiVanda stad:
Hälsostationernafinska _ svenska _ engelska
linkkiVanda stad:
Jourmottagningarfinska _ svenska _ engelska
Tandvård
Offentlig tandvård
Tidsbokningsnumret till Vanda tandvård (hammashoito) är (09) 8393 5300.
Om du inte behöver brådskande tandvård, ring efter kl. 10.00.
Om du behöver brådskande tandvård, ska du ringa tidsbokningen så fort den öppnar kl. 7.30.
Mottagningen för brådskande vård finns vid Dickursby hälsostation måndag till fredag kl. 8–14.
linkkiVanda stad:
Information om tandvårdenfinska _ svenska _ engelska
linkkiVanda stad:
Tandklinikerfinska _ svenska
Tandvårdens jourmottagning
Under kvällar och veckoslut finns tandvårdsjouren (hammashoidon päivystys) vid Haartmanska sjukhuset i Helsingfors.
Telefonnumret är 09 471 71110.
Tidsbokningen har öppet vardagar kl. 14–21 och på veckoslut kl. 8–21.
Tandvårdens nattjour (hammashoidon yöpäivystys) finns på Tölö sjukhus olycksfallsstation.
Tölö sjukhus olycksfallsstation, Oral och käkkirurgisk jourmottagning
Tfn 040 621 5699
Tandvårdens jourmottagning kvällar och veckoslutfinska _ svenska _ engelska
Barns tandvård
Om tandvården för barn under skolåldern får du information på barnrådgivningen (lastenneuvola) och vid tandklinikerna (hammashoitola).
Barn under 17 år kallas till tandkliniken för undersökning med cirka två års mellanrum.
linkkiVanda stad:
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad:
Information om tandvården för skolbarnfinska
Privata tandvårdstjänster
I Vanda finns också privata tandläkare.
Om du inte har rätt att använda de offentliga hälsovårdstjänsterna, kan du söka dig till en privat tandläkare.
Hos en privat tandläkare måste du betala samtliga kostnader själv.
I vissa fall ersätter Kela en liten del av kostnaderna för privat tandvård.
Läs mer: Tandvård.
Sök tandläkarefinska
Mental hälsa
Om du behöver psykisk hjälp eller stöd, ska du kontakta din hälsostation (terveysasema).
På hälsostationen behandlas de vanligaste psykiska problemen.
Från hälsostationen kan du remitteras vidare exempelvis till depressionsskötare.
Om hälsostationen inte har öppet och situationen är akut, ska du kontakta samjouren vid Pejas sjukhus (Peijaksen sairaalan yhteispäivystys).
Sjukhusgatan 1
Tfn 116 117
Om du behöver omedelbar krishjälp, kan du också ta kontakt med social- och krisjouren.
Den har öppet dygnet runt.
Social- och krisjouren
Tfn (09) 8392 4005
Läs mer: Mental hälsa.
linkkiVanda stad:
Information om mentalvårdstjänsternafinska _ svenska _ engelska
linkkiVanda stad:
Hälsostationernafinska _ svenska _ engelska
linkkiVanda stad:
Jourmottagningarfinska _ svenska _ engelska
linkkiVanda stad:
Social- och krisjourenfinska _ svenska _ engelska
Sexuell hälsa och prevention
Om du behöver preventivmedel eller abort eller misstänker att du har en könssjukdom, kan du kontakta preventivmedels- och familjeplaneringsrådgivningen.
Du kan boka tid per telefon.
Numret är 09 839 50030.
Om du har en könssjukdom kan du även besöka polikliniken för könssjukdomar i Helsingfors eller en hälsostation.
Vanda erbjuder ungdomar under 20 år gratis preventivmedel.
Även unga vuxna under 24 år kan få gratis preventivmedel om de använder långvariga preventivmedel såsom spiral eller p-stav.
Läs mer: Sexuell hälsa och prevention.
linkkiVanda stad:
Rådgivningarna för familjeplaneringfinska _ svenska.
linkkiVanda stad:
Hälsostationernafinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Polikliniken för könssjukdomarfinska _ svenska _ engelska
Graviditet och förlossning
Vid mödrarådgivningen (äitiysneuvola) följs moderns, fostrets och hela familjens hälsotillstånd under graviditeten.
Kontakta rådgivningsbyrån (neuvola) när du upptäcker att du är gravid.
Rådgivningarnas telefontjänst
Via rådgivningsbyråernas telefontjänst kan du boka tid på rådgivningsbyrån och fråga hälsovårdaren om råd beträffande graviditet och förlossning.
Läs mer: Graviditet och förlossning och När ett barn föds i Finland.
linkkiVanda stad:
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad:
Rådgivningarna för familjeplaneringfinska _ svenska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Förlossningfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Handikappade
Du kan få tjänster för handikappade (vammaispalvelut) om du eller en närstående till dig har en invaliditet eller en sjukdom som orsakar långvariga, betydande svårigheter att klara sig hemma och i livet utanför hemmet.
Tjänster för handikappade är till exempel personlig assistans, serviceboende, färdtjänst och ombyggnadsarbeten i bostaden.
Ta kontakt med handikapprådgivningen som utreder ditt behov av stöd, handledning och tjänster utifrån din situation.
Mån.-fre. kl. 9–15
Tfn: (09) 8392 4682
Läs mer: Handikappade personer.
linkkiVanda stad:
Information om handikapptjänsternafinska _ svenska _ engelska
Hälsotjänster i Vanda
Barns hälsa
Tandvård
Mental hälsa
Sexuell hälsa och prevention
Graviditet och förlossning
Handikappade
Hälsotjänsterna i Vanda
Det allmänna nödnumret är 112.
Ring nödnumret endast om det handlar om ett nödfall, till exempel en akut sjukdomsattack.
Om din hemkommun är Vanda kan du använda kommunens offentliga hälsovårdstjänster.
Offentliga hälsovårdstjänster tillhandahålls till exempel vid hälsostationer, tandkliniker, rådgivningsbyråer och sjukhus.
Om du insjuknar akut eller råkar ut för en olycka får du akut sjukvård även om din hemkommun inte är Vanda.
Om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna, kan du boka tid på en privat läkarstation.
Läs mer: Hälsovårdstjänster i Finland.
Offentliga hälsovårdstjänster
Telefonnumret till den gemensamma telefontjänsten för hälsostationerna i Vanda är 09 839 50 000.
Du kan ringa detta nummer om du behöver rådgivning i behandlingen av en sjukdom eller vill boka eller avboka en läkartid.
Tjänsten har öppet måndag till fredag kl. 8–16.
I Vanda finns sju hälsostationer som tillhandahåller offentliga hälsovårdstjänster.
På hälsostationerna finns läkarens, sjukskötarens och hälsovårdarens mottagningar.
Om du insjuknar akut kan du gå direkt till vilken som helst hälsostation.
Det är bäst att gå till hälsostationen direkt på morgonen.
Hälsostationerna har öppet vardagar kl. 8.00–16.00.
linkkiVanda stad:
Information om hälsorådgivningfinska _ svenska _ engelska
linkkiVanda stad:
Hälsostationernafinska _ svenska _ engelska
Privata hälsotjänster
I Vanda finns flera läkarstationer som erbjuder privata hälsovårdstjänster.
Du kan gå till en privat läkarstation även om du inte har rätt att använda den offentliga hälsovårdens tjänster i Finland.
På en privat läkarstation måste du betala samtliga kostnader själv.
I vissa fall ersätter Kela en liten del av kostnaderna för privat sjukvård.
Läs mer: Hälsovårdstjänster i Finland.
Privat läkarstationfinska _ svenska _ engelska
Privat läkarstationfinska _ svenska _ engelska _ ryska
Privat läkarstationfinska _ svenska _ engelska
linkkiAava:
Privat läkarstationfinska _ svenska _ engelska
Läkemedel
Information om köp av läkemedel hittar du på InfoFinlands sida Läkemedel.
linkkiApotekareförbundet:
Apotekens kontaktuppgifterfinska
Hälsovård för papperslösa
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärhälsovård.
Tjänsterna vid Global Clinic är avgiftsfria för kunderna.
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter.
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
Telefonnumret till Helsingfors Global Clinicin är 044 948 1698.
En sjuksköterska eller läkare svarar i telefonen.
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
På kvällar, helger och storhelger är hälsostationerna stängda.
Om du insjuknar akut eller råkar ut för en olycka och inte kan vänta tills hälsostationen öppnar, kontakta jourmottagningen.
I Vanda finns jourmottagningen på Pejas sjukhus (Peijaksen sairaala).
Adress:
Sjukhusgatan 1
Tfn 116 117
Om du blir akut sjuk, kan du även besöka någon annan jourmottagning i huvudstadsregionen.
Mer information om jourmottagningarna hittar du på Vanda stads webbplats om hälsovårdstjänster.
linkkiVanda stad:
Jourmottagningarfinska _ svenska _ engelska
Barns hälsa
I hälsovården av barn under skolåldern får man hjälp av rådgivningsbyråerna (neuvola).
Telefonnumret till rådgivningsbyråerna i Vanda är 09 8392 5900.
Du kan boka en tid på rådgivningen eller fråga om råd om du har frågor kring barnets hälsa.
Skolhälsovården har hand om skolbarns hälsa.
Mer information hittar du på Vanda stads webbplats.
Om ett barn insjuknar akut, ska du kontakta hälsostationen.
Hälsostationerna har öppet måndag till fredag kl. 8–16.
När hälsostationen har stängt ska du kontakta jourmottagningen vid Barnsjukhuset.
Jourmottagningen tar endast hand om barn med brådskande hjälpbehov.
Telefonnumret till jourmottagningen är 116 117.
Adress:
Barnsjukhuset
Stenbäcksgatan 9
Du kan även ta barnet till en privat läkarstation.
I Vanda finns många privata läkarstationer som även tar hand om barn.
Läs mer: Barns hälsa.
linkkiVanda stad:
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad:
Tidsbokning och rådgivningfinska _ svenska _ engelska
linkkiVanda stad:
Information om skolhälsovårdenfinska _ svenska _ engelska
linkkiVanda stad:
Hälsostationernafinska _ svenska _ engelska
linkkiVanda stad:
Jourmottagningarfinska _ svenska _ engelska
Tandvård
Offentlig tandvård
Tidsbokningsnumret till Vanda tandvård (hammashoito) är (09) 8393 5300.
Om du inte behöver brådskande tandvård, ring efter kl. 10.00.
Om du behöver brådskande tandvård, ska du ringa tidsbokningen så fort den öppnar kl. 7.30.
Mottagningen för brådskande vård finns vid Dickursby hälsostation måndag till fredag kl. 8–14.
linkkiVanda stad:
Information om tandvårdenfinska _ svenska _ engelska
linkkiVanda stad:
Tandklinikerfinska _ svenska
Tandvårdens jourmottagning
Under kvällar och veckoslut finns tandvårdsjouren (hammashoidon päivystys) vid Haartmanska sjukhuset i Helsingfors.
Telefonnumret är 09 471 71110.
Tidsbokningen har öppet vardagar kl. 14–21 och på veckoslut kl. 8–21.
Tandvårdens nattjour (hammashoidon yöpäivystys) finns på Tölö sjukhus olycksfallsstation.
Tölö sjukhus olycksfallsstation, Oral och käkkirurgisk jourmottagning
Tfn 040 621 5699
Tandvårdens jourmottagning kvällar och veckoslutfinska _ svenska _ engelska
Barns tandvård
Om tandvården för barn under skolåldern får du information på barnrådgivningen (lastenneuvola) och vid tandklinikerna (hammashoitola).
Barn under 17 år kallas till tandkliniken för undersökning med cirka två års mellanrum.
linkkiVanda stad:
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad:
Information om tandvården för skolbarnfinska
Privata tandvårdstjänster
I Vanda finns också privata tandläkare.
Om du inte har rätt att använda de offentliga hälsovårdstjänsterna, kan du söka dig till en privat tandläkare.
Hos en privat tandläkare måste du betala samtliga kostnader själv.
I vissa fall ersätter Kela en liten del av kostnaderna för privat tandvård.
Läs mer: Tandvård.
Sök tandläkarefinska
Mental hälsa
Om du behöver psykisk hjälp eller stöd, ska du kontakta din hälsostation (terveysasema).
På hälsostationen behandlas de vanligaste psykiska problemen.
Från hälsostationen kan du remitteras vidare exempelvis till depressionsskötare.
Om hälsostationen inte har öppet och situationen är akut, ska du kontakta samjouren vid Pejas sjukhus (Peijaksen sairaalan yhteispäivystys).
Sjukhusgatan 1
Tfn 116 117
Om du behöver omedelbar krishjälp, kan du också ta kontakt med social- och krisjouren.
Den har öppet dygnet runt.
Social- och krisjouren
Tfn (09) 8392 4005
Läs mer: Mental hälsa.
linkkiVanda stad:
Information om mentalvårdstjänsternafinska _ svenska _ engelska
linkkiVanda stad:
Hälsostationernafinska _ svenska _ engelska
linkkiVanda stad:
Jourmottagningarfinska _ svenska _ engelska
linkkiVanda stad:
Social- och krisjourenfinska _ svenska _ engelska
Sexuell hälsa och prevention
Om du behöver preventivmedel eller abort eller misstänker att du har en könssjukdom, kan du kontakta preventivmedels- och familjeplaneringsrådgivningen.
Du kan boka tid per telefon.
Numret är 09 839 50030.
Om du har en könssjukdom kan du även besöka polikliniken för könssjukdomar i Helsingfors eller en hälsostation.
Vanda erbjuder ungdomar under 20 år gratis preventivmedel.
Även unga vuxna under 24 år kan få gratis preventivmedel om de använder långvariga preventivmedel såsom spiral eller p-stav.
Läs mer: Sexuell hälsa och prevention.
linkkiVanda stad:
Rådgivningarna för familjeplaneringfinska _ svenska.
linkkiVanda stad:
Hälsostationernafinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Polikliniken för könssjukdomarfinska _ svenska _ engelska
Graviditet och förlossning
Vid mödrarådgivningen (äitiysneuvola) följs moderns, fostrets och hela familjens hälsotillstånd under graviditeten.
Kontakta rådgivningsbyrån (neuvola) när du upptäcker att du är gravid.
Rådgivningarnas telefontjänst
Via rådgivningsbyråernas telefontjänst kan du boka tid på rådgivningsbyrån och fråga hälsovårdaren om råd beträffande graviditet och förlossning.
Läs mer: Graviditet och förlossning och När ett barn föds i Finland.
linkkiVanda stad:
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad:
Rådgivningarna för familjeplaneringfinska _ svenska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Förlossningfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Handikappade
Du kan få tjänster för handikappade (vammaispalvelut) om du eller en närstående till dig har en invaliditet eller en sjukdom som orsakar långvariga, betydande svårigheter att klara sig hemma och i livet utanför hemmet.
Tjänster för handikappade är till exempel personlig assistans, serviceboende, färdtjänst och ombyggnadsarbeten i bostaden.
Ta kontakt med handikapprådgivningen som utreder ditt behov av stöd, handledning och tjänster utifrån din situation.
Mån.-fre. kl. 9–15
Tfn: (09) 8392 4682
Läs mer: Handikappade personer.
linkkiVanda stad:
Information om handikapptjänsternafinska _ svenska _ engelska
Dagvård
Förskoleundervisning
Grundläggande utbildning
Yrkesutbildning
Gymnasium
Stöd och handledning för unga
Högskoleutbildning
Övriga studiemöjligheter
Dagvård
I Vanda finns både kommunala och privata daghem.
Kommunen övervakar också den privata dagvården.
I Vanda ges dagvård på finska, svenska, ryska och engelska.
Inom dagvården ges även undervisning i finska som andra språk.
Dagvård ordnas också inom familjedagvården och i gruppfamiljedaghem.
Man ska ansöka om dagvårdsplats för sitt barn minst fyra månader innan barnet ska börja i dagvården.
Du kan ansöka om plats i den kommunala dagvården via Internet eller med en pappersblankett.
För en elektronisk ansökan behöver du egna nätbankskoder eller en elektronisk legitimation.
Pappersblanketter kan hämtas till exempel vid Vandainfo eller daghemmen.
Privata dagvårdsplatser söks direkt på daghemmet.
Frågor kring dagvård och ansökan om dagvårdsplats kan du ställa till daghemsföreståndaren eller skicka till adressen varhaiskasvatus(at)vantaa.fi.
Vanligtvis ansöker man om dagvårdsplats i den egna kommunen.
Om familjen bor nära gränsen till Helsingfors eller Esbo, kan du också söka dagvårdsplats i grannkommunen.
Du ska ändå lämna in din ansökan i den egna kommunen.
Mer information hittar du via tjänsten Helsingforsregionen.fi.
Läs mer: Dagvård
linkkiVanda stad:
Privat dagvårdfinska _ svenska _ engelska
linkkiVanda stad:
Privat dagvårdfinska
linkkiVanda stad:
Ansökan om dagvårdsplatsfinska _ svenska _ engelska
linkkiVanda stad:
Elektronisk ansökningsblankett för dagvårdenfinska _ svenska _ engelska
Information om dagvården finska _ svenska _ engelska
Förskoleundervisning
Förskoleundervisning (esiopetus) ordnas i både kommunala och privata daghem samt i förskoleenheter i skolornas lokaler.
I Vanda kan man få förskoleundervisning på finska, svenska och engelska.
Du måste ansöka om plats i förskoleundervisningen.
Ansökan kan göras elektroniskt via stadens webbplats eller med en pappersblankett.
Ansökningstiden är i januari, men ansökan kan även lämnas in övriga tider, om familjen till exempel flyttar till Vanda mitt under året.
Förberedande undervisning tillhandahålls för invandrarbarn som inte har tillräckliga kunskaper i finska för att klara sig i förskoleundervisningen.
Den förberedande undervisningen är avsedd för 6-åriga barn med invandrarbakgrund.
Den ordnas i daghemmens förskolegrupper.
Daghemmet anvisar barnet till den förberedande undervisningen i samband med ansökningen till förskoleundervisningen.
Du hittar mer information om förskoleundervisningen, ansökning till förskoleundervisningen och om undervisning som förbereder för förskoleundervisning på Vanda stads (Vantaan kaupunki) webbplats.
Du kan även fråga om mer information på daghemmen.
Läs mer: Förskoleundervisning
linkkiVanda stad:
Ansökan till förskoleundervisningfinska _ svenska _ engelska
linkkiVanda stad:
Information om den förberedande undervisningenfinska _ engelska
linkkiVanda stad:
Elektronisk ansökningsblankett för förskoleundervisningenfinska _ svenska _ engelska
linkkiVanda stad:
Daghem som ger förskoleundervisningfinska _ engelska
Grundläggande utbildning
I Vanda finns finskspråkiga och svenskspråkiga grundskolor (peruskoulu).
I Vanda finns även en internationell skola, där man kan avlägga grundskolan på engelska.
Mer information om skolorna i Vanda hittar du på Vanda stads (Vantaan kaupunki) webbplats.
Anmälan till grundskolan ska göras på förhand.
Anmälningstiden är vanligtvis i januari.
På stadens webbplats hittar du kontaktuppgifterna till skolorna och mer information om anmälan.
Läs mer: Grundläggande utbildning
linkkiVanda stad:
Anmälan till skolanfinska _ svenska _ engelska
linkkiVanda stad:
Skolornas kontaktuppgifterfinska
Eftermiddagsverksamhetfinska _ svenska
Förberedande utbildning inför grundskola
Om barnets kunskaper i det finska språket inte är tillräckligt bra för studier i den finskspråkiga grundskolan, kan barnet få förberedande utbildning (valmistava opetus).
I den förberedande utbildningen läser barnen det finska språket och grundskolans läroämnen.
Undervisningen pågår vanligtvis i ett år.
Om du har anlänt till Finland för en kort tid sedan och har barn under skolåldern ska du ta kontakt med områdeskoordinatorn för ditt bostadsområde (aluekoordinaattori).
Områdeskoordinatorn berättar om hur undervisningen ordnas och hjälper dig i frågor som rör barnets skolgång.
Information om den förberedande undervisningenfinska
linkkiVanda stad:
Områdeskoordinatorerfinska
Grundläggande utbildning för unga invandrare
Vid Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto) kan 17–24-åriga invandrarungdomar avlägga grundskolans avgångsbetyg.
Om man har hoppat av grundskolan, kan man avlägga grundskolans lärokurs också vid Eira vuxengymnasium (Eiran aikuislukio).
Grundläggande utbildning för invandrarefinska
linkkiEira vuxengymnasium:
Grundundervisning för vuxnafinska
Tionde klasserna
Du kan ansöka till den grundläggande utbildningens tilläggsundervisning, det vill säga till en tionde klass (kymppiluokka), om du fick grundskolans avgångsbetyg samma år eller året innan, men inte har fått en studieplats på andra stadiet.
På tionde klassen kan du höja dina betyg från grundskolan och du får en plan för fortsatta studier.
Tiondeklasserna i Vanda finns i östra och västra Vanda vid Varias verksamhetsställen och vid Lumo gymnasium (Lumon lukio).
linkkiVanda stad:
Tiondeklasserfinska _ svenska
Invandrare och grundläggande utbildning
I skolorna i Vanda ges hemspråksundervisning i flera olika språk.
I grundskolorna ges även utbildning i finska som andraspråk (suomi toisena kielenä) till elever som har ett annat modersmål än finska, svenska eller samiska, och vars kunskaper i det finska språket inte är i nivå med modersmålet.
När du anmäler dig till skolan, kan du samtidigt anmäla dig till hemspråksundervisning och undervisning i din egen religion.
Du kan även anmäla dig till undervisningen genom att fylla i en blankett, som du får från din egen skola.
Den ifyllda blanketten returneras till den egna skolan.
Undervisning i den egna religionen kan ordnas om gruppen består av minst tre elever.
Mer information om hemspråksundervisning och om undervisning i elevens egen religion hittar du på stadens webbplats och hos områdeskoordinatorerna (aluekoordinaattori).
linkkiVanda stad:
Information om hemspråksundervisningfinska
linkkiVanda stad:
Undervisning i den egna religionenfinska
Finska som andra språk i den grundläggande undervisningenfinska
linkkiVanda stad:
Områdeskoordinatorerfinska
Yrkesutbildning
I Vanda ordnas yrkesutbildning vid yrkesinstitutet Vantaan ammattiopisto Varia, handelsläroanstalten MERCURIA samt TTS Arbetseffektivitetsföreningen rf:s verksamhetsställe i Vanda.
I Varia ordnas även engelskspråkig undervisning samt finskspråkiga yrkesutbildningar särskilt avsedda för invandrare.
Edupoli ordnar yrkesutbildning för vuxna.
I Vanda finns även Finavia Avia College som ger utbildning för olika luftfartsyrken.
Läs mer: Yrkesutbildning.
linkkiVanda stad:
Yrkesutbildningfinska _ svenska
linkkiYrkesläroanstalten Varia i Vanda:
Yrkesutbildningfinska _ engelska
Yrkesutbildningfinska _ engelska
linkkiTTS Arbetseffektivitetsföreningen rf:s verksamhetsställe i Vanda:
Yrkesutbildningfinska
Utbildning som handleder för yrkesutbildning (VALMA)
Utbildning som handleder för grundläggande yrkesutbildning (Ammatilliseen peruskoulutukseen valmentava koulutus) d.v.s. VALMA är avsedd för dem som vill avlägga en grundläggande yrkesutbildning.
Under VALMA-utbildningen får du kunskap och färdigheter som hjälper dig i dina senare yrkesinriktade studier.
Du kan även förbättra din språkkunskap. Du kan också höja dina grundskolebetyg.
I Vanda ordnas VALMA-utbildning av Varia.
Läs mer om VALMA-utbildningen på InfoFinlands sida Utbildning som handleder för yrkesutbildning.
linkkiVanda stad:
Information om VALMA-utbildningarfinska
linkkiYrkesläroanstalten Varia i Vanda:
I Vanda kan du studera på gymnasiet (lukio) på finska, svenska eller engelska.
Undervisning på engelska erbjuds på IB-linjen vid gymnasieskolan Tikkurilan lukio.
I Vanda finns även ett vuxengymnasium.
Läs mer: Gymnasium.
linkkiVanda stad:
Information om gymnasieutbildningfinska _ svenska
linkkiVanda stad:
Gymnasierna och gymnasiernas hemsidorfinska
linkkiVanda stad:
Vuxengymnasiumfinska
linkkiVanda stad:
Distansgymnasiumfinska
linkkiVanda stad:
Steinergymnasietfinska
Förberedande gymnasieutbildning (LUVA)
Om du vill förbättra dina kunskaper i finska eller svenska innan du söker till ett gymnasium, kan du söka till en förberedande gymnasieutbildning.
Den är avsedd för invandrare.
I Vanda ordnas LUVA-utbildning av Lumon lukio.
Läs mer om LUVA-utbildningen på InfoFinlands sida Förberedande gymnasieutbildning.
linkkiVanda stad:
Förberedande gymnasieutbildningfinska
Stöd och handledning för unga
Om du är under 30 år gammal kan du få råd och handledning via Ohjaamo-tjänsten.
Ohjaamos personal hjälper dig om du inte har ett arbete eller en studieplats.
Du kan även fråga om andra saker, som till exempel boende eller ekonomiska frågor.
linkkiOhjaamo:
Stöd och handledning för ungafinska _ engelska
Vägledningscentret Kipinä
Om du är under 29 år gammal, bor i Vanda och inte har ett jobb eller en studieplats, kan du få råd och handledning i Kipinä.
Ring och boka en tid i förväg.
Utan tidsbokning kan du besöka Kipinä på tisdagar och onsdagar kl. 12.00–18.00.
Mer information hittar du på webbplatsen.
Kipinä
Banvägen 2, Dickursby
Tfn 050 312 4372
Vägledning och stöd för ungafinska _ svenska
Högskoleutbildning
I Vanda finns två yrkeshögskolor (ammattikorkeakoulu), Laurea och Metropolia.
De erbjuder utbildning inom många olika branscher.
Mer information om utbildningsprogram och om ansökan hittar du på läroanstalternas webbplats.
Också Helsingfors universitets öppna universitet (avoin yliopisto) har verksamhetsställen i Vanda. Där ges undervisning på högskolenivå och fortbildning.
Läs mer: Högskoleutbildning.
linkkiVanda stad:
Högskoleutbildningfinska
Yrkeshögskolafinska _ engelska
linkkiMetropolia:
Yrkeshögskolafinska _ engelska
Ubildning vid öppna universitetet i Vandafinska _ svenska _ engelska
Övriga studiemöjligheter
Vid Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto) kan du studera till exempel språk, handarbete och matlagning eller delta i ledd motion.
Kurserna är avgiftsbelagda och de ordnas både dag- och kvällstid.
Vuxenutbildningsinstitutet ordnar även kurser för invandrare.
Mer information hittar du på Vanda stads webbplats.
Läs mer: Andra studiemöjligheter.
linkkiVanda vuxenutbildningsinstitut:
Studiehandbokfinska
linkkiVanda vuxenutbildningsinstitut:
Kurser i finska och svenska språket för invandrarefinska
linkkiEdupoli:
Vuxenutbildningscenterfinska
Dagvård
Förskoleundervisning
Grundläggande utbildning
Yrkesutbildning
Gymnasium
Stöd och handledning för unga
Högskoleutbildning
Övriga studiemöjligheter
Dagvård
I Vanda finns både kommunala och privata daghem.
Kommunen övervakar också den privata dagvården.
I Vanda ges dagvård på finska, svenska, ryska och engelska.
Inom dagvården ges även undervisning i finska som andra språk.
Dagvård ordnas också inom familjedagvården och i gruppfamiljedaghem.
Man ska ansöka om dagvårdsplats för sitt barn minst fyra månader innan barnet ska börja i dagvården.
Du kan ansöka om plats i den kommunala dagvården via Internet eller med en pappersblankett.
För en elektronisk ansökan behöver du egna nätbankskoder eller en elektronisk legitimation.
Pappersblanketter kan hämtas till exempel vid Vandainfo eller daghemmen.
Privata dagvårdsplatser söks direkt på daghemmet.
Frågor kring dagvård och ansökan om dagvårdsplats kan du ställa till daghemsföreståndaren eller skicka till adressen varhaiskasvatus(at)vantaa.fi.
Vanligtvis ansöker man om dagvårdsplats i den egna kommunen.
Om familjen bor nära gränsen till Helsingfors eller Esbo, kan du också söka dagvårdsplats i grannkommunen.
Du ska ändå lämna in din ansökan i den egna kommunen.
Mer information hittar du via tjänsten Helsingforsregionen.fi.
Läs mer: Dagvård
linkkiVanda stad:
Privat dagvårdfinska _ svenska _ engelska
linkkiVanda stad:
Privat dagvårdfinska
linkkiVanda stad:
Ansökan om dagvårdsplatsfinska _ svenska _ engelska
linkkiVanda stad:
Elektronisk ansökningsblankett för dagvårdenfinska _ svenska _ engelska
Information om dagvården finska _ svenska _ engelska
Förskoleundervisning
Förskoleundervisning (esiopetus) ordnas i både kommunala och privata daghem samt i förskoleenheter i skolornas lokaler.
I Vanda kan man få förskoleundervisning på finska, svenska och engelska.
Du måste ansöka om plats i förskoleundervisningen.
Ansökan kan göras elektroniskt via stadens webbplats eller med en pappersblankett.
Ansökningstiden är i januari, men ansökan kan även lämnas in övriga tider, om familjen till exempel flyttar till Vanda mitt under året.
Förberedande undervisning tillhandahålls för invandrarbarn som inte har tillräckliga kunskaper i finska för att klara sig i förskoleundervisningen.
Den förberedande undervisningen är avsedd för 6-åriga barn med invandrarbakgrund.
Den ordnas i daghemmens förskolegrupper.
Daghemmet anvisar barnet till den förberedande undervisningen i samband med ansökningen till förskoleundervisningen.
Du hittar mer information om förskoleundervisningen, ansökning till förskoleundervisningen och om undervisning som förbereder för förskoleundervisning på Vanda stads (Vantaan kaupunki) webbplats.
Du kan även fråga om mer information på daghemmen.
Läs mer: Förskoleundervisning
linkkiVanda stad:
Ansökan till förskoleundervisningfinska _ svenska _ engelska
linkkiVanda stad:
Information om den förberedande undervisningenfinska _ engelska
linkkiVanda stad:
Elektronisk ansökningsblankett för förskoleundervisningenfinska _ svenska _ engelska
linkkiVanda stad:
Daghem som ger förskoleundervisningfinska _ engelska
Grundläggande utbildning
I Vanda finns finskspråkiga och svenskspråkiga grundskolor (peruskoulu).
I Vanda finns även en internationell skola, där man kan avlägga grundskolan på engelska.
Mer information om skolorna i Vanda hittar du på Vanda stads (Vantaan kaupunki) webbplats.
Anmälan till grundskolan ska göras på förhand.
Anmälningstiden är vanligtvis i januari.
På stadens webbplats hittar du kontaktuppgifterna till skolorna och mer information om anmälan.
Läs mer: Grundläggande utbildning
linkkiVanda stad:
Anmälan till skolanfinska _ svenska _ engelska
linkkiVanda stad:
Skolornas kontaktuppgifterfinska
Eftermiddagsverksamhetfinska _ svenska
Förberedande utbildning inför grundskola
Om barnets kunskaper i det finska språket inte är tillräckligt bra för studier i den finskspråkiga grundskolan, kan barnet få förberedande utbildning (valmistava opetus).
I den förberedande utbildningen läser barnen det finska språket och grundskolans läroämnen.
Undervisningen pågår vanligtvis i ett år.
Om du har anlänt till Finland för en kort tid sedan och har barn under skolåldern ska du ta kontakt med områdeskoordinatorn för ditt bostadsområde (aluekoordinaattori).
Områdeskoordinatorn berättar om hur undervisningen ordnas och hjälper dig i frågor som rör barnets skolgång.
Information om den förberedande undervisningenfinska
linkkiVanda stad:
Områdeskoordinatorerfinska
Grundläggande utbildning för unga invandrare
Vid Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto) kan 17–24-åriga invandrarungdomar avlägga grundskolans avgångsbetyg.
Om man har hoppat av grundskolan, kan man avlägga grundskolans lärokurs också vid Eira vuxengymnasium (Eiran aikuislukio).
Grundläggande utbildning för invandrarefinska
linkkiEira vuxengymnasium:
Grundundervisning för vuxnafinska
Tionde klasserna
Du kan ansöka till den grundläggande utbildningens tilläggsundervisning, det vill säga till en tionde klass (kymppiluokka), om du fick grundskolans avgångsbetyg samma år eller året innan, men inte har fått en studieplats på andra stadiet.
På tionde klassen kan du höja dina betyg från grundskolan och du får en plan för fortsatta studier.
Tiondeklasserna i Vanda finns i östra och västra Vanda vid Varias verksamhetsställen och vid Lumo gymnasium (Lumon lukio).
linkkiVanda stad:
Tiondeklasserfinska _ svenska
Invandrare och grundläggande utbildning
I skolorna i Vanda ges hemspråksundervisning i flera olika språk.
I grundskolorna ges även utbildning i finska som andraspråk (suomi toisena kielenä) till elever som har ett annat modersmål än finska, svenska eller samiska, och vars kunskaper i det finska språket inte är i nivå med modersmålet.
När du anmäler dig till skolan, kan du samtidigt anmäla dig till hemspråksundervisning och undervisning i din egen religion.
Du kan även anmäla dig till undervisningen genom att fylla i en blankett, som du får från din egen skola.
Den ifyllda blanketten returneras till den egna skolan.
Undervisning i den egna religionen kan ordnas om gruppen består av minst tre elever.
Mer information om hemspråksundervisning och om undervisning i elevens egen religion hittar du på stadens webbplats och hos områdeskoordinatorerna (aluekoordinaattori).
linkkiVanda stad:
Information om hemspråksundervisningfinska
linkkiVanda stad:
Undervisning i den egna religionenfinska
Finska som andra språk i den grundläggande undervisningenfinska
linkkiVanda stad:
Områdeskoordinatorerfinska
Yrkesutbildning
I Vanda ordnas yrkesutbildning vid yrkesinstitutet Vantaan ammattiopisto Varia, handelsläroanstalten MERCURIA samt TTS Arbetseffektivitetsföreningen rf:s verksamhetsställe i Vanda.
I Varia ordnas även engelskspråkig undervisning samt finskspråkiga yrkesutbildningar särskilt avsedda för invandrare.
Edupoli ordnar yrkesutbildning för vuxna.
I Vanda finns även Finavia Avia College som ger utbildning för olika luftfartsyrken.
Läs mer: Yrkesutbildning.
linkkiVanda stad:
Yrkesutbildningfinska _ svenska
linkkiYrkesläroanstalten Varia i Vanda:
Yrkesutbildningfinska _ engelska
Yrkesutbildningfinska _ engelska
linkkiTTS Arbetseffektivitetsföreningen rf:s verksamhetsställe i Vanda:
Yrkesutbildningfinska
Utbildning som handleder för yrkesutbildning (VALMA)
Utbildning som handleder för grundläggande yrkesutbildning (Ammatilliseen peruskoulutukseen valmentava koulutus) d.v.s. VALMA är avsedd för dem som vill avlägga en grundläggande yrkesutbildning.
Under VALMA-utbildningen får du kunskap och färdigheter som hjälper dig i dina senare yrkesinriktade studier.
Du kan även förbättra din språkkunskap. Du kan också höja dina grundskolebetyg.
I Vanda ordnas VALMA-utbildning av Varia.
Läs mer om VALMA-utbildningen på InfoFinlands sida Utbildning som handleder för yrkesutbildning.
linkkiVanda stad:
Information om VALMA-utbildningarfinska
linkkiYrkesläroanstalten Varia i Vanda:
I Vanda kan du studera på gymnasiet (lukio) på finska, svenska eller engelska.
Undervisning på engelska erbjuds på IB-linjen vid gymnasieskolan Tikkurilan lukio.
I Vanda finns även ett vuxengymnasium.
Läs mer: Gymnasium.
linkkiVanda stad:
Information om gymnasieutbildningfinska _ svenska
linkkiVanda stad:
Gymnasierna och gymnasiernas hemsidorfinska
linkkiVanda stad:
Vuxengymnasiumfinska
linkkiVanda stad:
Distansgymnasiumfinska
linkkiVanda stad:
Steinergymnasietfinska
Förberedande gymnasieutbildning (LUVA)
Om du vill förbättra dina kunskaper i finska eller svenska innan du söker till ett gymnasium, kan du söka till en förberedande gymnasieutbildning.
Den är avsedd för invandrare.
I Vanda ordnas LUVA-utbildning av Lumon lukio.
Läs mer om LUVA-utbildningen på InfoFinlands sida Förberedande gymnasieutbildning.
linkkiVanda stad:
Förberedande gymnasieutbildningfinska
Stöd och handledning för unga
Om du är under 30 år gammal kan du få råd och handledning via Ohjaamo-tjänsten.
Ohjaamos personal hjälper dig om du inte har ett arbete eller en studieplats.
Du kan även fråga om andra saker, som till exempel boende eller ekonomiska frågor.
linkkiOhjaamo:
Stöd och handledning för ungafinska _ engelska
Vägledningscentret Kipinä
Om du är under 29 år gammal, bor i Vanda och inte har ett jobb eller en studieplats, kan du få råd och handledning i Kipinä.
Ring och boka en tid i förväg.
Utan tidsbokning kan du besöka Kipinä på tisdagar och onsdagar kl. 12.00–18.00.
Mer information hittar du på webbplatsen.
Kipinä
Banvägen 2, Dickursby
Tfn 050 312 4372
Vägledning och stöd för ungafinska _ svenska
Högskoleutbildning
I Vanda finns två yrkeshögskolor (ammattikorkeakoulu), Laurea och Metropolia.
De erbjuder utbildning inom många olika branscher.
Mer information om utbildningsprogram och om ansökan hittar du på läroanstalternas webbplats.
Också Helsingfors universitets öppna universitet (avoin yliopisto) har verksamhetsställen i Vanda. Där ges undervisning på högskolenivå och fortbildning.
Läs mer: Högskoleutbildning.
linkkiVanda stad:
Högskoleutbildningfinska
Yrkeshögskolafinska _ engelska
linkkiMetropolia:
Yrkeshögskolafinska _ engelska
Ubildning vid öppna universitetet i Vandafinska _ svenska _ engelska
Övriga studiemöjligheter
Vid Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto) kan du studera till exempel språk, handarbete och matlagning eller delta i ledd motion.
Kurserna är avgiftsbelagda och de ordnas både dag- och kvällstid.
Vuxenutbildningsinstitutet ordnar även kurser för invandrare.
Mer information hittar du på Vanda stads webbplats.
Läs mer: Andra studiemöjligheter.
linkkiVanda vuxenutbildningsinstitut:
Studiehandbokfinska
linkkiVanda vuxenutbildningsinstitut:
Kurser i finska och svenska språket för invandrarefinska
linkkiEdupoli:
Vuxenutbildningscenterfinska
Dagvård
Förskoleundervisning
Grundläggande utbildning
Yrkesutbildning
Gymnasium
Stöd och handledning för unga
Högskoleutbildning
Övriga studiemöjligheter
Dagvård
I Vanda finns både kommunala och privata daghem.
Kommunen övervakar också den privata dagvården.
I Vanda ges dagvård på finska, svenska, ryska och engelska.
Inom dagvården ges även undervisning i finska som andra språk.
Dagvård ordnas också inom familjedagvården och i gruppfamiljedaghem.
Man ska ansöka om dagvårdsplats för sitt barn minst fyra månader innan barnet ska börja i dagvården.
Du kan ansöka om plats i den kommunala dagvården via Internet eller med en pappersblankett.
För en elektronisk ansökan behöver du egna nätbankskoder eller en elektronisk legitimation.
Pappersblanketter kan hämtas till exempel vid Vandainfo eller daghemmen.
Privata dagvårdsplatser söks direkt på daghemmet.
Frågor kring dagvård och ansökan om dagvårdsplats kan du ställa till daghemsföreståndaren eller skicka till adressen varhaiskasvatus(at)vantaa.fi.
Vanligtvis ansöker man om dagvårdsplats i den egna kommunen.
Om familjen bor nära gränsen till Helsingfors eller Esbo, kan du också söka dagvårdsplats i grannkommunen.
Du ska ändå lämna in din ansökan i den egna kommunen.
Mer information hittar du via tjänsten Helsingforsregionen.fi.
Läs mer: Dagvård
linkkiVanda stad:
Privat dagvårdfinska _ svenska _ engelska
linkkiVanda stad:
Privat dagvårdfinska
linkkiVanda stad:
Ansökan om dagvårdsplatsfinska _ svenska _ engelska
linkkiVanda stad:
Elektronisk ansökningsblankett för dagvårdenfinska _ svenska _ engelska
Information om dagvården finska _ svenska _ engelska
Förskoleundervisning
Förskoleundervisning (esiopetus) ordnas i både kommunala och privata daghem samt i förskoleenheter i skolornas lokaler.
I Vanda kan man få förskoleundervisning på finska, svenska och engelska.
Du måste ansöka om plats i förskoleundervisningen.
Ansökan kan göras elektroniskt via stadens webbplats eller med en pappersblankett.
Ansökningstiden är i januari, men ansökan kan även lämnas in övriga tider, om familjen till exempel flyttar till Vanda mitt under året.
Förberedande undervisning tillhandahålls för invandrarbarn som inte har tillräckliga kunskaper i finska för att klara sig i förskoleundervisningen.
Den förberedande undervisningen är avsedd för 6-åriga barn med invandrarbakgrund.
Den ordnas i daghemmens förskolegrupper.
Daghemmet anvisar barnet till den förberedande undervisningen i samband med ansökningen till förskoleundervisningen.
Du hittar mer information om förskoleundervisningen, ansökning till förskoleundervisningen och om undervisning som förbereder för förskoleundervisning på Vanda stads (Vantaan kaupunki) webbplats.
Du kan även fråga om mer information på daghemmen.
Läs mer: Förskoleundervisning
linkkiVanda stad:
Ansökan till förskoleundervisningfinska _ svenska _ engelska
linkkiVanda stad:
Information om den förberedande undervisningenfinska _ engelska
linkkiVanda stad:
Elektronisk ansökningsblankett för förskoleundervisningenfinska _ svenska _ engelska
linkkiVanda stad:
Daghem som ger förskoleundervisningfinska _ engelska
Grundläggande utbildning
I Vanda finns finskspråkiga och svenskspråkiga grundskolor (peruskoulu).
I Vanda finns även en internationell skola, där man kan avlägga grundskolan på engelska.
Mer information om skolorna i Vanda hittar du på Vanda stads (Vantaan kaupunki) webbplats.
Anmälan till grundskolan ska göras på förhand.
Anmälningstiden är vanligtvis i januari.
På stadens webbplats hittar du kontaktuppgifterna till skolorna och mer information om anmälan.
Läs mer: Grundläggande utbildning
linkkiVanda stad:
Anmälan till skolanfinska _ svenska _ engelska
linkkiVanda stad:
Skolornas kontaktuppgifterfinska
Eftermiddagsverksamhetfinska _ svenska
Förberedande utbildning inför grundskola
Om barnets kunskaper i det finska språket inte är tillräckligt bra för studier i den finskspråkiga grundskolan, kan barnet få förberedande utbildning (valmistava opetus).
I den förberedande utbildningen läser barnen det finska språket och grundskolans läroämnen.
Undervisningen pågår vanligtvis i ett år.
Om du har anlänt till Finland för en kort tid sedan och har barn under skolåldern ska du ta kontakt med områdeskoordinatorn för ditt bostadsområde (aluekoordinaattori).
Områdeskoordinatorn berättar om hur undervisningen ordnas och hjälper dig i frågor som rör barnets skolgång.
Information om den förberedande undervisningenfinska
linkkiVanda stad:
Områdeskoordinatorerfinska
Grundläggande utbildning för unga invandrare
Vid Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto) kan 17–24-åriga invandrarungdomar avlägga grundskolans avgångsbetyg.
Om man har hoppat av grundskolan, kan man avlägga grundskolans lärokurs också vid Eira vuxengymnasium (Eiran aikuislukio).
Grundläggande utbildning för invandrarefinska
linkkiEira vuxengymnasium:
Grundundervisning för vuxnafinska
Tionde klasserna
Du kan ansöka till den grundläggande utbildningens tilläggsundervisning, det vill säga till en tionde klass (kymppiluokka), om du fick grundskolans avgångsbetyg samma år eller året innan, men inte har fått en studieplats på andra stadiet.
På tionde klassen kan du höja dina betyg från grundskolan och du får en plan för fortsatta studier.
Tiondeklasserna i Vanda finns i östra och västra Vanda vid Varias verksamhetsställen och vid Lumo gymnasium (Lumon lukio).
linkkiVanda stad:
Tiondeklasserfinska _ svenska
Invandrare och grundläggande utbildning
I skolorna i Vanda ges hemspråksundervisning i flera olika språk.
I grundskolorna ges även utbildning i finska som andraspråk (suomi toisena kielenä) till elever som har ett annat modersmål än finska, svenska eller samiska, och vars kunskaper i det finska språket inte är i nivå med modersmålet.
När du anmäler dig till skolan, kan du samtidigt anmäla dig till hemspråksundervisning och undervisning i din egen religion.
Du kan även anmäla dig till undervisningen genom att fylla i en blankett, som du får från din egen skola.
Den ifyllda blanketten returneras till den egna skolan.
Undervisning i den egna religionen kan ordnas om gruppen består av minst tre elever.
Mer information om hemspråksundervisning och om undervisning i elevens egen religion hittar du på stadens webbplats och hos områdeskoordinatorerna (aluekoordinaattori).
linkkiVanda stad:
Information om hemspråksundervisningfinska
linkkiVanda stad:
Undervisning i den egna religionenfinska
Finska som andra språk i den grundläggande undervisningenfinska
linkkiVanda stad:
Områdeskoordinatorerfinska
Yrkesutbildning
I Vanda ordnas yrkesutbildning vid yrkesinstitutet Vantaan ammattiopisto Varia, handelsläroanstalten MERCURIA samt TTS Arbetseffektivitetsföreningen rf:s verksamhetsställe i Vanda.
I Varia ordnas även engelskspråkig undervisning samt finskspråkiga yrkesutbildningar särskilt avsedda för invandrare.
Edupoli ordnar yrkesutbildning för vuxna.
I Vanda finns även Finavia Avia College som ger utbildning för olika luftfartsyrken.
Läs mer: Yrkesutbildning.
linkkiVanda stad:
Yrkesutbildningfinska _ svenska
linkkiYrkesläroanstalten Varia i Vanda:
Yrkesutbildningfinska _ engelska
Yrkesutbildningfinska _ engelska
linkkiTTS Arbetseffektivitetsföreningen rf:s verksamhetsställe i Vanda:
Yrkesutbildningfinska
Utbildning som handleder för yrkesutbildning (VALMA)
Utbildning som handleder för grundläggande yrkesutbildning (Ammatilliseen peruskoulutukseen valmentava koulutus) d.v.s. VALMA är avsedd för dem som vill avlägga en grundläggande yrkesutbildning.
Under VALMA-utbildningen får du kunskap och färdigheter som hjälper dig i dina senare yrkesinriktade studier.
Du kan även förbättra din språkkunskap. Du kan också höja dina grundskolebetyg.
I Vanda ordnas VALMA-utbildning av Varia.
Läs mer om VALMA-utbildningen på InfoFinlands sida Utbildning som handleder för yrkesutbildning.
linkkiVanda stad:
Information om VALMA-utbildningarfinska
linkkiYrkesläroanstalten Varia i Vanda:
I Vanda kan du studera på gymnasiet (lukio) på finska, svenska eller engelska.
Undervisning på engelska erbjuds på IB-linjen vid gymnasieskolan Tikkurilan lukio.
I Vanda finns även ett vuxengymnasium.
Läs mer: Gymnasium.
linkkiVanda stad:
Information om gymnasieutbildningfinska _ svenska
linkkiVanda stad:
Gymnasierna och gymnasiernas hemsidorfinska
linkkiVanda stad:
Vuxengymnasiumfinska
linkkiVanda stad:
Distansgymnasiumfinska
linkkiVanda stad:
Steinergymnasietfinska
Förberedande gymnasieutbildning (LUVA)
Om du vill förbättra dina kunskaper i finska eller svenska innan du söker till ett gymnasium, kan du söka till en förberedande gymnasieutbildning.
Den är avsedd för invandrare.
I Vanda ordnas LUVA-utbildning av Lumon lukio.
Läs mer om LUVA-utbildningen på InfoFinlands sida Förberedande gymnasieutbildning.
linkkiVanda stad:
Förberedande gymnasieutbildningfinska
Stöd och handledning för unga
Om du är under 30 år gammal kan du få råd och handledning via Ohjaamo-tjänsten.
Ohjaamos personal hjälper dig om du inte har ett arbete eller en studieplats.
Du kan även fråga om andra saker, som till exempel boende eller ekonomiska frågor.
linkkiOhjaamo:
Stöd och handledning för ungafinska _ engelska
Vägledningscentret Kipinä
Om du är under 29 år gammal, bor i Vanda och inte har ett jobb eller en studieplats, kan du få råd och handledning i Kipinä.
Ring och boka en tid i förväg.
Utan tidsbokning kan du besöka Kipinä på tisdagar och onsdagar kl. 12.00–18.00.
Mer information hittar du på webbplatsen.
Kipinä
Banvägen 2, Dickursby
Tfn 050 312 4372
Vägledning och stöd för ungafinska _ svenska
Högskoleutbildning
I Vanda finns två yrkeshögskolor (ammattikorkeakoulu), Laurea och Metropolia.
De erbjuder utbildning inom många olika branscher.
Mer information om utbildningsprogram och om ansökan hittar du på läroanstalternas webbplats.
Också Helsingfors universitets öppna universitet (avoin yliopisto) har verksamhetsställen i Vanda. Där ges undervisning på högskolenivå och fortbildning.
Läs mer: Yrkeshögskolor, Universitet.
linkkiVanda stad:
Högskoleutbildningfinska
Yrkeshögskolafinska _ engelska
linkkiMetropolia:
Yrkeshögskolafinska _ engelska
Ubildning vid öppna universitetet i Vandafinska _ svenska _ engelska
Övriga studiemöjligheter
Vid Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto) kan du studera till exempel språk, handarbete och matlagning eller delta i ledd motion.
Kurserna är avgiftsbelagda och de ordnas både dag- och kvällstid.
Vuxenutbildningsinstitutet ordnar även kurser för invandrare.
Mer information hittar du på Vanda stads webbplats.
Läs mer: Studier som hobby.
linkkiVanda vuxenutbildningsinstitut:
Studiehandbokfinska
linkkiVanda vuxenutbildningsinstitut:
Kurser i finska och svenska språket för invandrarefinska
linkkiEdupoli:
Vuxenutbildningscenterfinska
Detta innehåll finns inte på det språk som du har valt.
Välj något annat språk.
Finska
Detta innehåll finns inte på det språk som du har valt.
Välj något annat språk.
Finska
Detta innehåll finns inte på det språk som du har valt.
Välj något annat språk.
Finska
Hyresbostad
Boende i en krissituation
Bostadslöshet
Stöd- och serviceboende
Bostadens avfallshantering
Hyresbostad
Hyresbostäderna är ofta dyra i huvudstadsregionen.
Du är själv ansvarig för att skaffa bostad åt dig själv.
Varken staden eller andra hyresvärdar har skyldighet att erbjuda dig bostad.
Läs mer: Hyresbostad.
Privata hyresbostäder
I Vanda finns också många andra hyresvärdar, varav de största är VVO, Sato och Avara.
Därtill ägs hyresbostäder i Vanda av många försäkringsbolag, Kuntien eläkevakuutus och Kunta-asunnot.
Det kan gå snabbt att få bostad via en privat hyresvärd.
Om du är studerande kan du ansöka om en hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS (Helsingin seudun Opiskelija-asuntosäätiö HOAS).
Om du är yngre än 30 år, kan du söka bostad hos Förbundet för ungdomsbostäder (Nuorisoasuntoliitto) och stiftelsen Nuorisosäätiö (Nuorisosäätiö).
linkkiSATO:
Hyresbostäderfinska _ engelska
linkkiAvara:
Hyresbostäderfinska
linkkiKommunbostäder:
Hyresbostäderfinska _ svenska _ engelska
linkkiFörbundet för ungdomsbostäder:
Hyresbostäder för personer under 30 årfinska _ engelska
Hyresbostäder för ungafinska _ engelska
linkkiHOAS:
Hyresbostäder för studerandefinska _ svenska _ engelska
Stadens hyresbostäder
Stadens hyresbostäder är vanligtvis förmånligare än de bostäder som hyrs ut av företag och privatpersoner.
Väntetiden för dessa bostäder kan dock vara lång och endast en liten del av de sökande får en bostad.
Vanda stads hyresbostäder ägs och hyrs ut av VAV Asunnot Oy.
Lokgränden 7
Tfn 010 235 1450 (kundtjänst)
Du kan göra en bostadsansökan på VAV Asunnot Oy:s webbplats.
Ansökan är giltig i fyra månader och måste sedan förnyas.
Vid val av invånare till stadens hyresbostäder prioriteras de sökande som har ett akut bostadsbehov.
Också sökandens inkomster beaktas, eftersom bostäderna främst är avsedda för personer med låga inkomster.
Information om stadens hyresbostäderfinska _ engelska
Ansökan om hyresbostad i stadenfinska _ engelska
Boende i en krissituation
Om din bostad har skadats till exempel till följd av brand eller vattenskada kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
Kontakta ditt försäkringsbolag direkt när skadan har inträffat.
I krissituationer får man även hjälp vid Vanda stads social- och krisjour (sosiaali- ja kriisipäivystys), som har öppet dygnet runt.
Telefonnumret till social- och krisjouren är (09) 8392 4005
linkkiVanda stad:
Social- och krisjourenfinska _ svenska _ engelska
Skyddshem
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta ett skyddshem (turvakoti).
Skyddshemmen har jourmottagning dygnet runt.
Skyddshemmet Mona är ett skyddshem avsett för invandrarkvinnor och deras barn.
Tfn 045 639 6274
Du kan även gå till Vanda skyddshem eller huvudstadsregionens skyddshem.
Tfn (09) 8392 0071
Steniusvägen 20
Tfn (09) 4777 180
linkkiTurvakoti Mona:
Skyddshemfinska
Skyddshemfinska _ engelska
Hjälp till offer för familjevåldfinska
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
De ungas skyddshus
Finlands Röda Kors De ungas skyddshus (Suomen Punaisen Ristin Nuorten turvatalo) ger stöd och hjälp i krissituationer för 12–19-åriga ungdomar.
Skyddshuset har öppet kl. 17–10, telefonjouren betjänar dygnet runt.
Sjukhusgatan 3 (Räckhals gård)
Tfn (09) 871 4043
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Bostadslöshet
Om du blir bostadslös ska du kontakta socialstationen (sosiaaliasema) för ditt eget område.
Kontaktuppgifterna hittar du på Vanda stads webbplats.
Om din hemkommun är Vanda, kan du få en bostad via Sininauha Oy eller Villenpirtti.
Läs mer: Bostadslöshet
linkkiVanda stad:
Socialtjänsterfinska _ svenska _ engelska
Bostäder för bostadslösafinska
Stödboende för personer med psykisk ohälsa och missbruksproblemfinska
Stöd- och serviceboende
Staden ordnar boendetjänster till exempel för åldringar och handikappade, som har svårt att klara av de dagliga sysslorna utan hjälp.
Åldringar och handikappade som inte klarar av att bo självständigt, kan bo i servicehus (palvelutalo) eller på en vårdinrättning (laitos).
Mer information om dessa tjänster får du från enheten för socialt arbete (sosiaalityön yksikkö) i ditt bostadsområde.
Läs mer: Stöd- och serviceboende.
linkkiVanda stad:
Information om hemvårdens stödtjänsterfinska
linkkiVanda stad:
Information om stadens servicebostäderfinska
linkkiVanda stad:
Privata servicehusfinska
linkkiVanda stad:
Socialtjänsterfinska _ svenska _ engelska
Bostadens avfallshantering
Information om var din närmaste återvinningsstation (kierrätyspiste) ligger hittar du på webbplatsen kierrätys.info.
Läs mer: Avfallshantering och återvinning.
linkkiAvfallsverksföreningen:
Återvinningsstationerfinska
linkkiHRM:
Återvinningsstationerfinska _ svenska _ engelska
Hyresbostad
Boende i en krissituation
Bostadslöshet
Stöd- och serviceboende
Bostadens avfallshantering
Hyresbostad
Hyresbostäderna är ofta dyra i huvudstadsregionen.
Du är själv ansvarig för att skaffa bostad åt dig själv.
Varken staden eller andra hyresvärdar har skyldighet att erbjuda dig bostad.
Läs mer: Hyresbostad.
Privata hyresbostäder
I Vanda finns också många andra hyresvärdar, varav de största är VVO, Sato och Avara.
Därtill ägs hyresbostäder i Vanda av många försäkringsbolag, Kuntien eläkevakuutus och Kunta-asunnot.
Det kan gå snabbt att få bostad via en privat hyresvärd.
Om du är studerande kan du ansöka om en hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS (Helsingin seudun Opiskelija-asuntosäätiö HOAS).
Om du är yngre än 30 år, kan du söka bostad hos Förbundet för ungdomsbostäder (Nuorisoasuntoliitto) och stiftelsen Nuorisosäätiö (Nuorisosäätiö).
linkkiSATO:
Hyresbostäderfinska _ engelska
linkkiAvara:
Hyresbostäderfinska
linkkiKommunbostäder:
Hyresbostäderfinska _ svenska _ engelska
linkkiFörbundet för ungdomsbostäder:
Hyresbostäder för personer under 30 årfinska _ engelska
Hyresbostäder för ungafinska _ engelska
linkkiHOAS:
Hyresbostäder för studerandefinska _ svenska _ engelska
Stadens hyresbostäder
Stadens hyresbostäder är vanligtvis förmånligare än de bostäder som hyrs ut av företag och privatpersoner.
Väntetiden för dessa bostäder kan dock vara lång och endast en liten del av de sökande får en bostad.
Vanda stads hyresbostäder ägs och hyrs ut av VAV Asunnot Oy.
Lokgränden 7
Tfn 010 235 1450 (kundtjänst)
Du kan göra en bostadsansökan på VAV Asunnot Oy:s webbplats.
Ansökan är giltig i fyra månader och måste sedan förnyas.
Vid val av invånare till stadens hyresbostäder prioriteras de sökande som har ett akut bostadsbehov.
Också sökandens inkomster beaktas, eftersom bostäderna främst är avsedda för personer med låga inkomster.
Information om stadens hyresbostäderfinska _ engelska
Ansökan om hyresbostad i stadenfinska _ engelska
Boende i en krissituation
Om din bostad har skadats till exempel till följd av brand eller vattenskada kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
Kontakta ditt försäkringsbolag direkt när skadan har inträffat.
I krissituationer får man även hjälp vid Vanda stads social- och krisjour (sosiaali- ja kriisipäivystys), som har öppet dygnet runt.
Telefonnumret till social- och krisjouren är (09) 8392 4005
linkkiVanda stad:
Social- och krisjourenfinska _ svenska _ engelska
Skyddshem
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta ett skyddshem (turvakoti).
Skyddshemmen har jourmottagning dygnet runt.
Skyddshemmet Mona är ett skyddshem avsett för invandrarkvinnor och deras barn.
Tfn 045 639 6274
Du kan även gå till Vanda skyddshem eller huvudstadsregionens skyddshem.
Tfn (09) 8392 0071
Steniusvägen 20
Tfn (09) 4777 180
linkkiTurvakoti Mona:
Skyddshemfinska
Skyddshemfinska _ engelska
Hjälp till offer för familjevåldfinska
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
De ungas skyddshus
Finlands Röda Kors De ungas skyddshus (Suomen Punaisen Ristin Nuorten turvatalo) ger stöd och hjälp i krissituationer för 12–19-åriga ungdomar.
Skyddshuset har öppet kl. 17–10, telefonjouren betjänar dygnet runt.
Sjukhusgatan 3 (Räckhals gård)
Tfn (09) 871 4043
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Bostadslöshet
Om du blir bostadslös ska du kontakta socialstationen (sosiaaliasema) för ditt eget område.
Kontaktuppgifterna hittar du på Vanda stads webbplats.
Om din hemkommun är Vanda, kan du få en bostad via Sininauha Oy eller Villenpirtti.
Läs mer: Bostadslöshet
linkkiVanda stad:
Socialtjänsterfinska _ svenska _ engelska
Bostäder för bostadslösafinska
Stödboende för personer med psykisk ohälsa och missbruksproblemfinska
Stöd- och serviceboende
Staden ordnar boendetjänster till exempel för åldringar och handikappade, som har svårt att klara av de dagliga sysslorna utan hjälp.
Åldringar och handikappade som inte klarar av att bo självständigt, kan bo i servicehus (palvelutalo) eller på en vårdinrättning (laitos).
Mer information om dessa tjänster får du från enheten för socialt arbete (sosiaalityön yksikkö) i ditt bostadsområde.
Läs mer: Stöd- och serviceboende.
linkkiVanda stad:
Information om hemvårdens stödtjänsterfinska
linkkiVanda stad:
Information om stadens servicebostäderfinska
linkkiVanda stad:
Privata servicehusfinska
linkkiVanda stad:
Socialtjänsterfinska _ svenska _ engelska
Bostadens avfallshantering
Information om var din närmaste återvinningsstation (kierrätyspiste) ligger hittar du på webbplatsen kierrätys.info.
Läs mer: Avfallshantering och återvinning.
linkkiAvfallsverksföreningen:
Återvinningsstationerfinska
linkkiHRM:
Återvinningsstationerfinska _ svenska _ engelska
Hyresbostad
Boende i en krissituation
Bostadslöshet
Stöd- och serviceboende
Bostadens avfallshantering
Hyresbostad
Hyresbostäderna är ofta dyra i huvudstadsregionen.
Du är själv ansvarig för att skaffa bostad åt dig själv.
Varken staden eller andra hyresvärdar har skyldighet att erbjuda dig bostad.
Läs mer: Hyresbostad.
Privata hyresbostäder
I Vanda finns också många andra hyresvärdar, varav de största är VVO, Sato och Avara.
Därtill ägs hyresbostäder i Vanda av många försäkringsbolag, Kuntien eläkevakuutus och Kunta-asunnot.
Det kan gå snabbt att få bostad via en privat hyresvärd.
Om du är studerande kan du ansöka om en hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS (Helsingin seudun Opiskelija-asuntosäätiö HOAS).
Om du är yngre än 30 år, kan du söka bostad hos Förbundet för ungdomsbostäder (Nuorisoasuntoliitto) och stiftelsen Nuorisosäätiö (Nuorisosäätiö).
linkkiSATO:
Hyresbostäderfinska _ engelska
linkkiAvara:
Hyresbostäderfinska
linkkiKommunbostäder:
Hyresbostäderfinska _ svenska _ engelska
linkkiFörbundet för ungdomsbostäder:
Hyresbostäder för personer under 30 årfinska _ engelska
Hyresbostäder för ungafinska _ engelska
linkkiHOAS:
Hyresbostäder för studerandefinska _ svenska _ engelska
Stadens hyresbostäder
Stadens hyresbostäder är vanligtvis förmånligare än de bostäder som hyrs ut av företag och privatpersoner.
Väntetiden för dessa bostäder kan dock vara lång och endast en liten del av de sökande får en bostad.
Vanda stads hyresbostäder ägs och hyrs ut av VAV Asunnot Oy.
Lokgränden 7
Tfn 010 235 1450 (kundtjänst)
Du kan göra en bostadsansökan på VAV Asunnot Oy:s webbplats.
Ansökan är giltig i fyra månader och måste sedan förnyas.
Vid val av invånare till stadens hyresbostäder prioriteras de sökande som har ett akut bostadsbehov.
Också sökandens inkomster beaktas, eftersom bostäderna främst är avsedda för personer med låga inkomster.
Information om stadens hyresbostäderfinska _ engelska
Ansökan om hyresbostad i stadenfinska _ engelska
Boende i en krissituation
Om din bostad har skadats till exempel till följd av brand eller vattenskada kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
Kontakta ditt försäkringsbolag direkt när skadan har inträffat.
I krissituationer får man även hjälp vid Vanda stads social- och krisjour (sosiaali- ja kriisipäivystys), som har öppet dygnet runt.
Telefonnumret till social- och krisjouren är (09) 8392 4005
linkkiVanda stad:
Social- och krisjourenfinska _ svenska _ engelska
Skyddshem
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta ett skyddshem (turvakoti).
Skyddshemmen har jourmottagning dygnet runt.
Skyddshemmet Mona är ett skyddshem avsett för invandrarkvinnor och deras barn.
Tfn 045 639 6274
Du kan även gå till Vanda skyddshem eller huvudstadsregionens skyddshem.
Tfn (09) 8392 0071
Steniusvägen 20
Tfn (09) 4777 180
linkkiTurvakoti Mona:
Skyddshemfinska
Skyddshemfinska _ engelska
Hjälp till offer för familjevåldfinska
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
De ungas skyddshus
Finlands Röda Kors De ungas skyddshus (Suomen Punaisen Ristin Nuorten turvatalo) ger stöd och hjälp i krissituationer för 12–19-åriga ungdomar.
Skyddshuset har öppet kl. 17–10, telefonjouren betjänar dygnet runt.
Sjukhusgatan 3 (Räckhals gård)
Tfn (09) 871 4043
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Bostadslöshet
Om du blir bostadslös ska du kontakta socialstationen (sosiaaliasema) för ditt eget område.
Kontaktuppgifterna hittar du på Vanda stads webbplats.
Om din hemkommun är Vanda, kan du få en bostad via Sininauha Oy eller Villenpirtti.
Läs mer: Bostadslöshet
linkkiVanda stad:
Socialtjänsterfinska _ svenska _ engelska
Bostäder för bostadslösafinska
Stödboende för personer med psykisk ohälsa och missbruksproblemfinska
Stöd- och serviceboende
Staden ordnar boendetjänster till exempel för åldringar och handikappade, som har svårt att klara av de dagliga sysslorna utan hjälp.
Åldringar och handikappade som inte klarar av att bo självständigt, kan bo i servicehus (palvelutalo) eller på en vårdinrättning (laitos).
Mer information om dessa tjänster får du från enheten för socialt arbete (sosiaalityön yksikkö) i ditt bostadsområde.
Läs mer: Stöd- och serviceboende.
linkkiVanda stad:
Information om hemvårdens stödtjänsterfinska
linkkiVanda stad:
Information om stadens servicebostäderfinska
linkkiVanda stad:
Privata servicehusfinska
linkkiVanda stad:
Socialtjänsterfinska _ svenska _ engelska
Bostadens avfallshantering
Information om var din närmaste återvinningsstation (kierrätyspiste) ligger hittar du på webbplatsen kierrätys.info.
Läs mer: Avfallshantering och återvinning.
linkkiAvfallsverksföreningen:
Återvinningsstationerfinska
linkkiHRM:
Återvinningsstationerfinska _ svenska _ engelska
Möjligheter att studera det finska eller svenska språket
Språkkurser
Med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors, Vanda, Esbo eller Grankulla.
Kurserna i svenska hittar du genom att klicka på länken på tjänstens startsida.
Kurserna i tjänsten finnishcourses.fi är öppna för alla.
Tjänsten omfattar inte arbets- och näringsbyråns kurser.
I Vanda anordnas kurser i finska och svenska språket för invandrare av Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto) Kurserna vid institutet är öppna för alla.
Vuxenutbildningsinstitutet ligger i Dickursby, men kurser ordnas runtom i Vanda.
Adress:
Näckrosvägen 5
Tfn (09) 8392 4342
Ytterligare information om kurser och anmälan hittar du på Vanda vuxenutbildningsinstituts webbplats och i studiehandboken.
Du får studiehandboken till exempel på bibliotek eller Vandainfo samt i elektroniskt format på Vanda stads webbplats.
Arbets- och näringsbyrån anvisar invandrare till kurser i finska språket som ingår i integrationsprocessen.
I samband med att en integrations- eller sysselsättningsplan upprättas för dig, kan du också få också en studieplats på en finskakurs reserverad eller också kan du ställas i kö för en studieplats.
Mer information hittar du vid arbets- och näringsbyrån.
Läs mer: Studier i finska och svenska
Kurser i finska och svenska språketfinska _ engelska _ ryska
linkkiVanda vuxenutbildningsinstitut:
Kurser i finska och svenska språket för invandrarefinska
linkkiArbets- och näringsministeriet:
Utbildning i finska och svenska språketfinska _ svenska _ engelska
linkkiVanda vuxenutbildningsinstitut:
Grundundervisning för vuxnafinska
Samtal på finska
På Vanda stadsbibliotek anordnas språkcaféer (kielikahvila), där man kan öva på att prata finska.
Alla som vill lära sig tala finska är välkomna till caféerna.
På språkcaféerna talar vi finska, så det är bra om du redan kan lite finska.
Språkcaféerna är avgiftsfria.
Mer information om språkcaféerna får du från biblioteken.
I Vanda anordnas samtalsklubbar på finska också på Silkesportens verksamhetscenter (Silkinportin toimintakeskus) och Kafnettis och Myyrinkis boendeträffpunkter (Kafnetin ja Myyringin asukastila).
Finskaklubbar avsedda för föräldrar som vårdar barn i hemmet anordnas i invånarparkerna (asukaspuisto) och i de öppna daghemmen (avoin päiväkoti).
Klubbarna för att lära sig tala finska är avgiftsfria.
Läsundervisning
Nätverket Vi läser tillsammans (Luetaan yhdessä-verkosto) erbjuder undervisning i läsning och det finska språket för invandrarkvinnor.
Flera olika Vi läser tillsammans-nätverk är verksamma på olika håll i Vanda.
Det är avgiftsfritt att delta i grupperna.
Språkkaféerfinska _ engelska _ ryska
linkkiVanda stad:
Invånarlokalfinska _ engelska
linkkiVanda stad:
Invånarlokalfinska _ engelska
linkkiVanda stad:
Parker för invånare och öppna daghemfinska _ svenska _ engelska
linkkiVi läser tillsammans-nätverket:
Vi läser tillsammans i Vandafinska _ svenska _ engelska
Allmän språkexamen
Du kan avlägga allmän språkexamen i finska eller svenska språket.
På utbildningsstyrelsens (Opetushallitus) webbplats finns en sökmotor med vilken du kan kontrollera var och när du kan avlägga examen.
I Vanda ordnas språkexamina till exempel vid Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto).
Läs mer: Officiellt intyg på språkkunskaper.
linkkiUtbildningsstyrelsen:
Att anmäla sig till en allmän språkexamen och examensavgifterfinska _ svenska _ engelska
linkkiVanda vuxenutbildningsinstitut:
Allmän språkexamenfinska
linkkiUtbildningsstyrelsen:
Examenssökningfinska
Möjligheter att studera det finska eller svenska språket
Språkkurser
Med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors, Vanda, Esbo eller Grankulla.
Kurserna i svenska hittar du genom att klicka på länken på tjänstens startsida.
Kurserna i tjänsten finnishcourses.fi är öppna för alla.
Tjänsten omfattar inte arbets- och näringsbyråns kurser.
I Vanda anordnas kurser i finska och svenska språket för invandrare av Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto) Kurserna vid institutet är öppna för alla.
Vuxenutbildningsinstitutet ligger i Dickursby, men kurser ordnas runtom i Vanda.
Adress:
Näckrosvägen 5
Tfn (09) 8392 4342
Ytterligare information om kurser och anmälan hittar du på Vanda vuxenutbildningsinstituts webbplats och i studiehandboken.
Du får studiehandboken till exempel på bibliotek eller Vandainfo samt i elektroniskt format på Vanda stads webbplats.
Arbets- och näringsbyrån anvisar invandrare till kurser i finska språket som ingår i integrationsprocessen.
I samband med att en integrations- eller sysselsättningsplan upprättas för dig, kan du också få också en studieplats på en finskakurs reserverad eller också kan du ställas i kö för en studieplats.
Mer information hittar du vid arbets- och näringsbyrån.
Läs mer: Studier i finska och svenska
Kurser i finska och svenska språketfinska _ engelska _ ryska
linkkiVanda vuxenutbildningsinstitut:
Kurser i finska och svenska språket för invandrarefinska
linkkiArbets- och näringsministeriet:
Utbildning i finska och svenska språketfinska _ svenska _ engelska
linkkiVanda vuxenutbildningsinstitut:
Grundundervisning för vuxnafinska
Samtal på finska
På Vanda stadsbibliotek anordnas språkcaféer (kielikahvila), där man kan öva på att prata finska.
Alla som vill lära sig tala finska är välkomna till caféerna.
På språkcaféerna talar vi finska, så det är bra om du redan kan lite finska.
Språkcaféerna är avgiftsfria.
Mer information om språkcaféerna får du från biblioteken.
I Vanda anordnas samtalsklubbar på finska också på Silkesportens verksamhetscenter (Silkinportin toimintakeskus) och Kafnettis och Myyrinkis boendeträffpunkter (Kafnetin ja Myyringin asukastila).
Finskaklubbar avsedda för föräldrar som vårdar barn i hemmet anordnas i invånarparkerna (asukaspuisto) och i de öppna daghemmen (avoin päiväkoti).
Klubbarna för att lära sig tala finska är avgiftsfria.
Läsundervisning
Nätverket Vi läser tillsammans (Luetaan yhdessä-verkosto) erbjuder undervisning i läsning och det finska språket för invandrarkvinnor.
Flera olika Vi läser tillsammans-nätverk är verksamma på olika håll i Vanda.
Det är avgiftsfritt att delta i grupperna.
Språkkaféerfinska _ engelska _ ryska
linkkiVanda stad:
Invånarlokalfinska _ engelska
linkkiVanda stad:
Invånarlokalfinska _ engelska
linkkiVanda stad:
Parker för invånare och öppna daghemfinska _ svenska _ engelska
linkkiVi läser tillsammans-nätverket:
Vi läser tillsammans i Vandafinska _ svenska _ engelska
Allmän språkexamen
Du kan avlägga allmän språkexamen i finska eller svenska språket.
På utbildningsstyrelsens (Opetushallitus) webbplats finns en sökmotor med vilken du kan kontrollera var och när du kan avlägga examen.
I Vanda ordnas språkexamina till exempel vid Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto).
Läs mer: Officiellt intyg på språkkunskaper.
linkkiUtbildningsstyrelsen:
Att anmäla sig till en allmän språkexamen och examensavgifterfinska _ svenska _ engelska
linkkiVanda vuxenutbildningsinstitut:
Allmän språkexamenfinska
linkkiUtbildningsstyrelsen:
Examenssökningfinska
Möjligheter att studera det finska eller svenska språket
Språkkurser
Med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors, Vanda, Esbo eller Grankulla.
Kurserna i svenska hittar du genom att klicka på länken på tjänstens startsida.
Kurserna i tjänsten finnishcourses.fi är öppna för alla.
Tjänsten omfattar inte arbets- och näringsbyråns kurser.
I Vanda anordnas kurser i finska och svenska språket för invandrare av Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto) Kurserna vid institutet är öppna för alla.
Vuxenutbildningsinstitutet ligger i Dickursby, men kurser ordnas runtom i Vanda.
Adress:
Näckrosvägen 5
Tfn (09) 8392 4342
Ytterligare information om kurser och anmälan hittar du på Vanda vuxenutbildningsinstituts webbplats och i studiehandboken.
Du får studiehandboken till exempel på bibliotek eller Vandainfo samt i elektroniskt format på Vanda stads webbplats.
Arbets- och näringsbyrån anvisar invandrare till kurser i finska språket som ingår i integrationsprocessen.
I samband med att en integrations- eller sysselsättningsplan upprättas för dig, kan du också få också en studieplats på en finskakurs reserverad eller också kan du ställas i kö för en studieplats.
Mer information hittar du vid arbets- och näringsbyrån.
Läs mer: Studier i finska och svenska
Kurser i finska och svenska språketfinska _ engelska _ ryska
linkkiVanda vuxenutbildningsinstitut:
Kurser i finska och svenska språket för invandrarefinska
linkkiArbets- och näringsministeriet:
Utbildning i finska och svenska språketfinska _ svenska _ engelska
linkkiVanda vuxenutbildningsinstitut:
Grundundervisning för vuxnafinska
Samtal på finska
På Vanda stadsbibliotek anordnas språkcaféer (kielikahvila), där man kan öva på att prata finska.
Alla som vill lära sig tala finska är välkomna till caféerna.
På språkcaféerna talar vi finska, så det är bra om du redan kan lite finska.
Språkcaféerna är avgiftsfria.
Mer information om språkcaféerna får du från biblioteken.
I Vanda anordnas samtalsklubbar på finska också på Silkesportens verksamhetscenter (Silkinportin toimintakeskus) och Kafnettis och Myyrinkis boendeträffpunkter (Kafnetin ja Myyringin asukastila).
Finskaklubbar avsedda för föräldrar som vårdar barn i hemmet anordnas i invånarparkerna (asukaspuisto) och i de öppna daghemmen (avoin päiväkoti).
Klubbarna för att lära sig tala finska är avgiftsfria.
Läsundervisning
Nätverket Vi läser tillsammans (Luetaan yhdessä-verkosto) erbjuder undervisning i läsning och det finska språket för invandrarkvinnor.
Flera olika Vi läser tillsammans-nätverk är verksamma på olika håll i Vanda.
Det är avgiftsfritt att delta i grupperna.
Språkkaféerfinska _ engelska _ ryska
linkkiVanda stad:
Invånarlokalfinska _ engelska
linkkiVanda stad:
Invånarlokalfinska _ engelska
linkkiVanda stad:
Parker för invånare och öppna daghemfinska _ svenska _ engelska
linkkiVi läser tillsammans-nätverket:
Vi läser tillsammans i Vandafinska _ svenska _ engelska
Allmän språkexamen
Du kan avlägga allmän språkexamen i finska eller svenska språket.
På utbildningsstyrelsens (Opetushallitus) webbplats finns en sökmotor med vilken du kan kontrollera var och när du kan avlägga examen.
I Vanda ordnas språkexamina till exempel vid Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto).
Läs mer: Officiellt intyg på språkkunskaper.
linkkiUtbildningsstyrelsen:
Att anmäla sig till en allmän språkexamen och examensavgifterfinska _ svenska _ engelska
linkkiVanda vuxenutbildningsinstitut:
Allmän språkexamenfinska
linkkiUtbildningsstyrelsen:
Examenssökningfinska
Var hittar jag jobb?
Hjälp med jobbsökningen
Att starta ett företag
Beskattning
Var hittar jag jobb?
TE-byrån (TE-toimisto) hjälper dig att söka arbete.
Om du är arbetslös och söker efter arbete, ska du anmäla dig som arbetssökande hos TE-byrån.
Du kan anmäla dig antingen via nättjänsten eller personligen hos TE-byrån.
Medborgare i EU-länderna, Island, Liechtenstein och Schweiz kan anmäla sig som arbetssökande via TE-byråns nättjänst.
Övriga länders medborgare måste anmäla sig personligen hos TE-byrån.
Ta med dig din legitimation och ditt uppehållstillstånd.
Kontaktuppgifter:
Information om TE-byråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös.
Information om att söka arbete i Finland hittar du på InfoFinlands sida: Var hittar jag jobb?
linkkiVanda arbets- och näringsbyrå:
Kontaktuppgifter och tjänsterfinska _ svenska
linkkiArbets- och näringsministeriet:
Lediga jobbfinska _ svenska
linkkiArbets- och näringsförvaltningen:
Länkar till jobbsajterfinska _ svenska _ engelska
linkkiVanda stad:
Stöd för att hitta sysselsättningfinska _ svenska _ engelska
Hjälp med jobbsökningen
Stadens tjänster för arbetssökande
Vanda stad tillhandahåller olika tjänster för arbetslösa som hjälper dem att få kontakt med arbetslivet och hitta jobb.
I Vanda ordnas även många rekryteringsevenemang där arbetsgivarna söker arbetstagare.
Du hittar mer information om stadens tjänster på Vanda stads webbplats.
linkkiVanda stad:
Stadens tjänster för arbetssökandefinska _ svenska _ engelska
Om du behöver hjälp med jobbsökningen eller med att hitta en studieplats kan du kontakta rådgivarna i Håkansböle internationella förenings Tsemppari-projekt.
Du hittar kontaktuppgifterna på Håkansböle internationella förenings webbplats.
Integrationscentret Kotoutumiskeskus Monika hjälper arbetslösa invandrarkvinnor att hitta jobb.
Du kan få hjälp med att skriva din CV eller en jobbansökan, studera vardagsfinska och digitala färdigheter.
Luckan integration
Luckan Integration är en rådgivningstjänst, som erbjuder personlig rådgivning för invandrare och anordnar bland annat evenemang och grupper relaterade till jobbsökning.
Språket som talas vid träffarna är engelska.
Råd om jobbsökningfinska _ svenska _ engelska _ spanska
Väestöliittos karriärmentorskap är avsett för utbildade invandrare.
Via programmet kan du få en mentor, som stödjer dig i sökningen efter arbete eller utbildningsplats eller i att starta eget företag.
Verksamheten sker på finska.
Mentorskap i fråga om arbetskarriärfinska _ engelska
Om du är under 30 år, kan du få råd och handledning via tjänsten Navigatorn.
Personalen vid Navigatorn hjälper dig om du inte har något arbete eller en studieplats.
Stödföreningen för unga invandrare R3 (R3 Maahanmuuttajanuorten tuki ry) hjälper ungdomar i frågor som rör utbildning och sysselsättning.
Mer information hittar du på föreningens webbplats.
Stöd för unga invandrarefinska
Att starta ett företag
Om du har ett företag i Vanda, kan du bli medlem i Vanda Företagare.
Vanda Företagare rf är företagarnas intressebevakningsorganisation som erbjuder sina medlemmar till exempel utbildning och rådgivning.
Mer information hittar du på föreningens webbplats.
NewCo Helsinki erbjuder rådgivning och hjälp med att starta eget företag på finska, svenska, engelska, ryska, arabiska, estniska, tyska och italienska.
Vid NewCo Helsinki ordnas informationsmöten om att starta eget för invandrare på finska, engelska, ryska, arabiska och estniska.
Infomötena är avgiftsfria.
NewCo Helsinki ordnar företagarutbildningar på finska, engelska och ryska.
En del av kurserna är avsedda för personer som ska starta eget företag och en del för dem som redan har eget företag.
Kurser hålls på finska, engelska och ryska.
Mer information och anmälan finns på NewCo Helsinki webbplats.
Nylands TE-byrå (TE-toimisto) erbjuder mångsidiga tjänster för personer som funderar på att starta eget och dem som är på väg att starta eget.
På Nylands TE-byrå kan du till exempel delta i företagarutbildning och söka startpeng för att starta eget företag.
Läs mer: Att grunda ett företag
Tjänster för företagare med invandrarbakgrundfinska _ engelska
linkkiFöretagsFinland:
Företagsrådgivningfinska _ svenska _ engelska
Företagsrådgivningfinska _ engelska
Företagarnas intressebevakningsorganisationfinska
Beskattning
Huvudstadsregionens skattebyrå betjänar kunderna i centrala Helsingfors.
Kontaktuppgifter:
Alexandersgatan 9 (Gloet)
Tfn: 029 512 000
Invandrare kan även sköta ärenden vid servicestället International House Helsinki.
På servicestället hjälper FPA:s och Skatteförvaltningens experter invandrare som kommer till Finland för att arbeta i frågor som rör beskattning och social trygghet
Kontaktuppgifter till servicestället International House Helsinki:
Albertinkatu 25
Läs mer: Beskattning
linkkiSkatteförvaltningen:
Kontaktuppgifterfinska _ svenska _ engelska
Rådgivning om social trygghet och beskattningfinska _ svenska _ engelska
IHH – serviceställe för dig som flyttar till Finland engelska
Var hittar jag jobb?
Hjälp med jobbsökningen
Att starta ett företag
Beskattning
Var hittar jag jobb?
TE-byrån (TE-toimisto) hjälper dig att söka arbete.
Om du är arbetslös och söker efter arbete, ska du anmäla dig som arbetssökande hos TE-byrån.
Du kan anmäla dig antingen via nättjänsten eller personligen hos TE-byrån.
Medborgare i EU-länderna, Island, Liechtenstein och Schweiz kan anmäla sig som arbetssökande via TE-byråns nättjänst.
Övriga länders medborgare måste anmäla sig personligen hos TE-byrån.
Ta med dig din legitimation och ditt uppehållstillstånd.
Kontaktuppgifter:
Information om TE-byråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös.
Information om att söka arbete i Finland hittar du på InfoFinlands sida: Var hittar jag jobb?
linkkiVanda arbets- och näringsbyrå:
Kontaktuppgifter och tjänsterfinska _ svenska
linkkiArbets- och näringsministeriet:
Lediga jobbfinska _ svenska
linkkiArbets- och näringsförvaltningen:
Länkar till jobbsajterfinska _ svenska _ engelska
linkkiVanda stad:
Stöd för att hitta sysselsättningfinska _ svenska _ engelska
Hjälp med jobbsökningen
Stadens tjänster för arbetssökande
Vanda stad tillhandahåller olika tjänster för arbetslösa som hjälper dem att få kontakt med arbetslivet och hitta jobb.
I Vanda ordnas även många rekryteringsevenemang där arbetsgivarna söker arbetstagare.
Du hittar mer information om stadens tjänster på Vanda stads webbplats.
linkkiVanda stad:
Stadens tjänster för arbetssökandefinska _ svenska _ engelska
Om du behöver hjälp med jobbsökningen eller med att hitta en studieplats kan du kontakta rådgivarna i Håkansböle internationella förenings Tsemppari-projekt.
Du hittar kontaktuppgifterna på Håkansböle internationella förenings webbplats.
Integrationscentret Kotoutumiskeskus Monika hjälper arbetslösa invandrarkvinnor att hitta jobb.
Du kan få hjälp med att skriva din CV eller en jobbansökan, studera vardagsfinska och digitala färdigheter.
Luckan integration
Luckan Integration är en rådgivningstjänst, som erbjuder personlig rådgivning för invandrare och anordnar bland annat evenemang och grupper relaterade till jobbsökning.
Språket som talas vid träffarna är engelska.
Råd om jobbsökningfinska _ svenska _ engelska _ spanska
Väestöliittos karriärmentorskap är avsett för utbildade invandrare.
Via programmet kan du få en mentor, som stödjer dig i sökningen efter arbete eller utbildningsplats eller i att starta eget företag.
Verksamheten sker på finska.
Mentorskap i fråga om arbetskarriärfinska _ engelska
Om du är under 30 år, kan du få råd och handledning via tjänsten Navigatorn.
Personalen vid Navigatorn hjälper dig om du inte har något arbete eller en studieplats.
Stödföreningen för unga invandrare R3 (R3 Maahanmuuttajanuorten tuki ry) hjälper ungdomar i frågor som rör utbildning och sysselsättning.
Mer information hittar du på föreningens webbplats.
Stöd för unga invandrarefinska
Att starta ett företag
Om du har ett företag i Vanda, kan du bli medlem i Vanda Företagare.
Vanda Företagare rf är företagarnas intressebevakningsorganisation som erbjuder sina medlemmar till exempel utbildning och rådgivning.
Mer information hittar du på föreningens webbplats.
NewCo Helsinki erbjuder rådgivning och hjälp med att starta eget företag på finska, svenska, engelska, ryska, arabiska, estniska, tyska och italienska.
Vid NewCo Helsinki ordnas informationsmöten om att starta eget för invandrare på finska, engelska, ryska, arabiska och estniska.
Infomötena är avgiftsfria.
NewCo Helsinki ordnar företagarutbildningar på finska, engelska och ryska.
En del av kurserna är avsedda för personer som ska starta eget företag och en del för dem som redan har eget företag.
Kurser hålls på finska, engelska och ryska.
Mer information och anmälan finns på NewCo Helsinki webbplats.
Nylands TE-byrå (TE-toimisto) erbjuder mångsidiga tjänster för personer som funderar på att starta eget och dem som är på väg att starta eget.
På Nylands TE-byrå kan du till exempel delta i företagarutbildning och söka startpeng för att starta eget företag.
Läs mer: Att grunda ett företag
Tjänster för företagare med invandrarbakgrundfinska _ engelska
linkkiFöretagsFinland:
Företagsrådgivningfinska _ svenska _ engelska
Företagsrådgivningfinska _ engelska
Företagarnas intressebevakningsorganisationfinska
Beskattning
Huvudstadsregionens skattebyrå betjänar kunderna i centrala Helsingfors.
Kontaktuppgifter:
Alexandersgatan 9 (Gloet)
Tfn: 029 512 000
Invandrare kan även sköta ärenden vid servicestället International House Helsinki.
På servicestället hjälper FPA:s och Skatteförvaltningens experter invandrare som kommer till Finland för att arbeta i frågor som rör beskattning och social trygghet
Kontaktuppgifter till servicestället International House Helsinki:
Albertinkatu 25
Läs mer: Beskattning
linkkiSkatteförvaltningen:
Kontaktuppgifterfinska _ svenska _ engelska
Rådgivning om social trygghet och beskattningfinska _ svenska _ engelska
IHH – serviceställe för dig som flyttar till Finland engelska
Var hittar jag jobb?
Hjälp med jobbsökningen
Att starta ett företag
Beskattning
Var hittar jag jobb?
TE-byrån (TE-toimisto) hjälper dig att söka arbete.
Om du är arbetslös och söker efter arbete, ska du anmäla dig som arbetssökande hos TE-byrån.
Du kan anmäla dig antingen via nättjänsten eller personligen hos TE-byrån.
Medborgare i EU-länderna, Island, Liechtenstein och Schweiz kan anmäla sig som arbetssökande via TE-byråns nättjänst.
Övriga länders medborgare måste anmäla sig personligen hos TE-byrån.
Ta med dig din legitimation och ditt uppehållstillstånd.
Kontaktuppgifter:
Information om TE-byråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös.
Information om att söka arbete i Finland hittar du på InfoFinlands sida: Var hittar jag jobb?
linkkiVanda arbets- och näringsbyrå:
Kontaktuppgifter och tjänsterfinska _ svenska
linkkiArbets- och näringsministeriet:
Lediga jobbfinska _ svenska
linkkiArbets- och näringsförvaltningen:
Länkar till jobbsajterfinska _ svenska _ engelska
linkkiVanda stad:
Stöd för att hitta sysselsättningfinska _ svenska _ engelska
Hjälp med jobbsökningen
Stadens tjänster för arbetssökande
Vanda stad tillhandahåller olika tjänster för arbetslösa som hjälper dem att få kontakt med arbetslivet och hitta jobb.
I Vanda ordnas även många rekryteringsevenemang där arbetsgivarna söker arbetstagare.
Du hittar mer information om stadens tjänster på Vanda stads webbplats.
linkkiVanda stad:
Stadens tjänster för arbetssökandefinska _ svenska _ engelska
Om du behöver hjälp med jobbsökningen eller med att hitta en studieplats kan du kontakta rådgivarna i Håkansböle internationella förenings Tsemppari-projekt.
Du hittar kontaktuppgifterna på Håkansböle internationella förenings webbplats.
Integrationscentret Kotoutumiskeskus Monika hjälper arbetslösa invandrarkvinnor att hitta jobb.
Du kan få hjälp med att skriva din CV eller en jobbansökan, studera vardagsfinska och digitala färdigheter.
Luckan integration
Luckan Integration är en rådgivningstjänst, som erbjuder personlig rådgivning för invandrare och anordnar bland annat evenemang och grupper relaterade till jobbsökning.
Språket som talas vid träffarna är engelska.
Råd om jobbsökningfinska _ svenska _ engelska _ spanska
Väestöliittos karriärmentorskap är avsett för utbildade invandrare.
Via programmet kan du få en mentor, som stödjer dig i sökningen efter arbete eller utbildningsplats eller i att starta eget företag.
Verksamheten sker på finska.
Mentorskap i fråga om arbetskarriärfinska _ engelska
Om du är under 30 år, kan du få råd och handledning via tjänsten Navigatorn.
Personalen vid Navigatorn hjälper dig om du inte har något arbete eller en studieplats.
Stödföreningen för unga invandrare R3 (R3 Maahanmuuttajanuorten tuki ry) hjälper ungdomar i frågor som rör utbildning och sysselsättning.
Mer information hittar du på föreningens webbplats.
Stöd för unga invandrarefinska
Att starta ett företag
Om du har ett företag i Vanda, kan du bli medlem i Vanda Företagare.
Vanda Företagare rf är företagarnas intressebevakningsorganisation som erbjuder sina medlemmar till exempel utbildning och rådgivning.
Mer information hittar du på föreningens webbplats.
NewCo Helsinki erbjuder rådgivning och hjälp med att starta eget företag på finska, svenska, engelska, ryska, arabiska, estniska, tyska och italienska.
Vid NewCo Helsinki ordnas informationsmöten om att starta eget för invandrare på finska, engelska, ryska, arabiska och estniska.
Infomötena är avgiftsfria.
NewCo Helsinki ordnar företagarutbildningar på finska, engelska och ryska.
En del av kurserna är avsedda för personer som ska starta eget företag och en del för dem som redan har eget företag.
Kurser hålls på finska, engelska och ryska.
Mer information och anmälan finns på NewCo Helsinki webbplats.
Nylands TE-byrå (TE-toimisto) erbjuder mångsidiga tjänster för personer som funderar på att starta eget och dem som är på väg att starta eget.
På Nylands TE-byrå kan du till exempel delta i företagarutbildning och söka startpeng för att starta eget företag.
Läs mer: Att grunda ett företag
Tjänster för företagare med invandrarbakgrundfinska _ engelska
linkkiFöretagsFinland:
Företagsrådgivningfinska _ svenska _ engelska
Företagsrådgivningfinska _ engelska
Företagarnas intressebevakningsorganisationfinska
Beskattning
Huvudstadsregionens skattebyrå betjänar kunderna i centrala Helsingfors.
Kontaktuppgifter:
Alexandersgatan 9 (Gloet)
Tfn: 029 512 000
Invandrare kan även sköta ärenden vid servicestället International House Helsinki.
På servicestället hjälper FPA:s och Skatteförvaltningens experter invandrare som kommer till Finland för att arbeta i frågor som rör beskattning och social trygghet
Kontaktuppgifter till servicestället International House Helsinki:
Albertinkatu 25
Läs mer: Beskattning
linkkiSkatteförvaltningen:
Kontaktuppgifterfinska _ svenska _ engelska
Rådgivning om social trygghet och beskattningfinska _ svenska _ engelska
IHH – serviceställe för dig som flyttar till Finland engelska
Rådgivning för och integration av invandrare
Inledande kartläggning
Behöver du en tolk?
Rådgivning för och integration av invandrare
Invandrartjänster
Vanda stads tjänster för invandrare omfattar
mottagningstjänster för invandrare
integrationstjänster
Vanda stads tjänster för invandrare (Vantaan maahanmuuttajapalvelut) ger dig information om integration, social- och hälsovårdstjänster och om stadens och olika organisationers tjänster.
Du kan bli klient om du flyttat till Finland på grund av familjeband, är flykting, offer för människohandel eller har rätt till en inledande kartläggning.
Tfn (09) 839 21074 och (09) 839 32042
linkkiVanda stad:
Invandrartjänsterfinska _ engelska
Verksamhetscentret Silkesporten (Silkinportin toimintakeskus) ger rådgivning för invandrare och där ordnas många slags aktiviteter.
dickursbyvägen 44 F, vån.
Tfn (09) 839 23651
linkkiSilkesportens verksamhetscenter:
Rådgivning och verksamhet för invandrarefinska _ engelska
Vandainfo ger dig information om såväl Vandas stads som statens tjänster.
Vandainfon finns i Dickursby, Korso och Myrbacka.
Adresserna är:
Dixi, Banvägen 11, 2:a vån.
tfn (09) 839 22133
Tfn (09) 839 22133
Tfn (09) 839 22133
Kontaktuppgifterna och öppettiderna hittar du på Vanda stads webbplats.
linkkiVanda stad:
Vandainfofinska _ svenska _ engelska
Den internationella föreningen i Håkansböle (Hakunilan kansainvälinen yhdistys) har en rådgivningspunkt som betjänar invandrare i Håkansböle, Björkby och andra områden i Vanda, som vill ha information om till exempel studier, språkkurser, arbete, hobbyverksamhet, krissituationer eller juridiska frågor.
Sporrgränden 2 A, vån. 3 (Håkansböle)
Tfn (09) 272 2775 och 040 501 3199.
linkkiInternationella föreningen i Håkansböle:
Rådgivning för invandrarefinska _ engelska _ ryska _ somaliska _ arabiska
På invandrarrådgivningen vid föreningen Vantaan Järjestörinki ry (Vantaan Järjestörinki ry:n Maahanmuuttajien neuvontapiste) kan du fråga om sådant som rör till exempel arbetslivet, social trygghet, hälsa, utbildning och uppehållstillstånd.
Adress:
Ranunkelvägen 22
Asukastila Myyrinki
Eldstadstorget 1 eller Kopparbergsvägen 10 B, vån.
Vanda Tfn (09) 839 35703 och 040 183 0930
Rautbergsgatan 3
Tfn 045 134 1711
Rådgivning för invandrarefinska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
IHH – serviceställe för dig som flyttar till Finland engelska
Inledande kartläggning
Den inledande kartläggningen (alkukartoitus) hjälper dig att hitta lämpliga tjänster i din hemstad.
Vanda stad eller Nylands TE-byrå ordnar en inledande kartläggning för varje ny invandrare i Vanda.
Du har rätt att få en inledande kartläggning om
din hemkommun är Vanda
du har flyttat till Vanda från ett annat land eller en annan ort i Finland
någon inledande kartläggning inte har gjorts för dig tidigare
du har haft hemkommun i Finland i högst tre år.
I den inledande kartläggningen får du information om utbildning i finska eller svenska, arbetssökning, utbildning och tjänster i Vanda.
Vid den inledande kartläggningen talas man vid med hjälp av tolk.
Den inledande kartläggningen är avgiftsfri.
Begäran om inledande kartläggning
Du kan begära en inledande kartläggning via e-post eller så kan du boka en tid per telefon.
Tfn 09 839 32622, 09 839 27525 eller 09 839 31766
Om du söker arbete, bör du anmäla dig till TE-byrån.
TE-byrån gör den inledande kartläggningen.
Läs mer om den inledande kartläggningen och integrationsplanen på InfoFinlands webbplats Integration i Finland
linkkiVanda stad:
Inledande kartläggningfinska _ engelska
Behöver du en tolk?
Om du måste sköta ärenden med myndigheter, men inte kan finska eller svenska och det inte heller finns något annat språk som både du och myndigheten talar, kan du använda en tolktjänst.
Meddela alltid myndigheten i förväg om du behöver en tolk.
Myndigheten bokar tolken och då får du tolkningstjänsten gratis.
Om du själv bokar tolken och betalar kostnaderna, kan du anlita en tolk när som helst.
Läs mer: Behöver du en tolk?
linkkiVanda stad:
Information om tolktjänsterfinska
linkkiFinlands översättar- och tolkförbund:
Sök tolk eller översättarefinska _ svenska _ engelska
Rådgivning för och integration av invandrare
Inledande kartläggning
Behöver du en tolk?
Rådgivning för och integration av invandrare
Invandrartjänster
Vanda stads tjänster för invandrare omfattar
mottagningstjänster för invandrare
integrationstjänster
Vanda stads tjänster för invandrare (Vantaan maahanmuuttajapalvelut) ger dig information om integration, social- och hälsovårdstjänster och om stadens och olika organisationers tjänster.
Du kan bli klient om du flyttat till Finland på grund av familjeband, är flykting, offer för människohandel eller har rätt till en inledande kartläggning.
Tfn (09) 839 21074 och (09) 839 32042
linkkiVanda stad:
Invandrartjänsterfinska _ engelska
Verksamhetscentret Silkesporten (Silkinportin toimintakeskus) ger rådgivning för invandrare och där ordnas många slags aktiviteter.
dickursbyvägen 44 F, vån.
Tfn (09) 839 23651
linkkiSilkesportens verksamhetscenter:
Rådgivning och verksamhet för invandrarefinska _ engelska
Vandainfo ger dig information om såväl Vandas stads som statens tjänster.
Vandainfon finns i Dickursby, Korso och Myrbacka.
Adresserna är:
Dixi, Banvägen 11, 2:a vån.
tfn (09) 839 22133
Tfn (09) 839 22133
Tfn (09) 839 22133
Kontaktuppgifterna och öppettiderna hittar du på Vanda stads webbplats.
linkkiVanda stad:
Vandainfofinska _ svenska _ engelska
Den internationella föreningen i Håkansböle (Hakunilan kansainvälinen yhdistys) har en rådgivningspunkt som betjänar invandrare i Håkansböle, Björkby och andra områden i Vanda, som vill ha information om till exempel studier, språkkurser, arbete, hobbyverksamhet, krissituationer eller juridiska frågor.
Sporrgränden 2 A, vån. 3 (Håkansböle)
Tfn (09) 272 2775 och 040 501 3199.
linkkiInternationella föreningen i Håkansböle:
Rådgivning för invandrarefinska _ engelska _ ryska _ somaliska _ arabiska
På invandrarrådgivningen vid föreningen Vantaan Järjestörinki ry (Vantaan Järjestörinki ry:n Maahanmuuttajien neuvontapiste) kan du fråga om sådant som rör till exempel arbetslivet, social trygghet, hälsa, utbildning och uppehållstillstånd.
Adress:
Ranunkelvägen 22
Asukastila Myyrinki
Eldstadstorget 1 eller Kopparbergsvägen 10 B, vån.
Vanda Tfn (09) 839 35703 och 040 183 0930
Rautbergsgatan 3
Tfn 045 134 1711
Rådgivning för invandrarefinska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
IHH – serviceställe för dig som flyttar till Finland engelska
Inledande kartläggning
Den inledande kartläggningen (alkukartoitus) hjälper dig att hitta lämpliga tjänster i din hemstad.
Vanda stad eller Nylands TE-byrå ordnar en inledande kartläggning för varje ny invandrare i Vanda.
Du har rätt att få en inledande kartläggning om
din hemkommun är Vanda
du har flyttat till Vanda från ett annat land eller en annan ort i Finland
någon inledande kartläggning inte har gjorts för dig tidigare
du har haft hemkommun i Finland i högst tre år.
I den inledande kartläggningen får du information om utbildning i finska eller svenska, arbetssökning, utbildning och tjänster i Vanda.
Vid den inledande kartläggningen talas man vid med hjälp av tolk.
Den inledande kartläggningen är avgiftsfri.
Begäran om inledande kartläggning
Du kan begära en inledande kartläggning via e-post eller så kan du boka en tid per telefon.
Tfn 09 839 32622, 09 839 27525 eller 09 839 31766
Om du söker arbete, bör du anmäla dig till TE-byrån.
TE-byrån gör den inledande kartläggningen.
Läs mer om den inledande kartläggningen och integrationsplanen på InfoFinlands webbplats Integration i Finland
linkkiVanda stad:
Inledande kartläggningfinska _ engelska
Behöver du en tolk?
Om du måste sköta ärenden med myndigheter, men inte kan finska eller svenska och det inte heller finns något annat språk som både du och myndigheten talar, kan du använda en tolktjänst.
Meddela alltid myndigheten i förväg om du behöver en tolk.
Myndigheten bokar tolken och då får du tolkningstjänsten gratis.
Om du själv bokar tolken och betalar kostnaderna, kan du anlita en tolk när som helst.
Läs mer: Behöver du en tolk?
linkkiVanda stad:
Information om tolktjänsterfinska
linkkiFinlands översättar- och tolkförbund:
Sök tolk eller översättarefinska _ svenska _ engelska
Rådgivning för och integration av invandrare
Inledande kartläggning
Behöver du en tolk?
Rådgivning för och integration av invandrare
Invandrartjänster
Vanda stads tjänster för invandrare omfattar
mottagningstjänster för invandrare
integrationstjänster
Vanda stads tjänster för invandrare (Vantaan maahanmuuttajapalvelut) ger dig information om integration, social- och hälsovårdstjänster och om stadens och olika organisationers tjänster.
Du kan bli klient om du flyttat till Finland på grund av familjeband, är flykting, offer för människohandel eller har rätt till en inledande kartläggning.
Tfn (09) 839 21074 och (09) 839 32042
linkkiVanda stad:
Invandrartjänsterfinska _ engelska
Vandainfo ger dig information om såväl Vandas stads som statens tjänster.
Vandainfon finns i Dickursby, Korso och Myrbacka.
Adresserna är:
Dixi, Banvägen 11, 2:a vån.
tfn (09) 839 22133
Tfn (09) 839 22133
Tfn (09) 839 22133
Kontaktuppgifterna och öppettiderna hittar du på Vanda stads webbplats.
linkkiVanda stad:
Vandainfofinska _ svenska _ engelska
Den internationella föreningen i Håkansböle (Hakunilan kansainvälinen yhdistys) har en rådgivningspunkt som betjänar invandrare i Håkansböle, Björkby och andra områden i Vanda, som vill ha information om till exempel studier, språkkurser, arbete, hobbyverksamhet, krissituationer eller juridiska frågor.
Sporrgränden 2 A, vån. 3 (Håkansböle)
Tfn (09) 272 2775 och 040 501 3199.
linkkiInternationella föreningen i Håkansböle:
Rådgivning för invandrarefinska _ engelska _ ryska _ somaliska _ arabiska
På invandrarrådgivningen vid föreningen Vantaan Järjestörinki ry (Vantaan Järjestörinki ry:n Maahanmuuttajien neuvontapiste) kan du fråga om sådant som rör till exempel arbetslivet, social trygghet, hälsa, utbildning och uppehållstillstånd.
Adress:
Ranunkelvägen 22
Asukastila Myyrinki
Eldstadstorget 1 eller Kopparbergsvägen 10 B, vån.
Vanda Tfn (09) 839 35703 och 040 183 0930
Rautbergsgatan 3
Tfn 045 134 1711
Rådgivning för invandrarefinska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
IHH – serviceställe för dig som flyttar till Finland engelska
Inledande kartläggning
Den inledande kartläggningen (alkukartoitus) hjälper dig att hitta lämpliga tjänster i din hemstad.
Vanda stad eller Nylands TE-byrå ordnar en inledande kartläggning för varje ny invandrare i Vanda.
Du har rätt att få en inledande kartläggning om
din hemkommun är Vanda
du har flyttat till Vanda från ett annat land eller en annan ort i Finland
någon inledande kartläggning inte har gjorts för dig tidigare
du har haft hemkommun i Finland i högst tre år.
I den inledande kartläggningen får du information om utbildning i finska eller svenska, arbetssökning, utbildning och tjänster i Vanda.
Vid den inledande kartläggningen talas man vid med hjälp av tolk.
Den inledande kartläggningen är avgiftsfri.
Begäran om inledande kartläggning
Du kan begära en inledande kartläggning via e-post eller så kan du boka en tid per telefon.
Tfn 09 839 32622, 09 839 27525 eller 09 839 31766
Om du söker arbete, bör du anmäla dig till TE-byrån.
TE-byrån gör den inledande kartläggningen.
Läs mer om den inledande kartläggningen och integrationsplanen på InfoFinlands webbplats Integration i Finland
linkkiVanda stad:
Inledande kartläggningfinska _ engelska
Behöver du en tolk?
Om du måste sköta ärenden med myndigheter, men inte kan finska eller svenska och det inte heller finns något annat språk som både du och myndigheten talar, kan du använda en tolktjänst.
Meddela alltid myndigheten i förväg om du behöver en tolk.
Myndigheten bokar tolken och då får du tolkningstjänsten gratis.
Om du själv bokar tolken och betalar kostnaderna, kan du anlita en tolk när som helst.
Läs mer: Behöver du en tolk?
linkkiVanda stad:
Information om tolktjänsterfinska
linkkiFinlands översättar- och tolkförbund:
Sök tolk eller översättarefinska _ svenska _ engelska
Tillståndsärenden
På Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU-medborgarens uppehållsrätt.
Migrationsverkets tjänsteställe i Helsingfors :
Göksgränd 3A
Du kan också ansöka om många slags uppehållstillstånd och EU-registrering på internet i tjänsten Enter Finland.
Om du inte är van vid att använda en dator, fyll i en ansökan på papper och lämna in den på Migrationsverkets tjänsteställe.
Dät är alltid bra att boka en tid i förväg på tjänstestället.
Du kan boka en tid på Migrationsverkets tidsbokningstjänst.
Observera att tjänstestället inte kan ge rådgivning om tillståndsärenden.
Läs mer: Flytta till Finland.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Registrering som invånare
Om du flyttar ditt stadigvarande boende till Vanda, ska du registrera dig som invånare i kommunen.
Du kan registrera dig vid magistraten.
Albertsgatan 25
Växel 029 55 39391
Registrering av utlänningar 029 55 36 300
När du går till magistraten ska du ta med dig
legitimation (till exempel pass)
uppehållstillstånd och uppehållskort (om du behöver uppehållstillstånd i Finland)
registreringsintyget över uppehållsrätten (oleskeluoikeuden rekisteröintitodistus) om du är EU-medborgare.
äktenskapsintyg
dina barns födelseattester.
Observera att utländska handlingar ska vara legaliserade.
Du får mer information om att legalisera officiella handlingar vid magistraten eller beskickningen för ditt eget land i Finland.
Läs mer: Registrering som invånare.
Registrering av utlänningarfinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
Du kan få:
kostnadsfri rådgivning och information kring att flytta på flera olika språk
en finländsk personbeteckning, registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1-intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
Adress
Albertsgatan 25
IHH – serviceställe för dig som flyttar till Finland engelska
Webbappen IHH Service Advisor App engelska
Tillståndsärenden
På Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU-medborgarens uppehållsrätt.
Migrationsverkets tjänsteställe i Helsingfors :
Göksgränd 3A
Du kan också ansöka om många slags uppehållstillstånd och EU-registrering på internet i tjänsten Enter Finland.
Om du inte är van vid att använda en dator, fyll i en ansökan på papper och lämna in den på Migrationsverkets tjänsteställe.
Dät är alltid bra att boka en tid i förväg på tjänstestället.
Du kan boka en tid på Migrationsverkets tidsbokningstjänst.
Observera att tjänstestället inte kan ge rådgivning om tillståndsärenden.
Läs mer: Flytta till Finland.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Registrering som invånare
Om du flyttar ditt stadigvarande boende till Vanda, ska du registrera dig som invånare i kommunen.
Du kan registrera dig vid magistraten.
Albertsgatan 25
Växel 029 55 39391
Registrering av utlänningar 029 55 36 300
När du går till magistraten ska du ta med dig
legitimation (till exempel pass)
uppehållstillstånd och uppehållskort (om du behöver uppehållstillstånd i Finland)
registreringsintyget över uppehållsrätten (oleskeluoikeuden rekisteröintitodistus) om du är EU-medborgare.
äktenskapsintyg
dina barns födelseattester.
Observera att utländska handlingar ska vara legaliserade.
Du får mer information om att legalisera officiella handlingar vid magistraten eller beskickningen för ditt eget land i Finland.
Läs mer: Registrering som invånare.
Registrering av utlänningarfinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
Du kan få:
kostnadsfri rådgivning och information kring att flytta på flera olika språk
en finländsk personbeteckning, registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1-intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
Adress
IHH – serviceställe för dig som flyttar till Finland engelska
Webbappen IHH Service Advisor App engelska
Tillståndsärenden
På Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU-medborgarens uppehållsrätt.
Migrationsverkets tjänsteställe i Helsingfors :
Göksgränd 3A
Du kan också ansöka om många slags uppehållstillstånd och EU-registrering på internet i tjänsten Enter Finland.
Om du inte är van vid att använda en dator, fyll i en ansökan på papper och lämna in den på Migrationsverkets tjänsteställe.
Dät är alltid bra att boka en tid i förväg på tjänstestället.
Du kan boka en tid på Migrationsverkets tidsbokningstjänst.
Observera att tjänstestället inte kan ge rådgivning om tillståndsärenden.
Läs mer: Flytta till Finland.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Registrering som invånare
Om du flyttar ditt stadigvarande boende till Vanda, ska du registrera dig som invånare i kommunen.
Du kan registrera dig vid magistraten.
Albertsgatan 25
Växel 029 55 39391
Registrering av utlänningar 029 55 36 300
När du går till magistraten ska du ta med dig
legitimation (till exempel pass)
uppehållstillstånd och uppehållskort (om du behöver uppehållstillstånd i Finland)
registreringsintyget över uppehållsrätten (oleskeluoikeuden rekisteröintitodistus) om du är EU-medborgare.
äktenskapsintyg
dina barns födelseattester.
Observera att utländska handlingar ska vara legaliserade.
Du får mer information om att legalisera officiella handlingar vid magistraten eller beskickningen för ditt eget land i Finland.
Läs mer: Registrering som invånare.
Registrering av utlänningarfinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
Du kan få:
kostnadsfri rådgivning och information kring att flytta på flera olika språk
en finländsk personbeteckning, registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1-intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
Adress
IHH – serviceställe för dig som flyttar till Finland engelska
Webbappen IHH Service Advisor App engelska
Trafik
Beslutsfattande och påverkan
Religion
Grundläggande information
Historia
Trafik
Kollektivtrafiken
Esbo och hela huvudstadsregionen har goda kollektivtrafikförbindelser.
I Esbo finns flera tåg- och metrostationer.
I staden finns flera busslinjer.
Information och råd till resenärerfinska _ svenska _ engelska
Esbo tillhör samkommunen Helsingforsregionens trafik HRT (HSL), som ordnar kollektivtrafiken i huvudstadsregionen.
Du kan söka information om rutterna i reseplanerartjänsten (Reittiopas).
Tjänsten ger dig råd om olika kollektivtrafikförbindelser från ett ställe till ett annat.
Reseplanerarefinska _ svenska _ engelska _ ryska
I kollektivtrafiken kan du betala med kontanter eller resekort.
I närtågen måste du köpa biljetten i förväg.
Mer information om resekorten och deras försäljningsställen i Esbo hittar du på HRT:s webbplats.
Du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat.
Biljetter och priserfinska _ svenska _ engelska
Att gå och cykla
Om du vill gå eller cykla i Esbo kan du söka en lämplig rutt i reseplaneraren för cykling och gång.
Resplan för cycling och gångfinska _ svenska _ engelska _ ryska
Cykelkartor för Helsingfors, Vanda och Esbo delas ut vid samservicekontoren och idrottsverkens serviceställen.
Cykelkartorna är kostnadsfria.
Friluftskartafinska
Bil och flyg
Du kan parkera bilen på många järnvägsstationer och fortsätta färden med kollektivtrafiken.
Helsingfors-Vanda flygplats ligger Esbos grannkommun Vanda.
Läs mer: Trafik.
linkkiEsbo stad:
Trafikfinska _ svenska _ engelska
linkkiEsbo stad:
Kartorfinska _ svenska _ engelska
Beslutsfattande och påverkan
I Esbo beslutas ärenden av stadsfullmäktige.
I stadsfullmäktige sitter 75 ledamöter som representerar olika politiska grupper.
Fullmäktige väljs var fjärde år genom kommunalval.
Invånarna i Esbo kan påverka beslutsfattandet och beredning av ärenden på många olika sätt.
Du kan ge respons till beslutsfattarna och tjänstemännen till exempel via det elektroniska responssystemet.
Du kan vara med i invånarverksamheten eller ta ett invånarinitiativ.
Läs mer om hur du kan påverka på Esbo stads webbplats.
I Esbo finns en delegation för mångkulturella frågor som utvecklar stadens mångkulturella politik.
I Esbo finns många politiska föreningar, invandrarföreningar och andra föreningar via vilka du också kan påverka beslutsfattandet.
Läs mer: Beslutsfattande och påverkan
linkkiEsbo stad:
Information om beslutsfattandefinska _ svenska _ engelska
linkkiEsbo stad:
Information om påverkanfinska _ svenska _ engelska
linkkiEsbo stad:
Elektroniskt responssystemfinska _ svenska _ engelska
linkkiEsbo stad:
Mångkulturella ärendenfinska _ svenska _ engelska
Religion
Många religiösa samfund är verksamma i Esbo och Helsingfors.
Via tjänsten Uskonnot Suomessa kan du söka information efter det religiösa samfundet och orten.
Läs mer: Kulturer och religioner i Finland.
Religiösa samfundfinska _ engelska
linkkiEsbo kyrkliga samfällighet:
Evangelisk-lutherska församlingarfinska _ svenska _ engelska
linkkiHelsingfors ortodoxa församling:
Ortodoxa församlingenfinska _ ryska
Grundläggande information
Esbo är en av huvudstadsregionens fyra kommuner.
Det ligger bredvid Helsingfors, väster om staden.
Utöver dessa finns det flera mindre tätorter, landsbygd och skogar i Esbo.
Esbo har cirka 280 000 invånare.
De flesta invånarna är finskspråkiga.
Ungefär 7 procent av invånarna är svenskspråkiga och 16 procent har andra modersmål.
Esbos areal är cirka 528 km2, varav cirka 216 km2 är vatten.
linkkiEsbo stad:
Information om Esbofinska _ svenska _ engelska
Historia
Esboområdet var bebott redan för ungefär 8 000 år sedan.
Då var södra Esbo fortfarande hav.
På 1200-talet flyttade många emigranter från Sverige till Esbo.
På 1400-talet blev Esbo en självständig socken med många byar.
I Esbo byggdes stora herrgårdar som hade stor betydelse för områdets utveckling.
När Finland blev en del av Ryssland blev Helsingfors huvudstad år 1812.
Även om Helsingfors växte snabbt, var Esbo ännu länge en fridfull landssocken.
Inflyttningen till Esbo blev livligare från och med 1940-talet.
År 1950 hade Esbo 25 000 invånare och 15 år senare redan 65 000 invånare.
Esbo blev en stad år 1972.
linkkiEsbo stad:
Historiafinska _ svenska
linkkiEsbo stad:
Museerfinska _ svenska _ engelska
Trafik
Beslutsfattande och påverkan
Religion
Grundläggande information
Historia
Trafik
Kollektivtrafiken
Esbo och hela huvudstadsregionen har goda kollektivtrafikförbindelser.
I Esbo finns flera tåg- och metrostationer.
I staden finns flera busslinjer.
Information och råd till resenärerfinska _ svenska _ engelska
Esbo tillhör samkommunen Helsingforsregionens trafik HRT (HSL), som ordnar kollektivtrafiken i huvudstadsregionen.
Du kan söka information om rutterna i reseplanerartjänsten (Reittiopas).
Tjänsten ger dig råd om olika kollektivtrafikförbindelser från ett ställe till ett annat.
Reseplanerarefinska _ svenska _ engelska _ ryska
I kollektivtrafiken kan du betala med kontanter eller resekort.
I närtågen måste du köpa biljetten i förväg.
Mer information om resekorten och deras försäljningsställen i Esbo hittar du på HRT:s webbplats.
Du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat.
Biljetter och priserfinska _ svenska _ engelska
Att gå och cykla
Om du vill gå eller cykla i Esbo kan du söka en lämplig rutt i reseplaneraren för cykling och gång.
Resplan för cycling och gångfinska _ svenska _ engelska _ ryska
Cykelkartor för Helsingfors, Vanda och Esbo delas ut vid samservicekontoren och idrottsverkens serviceställen.
Cykelkartorna är kostnadsfria.
Friluftskartafinska
Bil och flyg
Du kan parkera bilen på många järnvägsstationer och fortsätta färden med kollektivtrafiken.
Helsingfors-Vanda flygplats ligger Esbos grannkommun Vanda.
Läs mer: Trafik.
linkkiEsbo stad:
Trafikfinska _ svenska _ engelska
linkkiEsbo stad:
Kartorfinska _ svenska _ engelska
Beslutsfattande och påverkan
I Esbo beslutas ärenden av stadsfullmäktige.
I stadsfullmäktige sitter 75 ledamöter som representerar olika politiska grupper.
Fullmäktige väljs var fjärde år genom kommunalval.
Invånarna i Esbo kan påverka beslutsfattandet och beredning av ärenden på många olika sätt.
Du kan ge respons till beslutsfattarna och tjänstemännen till exempel via det elektroniska responssystemet.
Du kan vara med i invånarverksamheten eller ta ett invånarinitiativ.
Läs mer om hur du kan påverka på Esbo stads webbplats.
I Esbo finns en delegation för mångkulturella frågor som utvecklar stadens mångkulturella politik.
I Esbo finns många politiska föreningar, invandrarföreningar och andra föreningar via vilka du också kan påverka beslutsfattandet.
Läs mer: Beslutsfattande och påverkan
linkkiEsbo stad:
Information om beslutsfattandefinska _ svenska _ engelska
linkkiEsbo stad:
Information om påverkanfinska _ svenska _ engelska
linkkiEsbo stad:
Elektroniskt responssystemfinska _ svenska _ engelska
linkkiEsbo stad:
Mångkulturella ärendenfinska _ svenska _ engelska
Religion
Många religiösa samfund är verksamma i Esbo och Helsingfors.
Via tjänsten Uskonnot Suomessa kan du söka information efter det religiösa samfundet och orten.
Läs mer: Kulturer och religioner i Finland.
Religiösa samfundfinska _ engelska
linkkiEsbo kyrkliga samfällighet:
Evangelisk-lutherska församlingarfinska _ svenska _ engelska
linkkiHelsingfors ortodoxa församling:
Ortodoxa församlingenfinska _ ryska
Grundläggande information
Esbo är en av huvudstadsregionens fyra kommuner.
Det ligger bredvid Helsingfors, väster om staden.
Utöver dessa finns det flera mindre tätorter, landsbygd och skogar i Esbo.
Esbo har cirka 280 000 invånare.
De flesta invånarna är finskspråkiga.
Ungefär 7 procent av invånarna är svenskspråkiga och 16 procent har andra modersmål.
Esbos areal är cirka 528 km2, varav cirka 216 km2 är vatten.
linkkiEsbo stad:
Information om Esbofinska _ svenska _ engelska
Historia
Esboområdet var bebott redan för ungefär 8 000 år sedan.
Då var södra Esbo fortfarande hav.
På 1200-talet flyttade många emigranter från Sverige till Esbo.
På 1400-talet blev Esbo en självständig socken med många byar.
I Esbo byggdes stora herrgårdar som hade stor betydelse för områdets utveckling.
När Finland blev en del av Ryssland blev Helsingfors huvudstad år 1812.
Även om Helsingfors växte snabbt, var Esbo ännu länge en fridfull landssocken.
Inflyttningen till Esbo blev livligare från och med 1940-talet.
År 1950 hade Esbo 25 000 invånare och 15 år senare redan 65 000 invånare.
Esbo blev en stad år 1972.
linkkiEsbo stad:
Historiafinska _ svenska
linkkiEsbo stad:
Museerfinska _ svenska _ engelska
Trafik
Beslutsfattande och påverkan
Religion
Grundläggande information
Historia
Trafik
Kollektivtrafiken
Esbo och hela huvudstadsregionen har goda kollektivtrafikförbindelser.
I Esbo finns flera tåg- och metrostationer.
I staden finns flera busslinjer.
Information och råd till resenärerfinska _ svenska _ engelska
Esbo tillhör samkommunen Helsingforsregionens trafik HRT (HSL), som ordnar kollektivtrafiken i huvudstadsregionen.
Du kan söka information om rutterna i reseplanerartjänsten (Reittiopas).
Tjänsten ger dig råd om olika kollektivtrafikförbindelser från ett ställe till ett annat.
Reseplanerarefinska _ svenska _ engelska
I kollektivtrafiken kan du betala med kontanter eller resekort.
I närtågen måste du köpa biljetten i förväg.
Mer information om resekorten och deras försäljningsställen i Esbo hittar du på HRT:s webbplats.
Du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat.
Biljetter och priserfinska _ svenska _ engelska
Att gå och cykla
Om du vill gå eller cykla i Esbo kan du söka en lämplig rutt i reseplaneraren för cykling och gång.
Resplan för cycling och gångfinska _ svenska _ engelska _ ryska
Bil och flyg
Du kan parkera bilen på många järnvägsstationer och fortsätta färden med kollektivtrafiken.
Helsingfors-Vanda flygplats ligger Esbos grannkommun Vanda.
Läs mer: Trafik.
linkkiEsbo stad:
Trafikfinska _ svenska _ engelska
linkkiEsbo stad:
Kartorfinska _ svenska _ engelska
Beslutsfattande och påverkan
I Esbo beslutas ärenden av stadsfullmäktige.
I stadsfullmäktige sitter 75 ledamöter som representerar olika politiska grupper.
Fullmäktige väljs var fjärde år genom kommunalval.
Invånarna i Esbo kan påverka beslutsfattandet och beredning av ärenden på många olika sätt.
Du kan ge respons till beslutsfattarna och tjänstemännen till exempel via det elektroniska responssystemet.
Du kan vara med i invånarverksamheten eller ta ett invånarinitiativ.
Läs mer om hur du kan påverka på Esbo stads webbplats.
I Esbo finns en delegation för mångkulturella frågor som utvecklar stadens mångkulturella politik.
I Esbo finns många politiska föreningar, invandrarföreningar och andra föreningar via vilka du också kan påverka beslutsfattandet.
Läs mer: Beslutsfattande och påverkan
linkkiEsbo stad:
Information om beslutsfattandefinska _ svenska _ engelska
linkkiEsbo stad:
Information om påverkanfinska _ svenska _ engelska
linkkiEsbo stad:
Elektroniskt responssystemfinska _ svenska _ engelska
linkkiEsbo stad:
Mångkulturella ärendenfinska _ svenska _ engelska
Religion
Många religiösa samfund är verksamma i Esbo och Helsingfors.
Via tjänsten Uskonnot Suomessa kan du söka information efter det religiösa samfundet och orten.
Läs mer: Kulturer och religioner i Finland.
Religiösa samfundfinska _ engelska
linkkiEsbo kyrkliga samfällighet:
Evangelisk-lutherska församlingarfinska _ svenska _ engelska
linkkiHelsingfors ortodoxa församling:
Ortodoxa församlingenfinska _ ryska
Grundläggande information
Esbo är en av huvudstadsregionens fyra kommuner.
Det ligger bredvid Helsingfors, väster om staden.
Utöver dessa finns det flera mindre tätorter, landsbygd och skogar i Esbo.
Esbo har cirka 280 000 invånare.
De flesta invånarna är finskspråkiga.
Ungefär 7 procent av invånarna är svenskspråkiga och 16 procent har andra modersmål.
Esbos areal är cirka 528 km2, varav cirka 216 km2 är vatten.
linkkiEsbo stad:
Information om Esbofinska _ svenska _ engelska
Historia
Esboområdet var bebott redan för ungefär 8 000 år sedan.
Då var södra Esbo fortfarande hav.
På 1200-talet flyttade många emigranter från Sverige till Esbo.
På 1400-talet blev Esbo en självständig socken med många byar.
I Esbo byggdes stora herrgårdar som hade stor betydelse för områdets utveckling.
När Finland blev en del av Ryssland blev Helsingfors huvudstad år 1812.
Även om Helsingfors växte snabbt, var Esbo ännu länge en fridfull landssocken.
Inflyttningen till Esbo blev livligare från och med 1940-talet.
År 1950 hade Esbo 25 000 invånare och 15 år senare redan 65 000 invånare.
Esbo blev en stad år 1972.
linkkiEsbo stad:
Historiafinska _ svenska
linkkiEsbo stad:
Museerfinska _ svenska _ engelska
Evenemang
Bibliotek
Motion
Att röra sig i naturen
Teater och film
Museer
Fritidsverksamhet för barn och unga
Föreningar
I Esbo finns många hobbymöjligheter.
Invånarhusen Kivenkolo och Kylämaja är öppna för alla.
I invånarhusen kan områdets invånare vistas och samlas samt få anvisningar och råd.
Invånarhuset Kivenkolo
Sjöstöveln 1 A
linkkiEsbo stad:
Kivenkolo invånarhusfinska _ svenska _ engelska
Invånarhuset Kylämaja
Mattsgatan 7
linkkiEsbo stad:
Invånarhus Kylämajafinska
Vid Esbo arbetarinstitut (Espoon työväenopisto) kan man till exempel skapa konst, handarbeten, laga mat, dansa eller idka motion.
Där kan man även studera finska och andra språk.
linkkiEsbo stad:
Arbetarinstitutetfinska _ svenska _ engelska
I Esbo finns flera läroanstalter som ger grundundervisning i konstämnen speciellt för barn och unga.
Olika konstarter är musik, bildkonst, dans, teater och cirkus.
linkkiEsbo stad:
Konstundervisningfinska _ engelska.
Konsthuset Lilla Aurora ordnar kulturevenemang för barn.
linkkiEsbo stad:
Kulturevenemang för barnfinska _ svenska _ engelska
Läs mer: Fritid.
Evenemang
Evenemangfinska _ svenska _ engelska _ ryska _ kinesiska
linkkiEsbo stad:
Evenemangfinska
Bibliotek
I Esbo finns flera bibliotek på olika håll i staden.
På biblioteket kan du låna böcker, tidningar, musik, filmer, spel och mycket annat.
Biblioteken har böcker och annat material på flera olika språk.
I biblioteket kan du också använda dator.
Ofta hålls också utställningar och evenemang på biblioteken.
linkkiEsbo stad:
Bibliotekfinska _ svenska _ engelska
Flerspråkiga biblioteket
Flerspråkiga biblioteket ligger i Böle i Helsingfors
Här finns böcker, musik, tidningar och tidskrifter samt ljudböcker på flera olika språk.
Du kan åka till Böle eller beställa material till ditt eget närbibliotek.
linkkiHelsingfors stadsbibliotek:
Flerspråkiga biblioteketfinska _ svenska _ engelska
Huvudstadsregionens gemensamma bibliotekstjänstfinska _ svenska _ engelska _ somaliska _ persiska _ arabiska
Läs mer: Bibliotek.
Motion
I Esbo finns simhallar, flera idrottshallar, idrottsplaner och andra idrottsplatser för olika idrottsgrenar.
På motionsslingorna kan man springa på somrarna och åka skidor på vintrarna.
Läs mer: Motion.
linkkiEsbo stad:
Information om motionstjänsternafinska _ svenska _ engelska
linkkiEsbo stad:
Idrottsklubbarfinska _ svenska
Att röra sig i naturen
I Esbo finns flera friluftsområden där man kan vandra i naturen.
Till exempel Noux nationalpark ligger delvis på Esbos område.
linkkiEsbo stad:
Naturobjekt i Esbofinska _ svenska _ engelska
Webbsidorfinska _ svenska _ engelska _ ryska _ kinesiska
Hemstadsstigarfinska _ svenska _ engelska
I naturhuset Villa Elfvik ordnas utflykter, evenemang och utställningar.
Naturhuset är öppet för alla och ligger vid sidan av Bredvikens naturskyddsområde.
linkkiVilla Elfvik:
Naturens husfinska _ svenska _ engelska
I Esbo finns motionsslingor och friluftsleder på olika håll i staden.
På vintern är många motionsslingor skidspår.
En del rutter är belysta.
linkkiEsbo stad:
Friluftslivfinska _ svenska _ engelska
linkkiEsbo stad:
Friluftsområdenfinska _ svenska _ engelska
Vid insjöarna och på havskusten finns många badstränder.
Alla Esbobor får fritt fiska med metspö och pimpla.
Om du använder andra fiskeredskap ska du ha ett fisketillstånd.
linkkiEsbo stad:
Fiske och jaktfinska _ svenska _ engelska
Läs mer: Att röra sig i naturen.
Teater och film
I Esbo finns flera yrkes- och amatörteatrar.
I Esbo finns tre biografer.
Mer information om filmerna hittar du på biografernas webbplatser.
Därtill ordnar Esbo stad filmvisningar.
Läs mer: Teater och film.
linkkiFinnkino:
Filmerfinska _ engelska
Filmerfinska
Filmerfinska _ svenska _ engelska
linkkiEsbo stad:
Teatrar i Esbofinska _ svenska _ engelska
Museer
I Esbo finns flera museer.
Esbo moderna konstmuseum EMMA är ett av Finlands största konstmuseer.
Läs mer: Museer.
linkkiEsbo stad:
Museerfinska _ svenska _ engelska
linkkiEsbo stad:
Stadsmuseetfinska _ svenska _ engelska
linkkiEsbo stad:
Museet för modern konst EMMAfinska _ svenska _ engelska _ ryska
Fritidsverksamhet för barn och unga
I Esbo finns flera läroanstalter som ger grundundervisning i konstämnen speciellt för barn och unga.
Olika konstarter är musik, bildkonst, dans, teater och cirkuskonst.
I Esbo finns ungdomsgårdar med utbildade ledare som övervakar verksamheten.
Ungdomsgårdarna är öppna för alla ungdomar i åldrarna 9–17.
På ungdomsgårdarna kan de unga vistas på fritiden.
Där bedrivs det även hobbyklubbar och ordnas kurser och evenemang.
Också föreningar och idrottsklubbar ordnar mycket verksamhet för ungdomar.
Läs mer: Fritidsverksamhet för barn och unga.
linkkiEsbo stad:
Verksamhet för ungafinska _ svenska _ engelska
linkkiEsbo stad:
Ungdomsgårdarfinska _ svenska _ engelska
linkkiEsbo stad:
Rådgivning för ungafinska _ svenska _ engelska
linkkiEsbo stad:
Idrottsklubbarfinska _ svenska
Hobbysökningfinska
Föreningar
I Esbo finns många olika föreningar, till exempel kulturföreningar och idrottsklubbar.
Läs mer: Föreningar.
linkkiEsbo stad:
Idrottsklubbarfinska _ svenska
Föreningsverksamhetfinska
linkkiEsbo stad:
Föreningar för seniorerfinska _ svenska
Evenemang
Bibliotek
Motion
Att röra sig i naturen
Teater och film
Museer
Fritidsverksamhet för barn och unga
Föreningar
I Esbo finns många hobbymöjligheter.
Invånarhusen Kivenkolo och Kylämaja är öppna för alla.
I invånarhusen kan områdets invånare vistas och samlas samt få anvisningar och råd.
Invånarhuset Kivenkolo
Sjöstöveln 1 A
linkkiEsbo stad:
Kivenkolo invånarhusfinska _ svenska _ engelska
Invånarhuset Kylämaja
Mattsgatan 7
linkkiEsbo stad:
Invånarhus Kylämajafinska
Vid Esbo arbetarinstitut (Espoon työväenopisto) kan man till exempel skapa konst, handarbeten, laga mat, dansa eller idka motion.
Där kan man även studera finska och andra språk.
linkkiEsbo stad:
Arbetarinstitutetfinska _ svenska _ engelska
I Esbo finns flera läroanstalter som ger grundundervisning i konstämnen speciellt för barn och unga.
Olika konstarter är musik, bildkonst, dans, teater och cirkus.
linkkiEsbo stad:
Konstundervisningfinska _ engelska.
Konsthuset Lilla Aurora ordnar kulturevenemang för barn.
linkkiEsbo stad:
Kulturevenemang för barnfinska _ svenska _ engelska
Läs mer: Fritid.
Evenemang
Evenemangfinska _ svenska _ engelska _ ryska
linkkiEsbo stad:
Evenemangfinska
Bibliotek
I Esbo finns flera bibliotek på olika håll i staden.
På biblioteket kan du låna böcker, tidningar, musik, filmer, spel och mycket annat.
Biblioteken har böcker och annat material på flera olika språk.
I biblioteket kan du också använda dator.
Ofta hålls också utställningar och evenemang på biblioteken.
linkkiEsbo stad:
Bibliotekfinska _ svenska _ engelska
Flerspråkiga biblioteket
Flerspråkiga biblioteket ligger i Böle i Helsingfors
Här finns böcker, musik, tidningar och tidskrifter samt ljudböcker på flera olika språk.
Du kan åka till Böle eller beställa material till ditt eget närbibliotek.
linkkiHelsingfors stadsbibliotek:
Flerspråkiga biblioteketfinska _ svenska _ engelska
Huvudstadsregionens gemensamma bibliotekstjänstfinska _ svenska _ engelska _ somaliska _ persiska _ arabiska
Läs mer: Bibliotek.
Motion
I Esbo finns simhallar, flera idrottshallar, idrottsplaner och andra idrottsplatser för olika idrottsgrenar.
På motionsslingorna kan man springa på somrarna och åka skidor på vintrarna.
Läs mer: Motion.
linkkiEsbo stad:
Information om motionstjänsternafinska _ svenska _ engelska
linkkiEsbo stad:
Idrottsklubbarfinska _ svenska
Att röra sig i naturen
I Esbo finns flera friluftsområden där man kan vandra i naturen.
Till exempel Noux nationalpark ligger delvis på Esbos område.
linkkiEsbo stad:
Naturobjekt i Esbofinska _ svenska _ engelska
Webbsidorfinska _ svenska _ engelska _ ryska _ kinesiska
Hemstadsstigarfinska _ svenska _ engelska
I naturhuset Villa Elfvik ordnas utflykter, evenemang och utställningar.
Naturhuset är öppet för alla och ligger vid sidan av Bredvikens naturskyddsområde.
linkkiVilla Elfvik:
Naturens husfinska _ svenska _ engelska
I Esbo finns motionsslingor och friluftsleder på olika håll i staden.
På vintern är många motionsslingor skidspår.
En del rutter är belysta.
linkkiEsbo stad:
Friluftslivfinska _ svenska _ engelska
linkkiEsbo stad:
Friluftsområdenfinska _ svenska _ engelska
Vid insjöarna och på havskusten finns många badstränder.
Alla Esbobor får fritt fiska med metspö och pimpla.
Om du använder andra fiskeredskap ska du ha ett fisketillstånd.
linkkiEsbo stad:
Fiske och jaktfinska _ svenska _ engelska
Läs mer: Att röra sig i naturen.
Teater och film
I Esbo finns flera yrkes- och amatörteatrar.
I Esbo finns tre biografer.
Mer information om filmerna hittar du på biografernas webbplatser.
Därtill ordnar Esbo stad filmvisningar.
Läs mer: Teater och film.
linkkiFinnkino:
Filmerfinska _ engelska
Filmerfinska
Filmerfinska _ svenska _ engelska
linkkiEsbo stad:
Teatrar i Esbofinska _ svenska _ engelska
Museer
I Esbo finns flera museer.
Esbo moderna konstmuseum EMMA är ett av Finlands största konstmuseer.
Läs mer: Museer.
linkkiEsbo stad:
Museerfinska _ svenska _ engelska
linkkiEsbo stad:
Stadsmuseetfinska _ svenska _ engelska
linkkiEsbo stad:
Museet för modern konst EMMAfinska _ svenska _ engelska _ ryska
Fritidsverksamhet för barn och unga
I Esbo finns flera läroanstalter som ger grundundervisning i konstämnen speciellt för barn och unga.
Olika konstarter är musik, bildkonst, dans, teater och cirkuskonst.
I Esbo finns ungdomsgårdar med utbildade ledare som övervakar verksamheten.
Ungdomsgårdarna är öppna för alla ungdomar i åldrarna 9–17.
På ungdomsgårdarna kan de unga vistas på fritiden.
Där bedrivs det även hobbyklubbar och ordnas kurser och evenemang.
Också föreningar och idrottsklubbar ordnar mycket verksamhet för ungdomar.
Läs mer: Fritidsverksamhet för barn och unga.
linkkiEsbo stad:
Verksamhet för ungafinska _ svenska _ engelska
linkkiEsbo stad:
Ungdomsgårdarfinska _ svenska _ engelska
linkkiEsbo stad:
Rådgivning för ungafinska _ svenska _ engelska
linkkiEsbo stad:
Idrottsklubbarfinska _ svenska
Hobbysökningfinska
Föreningar
I Esbo finns många olika föreningar, till exempel kulturföreningar och idrottsklubbar.
Läs mer: Föreningar.
linkkiEsbo stad:
Idrottsklubbarfinska _ svenska
Föreningsverksamhetfinska
linkkiEsbo stad:
Föreningar för seniorerfinska _ svenska
Evenemang
Bibliotek
Motion
Att röra sig i naturen
Teater och film
Museer
Fritidsverksamhet för barn och unga
Föreningar
I Esbo finns många hobbymöjligheter.
Invånarhusen Kivenkolo och Kylämaja är öppna för alla.
I invånarhusen kan områdets invånare vistas och samlas samt få anvisningar och råd.
Invånarhuset Kivenkolo
Sjöstöveln 1 A
linkkiEsbo stad:
Kivenkolo invånarhusfinska _ svenska _ engelska
Invånarhuset Kylämaja
Mattsgatan 7
linkkiEsbo stad:
Invånarhus Kylämajafinska
Vid Esbo arbetarinstitut (Espoon työväenopisto) kan man till exempel skapa konst, handarbeten, laga mat, dansa eller idka motion.
Där kan man även studera finska och andra språk.
linkkiEsbo stad:
Arbetarinstitutetfinska _ svenska _ engelska
I Esbo finns flera läroanstalter som ger grundundervisning i konstämnen speciellt för barn och unga.
Olika konstarter är musik, bildkonst, dans, teater och cirkus.
linkkiEsbo stad:
Konstundervisningfinska _ engelska.
Konsthuset Lilla Aurora ordnar kulturevenemang för barn.
linkkiEsbo stad:
Kulturevenemang för barnfinska _ svenska _ engelska
Läs mer: Fritid.
Evenemang
Evenemangfinska _ svenska _ engelska _ ryska
linkkiEsbo stad:
Evenemangfinska
Bibliotek
I Esbo finns flera bibliotek på olika håll i staden.
På biblioteket kan du låna böcker, tidningar, musik, filmer, spel och mycket annat.
Biblioteken har böcker och annat material på flera olika språk.
I biblioteket kan du också använda dator.
Ofta hålls också utställningar och evenemang på biblioteken.
linkkiEsbo stad:
Bibliotekfinska _ svenska _ engelska
Flerspråkiga biblioteket
Flerspråkiga biblioteket ligger i Böle i Helsingfors
Här finns böcker, musik, tidningar och tidskrifter samt ljudböcker på flera olika språk.
Du kan åka till Böle eller beställa material till ditt eget närbibliotek.
linkkiHelsingfors stadsbibliotek:
Flerspråkiga biblioteketfinska _ svenska _ engelska
Huvudstadsregionens gemensamma bibliotekstjänstfinska _ svenska _ engelska _ somaliska _ persiska _ arabiska
Läs mer: Bibliotek.
Motion
I Esbo finns simhallar, flera idrottshallar, idrottsplaner och andra idrottsplatser för olika idrottsgrenar.
På motionsslingorna kan man springa på somrarna och åka skidor på vintrarna.
Läs mer: Motion.
linkkiEsbo stad:
Information om motionstjänsternafinska _ svenska _ engelska
linkkiEsbo stad:
Idrottsklubbarfinska _ svenska
Att röra sig i naturen
I Esbo finns flera friluftsområden där man kan vandra i naturen.
Till exempel Noux nationalpark ligger delvis på Esbos område.
linkkiEsbo stad:
Naturobjekt i Esbofinska _ svenska _ engelska
Webbsidorfinska _ svenska _ engelska _ ryska _ kinesiska
Hemstadsstigarfinska _ svenska _ engelska
I naturhuset Villa Elfvik ordnas utflykter, evenemang och utställningar.
Naturhuset är öppet för alla och ligger vid sidan av Bredvikens naturskyddsområde.
linkkiVilla Elfvik:
Naturens husfinska _ svenska _ engelska
I Esbo finns motionsslingor och friluftsleder på olika håll i staden.
På vintern är många motionsslingor skidspår.
En del rutter är belysta.
linkkiEsbo stad:
Friluftslivfinska _ svenska _ engelska
linkkiEsbo stad:
Friluftsområdenfinska _ svenska _ engelska
Vid insjöarna och på havskusten finns många badstränder.
Alla Esbobor får fritt fiska med metspö och pimpla.
Om du använder andra fiskeredskap ska du ha ett fisketillstånd.
linkkiEsbo stad:
Fiske och jaktfinska _ svenska _ engelska
Läs mer: Att röra sig i naturen.
Teater och film
I Esbo finns flera yrkes- och amatörteatrar.
I Esbo finns tre biografer.
Mer information om filmerna hittar du på biografernas webbplatser.
Därtill ordnar Esbo stad filmvisningar.
Läs mer: Teater och film.
linkkiFinnkino:
Filmerfinska _ engelska
Filmerfinska
Filmerfinska _ svenska _ engelska
linkkiEsbo stad:
Teatrar i Esbofinska _ svenska _ engelska
Museer
I Esbo finns flera museer.
Esbo moderna konstmuseum EMMA är ett av Finlands största konstmuseer.
Läs mer: Museer.
linkkiEsbo stad:
Museerfinska _ svenska _ engelska
linkkiEsbo stad:
Stadsmuseetfinska _ svenska _ engelska
linkkiEsbo stad:
Museet för modern konst EMMAfinska _ svenska _ engelska _ ryska
Fritidsverksamhet för barn och unga
I Esbo finns flera läroanstalter som ger grundundervisning i konstämnen speciellt för barn och unga.
Olika konstarter är musik, bildkonst, dans, teater och cirkuskonst.
I Esbo finns ungdomsgårdar med utbildade ledare som övervakar verksamheten.
Ungdomsgårdarna är öppna för alla ungdomar i åldrarna 9–17.
På ungdomsgårdarna kan de unga vistas på fritiden.
Där bedrivs det även hobbyklubbar och ordnas kurser och evenemang.
Också föreningar och idrottsklubbar ordnar mycket verksamhet för ungdomar.
Läs mer: Fritidsverksamhet för barn och unga.
linkkiEsbo stad:
Verksamhet för ungafinska _ svenska _ engelska
linkkiEsbo stad:
Ungdomsgårdarfinska _ svenska _ engelska
linkkiEsbo stad:
Rådgivning för ungafinska _ svenska _ engelska
linkkiEsbo stad:
Idrottsklubbarfinska _ svenska
Hobbysökningfinska
Föreningar
I Esbo finns många olika föreningar, till exempel kulturföreningar och idrottsklubbar.
Läs mer: Föreningar.
linkkiEsbo stad:
Idrottsklubbarfinska _ svenska
Föreningsverksamhetfinska
linkkiEsbo stad:
Föreningar för seniorerfinska _ svenska
Problem med uppehållstillståndet
Brott
Behöver du en jurist?
Våld Problem i äktenskap eller parförhållande
Barns och ungas problem
Missbruksproblem
Dödsfall
Ring nödnumret 112 om det är fråga om en nödsituation.
Via nödnumret kan du tillkalla polis, ambulans eller brandkår.
Ring inte nödnumret om det inte är en nödsituation.
Läs mer:Nödsituationer
linkkiEsbo stad:
Jourmottagningarfinska _ svenska _ engelska
Social- och krisjouren
Social- och krisjouren (sosiaali- ja kriisipäivystys) hjälper dygnet runt om du eller din familj behöver hjälp i en akut krissituation.
Krisen kan till exempel ha med våld, parförhållandet eller barnens problem att göra.
Du kan även kontakta social- och krisjouren om du har problem med din mentala hälsa, missbruksproblem eller om du råkat ut för en traumatisk händelse i livet.
Social- och krisjouren
Jorvs sjukhus
Åbovägen 150
Tfn (09) 816 42439
Öppet varje dag dygnet runt.
linkkiEsbo stad:
Social- och krisjourenfinska _ svenska _ engelska
Föreningen för mental hälsa i Finland (Suomen Mielenterveysseura) har en krismottagning för invandrare.
Kontoret ligger i Böle i Helsingfors.
Krismottagningen ger dig hjälp och stöd i svåra situationer.
Boka en tid per telefon på numret (09) 4135 0501.
linkkiFöreningen för mental hälsa i Finland:
Krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Problem med uppehållstillståndet
Om du har problem eller oklarheter med uppehållstillståndet, ska du ta kontakt med migrationsverket.
Läs mer: Problem med uppehållstillstånd
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Om du är flykting, asylsökande eller vistas i Finland av någon annan anledning kan du be om juridisk hjälp och rådgivning vid Flyktingrådgivningen rf.
Kontoret ligger i Helsingfors.
Adress: Kaisaniemigatan 4 A
Tfn 09 2313 9325
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Brott
Om du blir utsatt för ett brott, gör en brottsanmälan hos polisen.
Du kan göra brottsanmälan på internet.
Du kan även fylla i en blankett och lämna den till Esbo huvudpolisstation.
Esbo huvudpolisstation
Knektbrogränden 4
Läs mer: Brott
Kontaktuppgifterfinska _ svenska _ engelska
Elektronisk polisanmälanfinska _ svenska _ engelska
Behöver du en jurist?
Om du behöver juridisk hjälp, kan du kontakta Västra Nylands rättshjälpsbyrå.
Biskopsbron 9 B
Tfn 029 56 61820
Läs mer: Behöver du en jurist?
linkkiVästra Nylands rättshjälpsbyrå:
Rättshjälpfinska
Våld
Omatila (Omatila) hjälper dig om du har blivit utsatt för närståendevåld eller våld inom familjen.
Omatila ordnar vid behov boende för dig och dina barn.
Du kan ringa Omatila-tjänsten dygnet runt. Du behöver inte uppge ditt namn när du ringer.
Du kan också komma utan tidsbokning för att prata om din situation, måndag till fredag kl. 9–11 och onsdagar kl. 16–20.
Omatila
Enheten för familjeärenden
Kamrersvägen 6 A
Tfn 043 825 0535
Läs mer: Våld
linkkiEsbo stad:
Hjälp till offer för familjevåldfinska _ svenska _ engelska
Miehen Linja (Miehen Linja) är en tjänst som hjälper män, som har utsatt sina familjemedlemmar för våld. Tjänsten är avsedd för invandrarmän.
Målargränden 3 B
Tfn (09) 276 62899
Hjälp för invandrarmänfinska _ engelska
Problem i äktenskap eller parförhållande
Om du har problem i ditt äktenskap eller parförhållande kan du kontakta familjerådgivningen.
Familjerådgivningsbyråerna är i synnerhet avsedda för familjer med barn.
linkkiEsbo stad:
Familjerådgivningarfinska _ svenska _ engelska
Väestöliitto erbjuder rådgivning och terapi för par på finska och engelska.
linkkiBefolkningsförbundet:
Rådgivning till invandrare telefonledes och via e-postfinska _ svenska _ engelska
Familia Clubs projekt Duo erbjuder relationsrådgivning för par från två kulturer på finska och engelska.
Rådgivningen är avgiftsbelagd.
Relationsrådgivning för par från två kulturerfinska _ engelska
Också kyrkans familjerådgivningscentral erbjuder familjerådgivning vid problem i parförhållandet.
Kyrkans familjerådgivningfinska _ svenska _ engelska
Läs mer: Problem i äktenskap och parförhållande
Barns och ungas problem
Hälsovårdaren vid barnrådgivningen ger råd i frågor som rör hälsan och utvecklingen av barn under skolåldern.
I Esbo finns flera rådgivningsbyråer runtom i staden.
Rådgivningsbyråernas tidsbokning och rådgivning
Tfn (09) 816 22800
linkkiEsbo stad:
Rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
Vid problem som berör barn i skolåldern hjälper till exempel skolans hälsovårdare.
linkkiEsbo stad:
Information om hälsovården för skolbarnfinska _ svenska _ engelska
Om du behöver råd i frågor kring barns psykiska utveckling, kan du boka en tid hos familjerådgivningen.
linkkiEsbo stad:
Familjerådgivningarfinska _ svenska _ engelska
Väestöliitto ger råd till invandrarfamiljer i frågor rörande barnfostran och familjens välmående.
Rådgivningen på olika språk:
Tfn 050 325 7173 (ryska, engelska)
Unga kan prata om sina problem med hälsovårdaren på den egna skolan eller läroanstalten.
Det finns även andra ställen där man kan få hjälp.
En ung i åldern 13–22 år kan få hjälp vid Ungdomspolikliniken Nupoli om hen har problem till exempel med den mentala hälsan, rusmedelsbruk, spelande eller fritidsaktiviteterna.
Man kan ringa eller besöka Nupoli.
Besök på Nupoli är kostnadsfria och konfidentiella.
Tfn 09 816 31300
linkkiEsbo stad:
Nupoli - hjälp för ungafinska _ svenska
Om den unga inte är trygg i sitt eget hem, kan hen kontakta Finlands Röda Kors De ungas skyddshus.
Skyddshuset finns i Alberga.
De ungas skyddshus
Tfn (09) 8195 5360
linkkiFinlands Röda Kors:
De ungas skyddshusfinska
Läs mer: Barns och ungas problem
Om du har ekonomiska problem kan du fråga om råd hos kommunens socialarbetare.
Om du eller din familj inte har tillräckliga inkomster eller tillgångar för den nödvändiga dagliga försörjningen kan du söka grundläggande utkomststöd hos FPA.
Information om utkomststödfinska _ svenska _ engelska _ ryska _ estniska
Om du har problem med skulder, kontakta rättshjälpsbyråns ekonomi- och skuldrådgivning.
Tjänsten är kostnadsfri.
linkkiRättshjälpsbyrå:
Ekonomi- och skuldrådgivningfinska _ svenska _ engelska
Missbruksproblem
Kliniken för mental- och missbruksvård erbjuder vuxna Esbobor hjälp och vård vid problem med den mentala hälsan och missbruk.
Köpcentret Iso Omena
Telefon: 09 816 31300
linkkiEsbo stad:
Information om mentalvårdstjänsternafinska _ svenska _ engelska
Unga i åldern 13-22 med missbruksproblem kan få hjälp vid Ungdomspolikliniken Nupoli.
Tfn 09 816 31300
linkkiEsbo stad:
Nupoli - hjälp för ungafinska _ svenska
Läs mer: Missbruksproblem
Dödsfall
Begravningsbyråer hjälper med de praktiska arrangemangen vid en begravning.
Du kan söka begravningsbyråer till exempel på Finlands begravningsbyråers förbunds webbplats.
linkkiFinlands Begravningbyråers Förbund:
Begravningsbyråerfinska _ svenska _ engelska
I Esbo finns fem kristna begravningsplatser.
På Klockarmalmens begravningsplats finns ett gravområde för konfessionslösa.
Där kan de avlidna begravas som hade en annan religionstillhörighet eller inte hörde till något religionssamfund.
linkkiEsbo församlingar:
Begravningsplatserfinska _ svenska _ engelska
Om en närstående dör oväntat och du behöver stöd kan du kontakta social- och krisjouren i Esbo, telefon (09) 816 42439.
Läs mer: Dödsfall
Problem med uppehållstillståndet
Brott
Behöver du en jurist?
Våld Problem i äktenskap eller parförhållande
Barns och ungas problem
Missbruksproblem
Dödsfall
Ring nödnumret 112 om det är fråga om en nödsituation.
Via nödnumret kan du tillkalla polis, ambulans eller brandkår.
Ring inte nödnumret om det inte är en nödsituation.
Läs mer:Nödsituationer
linkkiEsbo stad:
Jourmottagningarfinska _ svenska _ engelska
Social- och krisjouren
Social- och krisjouren (sosiaali- ja kriisipäivystys) hjälper dygnet runt om du eller din familj behöver hjälp i en akut krissituation.
Krisen kan till exempel ha med våld, parförhållandet eller barnens problem att göra.
Du kan även kontakta social- och krisjouren om du har problem med din mentala hälsa, missbruksproblem eller om du råkat ut för en traumatisk händelse i livet.
Social- och krisjouren
Jorvs sjukhus
Åbovägen 150
Tfn (09) 816 42439
Öppet varje dag dygnet runt.
linkkiEsbo stad:
Social- och krisjourenfinska _ svenska _ engelska
Föreningen för mental hälsa i Finland (Suomen Mielenterveysseura) har en krismottagning för invandrare.
Kontoret ligger i Böle i Helsingfors.
Krismottagningen ger dig hjälp och stöd i svåra situationer.
Boka en tid per telefon på numret (09) 4135 0501.
linkkiFöreningen för mental hälsa i Finland:
Krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Problem med uppehållstillståndet
Om du har problem eller oklarheter med uppehållstillståndet, ska du ta kontakt med migrationsverket.
Läs mer: Problem med uppehållstillstånd
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Om du är flykting, asylsökande eller vistas i Finland av någon annan anledning kan du be om juridisk hjälp och rådgivning vid Flyktingrådgivningen rf.
Kontoret ligger i Helsingfors.
Adress: Kaisaniemigatan 4 A
Tfn 09 2313 9325
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Brott
Om du blir utsatt för ett brott, gör en brottsanmälan hos polisen.
Du kan göra brottsanmälan på internet.
Du kan även fylla i en blankett och lämna den till Esbo huvudpolisstation.
Esbo huvudpolisstation
Knektbrogränden 4
Läs mer: Brott
Kontaktuppgifterfinska _ svenska _ engelska
Elektronisk polisanmälanfinska _ svenska _ engelska
Behöver du en jurist?
Om du behöver juridisk hjälp, kan du kontakta Västra Nylands rättshjälpsbyrå.
Biskopsbron 9 B
Tfn 029 56 61820
Läs mer: Behöver du en jurist?
linkkiVästra Nylands rättshjälpsbyrå:
Rättshjälpfinska
Våld
Omatila (Omatila) hjälper dig om du har blivit utsatt för närståendevåld eller våld inom familjen.
Omatila ordnar vid behov boende för dig och dina barn.
Du kan ringa Omatila-tjänsten dygnet runt. Du behöver inte uppge ditt namn när du ringer.
Du kan också komma utan tidsbokning för att prata om din situation, måndag till fredag kl. 9–11 och onsdagar kl. 16–20.
Omatila
Enheten för familjeärenden
Kamrersvägen 6 A
Tfn 043 825 0535
Läs mer: Våld
linkkiEsbo stad:
Hjälp till offer för familjevåldfinska _ svenska _ engelska
Miehen Linja (Miehen Linja) är en tjänst som hjälper män, som har utsatt sina familjemedlemmar för våld. Tjänsten är avsedd för invandrarmän.
Målargränden 3 B
Tfn (09) 276 62899
Hjälp för invandrarmänfinska _ engelska
Problem i äktenskap eller parförhållande
Om du har problem i ditt äktenskap eller parförhållande kan du kontakta familjerådgivningen.
Familjerådgivningsbyråerna är i synnerhet avsedda för familjer med barn.
linkkiEsbo stad:
Familjerådgivningarfinska _ svenska _ engelska
Väestöliitto erbjuder rådgivning och terapi för par på finska och engelska.
linkkiBefolkningsförbundet:
Rådgivning till invandrare telefonledes och via e-postfinska _ svenska _ engelska
Familia Clubs projekt Duo erbjuder relationsrådgivning för par från två kulturer på finska och engelska.
Rådgivningen är avgiftsbelagd.
Relationsrådgivning för par från två kulturerfinska _ engelska
Också kyrkans familjerådgivningscentral erbjuder familjerådgivning vid problem i parförhållandet.
Kyrkans familjerådgivningfinska _ svenska _ engelska
Läs mer: Problem i äktenskap och parförhållande
Barns och ungas problem
Hälsovårdaren vid barnrådgivningen ger råd i frågor som rör hälsan och utvecklingen av barn under skolåldern.
I Esbo finns flera rådgivningsbyråer runtom i staden.
Rådgivningsbyråernas tidsbokning och rådgivning
Tfn (09) 816 22800
linkkiEsbo stad:
Rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
Vid problem som berör barn i skolåldern hjälper till exempel skolans hälsovårdare.
linkkiEsbo stad:
Information om hälsovården för skolbarnfinska _ svenska _ engelska
Om du behöver råd i frågor kring barns psykiska utveckling, kan du boka en tid hos familjerådgivningen.
linkkiEsbo stad:
Familjerådgivningarfinska _ svenska _ engelska
Väestöliitto ger råd till invandrarfamiljer i frågor rörande barnfostran och familjens välmående.
Rådgivningen på olika språk:
Tfn 050 325 7173 (ryska, engelska)
Unga kan prata om sina problem med hälsovårdaren på den egna skolan eller läroanstalten.
Det finns även andra ställen där man kan få hjälp.
En ung i åldern 13–22 år kan få hjälp vid Ungdomspolikliniken Nupoli om hen har problem till exempel med den mentala hälsan, rusmedelsbruk, spelande eller fritidsaktiviteterna.
Man kan ringa eller besöka Nupoli.
Besök på Nupoli är kostnadsfria och konfidentiella.
Tfn 09 816 31300
linkkiEsbo stad:
Nupoli - hjälp för ungafinska _ svenska
Om den unga inte är trygg i sitt eget hem, kan hen kontakta Finlands Röda Kors De ungas skyddshus.
Skyddshuset finns i Alberga.
De ungas skyddshus
Tfn (09) 8195 5360
linkkiFinlands Röda Kors:
De ungas skyddshusfinska
Läs mer: Barns och ungas problem
Om du har ekonomiska problem kan du fråga om råd hos kommunens socialarbetare.
Om du eller din familj inte har tillräckliga inkomster eller tillgångar för den nödvändiga dagliga försörjningen kan du söka grundläggande utkomststöd hos FPA.
Information om utkomststödfinska _ svenska _ engelska _ ryska _ estniska
Om du har problem med skulder, kontakta rättshjälpsbyråns ekonomi- och skuldrådgivning.
Tjänsten är kostnadsfri.
linkkiRättshjälpsbyrå:
Ekonomi- och skuldrådgivningfinska _ svenska _ engelska
Missbruksproblem
Kliniken för mental- och missbruksvård erbjuder vuxna Esbobor hjälp och vård vid problem med den mentala hälsan och missbruk.
Köpcentret Iso Omena
Telefon: 09 816 31300
linkkiEsbo stad:
Information om mentalvårdstjänsternafinska _ svenska _ engelska
Unga i åldern 13-22 med missbruksproblem kan få hjälp vid Ungdomspolikliniken Nupoli.
Tfn 09 816 31300
linkkiEsbo stad:
Nupoli - hjälp för ungafinska _ svenska
Läs mer: Missbruksproblem
Dödsfall
Begravningsbyråer hjälper med de praktiska arrangemangen vid en begravning.
Du kan söka begravningsbyråer till exempel på Finlands begravningsbyråers förbunds webbplats.
linkkiFinlands Begravningbyråers Förbund:
Begravningsbyråerfinska
I Esbo finns fem kristna begravningsplatser.
På Klockarmalmens begravningsplats finns ett gravområde för konfessionslösa.
Där kan de avlidna begravas som hade en annan religionstillhörighet eller inte hörde till något religionssamfund.
linkkiEsbo församlingar:
Begravningsplatserfinska _ svenska _ engelska
Om en närstående dör oväntat och du behöver stöd kan du kontakta social- och krisjouren i Esbo, telefon (09) 816 42439.
Läs mer: Dödsfall
Problem med uppehållstillståndet
Brott
Behöver du en jurist?
Våld Problem i äktenskap eller parförhållande
Barns och ungas problem
Missbruksproblem
Dödsfall
Ring nödnumret 112 om det är fråga om en nödsituation.
Via nödnumret kan du tillkalla polis, ambulans eller brandkår.
Ring inte nödnumret om det inte är en nödsituation.
Läs mer:Nödsituationer
linkkiEsbo stad:
Jourmottagningarfinska _ svenska _ engelska
Social- och krisjouren
Social- och krisjouren (sosiaali- ja kriisipäivystys) hjälper dygnet runt om du eller din familj behöver hjälp i en akut krissituation.
Krisen kan till exempel ha med våld, parförhållandet eller barnens problem att göra.
Du kan även kontakta social- och krisjouren om du har problem med din mentala hälsa, missbruksproblem eller om du råkat ut för en traumatisk händelse i livet.
Social- och krisjouren
Jorvs sjukhus
Åbovägen 150
Tfn (09) 816 42439
Öppet varje dag dygnet runt.
linkkiEsbo stad:
Social- och krisjourenfinska _ svenska _ engelska
Föreningen för mental hälsa i Finland (Suomen Mielenterveysseura) har en krismottagning för invandrare.
Kontoret ligger i Böle i Helsingfors.
Krismottagningen ger dig hjälp och stöd i svåra situationer.
Boka en tid per telefon på numret (09) 4135 0501.
linkkiFöreningen för mental hälsa i Finland:
Krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Problem med uppehållstillståndet
Om du har problem eller oklarheter med uppehållstillståndet, ska du ta kontakt med migrationsverket.
Läs mer: Problem med uppehållstillstånd
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Om du är flykting, asylsökande eller vistas i Finland av någon annan anledning kan du be om juridisk hjälp och rådgivning vid Flyktingrådgivningen rf.
Kontoret ligger i Helsingfors.
Adress: Kaisaniemigatan 4 A
Tfn 09 2313 9325
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Brott
Om du blir utsatt för ett brott, gör en brottsanmälan hos polisen.
Du kan göra brottsanmälan på internet.
Du kan även fylla i en blankett och lämna den till Esbo huvudpolisstation.
Esbo huvudpolisstation
Knektbrogränden 4
Läs mer: Brott
Kontaktuppgifterfinska _ svenska _ engelska
Elektronisk polisanmälanfinska _ svenska _ engelska
Behöver du en jurist?
Om du behöver juridisk hjälp, kan du kontakta Västra Nylands rättshjälpsbyrå.
Biskopsbron 9 B
Tfn 029 56 61820
Läs mer: Behöver du en jurist?
linkkiVästra Nylands rättshjälpsbyrå:
Rättshjälpfinska
Våld
Omatila (Omatila) hjälper dig om du har blivit utsatt för närståendevåld eller våld inom familjen.
Omatila ordnar vid behov boende för dig och dina barn.
Du kan ringa Omatila-tjänsten dygnet runt. Du behöver inte uppge ditt namn när du ringer.
Du kan också komma utan tidsbokning för att prata om din situation, måndag till fredag kl. 9–11 och onsdagar kl. 16–20.
Omatila
Enheten för familjeärenden
Kamrersvägen 6 A
Tfn 043 825 0535
Läs mer: Våld
linkkiEsbo stad:
Hjälp till offer för familjevåldfinska _ svenska _ engelska
Miehen Linja (Miehen Linja) är en tjänst som hjälper män, som har utsatt sina familjemedlemmar för våld. Tjänsten är avsedd för invandrarmän.
Målargränden 3 B
Tfn (09) 276 62899
Hjälp för invandrarmänfinska _ engelska
Problem i äktenskap eller parförhållande
Om du har problem i ditt äktenskap eller parförhållande kan du kontakta familjerådgivningen.
Familjerådgivningsbyråerna är i synnerhet avsedda för familjer med barn.
linkkiEsbo stad:
Familjerådgivningarfinska _ svenska _ engelska
Väestöliitto erbjuder rådgivning och terapi för par på finska och engelska.
linkkiBefolkningsförbundet:
Rådgivning till invandrare telefonledes och via e-postfinska _ svenska _ engelska
Familia Clubs projekt Duo erbjuder relationsrådgivning för par från två kulturer på finska och engelska.
Rådgivningen är avgiftsbelagd.
Relationsrådgivning för par från två kulturerfinska _ engelska
Också kyrkans familjerådgivningscentral erbjuder familjerådgivning vid problem i parförhållandet.
Kyrkans familjerådgivningfinska _ svenska _ engelska
Läs mer: Problem i äktenskap och parförhållande
Barns och ungas problem
Hälsovårdaren vid barnrådgivningen ger råd i frågor som rör hälsan och utvecklingen av barn under skolåldern.
I Esbo finns flera rådgivningsbyråer runtom i staden.
Rådgivningsbyråernas tidsbokning och rådgivning
Tfn (09) 816 22800
linkkiEsbo stad:
Rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
Vid problem som berör barn i skolåldern hjälper till exempel skolans hälsovårdare.
linkkiEsbo stad:
Information om hälsovården för skolbarnfinska _ svenska _ engelska
Om du behöver råd i frågor kring barns psykiska utveckling, kan du boka en tid hos familjerådgivningen.
linkkiEsbo stad:
Familjerådgivningarfinska _ svenska _ engelska
Väestöliitto ger råd till invandrarfamiljer i frågor rörande barnfostran och familjens välmående.
Rådgivningen på olika språk:
Tfn 050 325 7173 (ryska, engelska)
Unga kan prata om sina problem med hälsovårdaren på den egna skolan eller läroanstalten.
Det finns även andra ställen där man kan få hjälp.
En ung i åldern 13–22 år kan få hjälp vid Ungdomspolikliniken Nupoli om hen har problem till exempel med den mentala hälsan, rusmedelsbruk, spelande eller fritidsaktiviteterna.
Man kan ringa eller besöka Nupoli.
Besök på Nupoli är kostnadsfria och konfidentiella.
Tfn 09 816 31300
linkkiEsbo stad:
Nupoli - hjälp för ungafinska _ svenska
Om den unga inte är trygg i sitt eget hem, kan hen kontakta Finlands Röda Kors De ungas skyddshus.
Skyddshuset finns i Alberga.
De ungas skyddshus
Tfn (09) 8195 5360
linkkiFinlands Röda Kors:
De ungas skyddshusfinska
Läs mer: Barns och ungas problem
Om du har ekonomiska problem kan du fråga om råd hos kommunens socialarbetare.
Om du eller din familj inte har tillräckliga inkomster eller tillgångar för den nödvändiga dagliga försörjningen kan du söka grundläggande utkomststöd hos FPA.
Information om utkomststödfinska _ svenska _ engelska _ ryska _ estniska
Om du har problem med skulder, kontakta rättshjälpsbyråns ekonomi- och skuldrådgivning.
Tjänsten är kostnadsfri.
linkkiRättshjälpsbyrå:
Ekonomi- och skuldrådgivningfinska _ svenska _ engelska
Missbruksproblem
Kliniken för mental- och missbruksvård erbjuder vuxna Esbobor hjälp och vård vid problem med den mentala hälsan och missbruk.
Köpcentret Iso Omena
Telefon: 09 816 31300
linkkiEsbo stad:
Information om mentalvårdstjänsternafinska _ svenska _ engelska
Unga i åldern 13-22 med missbruksproblem kan få hjälp vid Ungdomspolikliniken Nupoli.
Tfn 09 816 31300
linkkiEsbo stad:
Nupoli - hjälp för ungafinska _ svenska
Läs mer: Missbruksproblem
Dödsfall
Begravningsbyråer hjälper med de praktiska arrangemangen vid en begravning.
Du kan söka begravningsbyråer till exempel på Finlands begravningsbyråers förbunds webbplats.
linkkiFinlands Begravningbyråers Förbund:
Begravningsbyråerfinska
I Esbo finns fem kristna begravningsplatser.
På Klockarmalmens begravningsplats finns ett gravområde för konfessionslösa.
Där kan de avlidna begravas som hade en annan religionstillhörighet eller inte hörde till något religionssamfund.
linkkiEsbo församlingar:
Begravningsplatserfinska _ svenska _ engelska
Om en närstående dör oväntat och du behöver stöd kan du kontakta social- och krisjouren i Esbo, telefon (09) 816 42439.
Läs mer: Dödsfall
Äktenskap
Skilsmässa
Registrerat parförhållande
Vård av barn Invånarparker och klubbar
Problem i familjen
Äktenskap
Före äktenskapet ska du skriftligt begära hindersprövning (avioliiton esteiden tutkiminen).
Hindersprövningen görs på magistraten (maistraatti).
Du kan begära hindersprövning på vilken magistrat som helst.
Magistraten i Nyland, Esbo enhet
Miestentie 3
Tfn 029 553 9391
Läs mer: Äktenskap.
Vigselfinska _ svenska _ engelska
Anhållan om prövning av hinder mot äktenskapfinska _ svenska
Skilsmässa
Kvinnan eller mannen kan lämna in skilsmässoansökan i Västra Nylands tingsrätts kansli.
Du kan också söka skilsmässa ensam, utan din makes eller makas samtycke.
Du kan skicka in ansökan till tingsrättens kansli per post, fax eller via e-post.
Tfn 029 564 4000
Läs mer: Skilsmässa.
linkkiVästra Nylands tingsrätt:
Kontaktuppgifterfinska _ svenska
Barn vid skilsmässa
Om du har barn under 13 år och överväger att skilja dig, ta kontakt med familjerådgivningen (perheneuvola).
På familjerådgivningen kan du diskutera familjens situation med de anställda.
Familjerådgivningarnas kontaktuppgifter finns på Esbo stads webbplats.
Om du planerar skilsmässa kan du också ta kontakt med barnatillsyningsmannen (lastenvalvoja) vid enheten för familjeärenden.
Med barnatillsyningsmannen kan du diskutera skilsmässan och barnens framtid.
Makarna ska ingå ett avtal om barnens boende, umgängesrätt och underhållsbidrag.
Barnatillsyningsmännen bekräftar avtalet.
Kontaktuppgifterna till barnatillsyningsmännen finns på Esbo stads webbplats.
Esbo stad har en rådgivningstelefon där man kan fråga om råd i frågor rörande barnen när föräldrarna skiljer sig.
Tfn 046 877 3267
Läs mer: Barn vid skilsmässa.
linkkiEsbo stad:
Kontaktuppgifter till barnatillsyningsmännenfinska _ svenska
linkkiEsbo stad:
Skilsmässa i en barnfamiljfinska _ svenska
Vård av barn
Information om dagvård av barn i Esbo finns på InfoFinlands sida Utbildning i Esbo.
Tillfällig vård av barn
Du kan föra barnet till en parktant för tillfällig vård.
Det innebär kortvarig (2–3 tim. per gång) vård av småbarn ute i en lekpark.
Du får närmare uppgifter av parktanterna per telefon.
Du hittar telefonnumren på Esbo stads webbplats.
linkkiEsbo stad:
Parktanterfinska
Om du behöver en tillfällig barnskötare hem, kan du kontakta Mannerheims Barnskyddsförbund eller Väestöliitto.
Barnavård och hemhjälpfinska
linkkiMannerheims Barnskyddsförbund:
Barnavårdfinska _ svenska _ engelska
Läs mer: Dagvård.
Hemvårdsstöd
Om familjens yngsta barn är under tre år, kan barnets förälder få hemvårdsstöd (kotihoidon tuki) när han eller hon vårdar barnet i hemmet.
Om du har rätt till hemvårdsstödet kan du ansöka om det hos FPA.
Du kan fylla i ansökan på Internet eller posta den till FPA.
Du kan också besöka FPA:s kontor.
Esbo stad betalar ett kommuntillägg till de familjer som vårdar ett under treårigt barn i hemmet.
Man kan ansöka om Esbotillägget om en förälder tar hand om familjens alla barn under skolåldern i hemmet.
linkkiEsbo stad:
Vård av barn i hemmetfinska _ svenska _ engelska
Information om hemvårdsstödfinska _ svenska _ engelska
Sköta ärenden på Internetfinska _ svenska _ engelska
Kontaktuppgifter till FPAfinska _ svenska _ engelska
Invånarparker och klubbar
Esbo stad ordnar mycket verksamhet för de föräldrar som vårdar barn i hemmet. Det finns till exempel invånarparker, öppna daghem och klubbar.
Läs mer: Stöd för vård av barn i hemmet
linkkiEsbo stad:
Invånarparker och klubbarfinska _ engelska
Problem i familjen
På InfoFinlands sida Problematiska situationer i Esbo hittar du uppgifter om vart du kan vända dig i Esbo för att få hjälp vid barns och ungas problem och problem i familjen.
Du hittar uppgifter om barns och ungas problem också på InfoFinlands sida Barns och ungas problem och Var hittar jag hjälp när barn eller unga har problem?
På InfoFinlands sida Problem i äktenskap och parförhållande finns uppgifter om vart du kan vända dig för att få hjälp vid problem i parförhållandet.
Äktenskap
Skilsmässa
Registrerat parförhållande
Vård av barn Invånarparker och klubbar
Problem i familjen
Äktenskap
Före äktenskapet ska du skriftligt begära hindersprövning (avioliiton esteiden tutkiminen).
Hindersprövningen görs på magistraten (maistraatti).
Du kan begära hindersprövning på vilken magistrat som helst.
Magistraten i Nyland, Esbo enhet
Miestentie 3
Tfn 029 553 9391
Läs mer: Äktenskap.
Vigselfinska _ svenska _ engelska
Anhållan om prövning av hinder mot äktenskapfinska _ svenska
Skilsmässa
Kvinnan eller mannen kan lämna in skilsmässoansökan i Västra Nylands tingsrätts kansli.
Du kan också söka skilsmässa ensam, utan din makes eller makas samtycke.
Du kan skicka in ansökan till tingsrättens kansli per post, fax eller via e-post.
Tfn 029 564 4000
Läs mer: Skilsmässa.
linkkiVästra Nylands tingsrätt:
Kontaktuppgifterfinska _ svenska
Barn vid skilsmässa
Om du har barn under 13 år och överväger att skilja dig, ta kontakt med familjerådgivningen (perheneuvola).
På familjerådgivningen kan du diskutera familjens situation med de anställda.
Familjerådgivningarnas kontaktuppgifter finns på Esbo stads webbplats.
Om du planerar skilsmässa kan du också ta kontakt med barnatillsyningsmannen (lastenvalvoja) vid enheten för familjeärenden.
Med barnatillsyningsmannen kan du diskutera skilsmässan och barnens framtid.
Makarna ska ingå ett avtal om barnens boende, umgängesrätt och underhållsbidrag.
Barnatillsyningsmännen bekräftar avtalet.
Kontaktuppgifterna till barnatillsyningsmännen finns på Esbo stads webbplats.
Esbo stad har en rådgivningstelefon där man kan fråga om råd i frågor rörande barnen när föräldrarna skiljer sig.
Tfn 046 877 3267
Läs mer: Barn vid skilsmässa.
linkkiEsbo stad:
Kontaktuppgifter till barnatillsyningsmännenfinska _ svenska
linkkiEsbo stad:
Skilsmässa i en barnfamiljfinska _ svenska
Vård av barn
Information om dagvård av barn i Esbo finns på InfoFinlands sida Utbildning i Esbo.
Tillfällig vård av barn
Du kan föra barnet till en parktant för tillfällig vård.
Det innebär kortvarig (2–3 tim. per gång) vård av småbarn ute i en lekpark.
Du får närmare uppgifter av parktanterna per telefon.
Du hittar telefonnumren på Esbo stads webbplats.
linkkiEsbo stad:
Parktanterfinska
Om du behöver en tillfällig barnskötare hem, kan du kontakta Mannerheims Barnskyddsförbund eller Väestöliitto.
Barnavård och hemhjälpfinska
linkkiMannerheims Barnskyddsförbund:
Barnavårdfinska _ svenska _ engelska
Läs mer: Dagvård.
Hemvårdsstöd
Om familjens yngsta barn är under tre år, kan barnets förälder få hemvårdsstöd (kotihoidon tuki) när han eller hon vårdar barnet i hemmet.
Om du har rätt till hemvårdsstödet kan du ansöka om det hos FPA.
Du kan fylla i ansökan på Internet eller posta den till FPA.
Du kan också besöka FPA:s kontor.
Esbo stad betalar ett kommuntillägg till de familjer som vårdar ett under treårigt barn i hemmet.
Man kan ansöka om Esbotillägget om en förälder tar hand om familjens alla barn under skolåldern i hemmet.
linkkiEsbo stad:
Vård av barn i hemmetfinska _ svenska _ engelska
Information om hemvårdsstödfinska _ svenska _ engelska
Sköta ärenden på Internetfinska _ svenska _ engelska
Kontaktuppgifter till FPAfinska _ svenska _ engelska
Invånarparker och klubbar
Esbo stad ordnar mycket verksamhet för de föräldrar som vårdar barn i hemmet. Det finns till exempel invånarparker, öppna daghem och klubbar.
Läs mer: Stöd för vård av barn i hemmet
linkkiEsbo stad:
Invånarparker och klubbarfinska _ engelska
Äldre människor
Åldringar kan använda tjänsterna vid de vanliga hälsostationerna.
Dessutom erbjuds åldringar i Esbo egna tjänster, till exempel hemvårdens tjänster.
Om du vill ha mer information om tjänster för äldre kan du kontakta seniorrådgivningen (seniorineuvonta).
tfn (09) 816 33333
linkkiEsbo stad:
Seniorrådgivningenfinska _ svenska _ engelska
När du tar hand om en anhörig i hemmet
Om du tar hand om en äldre, sjuk eller handikappad anhörig hemma så att hen ska kunna bo hemma, kan du ha rätt till stöd för närståendevård.
linkkiEsbo stad:
Stöd för närståendevårdfinska _ svenska
Äldre människor
Problem i familjen
På InfoFinlands sida Problematiska situationer i Esbo hittar du uppgifter om vart du kan vända dig i Esbo för att få hjälp vid barns och ungas problem och problem i familjen.
Du hittar uppgifter om barns och ungas problem också på InfoFinlands sida Barns och ungas problem och Var hittar jag hjälp när barn eller unga har problem?
På InfoFinlands sida Problem i äktenskap och parförhållande finns uppgifter om vart du kan vända dig för att få hjälp vid problem i parförhållandet.
Äktenskap
Skilsmässa
Registrerat parförhållande
Vård av barn Invånarparker och klubbar
Problem i familjen
Äktenskap
Före äktenskapet ska du skriftligt begära hindersprövning (avioliiton esteiden tutkiminen).
Hindersprövningen görs på magistraten (maistraatti).
Du kan begära hindersprövning på vilken magistrat som helst.
Magistraten i Nyland, Esbo enhet
Miestentie 3
Tfn 029 553 9391
Läs mer: Äktenskap.
Vigselfinska _ svenska _ engelska
Anhållan om prövning av hinder mot äktenskapfinska _ svenska
Skilsmässa
Kvinnan eller mannen kan lämna in skilsmässoansökan i Västra Nylands tingsrätts kansli.
Du kan också söka skilsmässa ensam, utan din makes eller makas samtycke.
Du kan skicka in ansökan till tingsrättens kansli per post, fax eller via e-post.
Tfn 029 564 4000
Läs mer: Skilsmässa.
linkkiVästra Nylands tingsrätt:
Kontaktuppgifterfinska _ svenska
Barn vid skilsmässa
Om du har barn under 13 år och överväger att skilja dig, ta kontakt med familjerådgivningen (perheneuvola).
På familjerådgivningen kan du diskutera familjens situation med de anställda.
Familjerådgivningarnas kontaktuppgifter finns på Esbo stads webbplats.
Om du planerar skilsmässa kan du också ta kontakt med barnatillsyningsmannen (lastenvalvoja) vid enheten för familjeärenden.
Med barnatillsyningsmannen kan du diskutera skilsmässan och barnens framtid.
Makarna ska ingå ett avtal om barnens boende, umgängesrätt och underhållsbidrag.
Barnatillsyningsmännen bekräftar avtalet.
Kontaktuppgifterna till barnatillsyningsmännen finns på Esbo stads webbplats.
Esbo stad har en rådgivningstelefon där man kan fråga om råd i frågor rörande barnen när föräldrarna skiljer sig.
Tfn 046 877 3267
Läs mer: Barn vid skilsmässa.
linkkiEsbo stad:
Kontaktuppgifter till barnatillsyningsmännenfinska _ svenska
linkkiEsbo stad:
Skilsmässa i en barnfamiljfinska _ svenska
Vård av barn
Information om dagvård av barn i Esbo finns på InfoFinlands sida Utbildning i Esbo.
Tillfällig vård av barn
Du kan föra barnet till en parktant för tillfällig vård.
Det innebär kortvarig (2–3 tim. per gång) vård av småbarn ute i en lekpark.
Du får närmare uppgifter av parktanterna per telefon.
Du hittar telefonnumren på Esbo stads webbplats.
linkkiEsbo stad:
Parktanterfinska _ svenska
Om du behöver en tillfällig barnskötare hem, kan du kontakta Mannerheims Barnskyddsförbund eller Väestöliitto.
Barnavård och hemhjälpfinska
linkkiMannerheims Barnskyddsförbund:
Barnavårdfinska _ svenska _ engelska
Läs mer: Dagvård.
Hemvårdsstöd
Om familjens yngsta barn är under tre år, kan barnets förälder få hemvårdsstöd (kotihoidon tuki) när han eller hon vårdar barnet i hemmet.
Om du har rätt till hemvårdsstödet kan du ansöka om det hos FPA.
Du kan fylla i ansökan på Internet eller posta den till FPA.
Du kan också besöka FPA:s kontor.
Esbo stad betalar ett kommuntillägg till de familjer som vårdar ett under treårigt barn i hemmet.
Man kan ansöka om Esbotillägget om en förälder tar hand om familjens alla barn under skolåldern i hemmet.
linkkiEsbo stad:
Vård av barn i hemmetfinska _ svenska _ engelska
Information om hemvårdsstödfinska _ svenska _ engelska
Sköta ärenden på Internetfinska _ svenska _ engelska
Kontaktuppgifter till FPAfinska _ svenska _ engelska
Invånarparker och klubbar
Esbo stad ordnar mycket verksamhet för de föräldrar som vårdar barn i hemmet. Det finns till exempel invånarparker, öppna daghem och klubbar.
Läs mer: Stöd för vård av barn i hemmet
linkkiEsbo stad:
Invånarparker och klubbarfinska _ engelska
Äldre människor
Åldringar kan använda tjänsterna vid de vanliga hälsostationerna.
Dessutom erbjuds åldringar i Esbo egna tjänster, till exempel hemvårdens tjänster.
Om du vill ha mer information om tjänster för äldre kan du kontakta seniorrådgivningen (seniorineuvonta).
tfn (09) 816 33333
linkkiEsbo stad:
Seniorrådgivningenfinska _ svenska _ engelska
När du tar hand om en anhörig i hemmet
Om du tar hand om en äldre, sjuk eller handikappad anhörig hemma så att hen ska kunna bo hemma, kan du ha rätt till stöd för närståendevård.
linkkiEsbo stad:
Stöd för närståendevårdfinska _ svenska
Äldre människor
Problem i familjen
På InfoFinlands sida Problematiska situationer i Esbo hittar du uppgifter om vart du kan vända dig i Esbo för att få hjälp vid barns och ungas problem och problem i familjen.
Du hittar uppgifter om barns och ungas problem också på InfoFinlands sida Barns och ungas problem och Var hittar jag hjälp när barn eller unga har problem?
På InfoFinlands sida Problem i äktenskap och parförhållande finns uppgifter om vart du kan vända dig för att få hjälp vid problem i parförhållandet.
Hälsovårdstjänsterna i Esbo
Äldre människors hälsa
Tandvården
Mental hälsa
Sexuell hälsa
När du väntar barn
Handikappade personer
Ring nödnumret 112 om det är fråga om en brådskande nödsituation.
Ring nödnumret till exempel vid en allvarlig olycka eller när någon drabbas av en sjukdomsattack.
Ring inte nödnumret om det inte är en nödsituation.
Om du har din hemkommun i Esbo kan du utnyttja de offentliga hälsovårdstjänsterna.
Offentliga hälsovårdstjänster tillhandahålls vid hälsostationer, tandkliniker, rådgivningsbyråer och sjukhus.
Om du inte har rätt till de offentliga hälsovårdstjänsterna, kan du söka hjälp på en privat läkarstation.
På en privat läkarstation måste du betala samtliga kostnader själv.
Läs mer: Hälsa.
Hälsovårdstjänsterna i Esbo
Offentliga hälsovårdstjänster tillhandahålls av hälsostationerna (terveysasema).
Hälsostationerna har öppet vardagar klockan 8–16.
På hälsostationerna finns vanligtvis läkarens, sjukskötarens och hälsovårdarens mottagningar.
Du kan boka tid på hälsostationen per telefon.
På Esbo stads webbplats finns kontaktuppgifterna och telefonnumren till hälsostationerna.
När du ringer hälsostationen, besvaras ditt samtal inte nödvändigtvis omedelbart.
Ditt nummer sparas dock i en automat och du blir uppringd.
Kom i tid till mottagningen.
Om du inte kan komma till mottagningen, kom ihåg att avboka din tid senast föregående vardag före klockan 14.
Om du behöver första hjälpen snabbt, kan du komma till hälsostationen utan tidsbeställning.
linkkiEsbo stad:
Hälsostationernafinska _ svenska _ engelska
linkkiEsbo stad:
Hälsovårdscentralsavgifterfinska _ svenska
Privata hälsovårdstjänster
Vem som helst kan gå till en privat hälsostation.
Också de personer som inte har rätt till den offentliga hälsovården i Finland kan besöka privata hälsostationer.
På en privat hälsostation måste kunden själv betala samtliga kostnader.
I Esbo finns flera privata läkarstationer.
Kontaktuppgifter till privata läkare hittar du till exempel på Internet.
linkkietsilaakari.fi:
Privata hälsovårdstjänsterfinska
Privat läkarstationfinska _ svenska _ engelska
Privat läkarstationfinska _ svenska _ engelska
Läkemedel
Information om köp av läkemedel hittar du på InfoFinlands sida Läkemedel.
Hälsovård för papperslösa
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärhälsovård.
Tjänsterna vid Global Clinic är avgiftsfria för kunderna.
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter.
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
Telefonnumret till Global Clinic i Helsingfors är 044 977 4547.
Samtalet besvaras av en sjukskötare eller en läkare.
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Läs mer: Hälsovårdstjänster i Finland
Kvällstid och under veckoslut har hälsostationen stängt.
Då vårdas akuta sjukfall och olycksfall på jourmottagningen (päivystys).
Den närmaste jourmottagningen för vuxna finns vid Jorv sjukhus.
Ring den kostnadsfria Jourhjälpen på tfn 116 117 innan du kommer till jourmottagningen.
Jourmottagningen vid Jorv sjukhus
Åbovägen 150
Tfn (09) 4711
Jourmottagningar för barn under 16 år finns i Jorv och på Barnkliniken i Helsingfors.
Du behöver inte boka tid på jourmottagningen.
linkkiEsbo stad:
Jourmottagningarfinska _ svenska _ engelska
Läs mer: Hälsovårdstjänster i Finland
Barns hälsa
I hälsovården av 1–6-åriga barn får man hjälp av rådgivningsbyråns (neuvola) hälsovårdare och läkare.
Dem kan du fråga om råd och få hjälp med fostran av barn.
På rådgivningsbyrån följs att barnet är friskt och växer som det ska.
I Esbo finns flera rådgivningsbyråer på olika håll i staden.
Rådgivningsbyråernas kontaktuppgifter finns på Esbo stads webbplats.
Du kan boka tid vid alla rådgivningsbyråer på samma nummer.
Om ett barn blir sjukt och behöver snabbt vård, ta kontakt med hälsostationen (terveysasema).
Skolhälsovårdaren har hand om skolbarns hälsa.
Under kvällar och veckoslut finns jourmottagningen för barn under 16 år vid Jorv sjukhus och på Barnkliniken i Helsingfors.
Du kan också ta ditt barn till en privat läkarstation.
Läs mer: Barns hälsa.
linkkiEsbo stad:
Barnrådgivningsbyråernas tjänsterfinska _ svenska _ engelska
linkkiEsbo stad:
Rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
linkkiEsbo stad:
Hälsostationernafinska _ svenska _ engelska
linkkiEsbo stad:
Information om hälsovården för skolbarnfinska _ svenska _ engelska
linkkiEsbo stad:
Jourmottagningarfinska _ svenska _ engelska
Äldre människors hälsa
Åldringar kan använda tjänsterna vid de vanliga hälsostationerna.
Dessutom erbjuds åldringar i Esbo egna tjänster, till exempel hemvårdens tjänster.
Om du vill ha mer information om tjänster för äldre kan du kontakta seniorrådgivningen (seniorineuvonta).
tfn (09) 816 33333
linkkiEsbo stad:
Seniorrådgivningenfinska _ svenska
När du tar hand om en anhörig i hemmet
Om du tar hand om en äldre, sjuk eller handikappad anhörig hemma så att hen ska kunna bo hemma, kan du ha rätt till stöd för närståendevård.
linkkiEsbo stad:
Stöd för närståendevårdfinska _ svenska
Äldre människors hälsa, Äldre människor
Tandvården
Offentlig tandvård
Du kan använda de kommunala tandläkartjänsterna om du har hemkommun i Esbo.
I nödfall kan du använda kommunala tjänster även om Esbo inte är din hemkommun.
Du kan boka tid hos en tandläkare på Esbo tandklinikers gemensamma nummer.
Tandklinikernas tidsbeställning
Tfn (09) 816 30300
Du kan ringa numret på vardagar.
Om du behöver besöka tandläkaren snabbt, ta kontakt med social- och hälsostationen i Kilo.
Social- och hälsostationen i Kilo
Trillagatan 5
Tfn (09) 816 35900
Tidsbeställning på vardagar.
Om du behöver akut tandläkarvård kvällstid eller under veckoslut, kan du kontakta Haartmanska sjukhuset i Helsingfors.
Jourmottagningen vid Haartmanska sjukhuset har öppet vardagar kl. 14–21 och lö-sö kl. 8–21.
Tfn (09) 310 49999.
linkkiEsbo stad:
Mun- och tandhälsovårdenfinska _ svenska _ engelska
Privat tandvård
I Esbo finns också privata tandläkare.
Du kan gå till en privat tandläkare även om du inte har rätt att använda den offentliga hälsovårdens tjänster.
Privat tandvård är dyrare än offentlig tandvård.
Läs mer: Tandvård.
Sök tandläkarefinska
Mental hälsa
Om du behöver hjälp eller stöd i mental- och/eller missbruksfrågor, boka tid till en psykiatriskötare.
Du kan boka tid vardagar kl. 8–16 på numret 09 816 31300.
linkkiEsbo stad:
Information om mentalvårdstjänsternafinska _ svenska _ engelska
Psykiatriskötarna har mottagning på hälsostationerna.
Mottagning för unga finns vid Nupoli.
Du kan även besöka mottagningen vid Kliniken för mental- och missbruksvård på servicetorget i Iso Omena utan tidsbokning måndag till fredag kl. 8.30–10.30 och dessutom måndag till torsdag kl. 13–14.30.
Adress: Finnviksvägen 1, Köpcentret Iso Omena.
Om du behöver krishjälp snabbt, ta kontakt med Esbo social- och krisjour (Espoon sosiaali- ja kriisipäivystys).
Social- och krisjouren
Åbovägen 150
Tfn (09) 816 42439
Öppet alla dagar dygnet runt.
linkkiEsbo stad:
Social- och krisjourenfinska _ svenska _ engelska
Läs mer: Mental hälsa.
linkkiFöreningen för mental hälsa i Finland:
Krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Information om mentalvårdstjänsternafinska _ svenska _ engelska
Sexuell hälsa
Vid hälsostationernas preventivrådgivning (ehkäisyneuvola) får du hjälp med graviditetsprevention och familjeplanering.
Ungdomar kan diskutera frågor kring sexuell hälsa med hälsovårdaren vid sin egen skola.
linkkiEsbo stad:
Preventivrådgivningsbyråerfinska _ svenska _ engelska
Om du behöver en gynekologisk undersökning, ta kontakt med hälsostationen.
Du kan också boka tid vid hälsostationen om du behöver ett recept för preventivmedel eller om du överväger abort.
Hälsostationernas kontaktuppgifter finns på Esbo stads webbplats.
linkkiEsbo stad:
Hälsostationernafinska _ svenska _ engelska
Könssjukdomar behandlas i huvudstadsregionen på polikliniken för könssjukdomar i Helsingfors.
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Polikliniken för könssjukdomarfinska _ svenska _ engelska
När du väntar barn
Kontakta rådgivningen (neuvola) när du upptäcker att du är gravid.
Vid rådgivningen följs moderns, fostrets och hela familjens hälsotillstånd under graviditeten.
I Esbo finns flera rådgivningsbyråer på olika håll i staden.
Du kan boka tid vid alla rådgivningsbyråer på samma nummer.
Rådgivning och tidsbeställning vid rådgivningsbyrån
Tfn (09) 816 22800
Läs mer: När du väntar barn.
linkkiEsbo stad:
Rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
Förlossning
I Esbo finns Jorv sjukhus där man kan föda barn.
Om du vill kan du även föda barnet på något annat sjukhus inom samkommunen Helsingfors och Nylands sjukvårdsdistrikt (HNS).
Mer information hittar du på HNS webbplats.
Läs mer: Förlossning.
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Förlossningfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Handikappade personer
Esbo stad ordnar olika tjänster för handikappade, till exempel dagverksamhet och färdtjänster.
Personer som har sin hemkommun i Esbo har rätt till dessa tjänster.
Du kan ansöka om tjänster och stödfunktioner hos stadens socialarbetare.
Mer information om tjänsterna för handikappade hittar du på Esbo stads handikappservice.
Esbo handikappservice
Kamrersvägen 2 A, vån. 4
Tfn (09) 816 45285
Läs mer: Handikappade personer
linkkiEsbo stad:
Kontaktuppgifter till socialarbetarefinska _ svenska _ engelska
linkkiEsbo stad:
Stödtjänster för handikappadefinska _ svenska _ engelska
Ett handikappat barn
Om du har ett handikappat barn kan du kontakta socialarbetaren vid handikappservicen för ditt eget område vammaispalvelut(at)espoo.fi.
Frågor som rör skolgången för ett handikappat barn kan du ställa till skolväsendet (opetustoimi) samt till servicehandledaren för skolelever (koululaisten palveluohjaaja).
Läs mer: Ett handikappat barn
linkkiEsbo stad:
Kontaktuppgifter till utbildningsväsendetfinska _ engelska
Hälsovårdstjänsterna i Esbo
Tandvården
Mental hälsa
Sexuell hälsa
När du väntar barn
Handikappade personer
Ring nödnumret 112 om det är fråga om en brådskande nödsituation.
Ring nödnumret till exempel vid en allvarlig olycka eller när någon drabbas av en sjukdomsattack.
Ring inte nödnumret om det inte är en nödsituation.
Om du har din hemkommun i Esbo kan du utnyttja de offentliga hälsovårdstjänsterna.
Offentliga hälsovårdstjänster tillhandahålls vid hälsostationer, tandkliniker, rådgivningsbyråer och sjukhus.
Om du inte har rätt till de offentliga hälsovårdstjänsterna, kan du söka hjälp på en privat läkarstation.
På en privat läkarstation måste du betala samtliga kostnader själv.
Läs mer: Hälsa.
Hälsovårdstjänsterna i Esbo
Offentliga hälsovårdstjänster tillhandahålls av hälsostationerna (terveysasema).
Hälsostationerna har öppet vardagar klockan 8–16.
På hälsostationerna finns vanligtvis läkarens, sjukskötarens och hälsovårdarens mottagningar.
Du kan boka tid på hälsostationen per telefon.
På Esbo stads webbplats finns kontaktuppgifterna och telefonnumren till hälsostationerna.
När du ringer hälsostationen, besvaras ditt samtal inte nödvändigtvis omedelbart.
Ditt nummer sparas dock i en automat och du blir uppringd.
Kom i tid till mottagningen.
Om du inte kan komma till mottagningen, kom ihåg att avboka din tid senast föregående vardag före klockan 14.
Om du behöver första hjälpen snabbt, kan du komma till hälsostationen utan tidsbeställning.
linkkiEsbo stad:
Hälsostationernafinska _ svenska _ engelska
linkkiEsbo stad:
Hälsovårdscentralsavgifterfinska _ svenska
Privata hälsovårdstjänster
Vem som helst kan gå till en privat hälsostation.
Också de personer som inte har rätt till den offentliga hälsovården i Finland kan besöka privata hälsostationer.
På en privat hälsostation måste kunden själv betala samtliga kostnader.
I Esbo finns flera privata läkarstationer.
Kontaktuppgifter till privata läkare hittar du till exempel på Internet.
linkkietsilaakari.fi:
Privata hälsovårdstjänsterfinska
Privat läkarstationfinska _ svenska _ engelska
Privat läkarstationfinska _ svenska _ engelska
Läkemedel
Information om köp av läkemedel hittar du på InfoFinlands sida Läkemedel.
Hälsovård för papperslösa
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärhälsovård.
Tjänsterna vid Global Clinic är avgiftsfria för kunderna.
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter.
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
Telefonnumret till Global Clinic i Helsingfors är 044 977 4547.
Samtalet besvaras av en sjukskötare eller en läkare.
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Läs mer: Hälsovårdstjänster i Finland
Kvällstid och under veckoslut har hälsostationen stängt.
Då vårdas akuta sjukfall och olycksfall på jourmottagningen (päivystys).
Den närmaste jourmottagningen för vuxna finns vid Jorv sjukhus.
Ring den kostnadsfria Jourhjälpen på tfn 116 117 innan du kommer till jourmottagningen.
Jourmottagningen vid Jorv sjukhus
Åbovägen 150
Tfn (09) 4711
Jourmottagningar för barn under 16 år finns i Jorv och på Barnkliniken i Helsingfors.
Du behöver inte boka tid på jourmottagningen.
linkkiEsbo stad:
Jourmottagningarfinska _ svenska _ engelska
Läs mer: Hälsovårdstjänster i Finland
Barns hälsa
I hälsovården av 1–6-åriga barn får man hjälp av rådgivningsbyråns (neuvola) hälsovårdare och läkare.
Dem kan du fråga om råd och få hjälp med fostran av barn.
På rådgivningsbyrån följs att barnet är friskt och växer som det ska.
I Esbo finns flera rådgivningsbyråer på olika håll i staden.
Rådgivningsbyråernas kontaktuppgifter finns på Esbo stads webbplats.
Du kan boka tid vid alla rådgivningsbyråer på samma nummer.
Om ett barn blir sjukt och behöver snabbt vård, ta kontakt med hälsostationen (terveysasema).
Skolhälsovårdaren har hand om skolbarns hälsa.
Under kvällar och veckoslut finns jourmottagningen för barn under 16 år vid Jorv sjukhus och på Barnkliniken i Helsingfors.
Du kan också ta ditt barn till en privat läkarstation.
Läs mer: Barns hälsa.
linkkiEsbo stad:
Barnrådgivningsbyråernas tjänsterfinska _ svenska _ engelska
linkkiEsbo stad:
Rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
linkkiEsbo stad:
Hälsostationernafinska _ svenska _ engelska
linkkiEsbo stad:
Information om hälsovården för skolbarnfinska _ svenska _ engelska
linkkiEsbo stad:
Jourmottagningarfinska _ svenska _ engelska
Tandvården
Offentlig tandvård
Du kan använda de kommunala tandläkartjänsterna om du har hemkommun i Esbo.
I nödfall kan du använda kommunala tjänster även om Esbo inte är din hemkommun.
Du kan boka tid hos en tandläkare på Esbo tandklinikers gemensamma nummer.
Tandklinikernas tidsbeställning
Tfn (09) 816 30300
Du kan ringa numret på vardagar.
Om du behöver besöka tandläkaren snabbt, ta kontakt med social- och hälsostationen i Kilo.
Social- och hälsostationen i Kilo
Trillagatan 5
Tfn (09) 816 35900
Tidsbeställning på vardagar.
Om du behöver akut tandläkarvård kvällstid eller under veckoslut, kan du kontakta Haartmanska sjukhuset i Helsingfors.
Jourmottagningen vid Haartmanska sjukhuset har öppet vardagar kl. 14–21 och lö-sö kl. 8–21.
Tfn (09) 310 49999.
linkkiEsbo stad:
Mun- och tandhälsovårdenfinska _ svenska _ engelska
Privat tandvård
I Esbo finns också privata tandläkare.
Du kan gå till en privat tandläkare även om du inte har rätt att använda den offentliga hälsovårdens tjänster.
Privat tandvård är dyrare än offentlig tandvård.
Läs mer: Tandvård.
Sök tandläkarefinska
Mental hälsa
Om du behöver hjälp eller stöd i mental- och/eller missbruksfrågor, boka tid till en psykiatriskötare.
Du kan boka tid vardagar kl. 8–16 på numret 09 816 31300.
linkkiEsbo stad:
Information om mentalvårdstjänsternafinska _ svenska _ engelska
Psykiatriskötarna har mottagning på hälsostationerna.
Mottagning för unga finns vid Nupoli.
Du kan även besöka mottagningen vid Kliniken för mental- och missbruksvård på servicetorget i Iso Omena utan tidsbokning måndag till fredag kl. 8.30–10.30 och dessutom måndag till torsdag kl. 13–14.30.
Adress: Finnviksvägen 1, Köpcentret Iso Omena.
Om du behöver krishjälp snabbt, ta kontakt med Esbo social- och krisjour (Espoon sosiaali- ja kriisipäivystys).
Social- och krisjouren
Åbovägen 150
Tfn (09) 816 42439
Öppet alla dagar dygnet runt.
linkkiEsbo stad:
Social- och krisjourenfinska _ svenska _ engelska
Läs mer: Mental hälsa.
linkkiFöreningen för mental hälsa i Finland:
Krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Information om mentalvårdstjänsternafinska _ svenska _ engelska
Sexuell hälsa
Vid hälsostationernas preventivrådgivning (ehkäisyneuvola) får du hjälp med graviditetsprevention och familjeplanering.
Ungdomar kan diskutera frågor kring sexuell hälsa med hälsovårdaren vid sin egen skola.
linkkiEsbo stad:
Preventivrådgivningsbyråerfinska _ svenska _ engelska
Om du behöver en gynekologisk undersökning, ta kontakt med hälsostationen.
Du kan också boka tid vid hälsostationen om du behöver ett recept för preventivmedel eller om du överväger abort.
Hälsostationernas kontaktuppgifter finns på Esbo stads webbplats.
linkkiEsbo stad:
Hälsostationernafinska _ svenska _ engelska
Könssjukdomar behandlas i huvudstadsregionen på polikliniken för könssjukdomar i Helsingfors.
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Polikliniken för könssjukdomarfinska _ svenska _ engelska
När du väntar barn
Kontakta rådgivningen (neuvola) när du upptäcker att du är gravid.
Vid rådgivningen följs moderns, fostrets och hela familjens hälsotillstånd under graviditeten.
I Esbo finns flera rådgivningsbyråer på olika håll i staden.
Du kan boka tid vid alla rådgivningsbyråer på samma nummer.
Rådgivning och tidsbeställning vid rådgivningsbyrån
Tfn (09) 816 22800
Läs mer: När du väntar barn.
linkkiEsbo stad:
Rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
Förlossning
I Esbo finns Jorv sjukhus där man kan föda barn.
Om du vill kan du även föda barnet på något annat sjukhus inom samkommunen Helsingfors och Nylands sjukvårdsdistrikt (HNS).
Mer information hittar du på HNS webbplats.
Läs mer: Förlossning.
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Förlossningfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Handikappade personer
Esbo stad ordnar olika tjänster för handikappade, till exempel dagverksamhet och färdtjänster.
Personer som har sin hemkommun i Esbo har rätt till dessa tjänster.
Du kan ansöka om tjänster och stödfunktioner hos stadens socialarbetare.
Mer information om tjänsterna för handikappade hittar du på Esbo stads handikappservice.
Esbo handikappservice
Kamrersvägen 2 A, vån. 4
Tfn (09) 816 45285
Handikappade personerlinkkiEsbo stad:
linkkiEsbo stad:
Stödtjänster för handikappadefinska _ svenska _ engelska
Ett handikappat barn
Om du har ett handikappat barn kan du kontakta socialarbetaren vid handikappservicen för ditt eget område vammaispalvelut(at)espoo.fi.
Frågor som rör skolgången för ett handikappat barn kan du ställa till skolväsendet (opetustoimi) samt till servicehandledaren för skolelever (koululaisten palveluohjaaja).
Läs mer: Ett handikappat barn
linkkiEsbo stad:
Kontaktuppgifter till utbildningsväsendetfinska _ engelska
Hälsovårdstjänsterna i Esbo
Tandvården
Mental hälsa
Sexuell hälsa
När du väntar barn
Handikappade personer
Ring nödnumret 112 om det är fråga om en brådskande nödsituation.
Ring nödnumret till exempel vid en allvarlig olycka eller när någon drabbas av en sjukdomsattack.
Ring inte nödnumret om det inte är en nödsituation.
Om du har din hemkommun i Esbo kan du utnyttja de offentliga hälsovårdstjänsterna.
Offentliga hälsovårdstjänster tillhandahålls vid hälsostationer, tandkliniker, rådgivningsbyråer och sjukhus.
Om du inte har rätt till de offentliga hälsovårdstjänsterna, kan du söka hjälp på en privat läkarstation.
På en privat läkarstation måste du betala samtliga kostnader själv.
Läs mer: Hälsa.
Hälsovårdstjänsterna i Esbo
Offentliga hälsovårdstjänster tillhandahålls av hälsostationerna (terveysasema).
Hälsostationerna har öppet vardagar klockan 8–16.
På hälsostationerna finns vanligtvis läkarens, sjukskötarens och hälsovårdarens mottagningar.
Du kan boka tid på hälsostationen per telefon.
På Esbo stads webbplats finns kontaktuppgifterna och telefonnumren till hälsostationerna.
När du ringer hälsostationen, besvaras ditt samtal inte nödvändigtvis omedelbart.
Ditt nummer sparas dock i en automat och du blir uppringd.
Kom i tid till mottagningen.
Om du inte kan komma till mottagningen, kom ihåg att avboka din tid senast föregående vardag före klockan 14.
Om du behöver första hjälpen snabbt, kan du komma till hälsostationen utan tidsbeställning.
linkkiEsbo stad:
Hälsostationernafinska _ svenska _ engelska
linkkiEsbo stad:
Hälsovårdscentralsavgifterfinska _ svenska
Privata hälsovårdstjänster
Vem som helst kan gå till en privat hälsostation.
Också de personer som inte har rätt till den offentliga hälsovården i Finland kan besöka privata hälsostationer.
På en privat hälsostation måste kunden själv betala samtliga kostnader.
I Esbo finns flera privata läkarstationer.
Kontaktuppgifter till privata läkare hittar du till exempel på Internet.
linkkietsilaakari.fi:
Privata hälsovårdstjänsterfinska
Privat läkarstationfinska _ svenska _ engelska
Privat läkarstationfinska _ svenska _ engelska
Läkemedel
Information om köp av läkemedel hittar du på InfoFinlands sida Läkemedel.
Hälsovård för papperslösa
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärhälsovård.
Tjänsterna vid Global Clinic är avgiftsfria för kunderna.
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter.
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
Telefonnumret till Global Clinic i Helsingfors är 044 977 4547.
Samtalet besvaras av en sjukskötare eller en läkare.
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Läs mer: Hälsovårdstjänster i Finland
Kvällstid och under veckoslut har hälsostationen stängt.
Då vårdas akuta sjukfall och olycksfall på jourmottagningen (päivystys).
Den närmaste jourmottagningen för vuxna finns vid Jorv sjukhus.
Ring den kostnadsfria Jourhjälpen på tfn 116 117 innan du kommer till jourmottagningen.
Jourmottagningen vid Jorv sjukhus
Åbovägen 150
Tfn (09) 4711
Jourmottagningar för barn under 16 år finns i Jorv och på Barnkliniken i Helsingfors.
Du behöver inte boka tid på jourmottagningen.
linkkiEsbo stad:
Jourmottagningarfinska _ svenska _ engelska
Läs mer: Hälsovårdstjänster i Finland
Barns hälsa
I hälsovården av 1–6-åriga barn får man hjälp av rådgivningsbyråns (neuvola) hälsovårdare och läkare.
Dem kan du fråga om råd och få hjälp med fostran av barn.
På rådgivningsbyrån följs att barnet är friskt och växer som det ska.
I Esbo finns flera rådgivningsbyråer på olika håll i staden.
Rådgivningsbyråernas kontaktuppgifter finns på Esbo stads webbplats.
Du kan boka tid vid alla rådgivningsbyråer på samma nummer.
Om ett barn blir sjukt och behöver snabbt vård, ta kontakt med hälsostationen (terveysasema).
Skolhälsovårdaren har hand om skolbarns hälsa.
Under kvällar och veckoslut finns jourmottagningen för barn under 16 år vid Jorv sjukhus och på Barnkliniken i Helsingfors.
Du kan också ta ditt barn till en privat läkarstation.
Läs mer: Barns hälsa.
linkkiEsbo stad:
Barnrådgivningsbyråernas tjänsterfinska _ svenska _ engelska
linkkiEsbo stad:
Rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
linkkiEsbo stad:
Hälsostationernafinska _ svenska _ engelska
linkkiEsbo stad:
Information om hälsovården för skolbarnfinska _ svenska _ engelska
linkkiEsbo stad:
Jourmottagningarfinska _ svenska _ engelska
Tandvården
Offentlig tandvård
Du kan använda de kommunala tandläkartjänsterna om du har hemkommun i Esbo.
I nödfall kan du använda kommunala tjänster även om Esbo inte är din hemkommun.
Du kan boka tid hos en tandläkare på Esbo tandklinikers gemensamma nummer.
Tandklinikernas tidsbeställning
Tfn (09) 816 30300
Du kan ringa numret på vardagar.
Om du behöver besöka tandläkaren snabbt, ta kontakt med social- och hälsostationen i Kilo.
Social- och hälsostationen i Kilo
Trillagatan 5
Tfn (09) 816 35900
Tidsbeställning på vardagar.
Om du behöver akut tandläkarvård kvällstid eller under veckoslut, kan du kontakta Haartmanska sjukhuset i Helsingfors.
Jourmottagningen vid Haartmanska sjukhuset har öppet vardagar kl. 14–21 och lö-sö kl. 8–21.
Tfn (09) 310 49999.
linkkiEsbo stad:
Mun- och tandhälsovårdenfinska _ svenska _ engelska
Privat tandvård
I Esbo finns också privata tandläkare.
Du kan gå till en privat tandläkare även om du inte har rätt att använda den offentliga hälsovårdens tjänster.
Privat tandvård är dyrare än offentlig tandvård.
Läs mer: Tandvård.
Sök tandläkarefinska
Mental hälsa
Om du behöver hjälp eller stöd i mental- och/eller missbruksfrågor, boka tid till en psykiatriskötare.
Du kan boka tid vardagar kl. 8–16 på numret 09 816 31300.
linkkiEsbo stad:
Information om mentalvårdstjänsternafinska _ svenska _ engelska
Psykiatriskötarna har mottagning på hälsostationerna.
Mottagning för unga finns vid Nupoli.
Du kan även besöka mottagningen vid Kliniken för mental- och missbruksvård på servicetorget i Iso Omena utan tidsbokning måndag till fredag kl. 8.30–10.30 och dessutom måndag till torsdag kl. 13–14.30.
Adress: Finnviksvägen 1, Köpcentret Iso Omena.
Om du behöver krishjälp snabbt, ta kontakt med Esbo social- och krisjour (Espoon sosiaali- ja kriisipäivystys).
Social- och krisjouren
Åbovägen 150
Tfn (09) 816 42439
Öppet alla dagar dygnet runt.
linkkiEsbo stad:
Social- och krisjourenfinska _ svenska _ engelska
Läs mer: Mental hälsa.
linkkiFöreningen för mental hälsa i Finland:
Krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Information om mentalvårdstjänsternafinska _ svenska _ engelska
Sexuell hälsa
Vid hälsostationernas preventivrådgivning (ehkäisyneuvola) får du hjälp med graviditetsprevention och familjeplanering.
Ungdomar kan diskutera frågor kring sexuell hälsa med hälsovårdaren vid sin egen skola.
linkkiEsbo stad:
Preventivrådgivningsbyråerfinska _ svenska _ engelska
Om du behöver en gynekologisk undersökning, ta kontakt med hälsostationen.
Du kan också boka tid vid hälsostationen om du behöver ett recept för preventivmedel eller om du överväger abort.
Hälsostationernas kontaktuppgifter finns på Esbo stads webbplats.
linkkiEsbo stad:
Hälsostationernafinska _ svenska _ engelska
Könssjukdomar behandlas i huvudstadsregionen på polikliniken för könssjukdomar i Helsingfors.
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Polikliniken för könssjukdomarfinska _ svenska _ engelska
Läs mer: Sexualhälsa
När du väntar barn
Kontakta rådgivningen (neuvola) när du upptäcker att du är gravid.
Vid rådgivningen följs moderns, fostrets och hela familjens hälsotillstånd under graviditeten.
I Esbo finns flera rådgivningsbyråer på olika håll i staden.
Du kan boka tid vid alla rådgivningsbyråer på samma nummer.
Rådgivning och tidsbeställning vid rådgivningsbyrån
Tfn (09) 816 22800
Läs mer: Graviditet och förlossning.
linkkiEsbo stad:
Rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
Förlossning
I Esbo finns Jorv sjukhus där man kan föda barn.
Om du vill kan du även föda barnet på något annat sjukhus inom samkommunen Helsingfors och Nylands sjukvårdsdistrikt (HNS).
Mer information hittar du på HNS webbplats.
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Förlossningfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Handikappade personer
Esbo stad ordnar olika tjänster för handikappade, till exempel dagverksamhet och färdtjänster.
Personer som har sin hemkommun i Esbo har rätt till dessa tjänster.
Du kan ansöka om tjänster och stödfunktioner hos stadens socialarbetare.
Mer information om tjänsterna för handikappade hittar du på Esbo stads handikappservice.
Esbo handikappservice
Kamrersvägen 2 A, vån. 4
Tfn (09) 816 45285
Läs mer: Handikappade personer
linkkiEsbo stad:
Stödtjänster för handikappadefinska _ svenska _ engelska
Ett handikappat barn
Om du har ett handikappat barn kan du kontakta socialarbetaren vid handikappservicen för ditt eget område vammaispalvelut(at)espoo.fi.
Frågor som rör skolgången för ett handikappat barn kan du ställa till skolväsendet (opetustoimi) samt till servicehandledaren för skolelever (koululaisten palveluohjaaja).
Läs mer: Ett handikappat barn
linkkiEsbo stad:
Kontaktuppgifter till utbildningsväsendetfinska _ engelska
Detta innehåll finns inte på det språk som du har valt.
Välj något annat språk.
Finska
Detta innehåll finns inte på det språk som du har valt.
Välj något annat språk.
Finska
Detta innehåll finns inte på det språk som du har valt.
Välj något annat språk.
Finska
Dagvård
Förskoleundervisning
Grundläggande utbildning
Hemspråksundervisning för invandrare
Yrkesutbildning
Gymnasium
Stöd och handledning för unga
Högskoleutbildning
Andra studiemöjligheter
Dagvård
I Esbo finns både kommunala och privata daghem.
I Esbo finns dessutom familjedagvårdare.
Dagvård fås på finska och på svenska.
Ansök om dagvårdsplats minst fyra månader innan barnet ska börja i dagvården.
Om du till exempel oväntat får arbete eller en studieplats kan du ansöka om vårdplats senare.
När du ansöker om vårdplats ska du fylla i en ansökningsblankett.
Du kan också söka dagvårdsplats via Internet.
Familjer som bor i Esbo kan också söka dagvårdsplats till sitt barn i Helsingfors, Vanda eller Grankulla.
Du ska ändå lämna in din ansökan i Esbo.
Mer information får du via tjänsten Helsingforsregionen.fi.
Läs mer: Dagvård.
linkkiEsbo stad:
Dagvårdfinska _ svenska _ engelska
linkkiEsbo stad:
Ansökan om dagvårdsplatsfinska
linkkiEsbo stad:
Servicepunktfinska _ svenska _ engelska
linkkiEsbo stad:
Dagvårdens samanvändningsområdefinska _ svenska _ engelska
Förskoleundervisning
I Esbo anordnas förskoleundervisningen (esiopetus) i daghemmen.
Förskoleundervisning ges på finska och på svenska.
Till förskoleundervisningen anmäler man sig via Esbo stads webbplats.
Förskoleundervisningen börjar i augusti.
Ansökningstiden är vanligtvis i januari.
I frågor kring barndagvård och förskoleundervisning kan du också kontakta daghemsföreståndarna eller stadens chef för småbarnsfostran (varhaiskasvatuspäällikkö).
Kontaktuppgifterna finns på stadens webbplats.
Läs mer: Förskoleundervisning.
linkkiEsbo stad:
Förskoleundervisningfinska _ svenska _ engelska
linkkiEsbo stad:
Ansökan till förskoleundervisningfinska _ svenska _ engelska
Grundläggande utbildning
I Esbo finns finskspråkiga och svenskspråkiga grundskolor (peruskoulu).
Undervisning kan även fås på engelska.
Skolan börjar vanligtvis det året då barnet fyller sju år.
Anmälan till grundskolan ska göras på förhand.
Anmälningstiden är vanligtvis i januari.
På stadens webbplats hittar du kontaktuppgifterna till skolorna och mer information om anmälan.
Om du har frågor om den grundläggande utbildningen kan du kontakta Resultatenheten för den finskspråkiga undervisningen (Suomenkielisen opetuksen tulosyksikkö).
Resultatenheten för den finskspråkiga undervisningen
Kamrersvägen 3 B
Tfn (09) 816 52044 och (09) 816 52043
Grundläggande utbildning.
linkkiEsbo stad:
Grundläggande utbildningfinska _ svenska _ engelska
linkkiEsbo stad:
Anmälan till skolanfinska _ svenska _ engelska
linkkiEsbo stad:
Espoo International Schoolfinska _ engelska
Internationella skolor i huvudstadsregionenfinska
linkkiExpatFinland.fi:
Internationella skolor i huvudstadsregionenengelska
linkkiEsbo stad:
Eftermiddagsverksamhetfinska _ engelska
Hemspråksundervisning för invandrare
Barn med invandrarbakgrund och barn från tvåspråkiga familjer kan få hemspråksundervisning (oman äidinkielen opetus) om tillräckligt många barn anmäler sig till gruppen för det egna språket.
Undervisning ges två timmar i veckan.
Anmälan till hemspråksundervisning görs varje år i mars.
Mer information hittar du på Esbo stads webbplats.
linkkiEsbo stad:
Förberedande undervisning för barn i förskoleåldern(pdf, 100 kb)finska _ engelska _ ryska _ estniska _ somaliska _ kinesiska _ arabiska _ kurdiska _ albanska
linkkiEsbo stad:
Förberedande undervisning för barn i förskoleåldernfinska _ engelska
linkkiEsbo stad:
Hemspråksundervisningfinska _ engelska
Yrkesutbildning
På Omnia kan man studera många olika yrken.
På Omnia ordnas för invandrare utbildning som förbereder dem på yrkesutbildning.
Den förberedande utbildningen är avsedd för unga och vuxna, som är intresserade av yrkesstudier och vill förbättra sina kunskaper i finska..
Esbobor kan också ansöka till yrkesskolorna i Helsingfors och Vanda.
Läs mer: Yrkesutbildning
Yrkesutbildningfinska _ engelska
linkkiEsbo stad:
Yrkesläroanstalterfinska _ engelska
Yrkesläroanstalterfinska _ svenska _ engelska
linkkiVanda stad:
Yrkesutbildningfinska _ svenska
Gymnasium
I Esbo finns elva finskspråkiga och ett svenskspråkigt gymnasium (lukio).
I två av gymnasierna i Esbo finns en engelskspråkig IB-linje.
Ungdomar från Esbo kan också söka till gymnasier i andra städer.
I Esbo finns ett vuxengymnasium (aikuislukio) där vuxna kan avlägga gymnasie- och studentexamen.
På gymnasiet kan man även höja vitsorden i sitt avgångsbetyg eller studera enskilda ämnen.
Invandrarungdomar kan dessutom studera finska och avlägga grundskolans lärokurs.
I gymnasiet Leppävaaran lukio ordnas för invandrare och utlänningar utbildning som förbereder dem på gymnasiet.
Utbildningen är avsedd för unga som vill studera på gymnasiet, men vars språkkunskaper inte är tillräckliga för gymnasiestudier.
Läs mer: Gymnasium
linkkiEsbo stad:
Gymnasierfinska _ svenska _ engelska
linkkiEsbo stad:
Vuxengymnasietfinska
linkkiEsbo stad:
Gymnasieförberedande utbildning för invandrarefinska _ engelska
linkkiEsbo vuxengymnasium Omnia:
Grundläggande utbildning för invandrarefinska
Om du är under 30 år gammal kan du få råd och handledning via Ohjaamo-tjänsten.
Ohjaamos personal hjälper dig om du inte har ett arbete eller en studieplats.
Du kan även fråga om andra saker, som till exempel boende eller ekonomiska frågor.
Kontaktuppgifter:
Fågelbergavägen 2 A
Puh. 040 126 7513
linkkiEsbo stad:
Ohjaamofinska _ svenska _ engelska
Högskoleutbildning
I Esbo finns tre högskolor:
yrkeshögskolan Laurea
yrkeshögskolan Metropolia.
Vid högskolorna kan du avlägga högskoleexamen.
Mer information finns på Aalto-universitetets, Laureas och Metropolias webbplatser.
Också i Helsingfors finns det universitet och yrkeshögskolor där man kan studera inom många områden.
Mer information hittar du på Helsingfors stads webbplats.
Läs mer: Högskoleutbildning
Universitet inom teknik, konst och ekonomifinska _ svenska _ engelska
Yrkeshögskolafinska _ engelska
linkkiMetropolia:
Yrkeshögskolafinska _ engelska
Högskolorfinska
Andra studiemöjligheter
Vid Esbo arbetarinstitut (Espoon työväenopisto) kan du studera till exempel språk, handarbete och matlagning eller delta i ledd motion.
Kurserna är avgiftsbelagda. Kurser anordnas både dagtid och kvällstid.
Vid arbetarinstitutet kan vem som helst studera.
Vid Esbo bildkonstskola (Espoon kuvataidekoulu) kan barn och unga studera bildkonst.
Studierna är avgiftsbelagda.
Vid Esbo musikinstitut (Espoon musiikkiopisto) kan barn och vuxna studera musik.
Läs mer: Andra studiemöjligheter
linkkiEsbo stad:
Arbetarinstitutetfinska _ svenska _ engelska
linkkiEsbo biIdkonstskola:
Bildkonst för barn och ungafinska _ svenska _ engelska
linkkiEsbo musikinstitut:
Musikundervisning för barn och vuxnafinska _ engelska
Dagvård
Förskoleundervisning
Grundläggande utbildning
Hemspråksundervisning för invandrare
Yrkesutbildning
Gymnasium
Stöd och handledning för unga
Högskoleutbildning
Andra studiemöjligheter
Dagvård
I Esbo finns både kommunala och privata daghem.
I Esbo finns dessutom familjedagvårdare.
Dagvård fås på finska och på svenska.
Ansök om dagvårdsplats minst fyra månader innan barnet ska börja i dagvården.
Om du till exempel oväntat får arbete eller en studieplats kan du ansöka om vårdplats senare.
När du ansöker om vårdplats ska du fylla i en ansökningsblankett.
Du kan också söka dagvårdsplats via Internet.
Familjer som bor i Esbo kan också söka dagvårdsplats till sitt barn i Helsingfors, Vanda eller Grankulla.
Du ska ändå lämna in din ansökan i Esbo.
Mer information får du via tjänsten Helsingforsregionen.fi.
Läs mer: Dagvård.
linkkiEsbo stad:
Dagvårdfinska _ svenska _ engelska
linkkiEsbo stad:
Ansökan om dagvårdsplatsfinska
linkkiEsbo stad:
Servicepunktfinska _ svenska _ engelska
linkkiEsbo stad:
Dagvårdens samanvändningsområdefinska _ svenska _ engelska
Förskoleundervisning
I Esbo anordnas förskoleundervisningen (esiopetus) i daghemmen.
Förskoleundervisning ges på finska och på svenska.
Till förskoleundervisningen anmäler man sig via Esbo stads webbplats.
Förskoleundervisningen börjar i augusti.
Ansökningstiden är vanligtvis i januari.
I frågor kring barndagvård och förskoleundervisning kan du också kontakta daghemsföreståndarna eller stadens chef för småbarnsfostran (varhaiskasvatuspäällikkö).
Kontaktuppgifterna finns på stadens webbplats.
Läs mer: Förskoleundervisning.
linkkiEsbo stad:
Förskoleundervisningfinska _ svenska _ engelska
linkkiEsbo stad:
Ansökan till förskoleundervisningfinska _ engelska
Grundläggande utbildning
I Esbo finns finskspråkiga och svenskspråkiga grundskolor (peruskoulu).
Undervisning kan även fås på engelska.
Skolan börjar vanligtvis det året då barnet fyller sju år.
Anmälan till grundskolan ska göras på förhand.
Anmälningstiden är vanligtvis i januari.
På stadens webbplats hittar du kontaktuppgifterna till skolorna och mer information om anmälan.
Om du har frågor om den grundläggande utbildningen kan du kontakta Resultatenheten för den finskspråkiga undervisningen (Suomenkielisen opetuksen tulosyksikkö).
Resultatenheten för den finskspråkiga undervisningen
Kamrersvägen 3 B
Tfn (09) 816 52044 och (09) 816 52043
Grundläggande utbildning.
linkkiEsbo stad:
Grundläggande utbildningfinska _ svenska _ engelska
linkkiEsbo stad:
Anmälan till skolanfinska _ svenska _ engelska
linkkiEsbo stad:
Espoo International Schoolfinska _ engelska
Internationella skolor i huvudstadsregionenfinska
linkkiExpatFinland.fi:
Internationella skolor i huvudstadsregionenengelska
linkkiEsbo stad:
Eftermiddagsverksamhetfinska _ engelska
Hemspråksundervisning för invandrare
Barn med invandrarbakgrund och barn från tvåspråkiga familjer kan få hemspråksundervisning (oman äidinkielen opetus) om tillräckligt många barn anmäler sig till gruppen för det egna språket.
Undervisning ges två timmar i veckan.
Anmälan till hemspråksundervisning görs varje år i mars.
Mer information hittar du på Esbo stads webbplats.
linkkiEsbo stad:
Förberedande undervisning för barn i förskoleåldern(pdf, 100 kb)finska _ engelska _ ryska _ estniska _ somaliska _ kinesiska _ arabiska _ kurdiska _ albanska
linkkiEsbo stad:
Förberedande undervisning för barn i förskoleåldernfinska _ engelska
linkkiEsbo stad:
Hemspråksundervisningfinska _ engelska
Yrkesutbildning
På Omnia kan man studera många olika yrken.
På Omnia ordnas för invandrare utbildning som förbereder dem på yrkesutbildning.
Den förberedande utbildningen är avsedd för unga och vuxna, som är intresserade av yrkesstudier och vill förbättra sina kunskaper i finska..
Esbobor kan också ansöka till yrkesskolorna i Helsingfors och Vanda.
Läs mer: Yrkesutbildning
Yrkesutbildningfinska _ engelska
linkkiEsbo stad:
Yrkesläroanstalterfinska _ engelska
Yrkesläroanstalterfinska _ svenska _ engelska
linkkiVanda stad:
Yrkesutbildningfinska _ svenska
Gymnasium
I Esbo finns elva finskspråkiga och ett svenskspråkigt gymnasium (lukio).
I två av gymnasierna i Esbo finns en engelskspråkig IB-linje.
Ungdomar från Esbo kan också söka till gymnasier i andra städer.
I Esbo finns ett vuxengymnasium (aikuislukio) där vuxna kan avlägga gymnasie- och studentexamen.
På gymnasiet kan man även höja vitsorden i sitt avgångsbetyg eller studera enskilda ämnen.
Invandrarungdomar kan dessutom studera finska och avlägga grundskolans lärokurs.
I gymnasiet Leppävaaran lukio ordnas för invandrare och utlänningar utbildning som förbereder dem på gymnasiet.
Utbildningen är avsedd för unga som vill studera på gymnasiet, men vars språkkunskaper inte är tillräckliga för gymnasiestudier.
Läs mer: Gymnasium
linkkiEsbo stad:
Gymnasierfinska _ svenska _ engelska
linkkiEsbo stad:
Vuxengymnasietfinska
linkkiEsbo stad:
Gymnasieförberedande utbildning för invandrarefinska _ engelska
linkkiEsbo vuxengymnasium Omnia:
Grundläggande utbildning för invandrarefinska
Om du är under 30 år gammal kan du få råd och handledning via Ohjaamo-tjänsten.
Ohjaamos personal hjälper dig om du inte har ett arbete eller en studieplats.
Du kan även fråga om andra saker, som till exempel boende eller ekonomiska frågor.
Kontaktuppgifter:
Fågelbergavägen 2 A
Puh. 040 126 7513
linkkiEsbo stad:
Ohjaamofinska _ svenska _ engelska
Högskoleutbildning
I Esbo finns tre högskolor:
yrkeshögskolan Laurea
yrkeshögskolan Metropolia.
Vid högskolorna kan du avlägga högskoleexamen.
Mer information finns på Aalto-universitetets, Laureas och Metropolias webbplatser.
Också i Helsingfors finns det universitet och yrkeshögskolor där man kan studera inom många områden.
Mer information hittar du på Helsingfors stads webbplats.
Läs mer: Högskoleutbildning
Universitet inom teknik, konst och ekonomifinska _ svenska _ engelska
Yrkeshögskolafinska _ engelska
linkkiMetropolia:
Yrkeshögskolafinska _ engelska
Högskolorfinska
Andra studiemöjligheter
Vid Esbo arbetarinstitut (Espoon työväenopisto) kan du studera till exempel språk, handarbete och matlagning eller delta i ledd motion.
Kurserna är avgiftsbelagda. Kurser anordnas både dagtid och kvällstid.
Vid arbetarinstitutet kan vem som helst studera.
Vid Esbo bildkonstskola (Espoon kuvataidekoulu) kan barn och unga studera bildkonst.
Studierna är avgiftsbelagda.
Vid Esbo musikinstitut (Espoon musiikkiopisto) kan barn och vuxna studera musik.
Läs mer: Andra studiemöjligheter
linkkiEsbo stad:
Arbetarinstitutetfinska _ svenska _ engelska
linkkiEsbo biIdkonstskola:
Bildkonst för barn och ungafinska _ svenska _ engelska
linkkiEsbo musikinstitut:
Musikundervisning för barn och vuxnafinska _ engelska
Dagvård
Förskoleundervisning
Grundläggande utbildning
Hemspråksundervisning för invandrare
Yrkesutbildning
Gymnasium
Stöd och handledning för unga
Högskoleutbildning
Andra studiemöjligheter
Dagvård
I Esbo finns både kommunala och privata daghem.
I Esbo finns dessutom familjedagvårdare.
Dagvård fås på finska och på svenska.
Ansök om dagvårdsplats minst fyra månader innan barnet ska börja i dagvården.
Om du till exempel oväntat får arbete eller en studieplats kan du ansöka om vårdplats senare.
När du ansöker om vårdplats ska du fylla i en ansökningsblankett.
Du kan också söka dagvårdsplats via Internet.
Familjer som bor i Esbo kan också söka dagvårdsplats till sitt barn i Helsingfors, Vanda eller Grankulla.
Du ska ändå lämna in din ansökan i Esbo.
Mer information får du via tjänsten Helsingforsregionen.fi.
Läs mer: Småbarnspedagogik
linkkiEsbo stad:
Dagvårdfinska _ svenska _ engelska
linkkiEsbo stad:
Ansökan om dagvårdsplatsfinska _ engelska
linkkiEsbo stad:
Servicepunktfinska _ svenska _ engelska
linkkiEsbo stad:
Dagvårdens samanvändningsområdefinska _ svenska _ engelska
Förskoleundervisning
I Esbo anordnas förskoleundervisningen (esiopetus) i daghemmen.
Förskoleundervisning ges på finska och på svenska.
Till förskoleundervisningen anmäler man sig via Esbo stads webbplats.
Förskoleundervisningen börjar i augusti.
Ansökningstiden är vanligtvis i januari.
I frågor kring barndagvård och förskoleundervisning kan du också kontakta daghemsföreståndarna eller stadens chef för småbarnsfostran (varhaiskasvatuspäällikkö).
Kontaktuppgifterna finns på stadens webbplats.
Läs mer: Förskoleundervisning.
linkkiEsbo stad:
Förskoleundervisningfinska _ svenska _ engelska
linkkiEsbo stad:
Ansökan till förskoleundervisningfinska _ engelska
Grundläggande utbildning
I Esbo finns finskspråkiga och svenskspråkiga grundskolor (peruskoulu).
Undervisning kan även fås på engelska.
Skolan börjar vanligtvis det året då barnet fyller sju år.
Anmälan till grundskolan ska göras på förhand.
Anmälningstiden är vanligtvis i januari.
På stadens webbplats hittar du kontaktuppgifterna till skolorna och mer information om anmälan.
Om du har frågor om den grundläggande utbildningen kan du kontakta Resultatenheten för den finskspråkiga undervisningen (Suomenkielisen opetuksen tulosyksikkö).
Resultatenheten för den finskspråkiga undervisningen
Kamrersvägen 3 B
Tfn (09) 816 52044 och (09) 816 52043
Grundläggande utbildning.
linkkiEsbo stad:
Grundläggande utbildningfinska _ svenska _ engelska
linkkiEsbo stad:
Anmälan till skolanfinska _ svenska _ engelska
linkkiEsbo stad:
Espoo International Schoolfinska _ engelska
Internationella skolor i huvudstadsregionenfinska
linkkiExpatFinland.fi:
Internationella skolor i huvudstadsregionenengelska
linkkiEsbo stad:
Eftermiddagsverksamhetfinska _ engelska
Hemspråksundervisning för invandrare
Barn med invandrarbakgrund och barn från tvåspråkiga familjer kan få hemspråksundervisning (oman äidinkielen opetus) om tillräckligt många barn anmäler sig till gruppen för det egna språket.
Undervisning ges två timmar i veckan.
Anmälan till hemspråksundervisning görs varje år i mars.
Mer information hittar du på Esbo stads webbplats.
linkkiEsbo stad:
Förberedande undervisning för barn i förskoleåldern(pdf, 100 kb)finska _ engelska _ ryska _ estniska _ somaliska _ kinesiska _ arabiska _ kurdiska _ albanska
linkkiEsbo stad:
Förberedande undervisning för barn i förskoleåldernfinska _ engelska
linkkiEsbo stad:
Hemspråksundervisningfinska _ engelska
Yrkesutbildning
På Omnia kan man studera många olika yrken.
På Omnia ordnas för invandrare utbildning som förbereder dem på yrkesutbildning.
Den förberedande utbildningen är avsedd för unga och vuxna, som är intresserade av yrkesstudier och vill förbättra sina kunskaper i finska..
Esbobor kan också ansöka till yrkesskolorna i Helsingfors och Vanda.
Läs mer: Yrkesutbildning
Yrkesutbildningfinska _ engelska
linkkiEsbo stad:
Yrkesläroanstalterfinska _ engelska
Yrkesläroanstalterfinska _ svenska _ engelska
linkkiVanda stad:
Yrkesutbildningfinska _ svenska
Gymnasium
I Esbo finns elva finskspråkiga och ett svenskspråkigt gymnasium (lukio).
I två av gymnasierna i Esbo finns en engelskspråkig IB-linje.
Ungdomar från Esbo kan också söka till gymnasier i andra städer.
I Esbo finns ett vuxengymnasium (aikuislukio) där vuxna kan avlägga gymnasie- och studentexamen.
På gymnasiet kan man även höja vitsorden i sitt avgångsbetyg eller studera enskilda ämnen.
Invandrarungdomar kan dessutom studera finska och avlägga grundskolans lärokurs.
I gymnasiet Leppävaaran lukio ordnas för invandrare och utlänningar utbildning som förbereder dem på gymnasiet.
Utbildningen är avsedd för unga som vill studera på gymnasiet, men vars språkkunskaper inte är tillräckliga för gymnasiestudier.
Läs mer: Gymnasium
linkkiEsbo stad:
Gymnasierfinska _ svenska _ engelska
linkkiEsbo stad:
Vuxengymnasietfinska
linkkiEsbo stad:
Gymnasieförberedande utbildning för invandrarefinska _ engelska
linkkiEsbo vuxengymnasium Omnia:
Grundläggande utbildning för invandrarefinska
Om du är under 30 år gammal kan du få råd och handledning via Ohjaamo-tjänsten.
Ohjaamos personal hjälper dig om du inte har ett arbete eller en studieplats.
Du kan även fråga om andra saker, som till exempel boende eller ekonomiska frågor.
Kontaktuppgifter:
Fågelbergavägen 2 A
Puh. 040 126 7513
linkkiEsbo stad:
Ohjaamofinska _ svenska _ engelska
Högskoleutbildning
I Esbo finns tre högskolor:
yrkeshögskolan Laurea
yrkeshögskolan Metropolia.
Vid högskolorna kan du avlägga högskoleexamen.
Mer information finns på Aalto-universitetets, Laureas och Metropolias webbplatser.
Också i Helsingfors finns det universitet och yrkeshögskolor där man kan studera inom många områden.
Mer information hittar du på Helsingfors stads webbplats.
Läs mer: Yrkeshögskolor
Universitet inom teknik, konst och ekonomifinska _ svenska _ engelska
Yrkeshögskolafinska _ engelska
linkkiMetropolia:
Yrkeshögskolafinska _ engelska
Högskolorfinska
Andra studiemöjligheter
Vid Esbo arbetarinstitut (Espoon työväenopisto) kan du studera till exempel språk, handarbete och matlagning eller delta i ledd motion.
Kurserna är avgiftsbelagda. Kurser anordnas både dagtid och kvällstid.
Vid arbetarinstitutet kan vem som helst studera.
Vid Esbo bildkonstskola (Espoon kuvataidekoulu) kan barn och unga studera bildkonst.
Studierna är avgiftsbelagda.
Vid Esbo musikinstitut (Espoon musiikkiopisto) kan barn och vuxna studera musik.
Läs mer: Studier som hobby
linkkiEsbo stad:
Arbetarinstitutetfinska _ svenska _ engelska
linkkiEsbo biIdkonstskola:
Bildkonst för barn och ungafinska _ svenska _ engelska
linkkiEsbo musikinstitut:
Musikundervisning för barn och vuxnafinska _ engelska
Hyresbostad
Ägarbostad
Bostadsrättsbostad
Delägarbostad
Tillfälligt boende
Boende i en krissituation
Stöd- och serviceboende
Bostadslöshet
Avfallshantering och återvinning
Hyresbostad
I Esbo och huvudstadsregionen är hyrorna ofta högre än i resten av Finland.
Det kan vara svårt att hitta en bostad med lämplig hyra.
Det lönar sig att avsätta tid för bostadssökandet och undersöka olika alternativ.
Privata hyresbostäder
Hos en privat hyresvärd kan det gå snabbt att få en bostad, men hyran kan vara högre än i stadens hyresbostäder.
Du kan söka privata hyresbostäder i Esbo via hyresvärdarnas webbplatser:
Sökning av hyresbostäderfinska
Sökning av hyresbostäderfinska _ engelska
Hyresbostäder för ungafinska _ engelska
Hyresbostäder för ungafinska _ engelska
Om du är studerande kan du få en hyresbostad för studerande i Esbo.
Hyresbostäder för studerande erbjuds av Helsingforsregionens studentbostadsstiftelse HOAS och Aalto-universitets studentkår AUS.
linkkiHOAS:
Hyresbostäder för studerandefinska _ svenska _ engelska
Hyresbostäder för studerandefinska _ svenska _ engelska
Stadens hyresbostäder
Stadens hyresbostäder är ofta billigare än bostäder som man hyr av företag eller privatpersoner.
Det är dock många som ansöker om stadens bostäder och endast en liten del av de sökande får en bostad.
Störst är bristen på små bostäder.
Stadens hyresbostäder förvaltas av Espoon Asunnot Oy (Espoon Asunnot Oy).
Om du vill ansöka om en hyresbostad, fyll i en ansökningsblankett för hyresbostad på Espoon Asunnot Oy:s webbplats.
Du kan även fylla i ansökningsblanketten på Espoon Asunnot Oy:s kontor.
Du kan också få blanketten hemskickad per post.
Dina möjligheter att få en bostad påverkas av ditt bostadsbehov och dina tillgångar och inkomster.
För att kunna ansöka om en hyresbostad hos staden, måste du ha uppehållstillstånd för minst ett år.
Tfn (09) 816 5800
Ansökan är giltig i tre månader.
Efter det måste du förnya din ansökan om du fortfarande letar efter bostad.
Läs mer: Hyresbostad
linkkiEsbo Bostäder Ab:
Ansökan om hyresbostad i stadenfinska _ engelska
linkkiEsbo stad:
Stadens hyresbostäderfinska _ svenska _ engelska
linkkiEsbo stad:
Seniorbostäderfinska _ svenska
Ägarbostad
På internet finns många bostadsförsäljningsannonser. Bostäderna i Esbo är tämligen dyra.
Information om köp av bostad hittar du på InfoFinlands sida Ägarbostad.
Bostadsrättsbostad
Om du ansöker om en bostadsrättsbostad, behöver du ett ordningsnummer. Du ansöker om ordningsnumret vid Esbo eller Helsingfors stad.
Läs mer: Bostadsrättsbostad.
linkkiEsbo stad:
Bostadsrättsbostäderfinska _ svenska _ engelska
Delägarbostad
Asuntosäätiö har delägarbostäder i Esbo.
Mer information hittar du på Asuntosäätiös webbplats.
Läs mer: Delägarbostad.
Delägarbostadfinska
Tillfälligt boende
I Esbo finns många olika hotell där man kan bo tillfälligt.
Läs mer: Tillfälligt boende.
linkkiVisitEspoo.fi:
Hotellfinska _ svenska _ engelska _ ryska _ kinesiska
Brand eller vattenskada
Om din bostad har skadats till exempel till följd av brand eller vattenskada kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
Kontakta ditt försäkringsbolag direkt när skadan har inträffat.
Våld i hemmet
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta tjänsten Omatila (Omatila).
Omatila ordnar vid behov boende för dig och dina barn.
Omatila-tjänsten
Kamrersvägen 6 A
Tfn 043 825 0535
Öppet
Lördag-söndag kl. 9-16
Social- och krisjouren 24 h
Tfn 09 816 42439
linkkiEsbo stad:
Hjälp till offer för familjevåldfinska _ svenska _ engelska
Om du är ung och har problem hemma, kan du kontakta Finlands Röda Kors De ungas skyddshus.
Skyddshuset finns i Alberga.
De ungas skyddshus
Tfn (09) 8195 5360
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Stöd- och serviceboende
En del människor, till exempel åldringar och handikappade, har svårt att klara av de dagliga sysslorna utan hjälp.
Personer som har sin hemkommun i Esbo kan få hemvårdens stödtjänster av Esbo stad, till exempel måltidstjänster eller färdtjänst.
Dessa tjänster hjälper människorna att klara sig bättre hemma.
Åldringar och handikappade som inte klarar av att bo självständigt, kan bo i ett servicehus eller på en vårdinrättning.
Läs mer: Stöd- och serviceboende
Om du har frågor kring stödtjänsterna för handikappade, kontakta handikappservicen vid Esbo stad.
Esbo stads handikappservice
Telefonrådgivning: (09) 816 45285
linkkiEsbo stad:
Stödtjänster för handikappadefinska _ svenska _ engelska
Om du har frågor kring stödtjänsterna för äldre, kontakta Esbo stads rådgivning för seniorer.
Esbo stads rådgivning för seniorer
tfn (09) 816 33333
linkkiEsbo stad:
Stödtjänster för äldrefinska _ svenska _ engelska
linkkiEsbo stad:
Information om hemvårdens stödtjänsterfinska _ svenska
linkkiEsbo stad:
Information om boende i servicehusfinska _ svenska
Bostadslöshet
Om du blir bostadslös, kontakta Esbo stads verksamhetsställe för vuxensocialarbete.
linkkiEsbo stad:
Kontaktuppgifter till vuxensocialarbetetfinska _ svenska _ engelska
Om läget är akut, kan du även kontakta social- och krisjouren i Esbo.
Social- och krisjouren
Jorvs sjukhus
Åbovägen 150
Tfn (09) 816 42439
linkkiEsbo stad:
Social- och krisjourenfinska _ svenska _ engelska
Läs mer: Bostadslöshet
Avfallshantering och återvinning
På InfoFinlands sida Avfallshantering och återvinning hittar du information om sopsortering.
linkkiHelsingforsregionens miljötjänster:
Sopsorteringsanvisningarfinska _ svenska _ engelska
linkkiHelsingforsregionens miljötjänster:
Återvinningsstationerfinska _ svenska _ engelska
Hyresbostad
Ägarbostad
Bostadsrättsbostad
Delägarbostad
Tillfälligt boende
Boende i en krissituation
Stöd- och serviceboende
Bostadslöshet
Avfallshantering och återvinning
Hyresbostad
I Esbo och huvudstadsregionen är hyrorna ofta högre än i resten av Finland.
Det kan vara svårt att hitta en bostad med lämplig hyra.
Det lönar sig att avsätta tid för bostadssökandet och undersöka olika alternativ.
Privata hyresbostäder
Hos en privat hyresvärd kan det gå snabbt att få en bostad, men hyran kan vara högre än i stadens hyresbostäder.
Du kan söka privata hyresbostäder i Esbo via hyresvärdarnas webbplatser:
Sökning av hyresbostäderfinska
Sökning av hyresbostäderfinska _ engelska
Hyresbostäder för ungafinska _ engelska
Hyresbostäder för ungafinska _ engelska
Om du är studerande kan du få en hyresbostad för studerande i Esbo.
Hyresbostäder för studerande erbjuds av Helsingforsregionens studentbostadsstiftelse HOAS och Aalto-universitets studentkår AUS.
linkkiHOAS:
Hyresbostäder för studerandefinska _ svenska _ engelska
Hyresbostäder för studerandefinska _ svenska _ engelska
Stadens hyresbostäder
Stadens hyresbostäder är ofta billigare än bostäder som man hyr av företag eller privatpersoner.
Det är dock många som ansöker om stadens bostäder och endast en liten del av de sökande får en bostad.
Störst är bristen på små bostäder.
Stadens hyresbostäder förvaltas av Espoon Asunnot Oy (Espoon Asunnot Oy).
Om du vill ansöka om en hyresbostad, fyll i en ansökningsblankett för hyresbostad på Espoon Asunnot Oy:s webbplats.
Du kan även fylla i ansökningsblanketten på Espoon Asunnot Oy:s kontor.
Du kan också få blanketten hemskickad per post.
Dina möjligheter att få en bostad påverkas av ditt bostadsbehov och dina tillgångar och inkomster.
För att kunna ansöka om en hyresbostad hos staden, måste du ha uppehållstillstånd för minst ett år.
Tfn (09) 816 5800
Ansökan är giltig i tre månader.
Efter det måste du förnya din ansökan om du fortfarande letar efter bostad.
Läs mer: Hyresbostad
linkkiEsbo Bostäder Ab:
Ansökan om hyresbostad i stadenfinska _ engelska
linkkiEsbo stad:
Stadens hyresbostäderfinska _ svenska _ engelska
linkkiEsbo stad:
Seniorbostäderfinska _ svenska
Ägarbostad
På internet finns många bostadsförsäljningsannonser.
Bostäderna i Esbo är tämligen dyra.
Information om köp av bostad hittar du på InfoFinlands sida Ägarbostad.
Bostadsrättsbostad
Om du ansöker om en bostadsrättsbostad, behöver du ett ordningsnummer. Du ansöker om ordningsnumret vid Esbo eller Helsingfors stad.
Läs mer: Bostadsrättsbostad.
linkkiEsbo stad:
Bostadsrättsbostäderfinska _ svenska _ engelska
Delägarbostad
Asuntosäätiö har delägarbostäder i Esbo.
Mer information hittar du på Asuntosäätiös webbplats.
Läs mer: Delägarbostad.
Delägarbostadfinska
Tillfälligt boende
I Esbo finns många olika hotell där man kan bo tillfälligt.
Läs mer: Tillfälligt boende.
linkkiVisitEspoo.fi:
Hotellfinska _ svenska _ engelska _ ryska
Brand eller vattenskada
Om din bostad har skadats till exempel till följd av brand eller vattenskada kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
Kontakta ditt försäkringsbolag direkt när skadan har inträffat.
Våld i hemmet
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta tjänsten Omatila (Omatila).
Omatila ordnar vid behov boende för dig och dina barn.
Omatila-tjänsten
Kamrersvägen 6 A
Tfn 043 825 0535
Öppet
Lördag-söndag kl. 9-16
Social- och krisjouren 24 h
Tfn 09 816 42439
linkkiEsbo stad:
Hjälp till offer för familjevåldfinska _ svenska _ engelska
Om du är ung och har problem hemma, kan du kontakta Finlands Röda Kors De ungas skyddshus.
Skyddshuset finns i Alberga.
De ungas skyddshus
Tfn (09) 8195 5360
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Stöd- och serviceboende
En del människor, till exempel åldringar och handikappade, har svårt att klara av de dagliga sysslorna utan hjälp.
Personer som har sin hemkommun i Esbo kan få hemvårdens stödtjänster av Esbo stad, till exempel måltidstjänster eller färdtjänst.
Dessa tjänster hjälper människorna att klara sig bättre hemma.
Åldringar och handikappade som inte klarar av att bo självständigt, kan bo i ett servicehus eller på en vårdinrättning.
Läs mer: Stöd- och serviceboende
Om du har frågor kring stödtjänsterna för handikappade, kontakta handikappservicen vid Esbo stad.
Esbo stads handikappservice
Telefonrådgivning: (09) 816 45285
linkkiEsbo stad:
Stödtjänster för handikappadefinska _ svenska _ engelska
Om du har frågor kring stödtjänsterna för äldre, kontakta Esbo stads rådgivning för seniorer.
Esbo stads rådgivning för seniorer
tfn (09) 816 33333
linkkiEsbo stad:
Stödtjänster för äldrefinska _ svenska _ engelska
linkkiEsbo stad:
Information om hemvårdens stödtjänsterfinska _ svenska
linkkiEsbo stad:
Information om boende i servicehusfinska _ svenska
Bostadslöshet
Om du blir bostadslös, kontakta Esbo stads verksamhetsställe för vuxensocialarbete.
linkkiEsbo stad:
Kontaktuppgifter till vuxensocialarbetetfinska _ svenska _ engelska
Om läget är akut, kan du även kontakta social- och krisjouren i Esbo.
Social- och krisjouren
Jorvs sjukhus
Åbovägen 150
Tfn (09) 816 42439
linkkiEsbo stad:
Social- och krisjourenfinska _ svenska _ engelska
Läs mer: Bostadslöshet
Avfallshantering och återvinning
På InfoFinlands sida Avfallshantering och återvinning hittar du information om sopsortering.
linkkiHelsingforsregionens miljötjänster:
Sopsorteringsanvisningarfinska _ svenska _ engelska
linkkiHelsingforsregionens miljötjänster:
Återvinningsstationerfinska _ svenska _ engelska
Hyresbostad
Ägarbostad
Bostadsrättsbostad
Delägarbostad
Tillfälligt boende
Boende i en krissituation
Stöd- och serviceboende
Bostadslöshet
Avfallshantering och återvinning
Hyresbostad
I Esbo och huvudstadsregionen är hyrorna ofta högre än i resten av Finland.
Det kan vara svårt att hitta en bostad med lämplig hyra.
Det lönar sig att avsätta tid för bostadssökandet och undersöka olika alternativ.
Privata hyresbostäder
Hos en privat hyresvärd kan det gå snabbt att få en bostad, men hyran kan vara högre än i stadens hyresbostäder.
Du kan söka privata hyresbostäder i Esbo via hyresvärdarnas webbplatser:
Sökning av hyresbostäderfinska
Sökning av hyresbostäderfinska _ engelska
Hyresbostäder för ungafinska _ engelska
Hyresbostäder för ungafinska _ engelska
Om du är studerande kan du få en hyresbostad för studerande i Esbo.
Hyresbostäder för studerande erbjuds av Helsingforsregionens studentbostadsstiftelse HOAS och Aalto-universitets studentkår AUS.
linkkiHOAS:
Hyresbostäder för studerandefinska _ svenska _ engelska
Hyresbostäder för studerandefinska _ svenska _ engelska
Stadens hyresbostäder
Stadens hyresbostäder är ofta billigare än bostäder som man hyr av företag eller privatpersoner.
Det är dock många som ansöker om stadens bostäder och endast en liten del av de sökande får en bostad.
Störst är bristen på små bostäder.
Stadens hyresbostäder förvaltas av Espoon Asunnot Oy (Espoon Asunnot Oy).
Om du vill ansöka om en hyresbostad, fyll i en ansökningsblankett för hyresbostad på Espoon Asunnot Oy:s webbplats.
Du kan även fylla i ansökningsblanketten på Espoon Asunnot Oy:s kontor.
Du kan också få blanketten hemskickad per post.
Dina möjligheter att få en bostad påverkas av ditt bostadsbehov och dina tillgångar och inkomster.
För att kunna ansöka om en hyresbostad hos staden, måste du ha uppehållstillstånd för minst ett år.
Tfn (09) 816 5800
Ansökan är giltig i tre månader.
Efter det måste du förnya din ansökan om du fortfarande letar efter bostad.
Läs mer: Hyresbostad
linkkiEsbo Bostäder Ab:
Ansökan om hyresbostad i stadenfinska _ engelska
linkkiEsbo stad:
Stadens hyresbostäderfinska _ svenska _ engelska
linkkiEsbo stad:
Seniorbostäderfinska _ svenska
Ägarbostad
På internet finns många bostadsförsäljningsannonser.
Bostäderna i Esbo är tämligen dyra.
Information om köp av bostad hittar du på InfoFinlands sida Ägarbostad.
Bostadsrättsbostad
Om du ansöker om en bostadsrättsbostad, behöver du ett ordningsnummer. Du ansöker om ordningsnumret vid Esbo eller Helsingfors stad.
Läs mer: Bostadsrättsbostad.
linkkiEsbo stad:
Bostadsrättsbostäderfinska _ svenska _ engelska
Delägarbostad
Asuntosäätiö har delägarbostäder i Esbo.
Mer information hittar du på Asuntosäätiös webbplats.
Läs mer: Delägarbostad.
Delägarbostadfinska
Tillfälligt boende
I Esbo finns många olika hotell där man kan bo tillfälligt.
Läs mer: Tillfälligt boende.
linkkiVisitEspoo.fi:
Hotellfinska _ svenska _ engelska _ ryska
Brand eller vattenskada
Om din bostad har skadats till exempel till följd av brand eller vattenskada kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
Kontakta ditt försäkringsbolag direkt när skadan har inträffat.
Våld i hemmet
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta tjänsten Omatila (Omatila).
Omatila ordnar vid behov boende för dig och dina barn.
Omatila-tjänsten
Kamrersvägen 6 A
Tfn 043 825 0535
Öppet
Lördag-söndag kl. 9-16
Social- och krisjouren 24 h
Tfn 09 816 42439
linkkiEsbo stad:
Hjälp till offer för familjevåldfinska _ svenska _ engelska
Om du är ung och har problem hemma, kan du kontakta Finlands Röda Kors De ungas skyddshus.
Skyddshuset finns i Alberga.
De ungas skyddshus
Tfn (09) 8195 5360
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Stöd- och serviceboende
En del människor, till exempel åldringar och handikappade, har svårt att klara av de dagliga sysslorna utan hjälp.
Personer som har sin hemkommun i Esbo kan få hemvårdens stödtjänster av Esbo stad, till exempel måltidstjänster eller färdtjänst.
Dessa tjänster hjälper människorna att klara sig bättre hemma.
Åldringar och handikappade som inte klarar av att bo självständigt, kan bo i ett servicehus eller på en vårdinrättning.
Läs mer: Stöd- och serviceboende
Om du har frågor kring stödtjänsterna för handikappade, kontakta handikappservicen vid Esbo stad.
Esbo stads handikappservice
Telefonrådgivning: (09) 816 45285
linkkiEsbo stad:
Stödtjänster för handikappadefinska _ svenska _ engelska
Om du har frågor kring stödtjänsterna för äldre, kontakta Esbo stads rådgivning för seniorer.
Esbo stads rådgivning för seniorer
tfn (09) 816 33333
linkkiEsbo stad:
Stödtjänster för äldrefinska _ svenska _ engelska
linkkiEsbo stad:
Information om hemvårdens stödtjänsterfinska _ svenska
linkkiEsbo stad:
Information om boende i servicehusfinska _ svenska
Bostadslöshet
Om du blir bostadslös, kontakta Esbo stads verksamhetsställe för vuxensocialarbete.
linkkiEsbo stad:
Kontaktuppgifter till vuxensocialarbetetfinska _ svenska _ engelska
Om läget är akut, kan du även kontakta social- och krisjouren i Esbo.
Social- och krisjouren
Jorvs sjukhus
Åbovägen 150
Tfn (09) 816 42439
linkkiEsbo stad:
Social- och krisjourenfinska _ svenska _ engelska
Läs mer: Bostadslöshet
Avfallshantering och återvinning
På InfoFinlands sida Avfallshantering och återvinning hittar du information om sopsortering.
linkkiHelsingforsregionens miljötjänster:
Sopsorteringsanvisningarfinska _ svenska _ engelska
linkkiHelsingforsregionens miljötjänster:
Återvinningsstationerfinska _ svenska _ engelska
Språkkurser
Med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors, Vanda, Esbo eller Grankulla.
I Esbo ordnas språkkurser i finska och svenska av Esbo arbetarinstitut, Esbo vuxengymnasium, Luksia och Axxell.
Kurser i finska och svenska språketfinska _ engelska _ ryska
Samtala på finska
På biblioteken i Esbo ordnas språkkaféer, där man kan öva sig i att prata finska.
På språkkaféerna samtalar man på finska, så det är bra om du redan kan lite finska.
Språkkaféerna är avgiftsfria.
Språkkaféer:
Entresse bibliotek, Iso Omena bibliotek, Stensvik bibliotek, Sello bibliotek och Hagalunds bibliotek.
Språkkaféerfinska _ engelska _ ryska
På den internationella träffpunkten Trapesa kan du delta i en samtals- och inlärningsgrupp på finska.
Gruppen är öppen för alla och den är avgiftsfri.
Diskussionsgrupp på finskafinska
Vi läser tillsammans för kvinnor
I Esbo finns även Vi läser tillsammans-grupper, där kvinnor kan studera finska språket.
linkkiVi läser tillsammans:
Finska för kvinnorfinska
Invånarlokalen i Kivenkolo
Man kan även träna sina finskakunskaper i invånarlokalen i Kivenkolo.
linkkiEsbo stad:
Kivenkolo invånarhusfinska _ svenska _ engelska
Om du är kund vid arbets- och näringsbyrån kan du fråga om språkkurser i finska och svenska vid arbets- och näringsbyrån.
Läs mer: Studier i finska och svenska
linkkiEsbo stad:
Kurser i finska och svenska språketfinska _ svenska _ engelska
linkkiEsbo stad:
Arbetarinstitutetfinska _ svenska _ engelska
linkkiEsbo stad:
Vuxengymnasietfinska
Kurser i finska och svenska språketfinska _ engelska
linkkiAxxell:
Kurser i finska och svenska språketfinska _ svenska
Allmän språkexamen
Du kan avlägga allmän språkexamen (yleinen kielitutkinto) i finska eller svenska i Esbo.
I Esbo ordnas språkexamina av Axxell och Esbo arbetarinstitut.
På utbildningsstyrelsens (opetushallitus) webbplats finns en sökmotor för språkexamina.
Med sökmotorn kan du kontrollera var och när du kan avlägga examen.
linkkiUtbildningsstyrelsen:
Examenssökningfinska
linkkiUtbildningsstyrelsen:
Allmänna språkexaminafinska _ svenska _ engelska
Språkkurser
Med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors, Vanda, Esbo eller Grankulla.
I Esbo ordnas språkkurser i finska och svenska av Esbo arbetarinstitut, Esbo vuxengymnasium, Luksia och Axxell.
Kurser i finska och svenska språketfinska _ engelska _ ryska
Samtala på finska
På biblioteken i Esbo ordnas språkkaféer, där man kan öva sig i att prata finska.
På språkkaféerna samtalar man på finska, så det är bra om du redan kan lite finska.
Språkkaféerna är avgiftsfria.
Språkkaféer:
Entresse bibliotek, Iso Omena bibliotek, Stensvik bibliotek, Sello bibliotek och Hagalunds bibliotek.
Språkkaféerfinska _ engelska _ ryska
På den internationella träffpunkten Trapesa kan du delta i en samtals- och inlärningsgrupp på finska.
Gruppen är öppen för alla och den är avgiftsfri.
Diskussionsgrupp på finskafinska
Vi läser tillsammans för kvinnor
I Esbo finns även Vi läser tillsammans-grupper, där kvinnor kan studera finska språket.
linkkiVi läser tillsammans:
Finska för kvinnorfinska
Invånarlokalen i Kivenkolo
Man kan även träna sina finskakunskaper i invånarlokalen i Kivenkolo.
linkkiEsbo stad:
Kivenkolo invånarhusfinska _ svenska _ engelska
Om du är kund vid arbets- och näringsbyrån kan du fråga om språkkurser i finska och svenska vid arbets- och näringsbyrån.
Läs mer: Studier i finska och svenska
linkkiEsbo stad:
Kurser i finska och svenska språketfinska _ svenska _ engelska
linkkiEsbo stad:
Arbetarinstitutetfinska _ svenska _ engelska
linkkiEsbo stad:
Vuxengymnasietfinska
Kurser i finska och svenska språketfinska _ engelska
linkkiAxxell:
Kurser i finska och svenska språketfinska _ svenska
Allmän språkexamen
Du kan avlägga allmän språkexamen (yleinen kielitutkinto) i finska eller svenska i Esbo.
I Esbo ordnas språkexamina av Axxell och Esbo arbetarinstitut.
På utbildningsstyrelsens (opetushallitus) webbplats finns en sökmotor för språkexamina.
Med sökmotorn kan du kontrollera var och när du kan avlägga examen.
linkkiUtbildningsstyrelsen:
Examenssökningfinska
linkkiUtbildningsstyrelsen:
Allmänna språkexaminafinska _ svenska _ engelska
Språkkurser
Med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors, Vanda, Esbo eller Grankulla.
I Esbo ordnas språkkurser i finska och svenska av Esbo arbetarinstitut, Esbo vuxengymnasium, Luksia och Axxell.
Kurser i finska och svenska språketfinska _ engelska _ ryska
Samtala på finska
På biblioteken i Esbo ordnas språkkaféer, där man kan öva sig i att prata finska.
På språkkaféerna samtalar man på finska, så det är bra om du redan kan lite finska.
Språkkaféerna är avgiftsfria.
Språkkaféer:
Entresse bibliotek, Iso Omena bibliotek, Stensvik bibliotek, Sello bibliotek och Hagalunds bibliotek.
Språkkaféerfinska _ engelska _ ryska
På den internationella träffpunkten Trapesa kan du delta i en samtals- och inlärningsgrupp på finska.
Gruppen är öppen för alla och den är avgiftsfri.
Diskussionsgrupp på finskafinska
Vi läser tillsammans för kvinnor
I Esbo finns även Vi läser tillsammans-grupper, där kvinnor kan studera finska språket.
linkkiVi läser tillsammans:
Finska för kvinnorfinska
Invånarlokalen i Kivenkolo
Man kan även träna sina finskakunskaper i invånarlokalen i Kivenkolo.
linkkiEsbo stad:
Kivenkolo invånarhusfinska _ svenska _ engelska
Om du är kund vid arbets- och näringsbyrån kan du fråga om språkkurser i finska och svenska vid arbets- och näringsbyrån.
Läs mer: Studier i finska och svenska
linkkiEsbo stad:
Kurser i finska och svenska språketfinska _ svenska _ engelska
linkkiEsbo stad:
Arbetarinstitutetfinska _ svenska _ engelska
linkkiEsbo stad:
Vuxengymnasietfinska
Kurser i finska och svenska språketfinska _ engelska
linkkiAxxell:
Kurser i finska och svenska språketfinska _ svenska
Allmän språkexamen
Du kan avlägga allmän språkexamen (yleinen kielitutkinto) i finska eller svenska i Esbo.
I Esbo ordnas språkexamina av Axxell och Esbo arbetarinstitut.
På utbildningsstyrelsens (opetushallitus) webbplats finns en sökmotor för språkexamina.
Med sökmotorn kan du kontrollera var och när du kan avlägga examen.
linkkiUtbildningsstyrelsen:
Examenssökningfinska
linkkiUtbildningsstyrelsen:
Allmänna språkexaminafinska _ svenska _ engelska
Var hittar jag jobb?
Hjälp med jobbsökningen
Att grunda ett företag
Beskattning
Var hittar jag jobb?
TE-byråns tjänster
Du kan få hjälp med jobbsökningen vid Nylands TE-byrå.
Verksamhetsstället i Esbo finns i Alberga.
linkkiArbets- och näringsministeriet:
Arbets- och näringsbyråerna i Nylandfinska _ svenska
TE-byrån betjänar på internet via sidan E-tjänster (Oma asiointi).
För att använda tjänsten behöver du nätbankskoder.
Medborgare i EU-länderna, Norge, Island, Liechtenstein och Schweiz kan anmäla sig som arbetssökande via TE-byråns E-tjänster.
Medborgare i andra länder måste anmäla sig personligen vid TE-byrån.
Ta med ett ID-kort och ditt uppehållstillstånd.
Information om TE-byråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös.
Information om jobbsökning i Finland hittar du på InfoFinlands sida Var hittar jag jobb?
linkkiTE-tjänster:
Anmälan utan nätbankskoderfinska _ svenska
linkkiArbets- och näringsministeriet:
Lediga jobbfinska _ svenska
linkkiArbets- och näringsförvaltningen:
Länkar till jobbsajterfinska _ svenska _ engelska
Lediga tjänster vid Esbo stad hittar du på stadens webbplats.
linkkiEsbo stad:
Arbetsplatser vid stadenfinska _ svenska _ engelska
Seure (Seure) är ett bemanningsbolag som erbjuder kortvariga jobb vid Helsingfors, Vanda, Esbo och Grankulla städer.
Jobben finns till exempel på skolor, daghem och sjukhus.
Arbetsplatser i kommunernafinska _ svenska
Hjälp med jobbsökningen
Råd om jobbsökningfinska _ svenska _ engelska _ spanska
Mentorskap i fråga om arbetskarriärfinska _ engelska
För unga under 30 år
linkkiEsbo stad:
Ohjaamofinska _ svenska _ engelska
Arbetslöshetsersättning
Information om att ansöka om arbetslöshetsersättning hittar du på InfoFinlands sida Arbetslöshetsförsäkring.
Att grunda ett företag
Om du vill grunda ett eget företag, kan du få hjälp vid FöretagsEsbo.
De hjälper dig att utveckla affärsidén och planera affärsverksamheten.
Tjänsterna är kostnadsfria.
linkkiFöretagsEsbo:
Företagsrådgivningfinska _ svenska _ engelska
Tjänster för företagarefinska _ svenska _ engelska
NewCo Yritys Helsinki erbjuder individuell rådgivning om grundande av företag samt ordnar informationsmöten och företagarutbildning på flera olika språk.
Tjänster för företagare med invandrarbakgrundfinska _ engelska
Guide om att grunda ett företagfinska _ engelska _ kinesiska
linkkiArbets- och näringsministeriet:
Tjänster för företagarefinska _ svenska _ engelska
Företagare i Esbo får även hjälp av Företagarna i Esbo rf.
Företagarna i Esbo rf är företagarnas egen organisation som erbjuder sina medlemmar till exempel utbildning, samarbete och rådgivning.
linkkiEsbo Företagare:
Företagarnas intressebevakningsorganisationfinska
Läs mer: Att grunda ett företag
Beskattning
Huvudstadsregionens skattebyrå ligger på Alexandersgatan 9 i Gloet i Helsingfors.
linkkiSkatteförvaltningen:
Kontaktuppgifter till skattebyråerfinska _ svenska _ engelska
Du kan även besöka servicestället In To Finland i Kampen i Helsingfors.
FPA:s och Skatteförvaltningens gemensamma rådgivning hjälper invandrare som har frågor om beskattningen eller den sociala tryggheten.
Här kan du hämta ett skattekort och ett inom byggbranschen obligatoriskt skattenummer.
Här kan dessutom utländska arbetstagare som ska arbeta i Finland tillfälligt få en finsk personbeteckning utan ett separat besök till magistraten.
Albertsgatan 25
Information om beskattningen hittar du på InfoFinlands sida Beskattning.
Var hittar jag jobb?
Hjälp med jobbsökningen
Att grunda ett företag
Beskattning
Var hittar jag jobb?
TE-byråns tjänster
Du kan få hjälp med jobbsökningen vid Nylands TE-byrå.
Verksamhetsstället i Esbo finns i Alberga.
linkkiArbets- och näringsministeriet:
Arbets- och näringsbyråerna i Nylandfinska _ svenska
TE-byrån betjänar på internet via sidan E-tjänster (Oma asiointi).
För att använda tjänsten behöver du nätbankskoder.
Medborgare i EU-länderna, Norge, Island, Liechtenstein och Schweiz kan anmäla sig som arbetssökande via TE-byråns E-tjänster.
Medborgare i andra länder måste anmäla sig personligen vid TE-byrån.
Ta med ett ID-kort och ditt uppehållstillstånd.
Information om TE-byråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös.
Information om jobbsökning i Finland hittar du på InfoFinlands sida Var hittar jag jobb?
linkkiTE-tjänster:
Anmälan utan nätbankskoderfinska _ svenska
linkkiArbets- och näringsministeriet:
Lediga jobbfinska _ svenska
linkkiArbets- och näringsförvaltningen:
Länkar till jobbsajterfinska _ svenska _ engelska
Lediga tjänster vid Esbo stad hittar du på stadens webbplats.
linkkiEsbo stad:
Arbetsplatser vid stadenfinska _ svenska _ engelska
Seure (Seure) är ett bemanningsbolag som erbjuder kortvariga jobb vid Helsingfors, Vanda, Esbo och Grankulla städer.
Jobben finns till exempel på skolor, daghem och sjukhus.
Arbetsplatser i kommunernafinska _ svenska
Hjälp med jobbsökningen
Råd om jobbsökningfinska _ svenska _ engelska _ spanska
Mentorskap i fråga om arbetskarriärfinska _ engelska
För unga under 30 år
linkkiEsbo stad:
Ohjaamofinska _ svenska _ engelska
Arbetslöshetsersättning
Information om att ansöka om arbetslöshetsersättning hittar du på InfoFinlands sida Arbetslöshetsförsäkring.
Att grunda ett företag
Om du vill grunda ett eget företag, kan du få hjälp vid FöretagsEsbo.
De hjälper dig att utveckla affärsidén och planera affärsverksamheten.
Tjänsterna är kostnadsfria.
linkkiFöretagsEsbo:
Företagsrådgivningfinska _ svenska _ engelska
Tjänster för företagarefinska _ svenska _ engelska
NewCo Yritys Helsinki erbjuder individuell rådgivning om grundande av företag samt ordnar informationsmöten och företagarutbildning på flera olika språk.
Tjänster för företagare med invandrarbakgrundfinska _ engelska
Guide om att grunda ett företagfinska _ engelska _ kinesiska
linkkiArbets- och näringsministeriet:
Tjänster för företagarefinska _ svenska _ engelska
Företagare i Esbo får även hjälp av Företagarna i Esbo rf.
Företagarna i Esbo rf är företagarnas egen organisation som erbjuder sina medlemmar till exempel utbildning, samarbete och rådgivning.
linkkiEsbo Företagare:
Företagarnas intressebevakningsorganisationfinska
Läs mer: Att grunda ett företag
Beskattning
Huvudstadsregionens skattebyrå ligger på Alexandersgatan 9 i Gloet i Helsingfors.
linkkiSkatteförvaltningen:
Kontaktuppgifter till skattebyråerfinska _ svenska _ engelska
Invandrare kan även sköta ärenden vid servicestället International House Helsinki.
På servicestället hjälper FPA:s och Skatteförvaltningens experter invandrare som kommer till Finland för att arbeta i frågor som rör beskattning och social trygghet.
Information om beskattningen hittar du på InfoFinlands sida Beskattning.
Var hittar jag jobb?
Hjälp med jobbsökningen
Att grunda ett företag
Beskattning
Var hittar jag jobb?
TE-byråns tjänster
Du kan få hjälp med jobbsökningen vid Nylands TE-byrå.
Verksamhetsstället i Esbo finns i Alberga.
linkkiArbets- och näringsministeriet:
Arbets- och näringsbyråerna i Nylandfinska _ svenska
TE-byrån betjänar på internet via sidan E-tjänster (Oma asiointi).
För att använda tjänsten behöver du nätbankskoder.
Medborgare i EU-länderna, Norge, Island, Liechtenstein och Schweiz kan anmäla sig som arbetssökande via TE-byråns E-tjänster.
Medborgare i andra länder måste anmäla sig personligen vid TE-byrån.
Ta med ett ID-kort och ditt uppehållstillstånd.
Information om TE-byråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös.
Information om jobbsökning i Finland hittar du på InfoFinlands sida Var hittar jag jobb?
linkkiTE-tjänster:
Anmälan utan nätbankskoderfinska _ svenska
linkkiArbets- och näringsministeriet:
Lediga jobbfinska _ svenska
linkkiArbets- och näringsförvaltningen:
Länkar till jobbsajterfinska _ svenska _ engelska
Lediga tjänster vid Esbo stad hittar du på stadens webbplats.
linkkiEsbo stad:
Arbetsplatser vid stadenfinska _ svenska _ engelska
Seure (Seure) är ett bemanningsbolag som erbjuder kortvariga jobb vid Helsingfors, Vanda, Esbo och Grankulla städer.
Jobben finns till exempel på skolor, daghem och sjukhus.
Arbetsplatser i kommunernafinska _ svenska _ engelska
Hjälp med jobbsökningen
Råd om jobbsökningfinska _ svenska _ engelska _ spanska
Mentorskap i fråga om arbetskarriärfinska _ engelska
För unga under 30 år
linkkiEsbo stad:
Ohjaamofinska _ svenska _ engelska
Arbetslöshetsersättning
Information om att ansöka om arbetslöshetsersättning hittar du på InfoFinlands sida Arbetslöshetsförsäkring.
Att grunda ett företag
Om du vill grunda ett eget företag, kan du få hjälp vid FöretagsEsbo.
De hjälper dig att utveckla affärsidén och planera affärsverksamheten.
Tjänsterna är kostnadsfria.
linkkiFöretagsEsbo:
Företagsrådgivningfinska _ svenska _ engelska
Tjänster för företagarefinska _ svenska _ engelska
NewCo Yritys Helsinki erbjuder individuell rådgivning om grundande av företag samt ordnar informationsmöten och företagarutbildning på flera olika språk.
Tjänster för företagare med invandrarbakgrundfinska _ engelska
Guide om att grunda ett företagfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ turkiska _ kinesiska _ arabiska
linkkiArbets- och näringsministeriet:
Tjänster för företagarefinska _ svenska _ engelska
Företagare i Esbo får även hjälp av Företagarna i Esbo rf.
Företagarna i Esbo rf är företagarnas egen organisation som erbjuder sina medlemmar till exempel utbildning, samarbete och rådgivning.
linkkiEsbo Företagare:
Företagarnas intressebevakningsorganisationfinska
Läs mer: Att grunda ett företag
Beskattning
Huvudstadsregionens skattebyrå ligger på Alexandersgatan 9 i Gloet i Helsingfors.
linkkiSkatteförvaltningen:
Kontaktuppgifter till skattebyråerfinska _ svenska _ engelska
Invandrare kan även sköta ärenden vid servicestället International House Helsinki.
På servicestället hjälper FPA:s och Skatteförvaltningens experter invandrare som kommer till Finland för att arbeta i frågor som rör beskattning och social trygghet.
Information om beskattningen hittar du på InfoFinlands sida Beskattning.
Rådgivning för och integration av invandrare
Inledande kartläggning och integrationsplan
Behöver du en tolk?
Rådgivning för och integration av invandrare
Servicepunkt
Vid Esbo stads servicepunkter (asiointipiste) får du mer information om stadens tjänster.
Servicepunkter finns på olika håll i staden.
Närmare kontaktuppgifter finns på Esbo stads webbplats.
Det gemensamma telefonnumret till servicepunkterna är (09) 816 57070 och e-postadressen är info(at)espoo.fi.
linkkiEsbo stad:
Servicepunktfinska _ svenska _ engelska
Kivenkolo
Invånarhuset Kivenkolo är ett öppet vardagsum där du kan få rådgivning och handledning på olika språk.
Kivenkolo
Sjöstöveln 1 A
Tfn 050 300 6093
linkkiEsbo stad:
Kivenkolo invånarhusfinska _ svenska _ engelska
Startpunkt för unga vuxna
Navigatorns Startpunkter erbjuder handledning och rådgivning utan tidsbokning till unga under 30 år.
Fågelbergavägen 2 A
Startpunkten i Iso Omena
linkkiEsbo stad:
Rådgivning för ungafinska _ svenska _ engelska
Den internationella mötesplatsen Trapesa erbjuder rådgivningstjänster.
Boka en tid i förväg.
Föreningen har även ett öppet vardagsrum, samtalsgrupper på finska och olika slags evenemang.
Stationsbron i Esbo
Tfn 010 583 7971
Invandrartjänster
Flyktingar kan även kontakta Esbo stads invandrartjänster (Maahanmuuttajapalvelut).
Vid servicerådgivningen får du råd och handledning utan tidsbeställning.
Rådgivningen ges på många olika språk.
Invandrartjänsterna
Fångstvägen 3
Tfn (09) 81621
linkkiEsbo stad:
Invandrartjänsterfinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
Du kan få:
kostnadsfri rådgivning och information kring att flytta på flera olika språk
en finländsk personbeteckning, registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1-intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
I tjänsten medverkar Helsingfors-info, magistraten i Nyland, skatteförvaltningens och FPA:s tjänst In To Finland, NTM-centralen i Nyland, Pensionsskyddscentralen och Helsingforsregionens handelskammare.
Adress
Albertsgatan 25
IHH – serviceställe för dig som flyttar till Finland engelska
Inledande kartläggning och integrationsplan
Inledande kartläggningar görs vid Esbo stads invandrartjänster eller enheten för vuxensocialarbete.
Invandrartjänsterna hjälper invandrare även i frågor som rör livet i Finland.
linkkiEsbo stad:
Invandrartjänsterfinska _ svenska _ engelska
linkkiEsbo stad:
Kontaktuppgifter till vuxensocialarbetetfinska _ svenska _ engelska
En anställd vid arbets- och näringsbyrån gör en inledande kartläggning tillsammans med dig, när du registrerar dig som arbetssökande.
Byrån i Esbo finns i Alberga.
Arbets- och näringsbyrån i Esbo
linkkiArbets- och näringsministeriet:
Arbets- och näringsbyråerna i Nylandfinska _ svenska
Behöver du en tolk?
Om du inte kan finska eller svenska kan du anlita en tolk när du sköter ärenden med myndigheter.
I vissa fall får du tolken via myndigheten.
Då är tolkningen kostnadsfri för dig.
Med myndigheter avses till exempel polisen, FPA, arbets- och näringsbyrån eller tjänstemän vid Esbo stad.
Myndigheten betalar dock inte alltid för en tolk.
Du ska alltså på förhand fråga om myndigheten betalar för tolktjänsterna.
Du kan använda en tolk när du vill, ifall du betalar och beställer tolken själv.
Du kan fråga om tolktjänsterna närmare till exempel vid Esbo stads invandrartjänster.
Läs mer: Behöver du en tolk?
linkkiEsbo stad:
Invandrartjänsterfinska _ svenska _ engelska
linkkiFinlands översättar- och tolkförbund:
Sök tolk eller översättarefinska _ svenska _ engelska
Rådgivning för och integration av invandrare
Inledande kartläggning och integrationsplan
Behöver du en tolk?
Rådgivning för och integration av invandrare
Servicepunkt
Vid Esbo stads servicepunkter (asiointipiste) får du mer information om stadens tjänster.
Servicepunkter finns på olika håll i staden.
Närmare kontaktuppgifter finns på Esbo stads webbplats.
Det gemensamma telefonnumret till servicepunkterna är (09) 816 57070 och e-postadressen är info(at)espoo.fi.
linkkiEsbo stad:
Servicepunktfinska _ svenska _ engelska
Kivenkolo
Invånarhuset Kivenkolo är ett öppet vardagsum där du kan få rådgivning och handledning på olika språk.
Kivenkolo
Sjöstöveln 1 A
Tfn 050 300 6093
linkkiEsbo stad:
Kivenkolo invånarhusfinska _ svenska _ engelska
Startpunkt för unga vuxna
Navigatorns Startpunkter erbjuder handledning och rådgivning utan tidsbokning till unga under 30 år.
Fågelbergavägen 2 A
Startpunkten i Iso Omena
linkkiEsbo stad:
Rådgivning för ungafinska _ svenska _ engelska
Den internationella mötesplatsen Trapesa erbjuder rådgivningstjänster.
Boka en tid i förväg.
Föreningen har även ett öppet vardagsrum, samtalsgrupper på finska och olika slags evenemang.
Stationsbron i Esbo
Tfn 010 583 7971
Invandrartjänster
Flyktingar kan även kontakta Esbo stads invandrartjänster (Maahanmuuttajapalvelut).
Vid servicerådgivningen får du råd och handledning utan tidsbeställning.
Rådgivningen ges på många olika språk.
Invandrartjänsterna
Fångstvägen 3
Tfn (09) 81621
linkkiEsbo stad:
Invandrartjänsterfinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
Du kan få:
kostnadsfri rådgivning och information kring att flytta på flera olika språk
en finländsk personbeteckning, registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1-intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
I tjänsten medverkar Helsingfors-info, magistraten i Nyland, skatteförvaltningens och FPA:s tjänst In To Finland, NTM-centralen i Nyland, Pensionsskyddscentralen och Helsingforsregionens handelskammare.
Adress
IHH – serviceställe för dig som flyttar till Finland engelska
Inledande kartläggning och integrationsplan
Inledande kartläggningar görs vid Esbo stads invandrartjänster eller enheten för vuxensocialarbete.
Invandrartjänsterna hjälper invandrare även i frågor som rör livet i Finland.
linkkiEsbo stad:
Invandrartjänsterfinska _ svenska _ engelska
linkkiEsbo stad:
Kontaktuppgifter till vuxensocialarbetetfinska _ svenska _ engelska
En anställd vid arbets- och näringsbyrån gör en inledande kartläggning tillsammans med dig, när du registrerar dig som arbetssökande.
Byrån i Esbo finns i Alberga.
Arbets- och näringsbyrån i Esbo
linkkiArbets- och näringsministeriet:
Arbets- och näringsbyråerna i Nylandfinska _ svenska
Behöver du en tolk?
Om du inte kan finska eller svenska kan du anlita en tolk när du sköter ärenden med myndigheter.
I vissa fall får du tolken via myndigheten.
Då är tolkningen kostnadsfri för dig.
Med myndigheter avses till exempel polisen, FPA, arbets- och näringsbyrån eller tjänstemän vid Esbo stad.
Myndigheten betalar dock inte alltid för en tolk.
Du ska alltså på förhand fråga om myndigheten betalar för tolktjänsterna.
Du kan använda en tolk när du vill, ifall du betalar och beställer tolken själv.
Du kan fråga om tolktjänsterna närmare till exempel vid Esbo stads invandrartjänster.
Läs mer: Behöver du en tolk?
linkkiEsbo stad:
Invandrartjänsterfinska _ svenska _ engelska
linkkiFinlands översättar- och tolkförbund:
Sök tolk eller översättarefinska _ svenska _ engelska
Rådgivning för och integration av invandrare
Inledande kartläggning och integrationsplan
Behöver du en tolk?
Rådgivning för och integration av invandrare
Servicepunkt
Vid Esbo stads servicepunkter (asiointipiste) får du mer information om stadens tjänster.
Servicepunkter finns på olika håll i staden.
Närmare kontaktuppgifter finns på Esbo stads webbplats.
Det gemensamma telefonnumret till servicepunkterna är (09) 816 57070 och e-postadressen är info(at)espoo.fi.
linkkiEsbo stad:
Servicepunktfinska _ svenska _ engelska
Kivenkolo
Invånarhuset Kivenkolo är ett öppet vardagsum där du kan få rådgivning och handledning på olika språk.
Kivenkolo
Sjöstöveln 1 A
Tfn 050 300 6093
linkkiEsbo stad:
Kivenkolo invånarhusfinska _ svenska _ engelska
Startpunkt för unga vuxna
Navigatorns Startpunkter erbjuder handledning och rådgivning utan tidsbokning till unga under 30 år.
Fågelbergavägen 2 A
Startpunkten i Iso Omena
linkkiEsbo stad:
Rådgivning för ungafinska _ svenska _ engelska
Den internationella mötesplatsen Trapesa erbjuder rådgivningstjänster.
Boka en tid i förväg.
Föreningen har även ett öppet vardagsrum, samtalsgrupper på finska och olika slags evenemang.
Stationsbron i Esbo
Tfn 010 583 7971
Invandrartjänster
Flyktingar kan även kontakta Esbo stads invandrartjänster (Maahanmuuttajapalvelut).
Vid servicerådgivningen får du råd och handledning utan tidsbeställning.
Rådgivningen ges på många olika språk.
Invandrartjänsterna
Fångstvägen 3
Tfn (09) 81621
linkkiEsbo stad:
Invandrartjänsterfinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
Du kan få:
kostnadsfri rådgivning och information kring att flytta på flera olika språk
en finländsk personbeteckning, registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1-intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
I tjänsten medverkar Helsingfors-info, Esbo stad, magistraten i Nyland, Migrationsverket, Skatteförvaltningen, FPA, NTM-centralen i Nyland, Pensionsskyddscentralen, Helsingforsregionens handelskammare och Finlands Fackförbunds Centralorganisation FFC.
Adress
IHH – serviceställe för dig som flyttar till Finland engelska
Inledande kartläggning och integrationsplan
Inledande kartläggningar görs vid Esbo stads invandrartjänster eller enheten för vuxensocialarbete.
Invandrartjänsterna hjälper invandrare även i frågor som rör livet i Finland.
linkkiEsbo stad:
Invandrartjänsterfinska _ svenska _ engelska
linkkiEsbo stad:
Kontaktuppgifter till vuxensocialarbetetfinska _ svenska _ engelska
En anställd vid arbets- och näringsbyrån gör en inledande kartläggning tillsammans med dig, när du registrerar dig som arbetssökande.
Byrån i Esbo finns i Alberga.
Arbets- och näringsbyrån i Esbo
linkkiArbets- och näringsministeriet:
Arbets- och näringsbyråerna i Nylandfinska _ svenska
Behöver du en tolk?
Om du inte kan finska eller svenska kan du anlita en tolk när du sköter ärenden med myndigheter.
I vissa fall får du tolken via myndigheten.
Då är tolkningen kostnadsfri för dig.
Med myndigheter avses till exempel polisen, FPA, arbets- och näringsbyrån eller tjänstemän vid Esbo stad.
Myndigheten betalar dock inte alltid för en tolk.
Du ska alltså på förhand fråga om myndigheten betalar för tolktjänsterna.
Du kan använda en tolk när du vill, ifall du betalar och beställer tolken själv.
Du kan fråga om tolktjänsterna närmare till exempel vid Esbo stads invandrartjänster.
Läs mer: Behöver du en tolk?
linkkiEsbo stad:
Invandrartjänsterfinska _ svenska _ engelska
linkkiFinlands översättar- och tolkförbund:
Sök tolk eller översättarefinska _ svenska _ engelska
Tillståndsärenden
På Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU-medborgarens uppehållsrätt.
Migrationsverkets tjänsteställe i Helsingfors :
Göksgränd 3A
Du kan också ansöka om många slags uppehållstillstånd och EU-registrering på internet i tjänsten Enter Finland.
Om du inte är van vid att använda en dator, fyll i en ansökan på papper och lämna in den på Migrationsverkets tjänsteställe.
Dät är alltid bra att boka en tid i förväg på tjänstestället.
Du kan boka en tid på Migrationsverkets tidsbokningstjänst.
Observera att tjänstestället inte kan ge rådgivning om tillståndsärenden.
Läs mer: Flytta till Finland.
Elektronisk tidsbokningfinska _ svenska _ engelska
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Registrering som invånare
Om du flyttar ditt stadigvarande boende till Esbo, ska du registrera dig som invånare i kommunen.
Du kan registrera dig vid magistraten i Nyland, Helsingfors enhet.
Magistraten i Nyland Helsingfors enhet
Albertsgatan 25
Tfn 029 55 39391
När du går till magistraten ska du ta med dig
legitimation (till exempel pass)
uppehållstillstånd och uppehållskort (om du behöver uppehållstillstånd i Finland)
registreringsintyget över uppehållsrätten (oleskeluoikeuden rekisteröintitodistus) om du är EU-medborgare.
äktenskapsintyg
dina barns födelseattester.
Observera att utländska handlingar ska vara legaliserade och översatta till finska, svenska eller engelska.
Du kan också ansöka om personbeteckning från magistraten.
Läs mer: Registrering som invånare, Hemkommun i Finland.
Registrering av utlänningarfinska _ svenska _ engelska
Kontaktuppgifter till magistratfinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
Du kan få:
kostnadsfri rådgivning och information kring att flytta på flera olika språk
en finländsk personbeteckning, registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1-intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
I tjänsten medverkar Helsingfors-info, magistraten i Nyland, skatteförvaltningens och FPA:s tjänst In To Finland, NTM-centralen i Nyland, Pensionsskyddscentralen och Helsingforsregionens handelskammare.
Adress
Albertsgatan 25
IHH – serviceställe för dig som flyttar till Finland engelska
Tillståndsärenden
På Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU-medborgarens uppehållsrätt.
Migrationsverkets tjänsteställe i Helsingfors :
Göksgränd 3A
Du kan också ansöka om många slags uppehållstillstånd och EU-registrering på internet i tjänsten Enter Finland.
Om du inte är van vid att använda en dator, fyll i en ansökan på papper och lämna in den på Migrationsverkets tjänsteställe.
Dät är alltid bra att boka en tid i förväg på tjänstestället.
Du kan boka en tid på Migrationsverkets tidsbokningstjänst.
Observera att tjänstestället inte kan ge rådgivning om tillståndsärenden.
Läs mer: Flytta till Finland.
Elektronisk tidsbokningfinska _ svenska _ engelska
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Registrering som invånare
Om du flyttar ditt stadigvarande boende till Esbo, ska du registrera dig som invånare i kommunen.
Du kan registrera dig vid magistraten i Nyland, Helsingfors enhet.
Magistraten i Nyland Helsingfors enhet
Tfn 029 55 39391
När du går till magistraten ska du ta med dig
legitimation (till exempel pass)
uppehållstillstånd och uppehållskort (om du behöver uppehållstillstånd i Finland)
registreringsintyget över uppehållsrätten (oleskeluoikeuden rekisteröintitodistus) om du är EU-medborgare.
äktenskapsintyg
dina barns födelseattester.
Observera att utländska handlingar ska vara legaliserade och översatta till finska, svenska eller engelska.
Du kan också ansöka om personbeteckning från magistraten.
Läs mer: Registrering som invånare, Hemkommun i Finland.
Registrering av utlänningarfinska _ svenska _ engelska
Kontaktuppgifter till magistratfinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
Du kan få:
kostnadsfri rådgivning och information kring att flytta på flera olika språk
en finländsk personbeteckning, registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1-intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
I tjänsten medverkar Helsingfors-info, magistraten i Nyland, skatteförvaltningens och FPA:s tjänst In To Finland, NTM-centralen i Nyland, Pensionsskyddscentralen och Helsingforsregionens handelskammare.
Adress
IHH – serviceställe för dig som flyttar till Finland engelska
Tillståndsärenden
På Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU-medborgarens uppehållsrätt.
Migrationsverkets tjänsteställe i Helsingfors :
Göksgränd 3A
Du kan också ansöka om många slags uppehållstillstånd och EU-registrering på internet i tjänsten Enter Finland.
Om du inte är van vid att använda en dator, fyll i en ansökan på papper och lämna in den på Migrationsverkets tjänsteställe.
Dät är alltid bra att boka en tid i förväg på tjänstestället.
Du kan boka en tid på Migrationsverkets tidsbokningstjänst.
Observera att tjänstestället inte kan ge rådgivning om tillståndsärenden.
Läs mer: Flytta till Finland.
Elektronisk tidsbokningfinska _ svenska _ engelska
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Registrering som invånare
Om du flyttar ditt stadigvarande boende till Esbo, ska du registrera dig som invånare i kommunen.
Du kan registrera dig vid magistraten i Nyland, Helsingfors enhet.
Magistraten i Nyland Helsingfors enhet
Tfn 029 55 39391
När du går till magistraten ska du ta med dig
legitimation (till exempel pass)
uppehållstillstånd och uppehållskort (om du behöver uppehållstillstånd i Finland)
registreringsintyget över uppehållsrätten (oleskeluoikeuden rekisteröintitodistus) om du är EU-medborgare.
äktenskapsintyg
dina barns födelseattester.
Observera att utländska handlingar ska vara legaliserade och översatta till finska, svenska eller engelska.
Du kan också ansöka om personbeteckning från magistraten.
Läs mer: Registrering som invånare, Hemkommun i Finland.
Registrering av utlänningarfinska _ svenska _ engelska
Kontaktuppgifter till magistratfinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
Du kan få:
kostnadsfri rådgivning och information kring att flytta på flera olika språk
en finländsk personbeteckning, registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1-intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
I tjänsten medverkar Helsingfors-info, magistraten i Nyland, skatteförvaltningens och FPA:s tjänst In To Finland, NTM-centralen i Nyland, Pensionsskyddscentralen och Helsingforsregionens handelskammare.
Adress
IHH – serviceställe för dig som flyttar till Finland engelska
Trafiken
Beslutsfattande och påverkan
Religion
Basfakta
Historia
Trafiken
Huvudstadsregionen har goda kollektivtrafikförbindelser.
I Helsingfors trafikerar tåg, bussar, spårvagnar, metron och Sveaborgsfärjorna.
Helsingfors är med i samkommunen Helsingforsregionens trafik (HRT) (Helsingin seudun liikenne -kuntayhtymä (HSL)) som sköter kollektivtrafiken i huvudstadsregionen.
I tjänsten Reseplaneraren (Reittiopas-palvelu) kan du söka information om kollektivtrafikens rutter i huvudstadsregionen.
Tjänsten ger dig förslag på olika kollektivtrafikförbindelser från ett ställe till ett annat.
I kollektivtrafikens färdmedel kan du betala med kontanter eller resekort (matkakortti).
Reseplanerarefinska _ svenska _ engelska _ ryska
Resekort
Med ett resekort (matkakortti) reser du förmånligare än med kontanter.
Resekortet gäller i lokaltrafikens bussar, närtågen, metron, spårvagnarna och Sveaborgsfärjorna.
Det finns två slags resekort.
Det är det billigaste sättet att resa.
Ett innehavarkort (haltijakohtainen kortti) kan användas av flera personer.
Innan du skaffar dig ett personligt kort ska du registrera dig som invånare i någon av kommunerna inom HRT-området.
Du kan köpa resekort vid HRT:s försäljningsställen (myyntipiste) eller serviceställen (palvelupiste).
De finns runtom i huvudstadsregionen.
Personligt resekort kan du köpa vid serviceställena.
Ta med dig identitetsbevis om du ska köpa personligt resekort.
Om du har finska nätbankskoder kan du även köpa personligt resekort på HRT:s webbplats.
Du kan resa med resekortet när du laddar kortet med period (kausi) eller värde (arvo).
En period betyder tid: till exempel en månad.
Värde betyder pengar.
Om du använder kollektivtrafiken ofta tjänar du på att ladda kortet med period.
Du kan ladda resekortet på vilket serviceställe för resekort (matkakortin latauspiste) som helst.
Du hittar mer information på HRT:s webbplats.
Ansökan om försäljningsplatserfinska _ svenska _ engelska
Information och råd till resenärerfinska _ svenska _ engelska
På cykel och till fots
I Helsingfors finns gott om cykelvägar.
I reseplaneraren för cykel- och gångtrafiken kan du söka en lämplig rutt om du vill gå eller cykla.
Bil och flyg
På många metrostationer kan du parkera din bil gratis för att fortsätta resan med kollektivtrafiken.
Helsingfors har goda landsvägsförbindelsermed resten av landet.
Den närmaste flygplatsen är Helsingfors-Vanda flygplats.
Läs mer: Trafiken.
Resplan för cycling och gångfinska _ svenska _ engelska _ ryska
linkkiVR:
Tågtidtabellerfinska _ svenska _ engelska _ ryska
Anslutningsparkeringfinska _ svenska _ engelska
Flygplatsenfinska _ svenska _ engelska _ ryska _ kinesiska
Beslutsfattande och påverkan
I Helsingfors beslutas ärenden av stadsfullmäktige.
Fullmäktigeledamöterna representerar olika politiska grupper.
Fullmäktige väljs vart fjärde år genom kommunalval.
Du kan följa fullmäktiges sammanträden och få mer information om beslutsfattandet på Helsingforskanalen eller på stadens webbplats.
Borgmästaren och stadens aktörer ordnar boendemöten runtom i Helsingfors för invånarna där man berättar om och diskuterar stadens ärenden.
Du kan även själv påverka beslutsfattande.
Att rösta i kommunalvalet är ett viktigt sätt att påverka.
Du kan även delta i utvecklingen av staden via olika slags elektroniska kanaler.
Till exempel på Helsingfors stads webbplats finns en färdig blankett, ett responssystem (palautejärjestelmä).
Via den kan du skicka frågor och förslag eller respons till staden.
I ditt bostadsområde arbetar dessutom stadens kontaktperson, stadslotsen (stadiluotsi), som kan hjälpa dig att föra vidare ditt förslag.
Stadslotsen har jour i områdets bibliotek vissa veckodagar och klockslag.
Mer information om stadslotsar och kontaktuppgifterna till dem hittar du på Helsingfors stads webbplats.
Stadsfullmäktigefinska _ svenska _ engelska
Stadsfullmäktiges sammanträden på Internetfinska _ svenska
Feedback till stadens ämbetsverk och inrättningarfinska _ svenska _ engelska
Delta och påverkafinska _ svenska _ engelska
Religion
I Helsingfors och Helsingforsregionen verkar många religiösa samfund.
I Helsingfors finns många olika religionssamfunds tempel och dessutom olika verksamhetscenter.
Via tjänsten Religionerna i Finland kan du söka information enligt religionssamfund och ort.
Läs mer: Kulturer och religioner i Finland.
Religiösa samfundfinska _ engelska
Basfakta
Helsingfors är Finlands huvudstad.
Staden ligger i södra Finland vid Finska viken.
Helsingfors är Finlands administrativa centrum: där sammanträder Finlands riksdag och där finns ministerierna.
Helsingfors är även ett viktigt centrum för affärs- och kulturlivet.
Helsingfors har cirka 600 000 invånare. 83 procent av invånarna har finska och 6 procent har svenska som modersmål.
11 procent har något annat modersmål.
Information om Helsingforsfinska _ svenska _ engelska
Helsingfors historia
Sveriges kung Gustav Vasa grundade Helsingfors på stranden av nuvarande Gammelstadsforsen genom att den 12 juni 1550 beordra invånare i andra städer att flytta till Helsingfors.
Finland var på den tiden en del av Sverige.
Gustav Vasa ville göra Helsingfors till en handelsstad som konkurrerar med Tallinn, och även holländska och tyska handelsmän flyttade till staden.
Inom kort erövrade Sverige Tallinn, och Helsingfors blev en krigsstad vars hamn användes för förflyttning av soldater först till Baltikum och på 1630-talet till tyska områden till trettioåriga kriget.
År 1640 flyttades Helsingfors till stadens nuvarande plats på Estnäs.
De första 200 åren var staden en anspråkslös småstad.
Under Stora nordiska kriget år 1710 föll två tredjedelar av Helsingfors befolkning offer till pesten.
Ryssland ockuperade Helsingfors två gånger på 1700-talet när Sverige och Ryssland var i krig.
År 1748 inleddes bygget av Sveaborgs sjöfästning på öarna utanför Helsingfors. (På finska Suomenlinna, "Finlands slott").
Bygget av fästningen förde med sig nya invånare till staden och också handeln blev livligare.
Helsingfors och Sveaborg erövrades av ryssarna 1808 och under kriget brann staden.
Ryssland gjorde området som erövrats till Finlands autonoma storfurstendöme.
År 1812 upphöjde kejsar Alexander I Helsingfors till Finlands huvudstad.
Samtidigt började man bygga Helsingfors innerstad i empirestil, vars byggnader inhyste storfurstendömets viktiga institutioner.
Också universitetet flyttades år 1828 från Åbo till Helsingfors.
När Finland blev självständigt år 1917 blev Helsingfors huvudstad i republiken Finland.
I januari 1918 tog det röda gardet, som representerade arbetarna, makten i HelsingforsHels.
Samtidigt organiserade sig de vita trupperna som representerade borgare och bönder i Österbotten och inbördeskriget bröt ut.
Tyska trupper som kom till Finland erövrade Helsingfors till de vita i april.
Under andra världskriget 1939–1944 bombade Sovjetunionen Helsingfors, men tack vare det duktiga luftvärnet vara skadorna i staden lindriga.
År 1946 inkorporerades nya områden till Helsingfors och staden yta mångfaldigades nästan åtta gånger.
Stadens befolkning växte snabbt och och på de inkorporerade områdena byggdes många nya förorter på 1950−1980-talen.
Helsingforsdagen firas varje år på dagen för stadens grundande, den 12 juni.
Då pågår många evenemang på olika håll i Helsingfors.
Helsingfors historiafinska _ svenska _ engelska
Trafiken
Beslutsfattande och påverkan
Religion
Basfakta
Historia
Trafiken
Huvudstadsregionen har goda kollektivtrafikförbindelser.
I Helsingfors trafikerar tåg, bussar, spårvagnar, metron och Sveaborgsfärjorna.
Helsingfors är med i samkommunen Helsingforsregionens trafik (HRT) (Helsingin seudun liikenne -kuntayhtymä (HSL)) som sköter kollektivtrafiken i huvudstadsregionen.
I tjänsten Reseplaneraren (Reittiopas-palvelu) kan du söka information om kollektivtrafikens rutter i huvudstadsregionen.
Tjänsten ger dig förslag på olika kollektivtrafikförbindelser från ett ställe till ett annat.
I kollektivtrafikens färdmedel kan du betala med kontanter eller resekort (matkakortti).
Reseplanerarefinska _ svenska _ engelska _ ryska
Resekort
Med ett resekort (matkakortti) reser du förmånligare än med kontanter.
Resekortet gäller i lokaltrafikens bussar, närtågen, metron, spårvagnarna och Sveaborgsfärjorna.
Det finns två slags resekort.
Det är det billigaste sättet att resa.
Ett innehavarkort (haltijakohtainen kortti) kan användas av flera personer.
Innan du skaffar dig ett personligt kort ska du registrera dig som invånare i någon av kommunerna inom HRT-området.
Du kan köpa resekort vid HRT:s försäljningsställen (myyntipiste) eller serviceställen (palvelupiste).
De finns runtom i huvudstadsregionen.
Personligt resekort kan du köpa vid serviceställena.
Ta med dig identitetsbevis om du ska köpa personligt resekort.
Om du har finska nätbankskoder kan du även köpa personligt resekort på HRT:s webbplats.
Du kan resa med resekortet när du laddar kortet med period (kausi) eller värde (arvo).
En period betyder tid: till exempel en månad.
Värde betyder pengar.
Om du använder kollektivtrafiken ofta tjänar du på att ladda kortet med period.
Du kan ladda resekortet på vilket serviceställe för resekort (matkakortin latauspiste) som helst.
Du hittar mer information på HRT:s webbplats.
Ansökan om försäljningsplatserfinska _ svenska _ engelska
Information och råd till resenärerfinska _ svenska _ engelska
På cykel och till fots
I Helsingfors finns gott om cykelvägar.
I reseplaneraren för cykel- och gångtrafiken kan du söka en lämplig rutt om du vill gå eller cykla.
Bil och flyg
På många metrostationer kan du parkera din bil gratis för att fortsätta resan med kollektivtrafiken.
Helsingfors har goda landsvägsförbindelsermed resten av landet.
Den närmaste flygplatsen är Helsingfors-Vanda flygplats.
Läs mer: Trafiken.
Resplan för cycling och gångfinska _ svenska _ engelska _ ryska
linkkiVR:
Tågtidtabellerfinska _ svenska _ engelska _ ryska
Anslutningsparkeringfinska _ svenska _ engelska
Flygplatsenfinska _ svenska _ engelska _ ryska _ kinesiska
Beslutsfattande och påverkan
I Helsingfors beslutas ärenden av stadsfullmäktige.
Fullmäktigeledamöterna representerar olika politiska grupper.
Fullmäktige väljs vart fjärde år genom kommunalval.
Du kan följa fullmäktiges sammanträden och få mer information om beslutsfattandet på Helsingforskanalen eller på stadens webbplats.
Borgmästaren och stadens aktörer ordnar boendemöten runtom i Helsingfors för invånarna där man berättar om och diskuterar stadens ärenden.
Du kan även själv påverka beslutsfattande.
Att rösta i kommunalvalet är ett viktigt sätt att påverka.
Du kan även delta i utvecklingen av staden via olika slags elektroniska kanaler.
Till exempel på Helsingfors stads webbplats finns en färdig blankett, ett responssystem (palautejärjestelmä).
Via den kan du skicka frågor och förslag eller respons till staden.
I ditt bostadsområde arbetar dessutom stadens kontaktperson, stadslotsen (stadiluotsi), som kan hjälpa dig att föra vidare ditt förslag.
Stadslotsen har jour i områdets bibliotek vissa veckodagar och klockslag.
Mer information om stadslotsar och kontaktuppgifterna till dem hittar du på Helsingfors stads webbplats.
Stadsfullmäktigefinska _ svenska _ engelska
Stadsfullmäktiges sammanträden på Internetfinska _ svenska
Feedback till stadens ämbetsverk och inrättningarfinska _ svenska _ engelska
Delta och påverkafinska _ svenska _ engelska
Religion
I Helsingfors och Helsingforsregionen verkar många religiösa samfund.
I Helsingfors finns många olika religionssamfunds tempel och dessutom olika verksamhetscenter.
Via tjänsten Religionerna i Finland kan du söka information enligt religionssamfund och ort.
Läs mer: Kulturer och religioner i Finland.
Religiösa samfundfinska _ engelska
Basfakta
Helsingfors är Finlands huvudstad.
Staden ligger i södra Finland vid Finska viken.
Helsingfors är Finlands administrativa centrum: där sammanträder Finlands riksdag och där finns ministerierna.
Helsingfors är även ett viktigt centrum för affärs- och kulturlivet.
Helsingfors har cirka 600 000 invånare. 83 procent av invånarna har finska och 6 procent har svenska som modersmål.
11 procent har något annat modersmål.
Information om Helsingforsfinska _ svenska _ engelska
Helsingfors historia
Sveriges kung Gustav Vasa grundade Helsingfors på stranden av nuvarande Gammelstadsforsen genom att den 12 juni 1550 beordra invånare i andra städer att flytta till Helsingfors.
Finland var på den tiden en del av Sverige.
Gustav Vasa ville göra Helsingfors till en handelsstad som konkurrerar med Tallinn, och även holländska och tyska handelsmän flyttade till staden.
Inom kort erövrade Sverige Tallinn, och Helsingfors blev en krigsstad vars hamn användes för förflyttning av soldater först till Baltikum och på 1630-talet till tyska områden till trettioåriga kriget.
År 1640 flyttades Helsingfors till stadens nuvarande plats på Estnäs.
De första 200 åren var staden en anspråkslös småstad.
Under Stora nordiska kriget år 1710 föll två tredjedelar av Helsingfors befolkning offer till pesten.
Ryssland ockuperade Helsingfors två gånger på 1700-talet när Sverige och Ryssland var i krig.
År 1748 inleddes bygget av Sveaborgs sjöfästning på öarna utanför Helsingfors. (På finska Suomenlinna, "Finlands slott").
Bygget av fästningen förde med sig nya invånare till staden och också handeln blev livligare.
Helsingfors och Sveaborg erövrades av ryssarna 1808 och under kriget brann staden.
Ryssland gjorde området som erövrats till Finlands autonoma storfurstendöme.
År 1812 upphöjde kejsar Alexander I Helsingfors till Finlands huvudstad.
Samtidigt började man bygga Helsingfors innerstad i empirestil, vars byggnader inhyste storfurstendömets viktiga institutioner.
Också universitetet flyttades år 1828 från Åbo till Helsingfors.
När Finland blev självständigt år 1917 blev Helsingfors huvudstad i republiken Finland.
I januari 1918 tog det röda gardet, som representerade arbetarna, makten i HelsingforsHels.
Samtidigt organiserade sig de vita trupperna som representerade borgare och bönder i Österbotten och inbördeskriget bröt ut.
Tyska trupper som kom till Finland erövrade Helsingfors till de vita i april.
Under andra världskriget 1939–1944 bombade Sovjetunionen Helsingfors, men tack vare det duktiga luftvärnet vara skadorna i staden lindriga.
År 1946 inkorporerades nya områden till Helsingfors och staden yta mångfaldigades nästan åtta gånger.
Stadens befolkning växte snabbt och och på de inkorporerade områdena byggdes många nya förorter på 1950−1980-talen.
Helsingforsdagen firas varje år på dagen för stadens grundande, den 12 juni.
Då pågår många evenemang på olika håll i Helsingfors.
Helsingfors historiafinska _ svenska _ engelska
Trafiken
Beslutsfattande och påverkan
Religion
Basfakta
Historia
Trafiken
Helsingfors är med i samkommunen Helsingforsregionens trafik (HRT) (Helsingin seudun liikenne -kuntayhtymä (HSL)) som sköter kollektivtrafiken i huvudstadsregionen.
Huvudstadsregionen har goda kollektivtrafikförbindelser.
I Helsingfors trafikerar tåg, bussar, spårvagnar, metron och Sveaborgsfärjorna.
I tjänsten Reseplaneraren (Reittiopas-palvelu) kan du söka information om kollektivtrafikens rutter i huvudstadsregionen.
Tjänsten ger dig förslag på olika kollektivtrafikförbindelser från ett ställe till ett annat.
I kollektivtrafikens färdmedel kan du betala med kontanter eller resekort (matkakortti).
Reseplanerarefinska _ svenska _ engelska
Resekort
Med ett resekort (matkakortti) reser du förmånligare än med kontanter.
Resekortet gäller i lokaltrafikens bussar, närtågen, metron, spårvagnarna och Sveaborgsfärjorna.
Det finns två slags resekort.
Det är det billigaste sättet att resa.
Ett innehavarkort (haltijakohtainen kortti) kan användas av flera personer.
Innan du skaffar dig ett personligt kort ska du registrera dig som invånare i någon av kommunerna inom HRT-området.
Du kan köpa resekort vid HRT:s försäljningsställen (myyntipiste) eller serviceställen (palvelupiste).
De finns runtom i huvudstadsregionen.
Personligt resekort kan du köpa vid serviceställena.
Ta med dig identitetsbevis om du ska köpa personligt resekort.
Om du har finska nätbankskoder kan du även köpa personligt resekort på HRT:s webbplats.
Du kan resa med resekortet när du laddar kortet med period (kausi) eller värde (arvo).
En period betyder tid: till exempel en månad.
Värde betyder pengar.
Om du använder kollektivtrafiken ofta tjänar du på att ladda kortet med period.
Du kan ladda resekortet på vilket serviceställe för resekort (matkakortin latauspiste) som helst.
Du hittar mer information på HRT:s webbplats.
Ansökan om försäljningsplatserfinska _ svenska _ engelska
Information och råd till resenärerfinska _ svenska _ engelska
På cykel och till fots
I Helsingfors finns gott om cykelvägar.
I reseplaneraren för cykel- och gångtrafiken kan du söka en lämplig rutt om du vill gå eller cykla.
Bil och flyg
På många metrostationer kan du parkera din bil gratis för att fortsätta resan med kollektivtrafiken.
Helsingfors har goda landsvägsförbindelsermed resten av landet.
Den närmaste flygplatsen är Helsingfors-Vanda flygplats.
Läs mer: Trafiken.
Resplan för cycling och gångfinska _ svenska _ engelska _ ryska
linkkiVR:
Tågtidtabellerfinska _ svenska _ engelska _ ryska
Anslutningsparkeringfinska _ svenska _ engelska
Flygplatsenfinska _ svenska _ engelska _ ryska _ kinesiska
Beslutsfattande och påverkan
I Helsingfors beslutas ärenden av stadsfullmäktige.
Fullmäktigeledamöterna representerar olika politiska grupper.
Fullmäktige väljs vart fjärde år genom kommunalval.
Du kan följa fullmäktiges sammanträden och få mer information om beslutsfattandet på Helsingforskanalen eller på stadens webbplats.
Borgmästaren och stadens aktörer ordnar boendemöten runtom i Helsingfors för invånarna där man berättar om och diskuterar stadens ärenden.
Du kan även själv påverka beslutsfattande.
Att rösta i kommunalvalet är ett viktigt sätt att påverka.
Du kan även delta i utvecklingen av staden via olika slags elektroniska kanaler.
Till exempel på Helsingfors stads webbplats finns en färdig blankett, ett responssystem (palautejärjestelmä).
Via den kan du skicka frågor och förslag eller respons till staden.
I ditt bostadsområde arbetar dessutom stadens kontaktperson, stadslotsen (stadiluotsi), som kan hjälpa dig att föra vidare ditt förslag.
Stadslotsen har jour i områdets bibliotek vissa veckodagar och klockslag.
Mer information om stadslotsar och kontaktuppgifterna till dem hittar du på Helsingfors stads webbplats.
Stadsfullmäktigefinska _ svenska _ engelska
Stadsfullmäktiges sammanträden på Internetfinska _ svenska
Feedback till stadens ämbetsverk och inrättningarfinska _ svenska _ engelska
Delta och påverkafinska _ svenska _ engelska
Religion
I Helsingfors och Helsingforsregionen verkar många religiösa samfund.
I Helsingfors finns många olika religionssamfunds tempel och dessutom olika verksamhetscenter.
Via tjänsten Religionerna i Finland kan du söka information enligt religionssamfund och ort.
Läs mer: Kulturer och religioner i Finland.
Religiösa samfundfinska _ engelska
Basfakta
Helsingfors är Finlands huvudstad.
Staden ligger i södra Finland vid Finska viken.
Helsingfors är Finlands administrativa centrum: där sammanträder Finlands riksdag och där finns ministerierna.
Helsingfors är även ett viktigt centrum för affärs- och kulturlivet.
Helsingfors har cirka 650 000 invånare. 78 procent av invånarna har finska och 6 procent har svenska som modersmål.
16 procent har något annat modersmål.
Information om Helsingfors(pdf, 5,9 MB)finska _ svenska _ engelska _ ryska _ franska _ kinesiska _ tyska
Helsingfors historia
Sveriges kung Gustav Vasa grundade Helsingfors på stranden av nuvarande Gammelstadsforsen genom att den 12 juni 1550 beordra invånare i andra städer att flytta till Helsingfors.
Finland var på den tiden en del av Sverige.
Gustav Vasa ville göra Helsingfors till en handelsstad som konkurrerar med Tallinn, och även holländska och tyska handelsmän flyttade till staden.
Inom kort erövrade Sverige Tallinn, och Helsingfors blev en krigsstad vars hamn användes för förflyttning av soldater först till Baltikum och på 1630-talet till tyska områden till trettioåriga kriget.
År 1640 flyttades Helsingfors till stadens nuvarande plats på Estnäs.
De första 200 åren var staden en anspråkslös småstad.
Under Stora nordiska kriget år 1710 föll två tredjedelar av Helsingfors befolkning offer till pesten.
Ryssland ockuperade Helsingfors två gånger på 1700-talet när Sverige och Ryssland var i krig.
År 1748 inleddes bygget av Sveaborgs sjöfästning på öarna utanför Helsingfors. (På finska Suomenlinna, "Finlands slott").
Bygget av fästningen förde med sig nya invånare till staden och också handeln blev livligare.
Helsingfors och Sveaborg erövrades av ryssarna 1808 och under kriget brann staden.
Ryssland gjorde området som erövrats till Finlands autonoma storfurstendöme.
År 1812 upphöjde kejsar Alexander I Helsingfors till Finlands huvudstad.
Samtidigt började man bygga Helsingfors innerstad i empirestil, vars byggnader inhyste storfurstendömets viktiga institutioner.
Också universitetet flyttades år 1828 från Åbo till Helsingfors.
När Finland blev självständigt år 1917 blev Helsingfors huvudstad i republiken Finland.
I januari 1918 tog det röda gardet, som representerade arbetarna, makten i HelsingforsHels.
Samtidigt organiserade sig de vita trupperna som representerade borgare och bönder i Österbotten och inbördeskriget bröt ut.
Tyska trupper som kom till Finland erövrade Helsingfors till de vita i april.
Under andra världskriget 1939–1944 bombade Sovjetunionen Helsingfors, men tack vare det duktiga luftvärnet vara skadorna i staden lindriga.
År 1946 inkorporerades nya områden till Helsingfors och staden yta mångfaldigades nästan åtta gånger.
Stadens befolkning växte snabbt och och på de inkorporerade områdena byggdes många nya förorter på 1950−1980-talen.
Helsingforsdagen firas varje år på dagen för stadens grundande, den 12 juni.
Då pågår många evenemang på olika håll i Helsingfors.
Helsingfors historiafinska _ svenska _ engelska
Bibliotek
Motion
Att röra sig i naturen
Teater och filmer
Museer
Hobbyer för barn och unga
Föreningar
Evenemang
Evenemang och sevärt i Helsingforsfinska _ svenska _ engelska _ ryska _ kinesiska _ tyska
Evenemangskalendrar och sökmaskinerfinska _ svenska _ engelska
Helsingfors evenemangskalenderfinska _ svenska _ engelska
Helsingfors evenemangskalenderfinska
Bibliotek
I Helsingfors finns många bibliotek på olika håll i staden.
I staden finns dessutom två bokbussar som åker runt.
Helsingfors stads bibliotek är en del av HelMet-biblioteket.
Till HelMet-biblioteket hör även biblioteken i Esbo, Vanda och Grankulla.
HelMet-biblioteken har en gemensam webbtjänst.
På webbtjänsten kan du söka och reservera material.
Du kan också förnya dina lån på Internet.
Nästan alla bibliotekstjänster är kostnadsfria.
För att kunna använda bibliotekstjänsterna behöver du ett bibliotekskort.
Du kan hämta ditt bibliotekskort vid vilket HelMet-bibliotek som helst.
Alla personer som har en adress i Finland kan få ett bibliotekskort.
Om du inte har en finländsk personbeteckning, är ditt bibliotekskort i kraft ett år i taget.
I biblioteken i Helsingfors finns mest böcker på finska, men du kan även låna böcker på många andra språk där.
I många bibliotek hittar du böcker på engelska, tyska, franska, italienska, spanska, estniska och ryska.
Flerspråkiga biblioteket
I huvudbiblioteket i Böle finns det flerspråkiga bibliotekets samling (monikielinen kirjasto).
Där finns böcker på fler än 60 olika språk.
Du kan också beställa böckerna till andra bibliotek.
Om du har ett bibliotekskort, kan du även läsa e-böcker och e-tidningar samt titta på filmer på din egen dator, läsplatta eller smarttelefon.
I Helsingfors finns även andra bibliotek, till exempel vid universiteten och högskolorna.
Läs mer: Bibliotek.
Bibliotek och öppettiderfinska _ svenska _ engelska
linkkiHelsingfors stadsbibliotek:
Flerspråkiga biblioteketfinska _ svenska _ engelska
Bibliotekets webbtjänstfinska _ svenska _ engelska
Motion
Du kan idka många slags motion på olika håll i Helsingfors.
I Helsingfors finns många simhallar, gym, idrottsplatser och motionsspår.
Helsingfors stad ordnar idrottskurser för stadsbor.
På sommaren ordnas avgiftsfri parkgympa på många håll i staden.
Läs mer: Motion.
Filmklipp om motionsalternativfinska _ engelska _ somaliska _ arabiska
Utomhusmotionfinska _ svenska _ engelska
Inomhusmotionfinska _ svenska _ engelska
Idrottsklubbarfinska _ svenska _ engelska
Handledd motionfinska _ svenska _ engelska
Att röra sig i naturen
I Helsingfors har man nära till naturen.
Du kan promenera eller cykla alternativt åka metro, buss, tåg spårvagn eller färja till parker, stränder, skogar eller naturskyddsområden.
På Helsingfors stads webbplats hittar du information om skogen i Helsingfors och i närheten av Helsingfors.
I Helsingfors finns även öar för friluftsliv som du når med ruttfärjor.
Sveaborg och Stora Räntan är också historiska sevärdheter.
Mer information om öarna och vattentrafiken får du på Helsingfors stads webbplats.
På sidan finns även information om båtliv i Helsingfors.
Du kan meta med metspö och pimpla på isen utan ett separat tillstånd.
Det är avgiftsfritt.
För annat fiske behöver du ett avgiftsbelagt tillstånd.
På Helsingfors stads webbplats finns mer information om var du kan köpa fisketillstånd.
Lämna inte linor eller annat fiskeavfall i naturen.
De kan orsaka stora plågor för fåglar och andra djur.
Läs mer: Att röra sig i naturen.
Friluftsområdenfinska _ svenska _ engelska
Friluftsliv i skärgårdenfinska _ svenska _ engelska
Båtlivfinska _ svenska _ engelska
Försäljningsställen för fisketillståndfinska _ svenska _ engelska
Teater och filmer
I Helsingfors finns många teatrar.
De flesta föreställningarna är finskspråkiga.
I Helsingfors finns även svenskspråkiga teatrar.
Du kan söka teaterföreställningar i evenemangskalendrarna på sidorna helsinki.fi och stadissa.fi.
I Helsingfors finns ett filmarkiv och flera biografer.
Information om vilka filmer som visas hittar du på biografernas webbplatser.
I evenemangskalendrarna hittar du information om filmfestivaler i Helsingfors.
Läs mer: Teater och filmer.
Information om filmer och filmvisningarfinska _ svenska _ engelska
Biograffinska
linkkiFinnkino:
Filmerfinska _ engelska
Museer
I Helsingfors finns många museer.
Mer information om museerna får du från Helsingfors turistbyrå.
Adress: Brunnsgatan 1 (Helsingfors huvudjärnvägsstation)
Tfn: 09 31013300
Läs mer: Museer.
Museer och utställningarfinska _ svenska _ engelska
linkkiAteneum:
Ateneumfinska _ svenska _ engelska
linkkiKiasma:
Museet för nutidskonst Kiasmafinska _ svenska _ engelska _ ryska
Designmuseetfinska _ svenska _ engelska
Sveaborgfinska _ svenska _ engelska
linkkiMuseiverket:
Fölisöns friluftsmuseumfinska _ svenska _ engelska _ franska _ tyska
linkkiMuseiverket:
Finlands nationalmuseumfinska _ svenska _ engelska
Naturhistoriska centralmuseetfinska _ svenska _ engelska _ ryska
Museer i Helsingforsfinska _ svenska _ engelska _ ryska _ kinesiska _ tyska
Hobbyer för barn och unga
Annegårdens konstcentrum är ett konsthus för barn och unga i centrala Helsingfors.
Adressen är Annegatan 30.
På Annegården ges konstundervisning och visas utställningar, dansföreställningar och teaterföreställningar.
Också i de andra konsthusen i Helsingfors ordnas kulturevenemang för barn och unga.
Barnkulturcentret Musikantit är ett aktivitetscenter med familjeevenemang, barnkonserter, utställningar och teater.
På centret kan barn studera musik, teater, bildkonst och dans på olika språk.
För barn finns även många idrottshobbyer.
Helsingfors stad ordnar till exempel gymnastik, simskolor och många andra idrottsaktiviteter för barn.
Också många privata företag erbjuder idrottshobbyer för barn.
Ungdomscentralen (Nuorisoasiainkeskus) erbjuder många idrottsmöjligheter till 9–18-åriga barn och unga.
På webbplatsen Munstadi.fi finns mycket information om aktiviteter och hobbyer för unga.
I tjänsten finns även Ruuti, som samlar de ungas egna idéer och initiativ.
I Helsingfors finns även många ungdomsgårdar, där de unga kan vistas på fritiden.
Läs mer: Hobbyer för barn och unga.
Verksamhet och evenemang för ungafinska _ svenska _ engelska
Information om medlemskortetfinska _ svenska _ engelska _ ryska _ franska _ somaliska
Idrottsklubbarfinska _ svenska _ engelska
Kulturcentralens verksamhetsställenfinska _ svenska _ engelska
Barnkulturcentralen Musikantitfinska _ engelska _ ryska
Ungdomsgårdarfinska
Hobbysökningfinska
Stöd och verksamhet för flickorfinska
Föreningar
I Helsingfors finns ett stort antal olika föreningar, till exempel kulturföreningar och idrottsorganisationer.
I Helsingfors finns även många invandrarföreningar.
Läs mer: Föreningar.
Föreningsverksamhetfinska _ svenska _ engelska
Bibliotek
Motion
Att röra sig i naturen
Teater och filmer
Museer
Hobbyer för barn och unga
Föreningar
Evenemang
Evenemang och sevärt i Helsingforsfinska _ svenska _ engelska _ ryska _ kinesiska _ tyska
Evenemangskalendrar och sökmaskinerfinska _ svenska _ engelska
Helsingfors evenemangskalenderfinska _ svenska _ engelska
Helsingfors evenemangskalenderfinska
Bibliotek
I Helsingfors finns många bibliotek på olika håll i staden.
I staden finns dessutom två bokbussar som åker runt.
Helsingfors stads bibliotek är en del av HelMet-biblioteket.
Till HelMet-biblioteket hör även biblioteken i Esbo, Vanda och Grankulla.
HelMet-biblioteken har en gemensam webbtjänst.
På webbtjänsten kan du söka och reservera material.
Du kan också förnya dina lån på Internet.
Nästan alla bibliotekstjänster är kostnadsfria.
För att kunna använda bibliotekstjänsterna behöver du ett bibliotekskort.
Du kan hämta ditt bibliotekskort vid vilket HelMet-bibliotek som helst.
Alla personer som har en adress i Finland kan få ett bibliotekskort.
Om du inte har en finländsk personbeteckning, är ditt bibliotekskort i kraft ett år i taget.
I biblioteken i Helsingfors finns mest böcker på finska, men du kan även låna böcker på många andra språk där.
I många bibliotek hittar du böcker på engelska, tyska, franska, italienska, spanska, estniska och ryska.
Flerspråkiga biblioteket
I huvudbiblioteket i Böle finns det flerspråkiga bibliotekets samling (monikielinen kirjasto).
Där finns böcker på fler än 60 olika språk.
Du kan också beställa böckerna till andra bibliotek.
Om du har ett bibliotekskort, kan du även läsa e-böcker och e-tidningar samt titta på filmer på din egen dator, läsplatta eller smarttelefon.
I Helsingfors finns även andra bibliotek, till exempel vid universiteten och högskolorna.
Läs mer: Bibliotek.
Bibliotek och öppettiderfinska _ svenska _ engelska
linkkiHelsingfors stadsbibliotek:
Flerspråkiga biblioteketfinska _ svenska _ engelska
Bibliotekets webbtjänstfinska _ svenska _ engelska
Motion
Du kan idka många slags motion på olika håll i Helsingfors.
I Helsingfors finns många simhallar, gym, idrottsplatser och motionsspår.
Helsingfors stad ordnar idrottskurser för stadsbor.
På sommaren ordnas avgiftsfri parkgympa på många håll i staden.
Läs mer: Motion.
Filmklipp om motionsalternativfinska _ engelska _ somaliska _ arabiska
Utomhusmotionfinska _ svenska _ engelska
Inomhusmotionfinska _ svenska _ engelska
Idrottsklubbarfinska _ svenska _ engelska
Handledd motionfinska _ svenska _ engelska
Att röra sig i naturen
I Helsingfors har man nära till naturen.
Du kan promenera eller cykla alternativt åka metro, buss, tåg spårvagn eller färja till parker, stränder, skogar eller naturskyddsområden.
På Helsingfors stads webbplats hittar du information om skogen i Helsingfors och i närheten av Helsingfors.
I Helsingfors finns även öar för friluftsliv som du når med ruttfärjor.
Sveaborg och Stora Räntan är också historiska sevärdheter.
Mer information om öarna och vattentrafiken får du på Helsingfors stads webbplats.
På sidan finns även information om båtliv i Helsingfors.
Du kan meta med metspö och pimpla på isen utan ett separat tillstånd.
Det är avgiftsfritt.
För annat fiske behöver du ett avgiftsbelagt tillstånd.
På Helsingfors stads webbplats finns mer information om var du kan köpa fisketillstånd.
Lämna inte linor eller annat fiskeavfall i naturen.
De kan orsaka stora plågor för fåglar och andra djur.
Läs mer: Att röra sig i naturen.
Friluftsområdenfinska _ svenska _ engelska
Friluftsliv i skärgårdenfinska _ svenska _ engelska
Båtlivfinska _ svenska _ engelska
Försäljningsställen för fisketillståndfinska _ svenska _ engelska
Teater och filmer
I Helsingfors finns många teatrar.
De flesta föreställningarna är finskspråkiga.
I Helsingfors finns även svenskspråkiga teatrar.
Du kan söka teaterföreställningar i evenemangskalendrarna på sidorna helsinki.fi och stadissa.fi.
I Helsingfors finns ett filmarkiv och flera biografer.
Information om vilka filmer som visas hittar du på biografernas webbplatser.
I evenemangskalendrarna hittar du information om filmfestivaler i Helsingfors.
Läs mer: Teater och filmer.
Information om filmer och filmvisningarfinska _ svenska _ engelska
Biograffinska
linkkiFinnkino:
Filmerfinska _ engelska
Museer
I Helsingfors finns många museer.
Mer information om museerna får du från Helsingfors turistbyrå.
Adress: Brunnsgatan 1 (Helsingfors huvudjärnvägsstation)
Tfn: 09 31013300
Läs mer: Museer.
Museer och utställningarfinska _ svenska _ engelska
linkkiAteneum:
Ateneumfinska _ svenska _ engelska
linkkiKiasma:
Museet för nutidskonst Kiasmafinska _ svenska _ engelska _ ryska
Designmuseetfinska _ svenska _ engelska
Sveaborgfinska _ svenska _ engelska
linkkiMuseiverket:
Fölisöns friluftsmuseumfinska _ svenska _ engelska _ franska _ tyska
linkkiMuseiverket:
Finlands nationalmuseumfinska _ svenska _ engelska
Naturhistoriska centralmuseetfinska _ svenska _ engelska _ ryska
Museer i Helsingforsfinska _ svenska _ engelska _ ryska _ kinesiska _ tyska
Hobbyer för barn och unga
Annegårdens konstcentrum är ett konsthus för barn och unga i centrala Helsingfors.
Adressen är Annegatan 30.
På Annegården ges konstundervisning och visas utställningar, dansföreställningar och teaterföreställningar.
Också i de andra konsthusen i Helsingfors ordnas kulturevenemang för barn och unga.
Barnkulturcentret Musikantit är ett aktivitetscenter med familjeevenemang, barnkonserter, utställningar och teater.
På centret kan barn studera musik, teater, bildkonst och dans på olika språk.
För barn finns även många idrottshobbyer.
Helsingfors stad ordnar till exempel gymnastik, simskolor och många andra idrottsaktiviteter för barn.
Också många privata företag erbjuder idrottshobbyer för barn.
Ungdomscentralen (Nuorisoasiainkeskus) erbjuder många idrottsmöjligheter till 9–18-åriga barn och unga.
På webbplatsen Munstadi.fi finns mycket information om aktiviteter och hobbyer för unga.
I tjänsten finns även Ruuti, som samlar de ungas egna idéer och initiativ.
I Helsingfors finns även många ungdomsgårdar, där de unga kan vistas på fritiden.
Läs mer: Hobbyer för barn och unga.
Verksamhet och evenemang för ungafinska _ svenska _ engelska
Information om medlemskortetfinska _ svenska _ engelska _ ryska _ franska _ somaliska
Idrottsklubbarfinska _ svenska _ engelska
Kulturcentralens verksamhetsställenfinska _ svenska _ engelska
Barnkulturcentralen Musikantitfinska _ engelska _ ryska
Ungdomsgårdarfinska
Hobbysökningfinska
Stöd och verksamhet för flickorfinska
Föreningar
I Helsingfors finns ett stort antal olika föreningar, till exempel kulturföreningar och idrottsorganisationer.
I Helsingfors finns även många invandrarföreningar.
Läs mer: Föreningar.
Föreningsverksamhetfinska _ svenska _ engelska
Bibliotek
Motion
Att röra sig i naturen
Teater och filmer
Museer
Hobbyer för barn och unga
Föreningar
Evenemang
Evenemang och sevärt i Helsingforsfinska _ svenska _ engelska _ ryska _ kinesiska _ tyska
Evenemang vid Helsingfors universitetfinska _ svenska _ engelska
Helsingfors evenemangskalenderfinska _ svenska _ engelska
Evenemang och platser i Helsingforsfinska
Bibliotek
I Helsingfors finns många bibliotek på olika håll i staden.
I staden finns dessutom två bokbussar som åker runt.
Helsingfors stads bibliotek är en del av HelMet-biblioteket.
Till HelMet-biblioteket hör även biblioteken i Esbo, Vanda och Grankulla.
HelMet-biblioteken har en gemensam webbtjänst.
På webbtjänsten kan du söka och reservera material.
Du kan också förnya dina lån på Internet.
Nästan alla bibliotekstjänster är kostnadsfria.
För att kunna använda bibliotekstjänsterna behöver du ett bibliotekskort.
Du kan hämta ditt bibliotekskort vid vilket HelMet-bibliotek som helst.
Alla personer som har en adress i Finland kan få ett bibliotekskort.
Om du inte har en finländsk personbeteckning, är ditt bibliotekskort i kraft ett år i taget.
I biblioteken i Helsingfors finns mest böcker på finska, men du kan även låna böcker på många andra språk där.
I många bibliotek hittar du böcker på engelska, tyska, franska, italienska, spanska, estniska och ryska.
Flerspråkiga biblioteket
I huvudbiblioteket i Böle finns det flerspråkiga bibliotekets samling (monikielinen kirjasto).
Där finns böcker på fler än 60 olika språk.
Du kan också beställa böckerna till andra bibliotek.
Om du har ett bibliotekskort, kan du även läsa e-böcker och e-tidningar samt titta på filmer på din egen dator, läsplatta eller smarttelefon.
I Helsingfors finns även andra bibliotek, till exempel vid universiteten och högskolorna.
Läs mer: Bibliotek.
Huvudstadsregionens gemensamma bibliotekstjänstfinska _ svenska _ engelska _ ryska _ somaliska _ persiska _ arabiska
Bibliotek och öppettiderfinska _ svenska _ engelska _ ryska
linkkiHelsingfors stadsbibliotek:
Flerspråkiga biblioteketfinska _ svenska _ engelska _ ryska
Motion
Du kan idka många slags motion på olika håll i Helsingfors.
I Helsingfors finns många simhallar, gym, idrottsplatser och motionsspår.
Helsingfors stad ordnar idrottskurser för stadsbor.
På sommaren ordnas avgiftsfri parkgympa på många håll i staden.
Läs mer: Motion.
Motion och friluftsliv i Helsingforsfinska _ svenska _ engelska
Inomhusmotionfinska _ svenska _ engelska
Idrottsklubbarfinska _ svenska _ engelska
Handledd motionfinska _ svenska _ engelska
Att röra sig i naturen
I Helsingfors har man nära till naturen.
Du kan promenera eller cykla alternativt åka metro, buss, tåg spårvagn eller färja till parker, stränder, skogar eller naturskyddsområden.
På Helsingfors stads webbplats hittar du information om skogen i Helsingfors och i närheten av Helsingfors.
I Helsingfors finns även öar för friluftsliv som du når med ruttfärjor.
Sveaborg och Stora Räntan är också historiska sevärdheter.
Mer information om öarna och vattentrafiken får du på Helsingfors stads webbplats.
På sidan finns även information om båtliv i Helsingfors.
Du kan meta med metspö och pimpla på isen utan ett separat tillstånd.
Det är avgiftsfritt.
För annat fiske behöver du ett avgiftsbelagt tillstånd.
På Helsingfors stads webbplats finns mer information om var du kan köpa fisketillstånd.
Lämna inte linor eller annat fiskeavfall i naturen.
De kan orsaka stora plågor för fåglar och andra djur.
Läs mer: Att röra sig i naturen.
Friluftsområdenfinska _ svenska _ engelska
Friluftsliv i skärgårdenfinska _ svenska _ engelska
Båtlivfinska _ svenska _ engelska
Försäljningsställen för fisketillståndfinska _ svenska _ engelska
Teater och filmer
I Helsingfors finns många teatrar.
De flesta föreställningarna är finskspråkiga.
I Helsingfors finns även svenskspråkiga teatrar.
Du kan söka teaterföreställningar i evenemangskalendrarna på sidorna myhelsinki.fi och stadissa.fi.
I Helsingfors finns ett filmarkiv och flera biografer.
Information om vilka filmer som visas hittar du på biografernas webbplatser.
I evenemangskalendrarna hittar du information om filmfestivaler i Helsingfors.
Läs mer: Teater och filmer.
Information om filmer och filmvisningarfinska _ svenska _ engelska
Biograffinska _ engelska _ ryska _ estniska
Biograffinska
linkkiFinnkino:
Filmerfinska _ engelska
Museer
I Helsingfors finns många museer.
Mer information om museerna får du från Helsingfors turistbyrå.
Adress: Brunnsgatan 1 (Helsingfors huvudjärnvägsstation)
Tfn: 09 31013300
Läs mer: Museer.
Museer och utställningarfinska _ svenska _ engelska
linkkiAteneum:
Ateneumfinska _ svenska _ engelska
linkkiKiasma:
Museet för nutidskonst Kiasmafinska _ svenska _ engelska _ ryska
Designmuseetfinska _ svenska _ engelska
Sveaborgfinska _ svenska _ engelska
linkkiMuseiverket:
Fölisöns friluftsmuseumfinska _ svenska _ engelska _ franska _ tyska
linkkiMuseiverket:
Finlands nationalmuseumfinska _ svenska _ engelska
Naturhistoriska centralmuseetfinska _ svenska _ engelska _ ryska
Museer i Helsingforsfinska _ svenska _ engelska _ ryska _ kinesiska _ tyska
Hobbyer för barn och unga
Annegårdens konstcentrum är ett konsthus för barn och unga i centrala Helsingfors.
Adressen är Annegatan 30.
På Annegården ges konstundervisning och visas utställningar, dansföreställningar och teaterföreställningar.
Också i de andra konsthusen i Helsingfors ordnas kulturevenemang för barn och unga.
Barnkulturcentret Musikantit är ett aktivitetscenter med familjeevenemang, barnkonserter, utställningar och teater.
På centret kan barn studera musik, teater, bildkonst och dans på olika språk.
För barn finns även många idrottshobbyer.
Helsingfors stad ordnar till exempel gymnastik, simskolor och många andra idrottsaktiviteter för barn.
Också många privata företag erbjuder idrottshobbyer för barn.
Ungdomscentralen (Nuorisoasiainkeskus) erbjuder många idrottsmöjligheter till 9–18-åriga barn och unga.
På webbplatsen Munstadi.fi finns mycket information om aktiviteter och hobbyer för unga.
I tjänsten finns även Ruuti, som samlar de ungas egna idéer och initiativ.
I Helsingfors finns även många ungdomsgårdar, där de unga kan vistas på fritiden.
Läs mer: Hobbyer för barn och unga.
Verksamhet och evenemang för ungafinska _ svenska _ engelska
Information om medlemskortetfinska _ svenska _ engelska _ ryska _ franska _ somaliska
Idrottsklubbarfinska _ svenska _ engelska
Kulturcentralens verksamhetsställenfinska _ svenska _ engelska
Barnkulturcentralen Musikantitfinska _ engelska _ ryska
Ungdomsgårdarfinska _ svenska _ engelska
Hobbysökningfinska _ svenska _ engelska
Stöd och verksamhet för flickorfinska
Föreningar
I Helsingfors finns ett stort antal olika föreningar, till exempel kulturföreningar och idrottsorganisationer.
I Helsingfors finns även många invandrarföreningar.
Läs mer: Föreningar.
Föreningsverksamhetfinska _ svenska _ engelska
Problem med uppehållstillståndet
Brott
Behöver du en jurist?
Våld
Problem i äktenskap eller parförhållande
Barns och ungas problem
Missbruksproblem
Dödsfall
Ring nödnumret 112 om det är fråga om en nödsituation.
Via nödnumret kan du tillkalla polis, ambulans eller brandkår.
Ring inte nödnumret om det inte är en nödsituation.
Socialjouren
Socialjouren (sosiaalipäivystys) hjälper kvällstid och under veckoslut om du är i akut behov av hjälp av en socialarbetare.
Socialjouren
Tfn 020 696 006
Krisjouren
På Krisjouren (kriisipäivystys) kan du få psykisk första hjälpen och stöd om du hamnar i en plötslig krissituation.
Plötsliga krissituationer kan till exempel vara en allvarlig olycka, att en närstående avlider eller att du blir offer för våld.
Du kan ringa jourtelefonen dygnet runt.
Telefonnumret är (09) 310 44222
Per telefon betjänar socialjouren och krisjouren på finska, svenska och i mån av möjlighet även på engelska.
Vid möten kan tolk användas.
Social- och krisjourenfinska _ svenska _ engelska
Problem med uppehållstillståndet
Om du har problem eller oklarheter med uppehållstillståndet, kan du ta kontakt med migrationsverket.
Du kan även fråga om råd vid Helsinki-info.
Telefon: 09 310 11111, mån.–tors. kl. 9–16, fre. kl. 10–15
Serviceställen:
Centrumbiblioteket Oodi, adress: Tölöviksgatan 1
Elektroniskt:
Rådgivning på chattenfinska _ svenska _ engelska
Skicka en fråga eller ge oss responsfinska _ svenska _ engelska
Flyktingar och asylsökande samt andra utlänningar kan söka hjälp och råd i frågor kring uppehållstillståndet hos Flyktingrådgivningen rf.
Adress: Kaisaniemigatan 4 A, vån. 6
Tfn 075 7575 100
Läs mer: Problem med uppehållstillstånd.
Brott
Om du behöver brådskande hjälp av polisen i en nödsituation, ring nödnumret 112.
Ring inte nödnumret om det inte är fråga om en nödsituation.
En brottsanmälan kan du göra på polisstationen.
Om det inte är fråga om ett allvarligt brott, kan du även göra brottsanmälan elektroniskt via polisens webbplats.
Läs mer: Brott.
Kontaktuppgifter till polisstationernafinska _ svenska _ engelska
Elektronisk polisanmälanfinska _ svenska _ engelska
Om du behöver rättshjälp, kan du kontakta Helsingfors rättshjälpsbyrå (Helsingin oikeusaputoimisto).
Adress: Porkalagatan 13 G, vån 2
Tfn 029 56 60120
Du kan även söka fram en privat advokat via Finlands Juristförbunds webbplats.
Läs mer: Behöver du en jurist?
linkkiFinlands Advokatförbund:
Advokaterfinska _ svenska _ engelska
Våld
Hjälp till invandrarkvinnor
Om du har blivit utsatt för våld eller hot, kan du få hjälp och stöd hos Kriscentret Monika.
Diu kan boka en tid genom att ringa hjälptelefonen i förväg eller besöka centret.
Tjänsten är helt konfidentiell och du behöver inte uppge ditt namn.
Du kan få hjälp på flera olika språk.
Hjälptelefon 0800 05058, mån.–fre. klockan 9–16
Adress: Hermanstads Strandväg 12 A, vån. 4
Öppettider: mån-fre 9-17
Skyddshem
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du ta dig till ett skyddshem (turvakoti).
Skyddshemmet Mona är ett skyddshem avsett för invandrarkvinnor och deras barn.
Du kan ta dig till ett skyddshem om det på grund av våld är för farligt att vistas hemma.
Skyddshemmets adress är hemlig.
Tfn 045 639 6274
Du kan även ta dig till Huvudstadens Skyddshem.
Adress: Steniusvägen 20
Tfn (09) 4777 180
Hjälp för män
Tjänsten Miehen Linja (Miehen Linja) är en tjänst som hjälper män, som har utsatt sin partner för våld.
Tjänsten är avsedd för män som flyttat till Finland, oberoende av bostadsort.
Tfn 09 276 62 8 99
På Miehen Linja kan du prata på finska, svenska, engelska, franska och grekiska eller medelst en tolk på ditt modersmål.
Läs mer: Våld.
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Hjälp till offer för familjevåldfinska
Hjälp för män för att sluta med våldsamt beteendefinska _ engelska
Problem i äktenskap eller parförhållande
Duo erbjuder relationsrådgivning för par från två kulturer på finska och engelska.
Rådgivningen är avgiftsbelagd.
Väestöliitto erbjuder parrådgivning och parterapi på finska och engelska.
Läs mer: Problem i äktenskap och parförhållande.
Relationsrådgivning för par från två kulturerfinska _ engelska
Sökning av relationsrådgivningstjänsterfinska _ svenska _ engelska
Barns och ungas problem
Hälsovårdaren vid barnrådgivningen ger råd i frågor som rör små barns hälsa, uppväxt och utveckling.
Om du behöver råd i sådant som rör fostran av barn eller barns utveckling, kan du boka en tid hos familjerådgivningen (perheneuvola).
Familjerådgivningen betjänar barn under 18 år och deras föräldrar.
Väestöliitto ger råd till invandrarfamiljer i frågor rörande barnfostran och familjens välmående.
Rådgivningen på olika språk:
Tfn 09-228 05 245 och 050 325 6450 (sorani, dari, persiska)
Tfn 09-228 05141, mobil 050 325 7173 (ryska, engelska)
Helsingfors ungdomsstation (Helsingin nuorisoasema) erbjuder hjälp till 13–23-åriga unga Helsingforsbor.
Du kan till exempel få hjälp med psykiska problem och missbruksproblem samt hjälp att sluta spela.
Också den ungas föräldrar kan kontakta ungdomsstationen.
Flickor kan få stöd och råd i Flickornas hus (Tyttöjen talo) och pojkar i Pojkarnas hus (Poikien talo).
Röda Korset har ett skyddshus för 12–19-åriga unga.
På De ungas skyddshus kan du få samtalshjälp och tillfällig logi.
Kontaktuppgifter till De ungas skyddshus:
Öppettider: varje dag kl. 17.00–10.00
Tfn (09) 622 4322
Information om rådgivningsbyråernas tjänsterfinska _ svenska _ engelska
Familjerådgivningfinska _ svenska _ engelska
linkkiFinlands Röda Kors:
De ungas skyddshus i Helsingforsfinska _ svenska
Stöd och verksamhet för flickorfinska
Om du har ekonomiska problem kan du fråga om råd hos en socialarbetare i din hemkommun eller hos FPA.I vissa situationer har du rätt till utkomststöd.
Du kan ansöka om utkomststöd hos FPA.
Information om utkomststödfinska _ svenska _ engelska _ ryska _ estniska
Ekonomi- och skuldrådgivning
Om du har problem med skulder, kontakta rättshjälpsbyråns ekonomi- och skuldrådgivning.
Tjänsten är kostnadsfri.
Helsingfors rättshjälpsbyrå
Ekonomi- och skuldrådgivning
Tfn 029 56 60123 mån–fre kl. 8–16.15
linkkiRättshjälpsbyrå:
Ekonomi- och skuldrådgivningfinska _ svenska _ engelska
Missbruks​problem
Om du behöver hjälp med ett missbruksproblem (såsom alkohol- eller drogmissbruk), kan du kontakta din närmaste hälsostation.
Du kan också kontakta A-kliniken.
Unga i åldern 13–23 med missbruksproblem kan få hjälp vid ungdomsstationen.
Läs mer: Missbruksproblem.
Missbrukarvårdfinska _ engelska
Dödsfall
Begravningsbyråer hjälper med de praktiska arrangemangen vid en begravning.
Du kan söka begravningsbyråer till exempel på Finlands begravningsbyråers förbunds webbplats.
I Helsingfors finns flera begravningsplatser.
Den evangelisk-lutherska kyrkan sköter om de flesta av dem.
I Sandudd finns dessutom Helsingfors ortodoxa begravningsplats, Helsingfors judiska begravningsplats och Helsingfors muslimska begravningsplats för tatarer.
Muslimerna i Helsingfors har sitt eget gravkvarter på Furumo begravningsplats i Vanda.
På Furumo begravningsplats finns även ett gravområde för konfessionslösa. Där kan de avlidna begravas som inte hörde till ett religionssamfund.
Om en närstående har avlidit och du behöver psykiskt stöd, kan du ringa krisjouren (kriisipäivystys).
Du kan ringa jourtelefonen dygnet runt.
Telefonnumret är (09) 310 44222
Läs mer: Dödsfall.
linkkiFinlands Begravningbyråers Förbund:
Begravningsbyråerfinska _ svenska _ engelska
linkkiHelsingfors kyrkliga samfällighet:
Begravningsplatserfinska _ svenska
linkkiHelsingfors kyrkliga samfällighet:
Muslimernas gravkvarterfinska
linkkiHelsingfors kyrkliga samfällighet:
Konfessionslös begravningsplatsfinska
Problem med uppehållstillståndet
Brott
Behöver du en jurist?
Våld
Problem i äktenskap eller parförhållande
Barns och ungas problem
Missbruksproblem
Dödsfall
Ring nödnumret 112 om det är fråga om en nödsituation.
Via nödnumret kan du tillkalla polis, ambulans eller brandkår.
Ring inte nödnumret om det inte är en nödsituation.
Socialjouren
Socialjouren (sosiaalipäivystys) hjälper kvällstid och under veckoslut om du är i akut behov av hjälp av en socialarbetare.
Socialjouren
Tfn 020 696 006
Krisjouren
På Krisjouren (kriisipäivystys) kan du få psykisk första hjälpen och stöd om du hamnar i en plötslig krissituation.
Plötsliga krissituationer kan till exempel vara en allvarlig olycka, att en närstående avlider eller att du blir offer för våld.
Du kan ringa jourtelefonen dygnet runt.
Telefonnumret är (09) 310 44222
Per telefon betjänar socialjouren och krisjouren på finska, svenska och i mån av möjlighet även på engelska.
Vid möten kan tolk användas.
Social- och krisjourenfinska _ svenska _ engelska
Problem med uppehållstillståndet
Om du har problem eller oklarheter med uppehållstillståndet, kan du ta kontakt med migrationsverket.
Du kan även fråga om råd vid Helsinki-info.
Telefon: 09 310 11111, mån.–tors. kl. 9–16, fre. kl. 10–15
Serviceställen:
Centrumbiblioteket Oodi, adress: Tölöviksgatan 1
Elektroniskt:
Rådgivning på chattenfinska _ svenska _ engelska
Skicka en fråga eller ge oss responsfinska _ svenska _ engelska
Flyktingar och asylsökande samt andra utlänningar kan söka hjälp och råd i frågor kring uppehållstillståndet hos Flyktingrådgivningen rf.
Adress: Kaisaniemigatan 4 A, vån. 6
Tfn 075 7575 100
Läs mer: Problem med uppehållstillstånd.
Brott
Om du behöver brådskande hjälp av polisen i en nödsituation, ring nödnumret 112.
Ring inte nödnumret om det inte är fråga om en nödsituation.
En brottsanmälan kan du göra på polisstationen.
Om det inte är fråga om ett allvarligt brott, kan du även göra brottsanmälan elektroniskt via polisens webbplats.
Läs mer: Brott.
Kontaktuppgifter till polisstationernafinska _ svenska _ engelska
Elektronisk polisanmälanfinska _ svenska _ engelska
Om du behöver rättshjälp, kan du kontakta Helsingfors rättshjälpsbyrå (Helsingin oikeusaputoimisto).
Adress: Porkalagatan 13 G, vån 2
Tfn 029 56 60120
Du kan även söka fram en privat advokat via Finlands Juristförbunds webbplats.
Läs mer: Behöver du en jurist?
linkkiFinlands Advokatförbund:
Advokaterfinska _ svenska _ engelska
Våld
Hjälp till invandrarkvinnor
Om du har blivit utsatt för våld eller hot, kan du få hjälp och stöd hos Kriscentret Monika.
Diu kan boka en tid genom att ringa hjälptelefonen i förväg eller besöka centret.
Tjänsten är helt konfidentiell och du behöver inte uppge ditt namn.
Du kan få hjälp på flera olika språk.
Hjälptelefon 0800 05058, mån.–fre. klockan 9–16
Adress: Hermanstads Strandväg 12 A, vån. 4
Öppettider: mån-fre 9-17
Skyddshem
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du ta dig till ett skyddshem (turvakoti).
Skyddshemmet Mona är ett skyddshem avsett för invandrarkvinnor och deras barn.
Du kan ta dig till ett skyddshem om det på grund av våld är för farligt att vistas hemma.
Skyddshemmets adress är hemlig.
Tfn 045 639 6274
Du kan även ta dig till Huvudstadens Skyddshem.
Adress: Steniusvägen 20
Tfn (09) 4777 180
Hjälp för män
Tjänsten Miehen Linja (Miehen Linja) är en tjänst som hjälper män, som har utsatt sin partner för våld.
Tjänsten är avsedd för män som flyttat till Finland, oberoende av bostadsort.
Tfn 09 276 62 8 99
På Miehen Linja kan du prata på finska, svenska, engelska, franska och grekiska eller medelst en tolk på ditt modersmål.
Läs mer: Våld.
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Hjälp till offer för familjevåldfinska
Hjälp för män för att sluta med våldsamt beteendefinska _ engelska
Problem i äktenskap eller parförhållande
Duo erbjuder relationsrådgivning för par från två kulturer på finska och engelska.
Rådgivningen är avgiftsbelagd.
Väestöliitto erbjuder parrådgivning och parterapi på finska och engelska.
Läs mer: Problem i äktenskap och parförhållande.
Relationsrådgivning för par från två kulturerfinska _ engelska
Sökning av relationsrådgivningstjänsterfinska _ svenska _ engelska
Barns och ungas problem
Hälsovårdaren vid barnrådgivningen ger råd i frågor som rör små barns hälsa, uppväxt och utveckling.
Om du behöver råd i sådant som rör fostran av barn eller barns utveckling, kan du boka en tid hos familjerådgivningen (perheneuvola).
Familjerådgivningen betjänar barn under 18 år och deras föräldrar.
Väestöliitto ger råd till invandrarfamiljer i frågor rörande barnfostran och familjens välmående.
Rådgivningen på olika språk:
Tfn 09-228 05 245 och 050 325 6450 (sorani, dari, persiska)
Tfn 09-228 05141, mobil 050 325 7173 (ryska, engelska)
Helsingfors ungdomsstation (Helsingin nuorisoasema) erbjuder hjälp till 13–23-åriga unga Helsingforsbor.
Du kan till exempel få hjälp med psykiska problem och missbruksproblem samt hjälp att sluta spela.
Också den ungas föräldrar kan kontakta ungdomsstationen.
Flickor kan få stöd och råd i Flickornas hus (Tyttöjen talo) och pojkar i Pojkarnas hus (Poikien talo).
Röda Korset har ett skyddshus för 12–19-åriga unga.
På De ungas skyddshus kan du få samtalshjälp och tillfällig logi.
Kontaktuppgifter till De ungas skyddshus:
Öppettider: varje dag kl. 17.00–10.00
Tfn (09) 622 4322
Information om rådgivningsbyråernas tjänsterfinska _ svenska _ engelska
Familjerådgivningfinska _ svenska _ engelska
linkkiFinlands Röda Kors:
De ungas skyddshus i Helsingforsfinska _ svenska
Stöd och verksamhet för flickorfinska
Om du har ekonomiska problem kan du fråga om råd hos en socialarbetare i din hemkommun eller hos FPA.I vissa situationer har du rätt till utkomststöd.
Du kan ansöka om utkomststöd hos FPA.
Information om utkomststödfinska _ svenska _ engelska _ ryska _ estniska
Ekonomi- och skuldrådgivning
Om du har problem med skulder, kontakta rättshjälpsbyråns ekonomi- och skuldrådgivning.
Tjänsten är kostnadsfri.
Helsingfors rättshjälpsbyrå
Ekonomi- och skuldrådgivning
Tfn 029 56 60123 mån–fre kl. 8–16.15
linkkiRättshjälpsbyrå:
Ekonomi- och skuldrådgivningfinska _ svenska _ engelska
Missbruks​problem
Om du behöver hjälp med ett missbruksproblem (såsom alkohol- eller drogmissbruk), kan du kontakta din närmaste hälsostation.
Du kan också kontakta A-kliniken.
Unga i åldern 13–23 med missbruksproblem kan få hjälp vid ungdomsstationen.
Läs mer: Missbruksproblem.
Missbrukarvårdfinska _ engelska
Dödsfall
Begravningsbyråer hjälper med de praktiska arrangemangen vid en begravning.
Du kan söka begravningsbyråer till exempel på Finlands begravningsbyråers förbunds webbplats.
I Helsingfors finns flera begravningsplatser.
Den evangelisk-lutherska kyrkan sköter om de flesta av dem.
I Sandudd finns dessutom Helsingfors ortodoxa begravningsplats, Helsingfors judiska begravningsplats och Helsingfors muslimska begravningsplats för tatarer.
Muslimerna i Helsingfors har sitt eget gravkvarter på Furumo begravningsplats i Vanda.
På Furumo begravningsplats finns även ett gravområde för konfessionslösa. Där kan de avlidna begravas som inte hörde till ett religionssamfund.
Om en närstående har avlidit och du behöver psykiskt stöd, kan du ringa krisjouren (kriisipäivystys).
Du kan ringa jourtelefonen dygnet runt.
Telefonnumret är (09) 310 44222
Läs mer: Dödsfall.
linkkiFinlands Begravningbyråers Förbund:
Begravningsbyråerfinska
linkkiHelsingfors kyrkliga samfällighet:
Begravningsplatserfinska _ svenska
linkkiHelsingfors kyrkliga samfällighet:
Muslimernas gravkvarterfinska
linkkiHelsingfors kyrkliga samfällighet:
Konfessionslös begravningsplatsfinska
Problem med uppehållstillståndet
Brott
Behöver du en jurist?
Våld
Problem i äktenskap eller parförhållande
Barns och ungas problem
Missbruksproblem
Dödsfall
Ring nödnumret 112 om det är fråga om en nödsituation.
Via nödnumret kan du tillkalla polis, ambulans eller brandkår.
Ring inte nödnumret om det inte är en nödsituation.
Socialjouren
Socialjouren (sosiaalipäivystys) hjälper kvällstid och under veckoslut om du är i akut behov av hjälp av en socialarbetare.
Socialjouren
Tfn 020 696 006
Krisjouren
På Krisjouren (kriisipäivystys) kan du få psykisk första hjälpen och stöd om du hamnar i en plötslig krissituation.
Plötsliga krissituationer kan till exempel vara en allvarlig olycka, att en närstående avlider eller att du blir offer för våld.
Du kan ringa jourtelefonen dygnet runt.
Telefonnumret är (09) 310 44222
Per telefon betjänar socialjouren och krisjouren på finska, svenska och i mån av möjlighet även på engelska.
Vid möten kan tolk användas.
Social- och krisjourenfinska _ svenska _ engelska
Problem med uppehållstillståndet
Om du har problem eller oklarheter med uppehållstillståndet, kan du ta kontakt med migrationsverket.
Du kan även fråga om råd vid Helsinki-info.
Telefon: 09 310 11111, mån.–tors. kl. 9–16, fre. kl. 10–15
Serviceställen:
Centrumbiblioteket Oodi, adress: Tölöviksgatan 4
Elektroniskt:
Rådgivning på chattenfinska _ svenska _ engelska
Skicka en fråga eller ge oss responsfinska _ svenska _ engelska
Flyktingar och asylsökande samt andra utlänningar kan söka hjälp och råd i frågor kring uppehållstillståndet hos Flyktingrådgivningen rf.
Adress: Kaisaniemigatan 4 A, vån. 6
Tfn 075 7575 100
Läs mer: Problem med uppehållstillstånd.
Brott
Om du behöver brådskande hjälp av polisen i en nödsituation, ring nödnumret 112.
Ring inte nödnumret om det inte är fråga om en nödsituation.
En brottsanmälan kan du göra på polisstationen.
Om det inte är fråga om ett allvarligt brott, kan du även göra brottsanmälan elektroniskt via polisens webbplats.
Läs mer: Brott.
Kontaktuppgifter till polisstationernafinska _ svenska _ engelska
Elektronisk polisanmälanfinska _ svenska _ engelska
Om du behöver rättshjälp, kan du kontakta Helsingfors rättshjälpsbyrå (Helsingin oikeusaputoimisto).
Adress: Porkalagatan 13 G, vån 2
Tfn 029 56 60120
Du kan även söka fram en privat advokat via Finlands Juristförbunds webbplats.
Läs mer: Behöver du en jurist?
linkkiFinlands Advokatförbund:
Advokaterfinska _ svenska _ engelska
Våld
Hjälp till invandrarkvinnor
Om du har blivit utsatt för våld eller hot, kan du få hjälp och stöd hos Kriscentret Monika.
Diu kan boka en tid genom att ringa hjälptelefonen i förväg eller besöka centret.
Tjänsten är helt konfidentiell och du behöver inte uppge ditt namn.
Du kan få hjälp på flera olika språk.
Hjälptelefon 0800 05058, mån.–fre. klockan 9–16
Adress: Hermanstads Strandväg 12 A, vån. 4
Öppettider: mån-fre 9-17
Skyddshem
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du ta dig till ett skyddshem (turvakoti).
Skyddshemmet Mona är ett skyddshem avsett för invandrarkvinnor och deras barn.
Du kan ta dig till ett skyddshem om det på grund av våld är för farligt att vistas hemma.
Skyddshemmets adress är hemlig.
Tfn 045 639 6274
Du kan även ta dig till Huvudstadens Skyddshem.
Adress: Steniusvägen 20
Tfn (09) 4777 180
Hjälp för män
Tjänsten Miehen Linja (Miehen Linja) är en tjänst som hjälper män, som har utsatt sin partner för våld.
Tjänsten är avsedd för män som flyttat till Finland, oberoende av bostadsort.
Tfn 09 276 62 8 99
På Miehen Linja kan du prata på finska, svenska, engelska, franska och grekiska eller medelst en tolk på ditt modersmål.
Läs mer: Våld.
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Hjälp till offer för familjevåldfinska
Hjälp för män för att sluta med våldsamt beteendefinska _ engelska
Problem i äktenskap eller parförhållande
Duo erbjuder relationsrådgivning för par från två kulturer på finska och engelska.
Rådgivningen är avgiftsbelagd.
Väestöliitto erbjuder parrådgivning och parterapi på finska och engelska.
Läs mer: Problem i äktenskap och parförhållande.
Relationsrådgivning för par från två kulturerfinska _ engelska
Sökning av relationsrådgivningstjänsterfinska _ svenska _ engelska
Barns och ungas problem
Hälsovårdaren vid barnrådgivningen ger råd i frågor som rör små barns hälsa, uppväxt och utveckling.
Om du behöver råd i sådant som rör fostran av barn eller barns utveckling, kan du boka en tid hos familjerådgivningen (perheneuvola).
Familjerådgivningen betjänar barn under 18 år och deras föräldrar.
Väestöliitto ger råd till invandrarfamiljer i frågor rörande barnfostran och familjens välmående.
Rådgivningen på olika språk:
Tfn 09-228 05 245 och 050 325 6450 (sorani, dari, persiska)
Tfn 09-228 05141, mobil 050 325 7173 (ryska, engelska)
Helsingfors ungdomsstation (Helsingin nuorisoasema) erbjuder hjälp till 13–23-åriga unga Helsingforsbor.
Du kan till exempel få hjälp med psykiska problem och missbruksproblem samt hjälp att sluta spela.
Också den ungas föräldrar kan kontakta ungdomsstationen.
Flickor kan få stöd och råd i Flickornas hus (Tyttöjen talo) och pojkar i Pojkarnas hus (Poikien talo).
Röda Korset har ett skyddshus för 12–19-åriga unga.
På De ungas skyddshus kan du få samtalshjälp och tillfällig logi.
Kontaktuppgifter till De ungas skyddshus:
Öppettider: varje dag kl. 17.00–10.00
Tfn (09) 622 4322
Information om rådgivningsbyråernas tjänsterfinska _ svenska _ engelska
Familjerådgivningfinska _ svenska _ engelska
linkkiFinlands Röda Kors:
De ungas skyddshus i Helsingforsfinska _ svenska
Stöd och verksamhet för flickorfinska
Om du har ekonomiska problem kan du fråga om råd hos en socialarbetare i din hemkommun eller hos FPA.I vissa situationer har du rätt till utkomststöd.
Du kan ansöka om utkomststöd hos FPA.
Information om utkomststödfinska _ svenska _ engelska _ ryska _ estniska
Ekonomi- och skuldrådgivning
Om du har problem med skulder, kontakta rättshjälpsbyråns ekonomi- och skuldrådgivning.
Tjänsten är kostnadsfri.
Helsingfors rättshjälpsbyrå
Ekonomi- och skuldrådgivning
Tfn 029 56 60123 mån–fre kl. 8–16.15
linkkiRättshjälpsbyrå:
Ekonomi- och skuldrådgivningfinska _ svenska _ engelska
Missbruks​problem
Om du behöver hjälp med ett missbruksproblem (såsom alkohol- eller drogmissbruk), kan du kontakta din närmaste hälsostation.
Du kan också kontakta A-kliniken.
Unga i åldern 13–23 med missbruksproblem kan få hjälp vid ungdomsstationen.
Läs mer: Missbruksproblem.
Missbrukarvårdfinska _ engelska
Dödsfall
Begravningsbyråer hjälper med de praktiska arrangemangen vid en begravning.
Du kan söka begravningsbyråer till exempel på Finlands begravningsbyråers förbunds webbplats.
I Helsingfors finns flera begravningsplatser.
Den evangelisk-lutherska kyrkan sköter om de flesta av dem.
I Sandudd finns dessutom Helsingfors ortodoxa begravningsplats, Helsingfors judiska begravningsplats och Helsingfors muslimska begravningsplats för tatarer.
Muslimerna i Helsingfors har sitt eget gravkvarter på Furumo begravningsplats i Vanda.
På Furumo begravningsplats finns även ett gravområde för konfessionslösa. Där kan de avlidna begravas som inte hörde till ett religionssamfund.
Om en närstående har avlidit och du behöver psykiskt stöd, kan du ringa krisjouren (kriisipäivystys).
Du kan ringa jourtelefonen dygnet runt.
Telefonnumret är (09) 310 44222
Läs mer: Dödsfall.
linkkiFinlands Begravningbyråers Förbund:
Begravningsbyråerfinska
linkkiHelsingfors kyrkliga samfällighet:
Begravningsplatserfinska _ svenska
linkkiHelsingfors kyrkliga samfällighet:
Muslimernas gravkvarterfinska
linkkiHelsingfors kyrkliga samfällighet:
Konfessionslös begravningsplatsfinska
Äktenskap
Skilsmässa
Barnets födelse
Vård av barnet
Lekparker och klubbar
Problem i familjen
Äktenskap
Före äktenskapet måste du begära prövning av äktenskapshinder.
Hindersprövningen görs på magistraten (maistraatti).
Begär hindersprövning på magistraten i god tid före bröllopsdagen.
Borgerliga vigslar förrättas på magistraten.
Boka tid för vigseln hos magistraten.
Magistraten i Helsingfors
Adress: Albertsgatan 25
Tfn 029 55 39391
Läs mer:
Äktenskap.
Vigselfinska _ svenska _ engelska
Skilsmässa
Kvinnan eller mannen kan lämna skilsmässoansökan i Helsingfors tingsrätts kansli.
Man kan också söka skilsmässa ensam.
Du kan skicka in ansökan till tingsrättens kansli per post eller via e-post.
Tfn 029 56 44200
När ni överväger att skiljas och behöver hjälp med att komma överens om saker, kan ni ansöka om medling i familjeärenden (perheasioiden sovittelu).
Läs mer: Skilsmässa.
Skilsmässoansökan(pdf, 100 kb)finska _ svenska
linkkiRättsväsendet:
Helsingfors tingsrättfinska _ svenska _ engelska
Förmedling i familjefrågorfinska _ svenska _ engelska
Barn vid skilsmässa
Om ni har barn och beslutar er för att skiljas ska ni boka en tid hos barnatillsyningsmannen (lastenvalvoja).
Barnatillsyningsmannen bekräftar överenskommelsen om var barnen ska bo, vården av barnen, umgängesrätt och underhållsbidrag.
Bokning av tid till barnatillsynsmannen:
Tfn (09) 310 44999
Tfn (09) 310 43447
Om ni behöver hjälp med att komma överens om sådant som rör barnen kan ni ansöka om medling i familjeärenden.
Läs mer: Barn vid skilsmässa.
Barnatillsyningsmännenfinska _ svenska _ engelska
Barnets födelse
Uppgifterna om barnets födelse skickas från sjukhuset till befolkningsdataregistret i Finland.
Du ska meddela barnets namn, modersmål och andra erforderliga uppgifter till magistraten (Maistraatti) med en separat blankett som skickas hem till dig.
Du kan läsa mer om registrering av barnets födelse, faderskapserkännande och vårdnaden om barnet på InfoFinlands sida: När ett barn föds i Finland.
Vård av barnet
På InfoFinlands sida Utbildning i Helsingfors hittar du information om dagvården av barn i Helsingfors.
Tillfällig vård av barn
I lekparkerna i Helsingfors stad finns parktanter (puistotäti).
Parktanterna erbjuder tillfällig hjälp med skötsel av barn på förmiddagar.
Parktanten övervakar och leder barnen som leker i parken.
Parktanterna sköter barnen mot en avgift.
Om du behöver en tillfällig barnskötare hem, kan du kontakta Mannerheims Barnskyddsförbund (Mannerheimin Lastensuojeluliitto) eller Väestöliitto (Väestöliitto).
Parktanterfinska _ svenska _ engelska
Barnavård och hemhjälpfinska
linkkiMannerheims barnskyddsförbund:
Barnvaktshjälpfinska
Läs mer:Vård av barnet.
Hemvårdsstöd
Om du sköter ett barn som är yngre än tre år hemma kan du ansöka om hemvårdsstöd (kotihoidon tuki).
Du ansöker om stödet från FPA.
Helsingfors stad betalar dessutom ett kommuntillägg vid hemvårdsstöd till familjer som hemma sköter ett barn som är yngre än tre år.
Hemvårdsstöd för barn och Helsingforstilläggetfinska _ svenska _ engelska
Lekparker och klubbar
I Helsingfors finns det lekparker och familjehus, där det ordnas verksamhet för barn och föräldrar som sköter barnen hemma.
Verksamheten kan till exempel bestå av handledd motion, sång eller sysselsättning.
Stadin aikuisopisto ordnar i vissa lekparker och familjehus kurser i finska för invandrarföräldrar.
Lekparkerna och familjehusen ordnar vården av barnen under den tid kursen varar.
I daghem, familjehus och lekparker ordnas klubbar på deltid för barn i åldern 2–5, som inte är i dagvård.
Också Helsingfors församlingar har klubbverksamhet.
Lekparkerfinska _ svenska _ engelska
Verksamhet för barnfamiljerfinska _ svenska _ engelska
Filmklipp om lekparksverksamhetfinska _ svenska _ engelska _ somaliska _ persiska _ arabiska
Familjehusfinska _ svenska _ engelska
Klubbar för barnfinska _ svenska _ engelska
Problem i familjen
På InfoFinlands sida Problematiska situationer i Helsingfors får du information om var i Helsingfors man kan få hjälp med barns och ungas problem, eller vid problem i familjen.
Information om barns och ungas problem finns också på InfoFinlands sida Barns och ungas problem.
På InfoFinlands sida Problem i äktenskap eller parförhållande, får du information om var du kan få råd vid problem i äktenskapet eller i parförhållandet.
Äktenskap
Skilsmässa
Barnets födelse
Vård av barnet
Lekparker och klubbar
Problem i familjen
Äldre människor
Äktenskap
Före äktenskapet måste du begära prövning av äktenskapshinder.
Hindersprövningen görs på magistraten (maistraatti).
Begär hindersprövning på magistraten i god tid före bröllopsdagen.
Borgerliga vigslar förrättas på magistraten.
Boka tid för vigseln hos magistraten.
Magistraten i Helsingfors
Adress: Fågelviksgränden 2
Tfn 029 55 39391
Läs mer:
Äktenskap.
Vigselfinska _ svenska _ engelska
Skilsmässa
Kvinnan eller mannen kan lämna skilsmässoansökan i Helsingfors tingsrätts kansli.
Man kan också söka skilsmässa ensam.
Du kan skicka in ansökan till tingsrättens kansli per post eller via e-post.
Tfn 029 56 44200
När ni överväger att skiljas och behöver hjälp med att komma överens om saker, kan ni ansöka om medling i familjeärenden (perheasioiden sovittelu).
Läs mer: Skilsmässa.
Skilsmässoansökan(pdf, 100 kb)finska _ svenska
linkkiRättsväsendet:
Helsingfors tingsrättfinska _ svenska _ engelska
Förmedling i familjefrågorfinska _ svenska _ engelska
Barn vid skilsmässa
Om ni har barn och beslutar er för att skiljas ska ni boka en tid hos barnatillsyningsmannen (lastenvalvoja).
Barnatillsyningsmannen bekräftar överenskommelsen om var barnen ska bo, vården av barnen, umgängesrätt och underhållsbidrag.
Bokning av tid till barnatillsynsmannen:
Tfn (09) 310 44999
Tfn (09) 310 43447
Om ni behöver hjälp med att komma överens om sådant som rör barnen kan ni ansöka om medling i familjeärenden.
Läs mer: Barn vid skilsmässa.
Barnatillsyningsmännenfinska _ svenska _ engelska
Barnets födelse
Uppgifterna om barnets födelse skickas från sjukhuset till befolkningsdataregistret i Finland.
Du ska meddela barnets namn, modersmål och andra erforderliga uppgifter till magistraten (Maistraatti) med en separat blankett som skickas hem till dig.
Du kan läsa mer om registrering av barnets födelse, faderskapserkännande och vårdnaden om barnet på InfoFinlands sida: När ett barn föds i Finland.
Vård av barnet
På InfoFinlands sida Utbildning i Helsingfors hittar du information om dagvården av barn i Helsingfors.
Tillfällig vård av barn
I lekparkerna i Helsingfors stad finns parktanter (puistotäti).
Parktanterna erbjuder tillfällig hjälp med skötsel av barn på förmiddagar.
Parktanten övervakar och leder barnen som leker i parken.
Parktanterna sköter barnen mot en avgift.
Om du behöver en tillfällig barnskötare hem, kan du kontakta Mannerheims Barnskyddsförbund (Mannerheimin Lastensuojeluliitto) eller Väestöliitto (Väestöliitto).
Parktanterfinska _ svenska _ engelska
Barnavård och hemhjälpfinska
linkkiMannerheims barnskyddsförbund:
Barnvaktshjälpfinska
Läs mer:Vård av barnet.
Hemvårdsstöd
Om du sköter ett barn som är yngre än tre år hemma kan du ansöka om hemvårdsstöd (kotihoidon tuki).
Du ansöker om stödet från FPA.
Helsingfors stad betalar dessutom ett kommuntillägg vid hemvårdsstöd till familjer som hemma sköter ett barn som är yngre än tre år.
Hemvårdsstöd för barn och Helsingforstilläggetfinska _ svenska _ engelska
Lekparker och klubbar
I Helsingfors finns det lekparker och familjehus, där det ordnas verksamhet för barn och föräldrar som sköter barnen hemma.
Verksamheten kan till exempel bestå av handledd motion, sång eller sysselsättning.
Stadin aikuisopisto ordnar i vissa lekparker och familjehus kurser i finska för invandrarföräldrar.
Lekparkerna och familjehusen ordnar vården av barnen under den tid kursen varar.
I daghem, familjehus och lekparker ordnas klubbar på deltid för barn i åldern 2–5, som inte är i dagvård.
Också Helsingfors församlingar har klubbverksamhet.
Lekparkerfinska _ svenska _ engelska
Verksamhet för barnfamiljerfinska _ svenska _ engelska
Filmklipp om lekparksverksamhetfinska _ svenska _ engelska _ somaliska _ persiska _ arabiska
Familjehusfinska _ svenska _ engelska
Klubbar för barnfinska _ svenska _ engelska
Problem i familjen
På InfoFinlands sida Problematiska situationer i Helsingfors får du information om var i Helsingfors man kan få hjälp med barns och ungas problem, eller vid problem i familjen.
Information om barns och ungas problem finns också på InfoFinlands sida Barns och ungas problem.
På InfoFinlands sida Problem i äktenskap eller parförhållande, får du information om var du kan få råd vid problem i äktenskapet eller i parförhållandet.
Äldre människor
Helsingfors stads Seniorinfo ger råd om tjänster för äldre i Helsingfors.
Äldre i Helsingfors och deras anhöriga kan kontakta Seniorinfo.
Seniorinfo betjänar på finska och svenska.
Seniori-info
Tfn 09 3104 4556 (mån–fre kl. 9–15)
Seniorinfofinska _ svenska _ engelska
När du tar hand om en anhörig i hemmet
När du tar hand om en gammal eller sjuk anhörig eller en anhörig med funktionsnedsättning för att han eller hon ska kunna bo kvar i sitt hem, kan du ha rätt till stöd för närståendevård.
Du får närmare uppgifter vid social- och närarbetets verksamhetsställe i ditt bostadsområde (sosiaali- ja lähityön toimipiste).
Läs mer: Äldre människor.
Enheterna för socialt arbete och närarbetefinska _ svenska _ engelska
Stöd för närståendevårdfinska _ svenska _ engelska
Äktenskap
Skilsmässa
Barnets födelse
Vård av barnet
Lekparker och klubbar
Problem i familjen
Äldre människor
Äktenskap
Före äktenskapet måste du begära prövning av äktenskapshinder.
Hindersprövningen görs på magistraten (maistraatti).
Begär hindersprövning på magistraten i god tid före bröllopsdagen.
Borgerliga vigslar förrättas på magistraten.
Boka tid för vigseln hos magistraten.
Magistraten i Helsingfors
Adress: Fågelviksgränden 2
Tfn 029 55 39391
Läs mer:
Äktenskap.
Vigselfinska _ svenska _ engelska
Skilsmässa
Kvinnan eller mannen kan lämna skilsmässoansökan i Helsingfors tingsrätts kansli.
Man kan också söka skilsmässa ensam.
Du kan skicka in ansökan till tingsrättens kansli per post eller via e-post.
Tfn 029 56 44200
När ni överväger att skiljas och behöver hjälp med att komma överens om saker, kan ni ansöka om medling i familjeärenden (perheasioiden sovittelu).
Läs mer: Skilsmässa.
Skilsmässoansökan(pdf, 100 kb)finska _ svenska
linkkiRättsväsendet:
Helsingfors tingsrättfinska _ svenska _ engelska
Förmedling i familjefrågorfinska _ svenska _ engelska
Barn vid skilsmässa
Om ni har barn och beslutar er för att skiljas ska ni boka en tid hos barnatillsyningsmannen (lastenvalvoja).
Barnatillsyningsmannen bekräftar överenskommelsen om var barnen ska bo, vården av barnen, umgängesrätt och underhållsbidrag.
Bokning av tid till barnatillsynsmannen:
Tfn (09) 310 44999
Tfn (09) 310 43447
Om ni behöver hjälp med att komma överens om sådant som rör barnen kan ni ansöka om medling i familjeärenden.
Läs mer: Barn vid skilsmässa.
Barnatillsyningsmännenfinska _ svenska _ engelska
Barnets födelse
Uppgifterna om barnets födelse skickas från sjukhuset till befolkningsdataregistret i Finland.
Du ska meddela barnets namn, modersmål och andra erforderliga uppgifter till magistraten (Maistraatti) med en separat blankett som skickas hem till dig.
Du kan läsa mer om registrering av barnets födelse, faderskapserkännande och vårdnaden om barnet på InfoFinlands sida: När ett barn föds i Finland.
linkkiHUS (Helsingfors och Nylands sjukvårdsdistrikt):
På babyresa - För dig som har fött barnfinska _ svenska _ engelska
Vård av barnet
På InfoFinlands sida Utbildning i Helsingfors hittar du information om dagvården av barn i Helsingfors.
Tillfällig vård av barn
I lekparkerna i Helsingfors stad finns parktanter (puistotäti).
Parktanterna erbjuder tillfällig hjälp med skötsel av barn på förmiddagar.
Parktanten övervakar och leder barnen som leker i parken.
Parktanterna sköter barnen mot en avgift.
Om du behöver en tillfällig barnskötare hem, kan du kontakta Mannerheims Barnskyddsförbund (Mannerheimin Lastensuojeluliitto) eller Väestöliitto (Väestöliitto).
Parktanterfinska _ svenska _ engelska
Barnavård och hemhjälpfinska
linkkiMannerheims barnskyddsförbund:
Barnvaktshjälpfinska
Läs mer:Vård av barnet.
Hemvårdsstöd
Om du sköter ett barn som är yngre än tre år hemma kan du ansöka om hemvårdsstöd (kotihoidon tuki).
Du ansöker om stödet från FPA.
Helsingfors stad betalar dessutom ett kommuntillägg vid hemvårdsstöd till familjer som hemma sköter ett barn som är yngre än två år.
Hemvårdsstöd för barn och Helsingforstilläggetfinska _ svenska _ engelska
Lekparker och klubbar
I Helsingfors finns det lekparker och familjehus, där det ordnas verksamhet för barn och föräldrar som sköter barnen hemma.
Verksamheten kan till exempel bestå av handledd motion, sång eller sysselsättning.
Stadin aikuisopisto ordnar i vissa lekparker och familjehus kurser i finska för invandrarföräldrar.
Lekparkerna och familjehusen ordnar vården av barnen under den tid kursen varar.
I daghem, familjehus och lekparker ordnas klubbar på deltid för barn i åldern 2–5, som inte är i dagvård.
Också Helsingfors församlingar har klubbverksamhet.
Lekparkerfinska _ svenska _ engelska
Verksamhet för barnfamiljerfinska _ svenska _ engelska
Filmklipp om lekparksverksamhetfinska _ svenska _ engelska _ somaliska _ persiska _ arabiska
Familjehusfinska _ svenska _ engelska
Klubbar för barnfinska _ svenska _ engelska
Problem i familjen
På InfoFinlands sida Problematiska situationer i Helsingfors får du information om var i Helsingfors man kan få hjälp med barns och ungas problem, eller vid problem i familjen.
Information om barns och ungas problem finns också på InfoFinlands sida Barns och ungas problem.
På InfoFinlands sida Problem i äktenskap eller parförhållande, får du information om var du kan få råd vid problem i äktenskapet eller i parförhållandet.
Äldre människor
Helsingfors stads Seniorinfo ger råd om tjänster för äldre i Helsingfors.
Äldre i Helsingfors och deras anhöriga kan kontakta Seniorinfo.
Seniorinfo betjänar på finska och svenska.
Seniori-info
Tfn 09 3104 4556 (mån–fre kl. 9–15)
Seniorinfofinska _ svenska _ engelska
När du tar hand om en anhörig i hemmet
När du tar hand om en gammal eller sjuk anhörig eller en anhörig med funktionsnedsättning för att han eller hon ska kunna bo kvar i sitt hem, kan du ha rätt till stöd för närståendevård.
Du får närmare uppgifter vid social- och närarbetets verksamhetsställe i ditt bostadsområde (sosiaali- ja lähityön toimipiste).
Läs mer: Äldre människor.
Enheterna för socialt arbete och närarbetefinska _ svenska _ engelska
Stöd för närståendevårdfinska _ svenska _ engelska
InfoFinland är en mångsidig webbplats som sammanställer viktig information för personer som planerar att flytta till Finland eller som redan bor här.
Webbplatsen betjänar även myndigheter i deras flerspråkiga informationsverksamhet.
I InfoFinland hittar användaren pålitlig information på sitt eget språk om flytten till Finland, arbete, studier, boende, utbildning, hälsa, familj, problematiska situationer och fritid.
InfoFinlands webbplats är responsiv.
Sidorna är enkla att använda med olika enheter, till exempel smarttelefonen eller surfplattan.
Språken i InfoFinland
Tjänsten finns på finska, svenska, engelska, ryska, estniska, franska, somaliska, spanska, turkiska, kinesiska, persiska och arabiska. De olika språkversionerna är identiska.
Översättningarna i tjänsten görs av en översättningsbyrå.
Mer information finns på InfoFinlands sida Översättningar
Dessutom innehåller InfoFinland länkar till material som publicerats på andra språk.
Information om lokala tjänster
I InfoFinland finns information om tjänsterna i många kommuner.
Länkar till kommunsidorna hittar du med hjälp av Menyn Städer i höger spalt.
När användaren är på en kommunsida, visas länkar till den grundläggande informationen om ämnet.
På sidan Städer hittar du kommunerna som finns i InfoFinland på en karta.
Sidunderhåll
InfoFinlands webbplats upprätthålls av Helsingfors stad.
InfoFinland-redaktionen sköter uppdateringen av uppgifterna i avsnitten Flytta till Finland, Livet i Finland och Information om Finland samt uppgifterna om Helsingfors, Esbo, Vanda och Grankulla.
De övriga medlemskommunernas egna redaktioner upprätthåller sina egna kommunsidor.
Kurssökningen för kurser i finska och svenska, Finnishcourses.fi, är en del av InfoFinland.
Kurser i finska och svenska språketfinska _ engelska _ ryska
InfoFinland finansieras av staten och samarbetskommunerna.
InfoFinlands chefredaktör och ansvariga redaktör är Eija Kyllönen-Saarnio.
Historia
Webbtjänsten InfoFinland hette tidigare Infobanken.
Namnet ändrades i november 2018.
Webbtjänsten Infopankki.fi publicerades vid Helsingfors kulturcentral 2003 som ett samarbete mellan Internationella kulturcentret Caisa och Helsingfors stadsbibliotek.
Caisafinska _ svenska _ engelska
Idag drivs InfoFinland vid Helsingfors stadskanslis kommunikationsavdelning.
InfoFinland är en mångsidig webbplats som sammanställer viktig information för personer som planerar att flytta till Finland eller som redan bor här.
Webbplatsen betjänar även myndigheter i deras flerspråkiga informationsverksamhet.
I InfoFinland hittar användaren pålitlig information på sitt eget språk om flytten till Finland, arbete, studier, boende, utbildning, hälsa, familj, problematiska situationer och fritid.
InfoFinlands webbplats är responsiv.
Sidorna är enkla att använda med olika enheter, till exempel smarttelefonen eller surfplattan.
Språken i InfoFinland
Tjänsten finns på finska, svenska, engelska, ryska, estniska, franska, somaliska, spanska, turkiska, kinesiska, persiska och arabiska. De olika språkversionerna är identiska.
Översättningarna i tjänsten görs av en översättningsbyrå.
Mer information finns på InfoFinlands sida Översättningar
Dessutom innehåller InfoFinland länkar till material som publicerats på andra språk.
Information om lokala tjänster
I InfoFinland finns information om tjänsterna i många kommuner.
Länkar till kommunsidorna hittar du med hjälp av Menyn Städer i höger spalt.
När användaren är på en kommunsida, visas länkar till den grundläggande informationen om ämnet.
På sidan Städer hittar du kommunerna som finns i InfoFinland på en karta.
Sidunderhåll
InfoFinlands webbplats upprätthålls av Helsingfors stad.
InfoFinland-redaktionen sköter uppdateringen av uppgifterna i avsnitten Flytta till Finland, Livet i Finland och Information om Finland samt uppgifterna om Helsingfors, Esbo, Vanda och Grankulla.
De övriga medlemskommunernas egna redaktioner upprätthåller sina egna kommunsidor.
Kurssökningen för kurser i finska och svenska, Finnishcourses.fi, är en del av InfoFinland.
Kurser i finska och svenska språketfinska _ engelska _ ryska
InfoFinland finansieras av staten och samarbetskommunerna.
InfoFinlands chefredaktör och ansvariga redaktör är Eija Kyllönen-Saarnio.
Historia
Webbtjänsten InfoFinland hette tidigare Infobanken.
Namnet ändrades i november 2018.
Webbtjänsten Infopankki.fi publicerades vid Helsingfors kulturcentral 2003 som ett samarbete mellan Internationella kulturcentret Caisa och Helsingfors stadsbibliotek.
Caisafinska _ svenska _ engelska
Idag drivs InfoFinland vid Helsingfors stadskanslis kommunikationsavdelning.
InfoFinland är en mångsidig webbplats som sammanställer viktig information för personer som planerar att flytta till Finland eller som redan bor här.
Webbplatsen betjänar även myndigheter i deras flerspråkiga informationsverksamhet.
I InfoFinland hittar användaren pålitlig information på sitt eget språk om flytten till Finland, arbete, studier, boende, utbildning, hälsa, familj, problematiska situationer och fritid.
InfoFinlands webbplats är responsiv.
Sidorna är enkla att använda med olika enheter, till exempel smarttelefonen eller surfplattan.
Språken i InfoFinland
Tjänsten finns på finska, svenska, engelska, ryska, estniska, franska, somaliska, spanska, turkiska, kinesiska, persiska och arabiska. De olika språkversionerna är identiska.
Översättningarna i tjänsten görs av en översättningsbyrå.
Mer information finns på InfoFinlands sida Översättningar
Dessutom innehåller InfoFinland länkar till material som publicerats på andra språk.
Information om lokala tjänster
I InfoFinland finns information om tjänsterna i många kommuner.
Länkar till kommunsidorna hittar du med hjälp av Menyn Städer i höger spalt.
När användaren är på en kommunsida, visas länkar till den grundläggande informationen om ämnet.
På sidan Städer hittar du kommunerna som finns i InfoFinland på en karta.
Sidunderhåll
InfoFinlands webbplats upprätthålls av Helsingfors stad.
InfoFinland-redaktionen sköter uppdateringen av uppgifterna i avsnitten Flytta till Finland, Livet i Finland och Information om Finland samt uppgifterna om Helsingfors, Esbo, Vanda och Grankulla.
De övriga medlemskommunernas egna redaktioner upprätthåller sina egna kommunsidor.
Kurssökningen för kurser i finska och svenska, Finnishcourses.fi, är en del av InfoFinland.
Kurser i finska och svenska språketfinska _ engelska _ ryska
InfoFinland finansieras av staten och samarbetskommunerna.
InfoFinlands chefredaktör och ansvariga redaktör är Eija Kyllönen-Saarnio.
Historia
Webbtjänsten InfoFinland hette tidigare Infobanken.
Namnet ändrades i november 2018.
Webbtjänsten Infopankki.fi publicerades vid Helsingfors kulturcentral 2003 som ett samarbete mellan Internationella kulturcentret Caisa och Helsingfors stadsbibliotek.
Caisafinska _ svenska _ engelska
Idag drivs InfoFinland vid Helsingfors stadskanslis kommunikationsavdelning.
Hälsotjänsterna i Helsingfors
Barns hälsa
Äldre människors hälsa
Tandvård
Mental hälsa
Sexuell hälsa
När du väntar barn
Patientens rättigheter
Handikappade personer
I brådskande nödsituationer ska du ringa nödnumret 112.
Ring nödnumret till exempel vid allvarliga olyckor eller om någon får en sjukdomsattack.
Ring inte nödnumret om det inte är fråga om en nödsituation.
Om du har hemkommun i Helsingfors, kan du använda de offentliga hälsotjänsterna.
Offentliga hälsotjänster tillhandahålls vid hälsostationer, tandkliniker, rådgivningsbyråer och sjukhus.
Om du inte har rätt att använda de offentliga hälsotjänsterna kan du söka hjälp på en privat läkarstation.
På en privat läkarstation måste du betala samtliga kostnader själv.
Om du behöver information om hälsotjänsterna, kan du ringa hälsorådgivningen: (09) 310 100 23.
Via tjänsten kan du också fråga om anvisningar för vård av sjukdomar.
Du kan tala finska, svenska eller engelska.
Läs mer: Hälsovårdstjänster i Finland.
Hälsotjänsterna i Helsingfors
När du kontaktar hälsostationen (terveysasema), bedömer en sjukskötare först din situation.
Utgående från bedömningen kan du få en tid hos läkare, hälsovårdare eller sjukskötare.
Hälsostationerna har öppet mån–fre kl. 8.00–16.00.
Om du behöver vård under samma dag ska du kontakta hälsostationen direkt på morgonen när den öppnar.
På Helsingfors stads hälsovårdscentrals webbplats hittar du kontaktuppgifterna till hälsostationerna.
linkkiHälsorådgivning:
Information om hälsorådgivningfinska
Hälsostationerna enligt stadsdelfinska _ svenska _ engelska
Patientavgifterfinska _ svenska _ engelska
Privata hälsovårdstjänster
Du kan gå till en privat läkarstation även om du inte har rätt att använda den offentliga hälso- och sjukvården i Finland.
På en privat läkarstation måste du betala samtliga kostnader själv.
Privat läkarstationfinska _ svenska _ engelska
Privat läkarstationfinska _ svenska _ engelska
Läkemedel
Du får information om hur du köper läkemedel på InfoFinlands sida Läkemedel.
Hälsovård för papperslösa
Med papperslösa avses invandrare som inte har uppehållstillstånd eller invandrare som inte har sjukförsäkring.
I Helsingfors har papperslösa invandrare rätt att få brådskande och nödvändig vård inom de offentliga hälsovårdstjänsterna.
Personer under 18 år och gravida har rätt att få alla de hälsovårdstjänster som övriga helsingforsare får.
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärhälsovård.
Tjänsterna vid Global Clinic är avgiftsfria för kunderna.
Global Clinic anmäler inte sina kunder till polisen eller andra myndigheter.
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
Telefonnumret till Global Clinic i Helsingfors är 044 977 4547.
Samtalet besvaras av en sjukskötare eller en läkare.
E-postadressen är globalclinic.finland(snabel-a)gmail.com.
Kontaktuppgifterfinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Under kvällar och helger är hälsostationerna stängda.
Om du behöver brådskande vård på kvällen eller veckoslutet, kontakta då jourmottagningen (päivystys).
Ring den kostnadsfria Jourhjälpen på tfn 116 117 innan du kommer till jourmottagningen.
Jourhjälpen (Päivystysapu) betjänar dygnet runt.
Om du bor i östra Helsingfors, sydöstra Helsingfors, nordöstra Helsingfors eller norra Helsingfors hittar du hälsovårdscentraljouren vid Malms sjukhus.
Malms sjukhus
Talvelavägen 6, J-trappan
Tfn (09) 310 6611 / 116 117
Om du bor i södra, mellersta eller västra Helsingfors finns hälsocentralsjouren vid Haartmanska sjukhuset.
Haartmanska sjukhuset
Haartmansgatan 4
Byggnad 12
Tfn (09) 310 5018 / 116 117
Hälsocentralsjourenfinska _ svenska _ engelska
Barns hälsa
På rådgivningsbyrån (neuvola) följs hälsa och uppväxt bland barn under skolåldern.
I Helsingfors kan du bli kund hos rådgivningen om du har ett FPA-kort.
Du kan boka tid på rådgivningsbyrån via din hälsostation.
Skolhälsovårdaren tar hand om skolbarns hälsa.
Du får mer information i skolan.
Om ditt barn plötsligt blir sjukt, ta kontakt med din hälsostation.
Ring hälsostationen direkt på morgonen när den öppnar.
Hälsostationerna har öppet mån–fre kl. 8.00–16.00.
När hälsostationen är stängd, kontakta jourmottagningen på Barnsjukhuset.
På jourmottagningen vårdas endast barn som är i akut behov av hjälp.
Barnsjukhuset (Lastensairaala)
Stenbäcksgatan 9
Tfn (09) 87 100 23
Du kan även föra barnet till en privat läkarstation.
I Helsingfors finns många privata läkarstationer som även tar hand om barn.
Läs mer: Barns hälsa.
Rådgivningsbyråernas kontaktuppgifterfinska _ engelska
Skolhälsovårdfinska _ svenska _ engelska
Hälsostationerna enligt stadsdelfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
Jourpolikliniken vid Barnklinikenfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
När ett barn insjuknar - råd till föräldrarnasvenska _ engelska
Äldre människors hälsa
Äldre människor kan anlita tjänster som tillhandahålls av vanliga hälsostationer.
Därtill är det möjligt att i vissa fall få tjänster som är särskilt avsedda för äldre.
Helsingfors stads Seniorinfo ger råd om tjänster för äldre i Helsingfors.
Äldre i Helsingfors och deras anhöriga kan kontakta Seniorinfo.
Seniorinfo betjänar på finska och svenska.
Seniori-info
Tfn 09 3104 4556 (mån–fre kl. 9–15)
Läs mer:
Äldre människors hälsa.
Hälsostationerna enligt stadsdelfinska _ svenska _ engelska
Seniorinfofinska _ svenska _ engelska
När du tar hand om en anhörig i hemmet
När du tar hand om en gammal eller sjuk anhörig eller en anhörig med funktionsnedsättning för att han eller hon ska kunna bo kvar i sitt hem, kan du ha rätt till stöd för närståendevård.
Du får närmare uppgifter vid social- och närarbetets verksamhetsställe i ditt bostadsområde (sosiaali- ja lähityön toimipiste).
Läs mer: Äldre människor.
Enheterna för socialt arbete och närarbetefinska _ svenska _ engelska
Stöd för närståendevårdfinska
Tandvård
Offentlig tandvård
Tidsbeställningsnumret till tandvården i Helsingfors är (09) 310 51400.
Du kan ringa tidsbeställningen mån–fre kl. 7–15.
Om du är i akut behov av vård, ring tidsbeställningen direkt på morgonen.
Om du behöver akut hjälp av tandläkaren på kvällen eller veckoslutet, ring jouren på tfn 09 471 71110.
Information om tandvårdenfinska _ svenska _ engelska
Information om tandvårdsjourenfinska _ svenska _ engelska
Film om munhälsovårdfinska _ engelska _ somaliska _ arabiska
Privat tandvård
I Helsingfors finns det också många privata tandläkare.
Du kan besöka en privat tandläkare även om du inte har rätt att anlita tjänster inom den offentliga hälso- och sjukvården.
Privat tandvård är dyrare än offentlig tandvård.
Läs mer: Tandvård.
Mental hälsa
Om du behöver psykiatrisk vård kan du kontakta din hälsocentral.
Vid behov skriver läkaren en remiss till den psykiatriska polikliniken för dig.
Föreningen för mental hälsa i Finland (Suomen Mielenterveysseura) har en krismottagning för invandrare som bor i Helsingforsregionen.
Vid krismottagningen får du hjälp och stöd i svåra situationer.
Du kan ringa och boka tid.
Krismottagningen betjänar på finska, svenska och engelska samt på andra språk med hjälp av tolk.
Boka tid per telefon på nummer (09) 413 50 510.
Läs mer: Mental hälsa.
Mentalvårdstjänsterfinska _ svenska _ engelska
Filmklipp om tjänster inom mental hälsafinska _ engelska _ somaliska _ arabiska
linkkiFöreningen för mental hälsa i Finland:
Krismottagningfinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Sexuell hälsa
Om du behöver ett recept för preventivmedel eller om du överväger abort, ta kontakt med din hälsostation (terveysasema).
Om du är under 16 år och behöver preventivmedel, ta kontakt med hälsovårdaren vid din läroinrättning.
Om du misstänker att du har en könssjukdom, men har inga symtom, ska du kontakta din hälsostation.
Om du har symtom kan du utan remiss besöka Helsingfors poliklinik för könssjukdomar mån–fre kl. 8–12.
Adressen är Mejlansvägen 2.
Läs mer: Sexuell hälsa.
Hälsostationerna enligt stadsdelfinska _ svenska _ engelska
Preventivrådgivningfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Polikliniken för könssjukdomarfinska _ svenska _ engelska
När du väntar barn
På rådgivningen (äitiysneuvola) följer man moderns, barnets och hela familjens välmående under graviditeten.
Kontakta rådgivningsbyrån i ditt område genast när du upptäcker att du väntar barn.
Förlossningssjukhusen i Helsingforsregionen är Kvinnokliniken (Helsingfors) och Jorv sjukhus (Esbo).
Du hittar kontaktuppgifterna på HNS webbplats.
Läs mer: När du väntar barn.
Rådgivningsbyråernas kontaktuppgifterfinska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Förlossningfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Patientens rättigheter
Om du upplever att du behandlats fel inom hälsovårdstjänsterna ska du först reda ut situationen vid din egen vårdenhet.
Om situationen inte löser sig, kontakta överläkaren eller överskötaren vid vårdenheten.
Därefter kan du vid behov kontakta patientombudsmannen (potilasasiamies).
Patientombudsmannens verksamhetfinska _ svenska _ engelska
Handikappade personer
Helsingfors stad ordnar tjänster för personer med funktionsnedsättning, till exempel hjälpmedel, färdtjänst och dagverksamhet.
Även barn med funktionsnedsättning kan få tjänster för personer med funktionsnedsättning.
Om du har en funktionsnedsättning, ta då först kontakt med hälsostationen (terveysasema).
På hälsostationen bedöms din situation.
Närmare information om tjänster för personer med funktionsnedsättning i Helsingfors får du av socialarbetarna vid stadens tjänster för personer med funktionsnedsättning.
Läs mer: Handikappade personer.
Läs mer: Ett handikappat barn.
Tjänster för handikappadefinska
Verksamhetsställen för handikappservicefinska
Hälsotjänsterna i Helsingfors
Barns hälsa
Tandvård
Mental hälsa
Sexuell hälsa och prevention
Graviditet och förlossning
Patientens rättigheter
Handikappade personer
I brådskande nödsituationer ska du ringa nödnumret 112.
Ring nödnumret till exempel vid allvarliga olyckor eller om någon får en sjukdomsattack.
Ring inte nödnumret om det inte är fråga om en nödsituation.
Om du har hemkommun i Helsingfors, kan du använda de offentliga hälsotjänsterna.
Offentliga hälsotjänster tillhandahålls vid hälsostationer, tandkliniker, rådgivningsbyråer och sjukhus.
Om du inte har rätt att använda de offentliga hälsotjänsterna kan du söka hjälp på en privat läkarstation.
På en privat läkarstation måste du betala samtliga kostnader själv.
Om du behöver information om hälsotjänsterna, kan du ringa hälsorådgivningen: (09) 310 100 23.
Via tjänsten kan du också fråga om anvisningar för vård av sjukdomar.
Du kan tala finska, svenska eller engelska.
Läs mer: Hälsovårdstjänster i Finland.
Hälsotjänsterna i Helsingfors
När du kontaktar hälsostationen (terveysasema), bedömer en sjukskötare först din situation.
Utgående från bedömningen kan du få en tid hos läkare, hälsovårdare eller sjukskötare.
Hälsostationerna har öppet mån–fre kl. 8.00–16.00.
Om du behöver vård under samma dag ska du kontakta hälsostationen direkt på morgonen när den öppnar.
På Helsingfors stads hälsovårdscentrals webbplats hittar du kontaktuppgifterna till hälsostationerna.
linkkiHälsorådgivning:
Information om hälsorådgivningfinska
Hälsostationerna enligt stadsdelfinska _ svenska _ engelska
Patientavgifterfinska _ svenska _ engelska
Privata hälsovårdstjänster
Du kan gå till en privat läkarstation även om du inte har rätt att använda den offentliga hälso- och sjukvården i Finland.
På en privat läkarstation måste du betala samtliga kostnader själv.
Privat läkarstationfinska _ svenska _ engelska
Privat läkarstationfinska _ svenska _ engelska
Läkemedel
Du får information om hur du köper läkemedel på InfoFinlands sida Läkemedel.
Hälsovård för papperslösa
Med papperslösa avses invandrare som inte har uppehållstillstånd eller invandrare som inte har sjukförsäkring.
I Helsingfors har papperslösa invandrare rätt att få brådskande och nödvändig vård inom de offentliga hälsovårdstjänsterna.
Personer under 18 år och gravida har rätt att få alla de hälsovårdstjänster som övriga helsingforsare får.
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärhälsovård.
Tjänsterna vid Global Clinic är avgiftsfria för kunderna.
Global Clinic anmäler inte sina kunder till polisen eller andra myndigheter.
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
Telefonnumret till Global Clinic i Helsingfors är 044 977 4547.
Samtalet besvaras av en sjukskötare eller en läkare.
E-postadressen är globalclinic.finland(snabel-a)gmail.com.
Kontaktuppgifterfinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Under kvällar och helger är hälsostationerna stängda.
Om du behöver brådskande vård på kvällen eller veckoslutet, kontakta då jourmottagningen (päivystys).
Ring den kostnadsfria Jourhjälpen på tfn 116 117 innan du kommer till jourmottagningen.
Jourhjälpen (Päivystysapu) betjänar dygnet runt.
Om du bor i östra Helsingfors, sydöstra Helsingfors, nordöstra Helsingfors eller norra Helsingfors hittar du hälsovårdscentraljouren vid Malms sjukhus.
Malms sjukhus
Talvelavägen 6, J-trappan
Tfn (09) 310 6611 / 116 117
Om du bor i södra, mellersta eller västra Helsingfors finns hälsocentralsjouren vid Haartmanska sjukhuset.
Haartmanska sjukhuset
Haartmansgatan 4
Byggnad 12
Tfn (09) 310 5018 / 116 117
Hälsocentralsjourenfinska _ svenska _ engelska
Barns hälsa
På rådgivningsbyrån (neuvola) följs hälsa och uppväxt bland barn under skolåldern.
I Helsingfors kan du bli kund hos rådgivningen om du har ett FPA-kort.
Du kan boka tid på rådgivningsbyrån via din hälsostation.
Skolhälsovårdaren tar hand om skolbarns hälsa.
Du får mer information i skolan.
Om ditt barn plötsligt blir sjukt, ta kontakt med din hälsostation.
Ring hälsostationen direkt på morgonen när den öppnar.
Hälsostationerna har öppet mån–fre kl. 8.00–16.00.
När hälsostationen är stängd, kontakta jourmottagningen på Barnsjukhuset.
På jourmottagningen vårdas endast barn som är i akut behov av hjälp.
Barnsjukhuset (Lastensairaala)
Stenbäcksgatan 9
Tfn (09) 87 100 23
Du kan även föra barnet till en privat läkarstation.
I Helsingfors finns många privata läkarstationer som även tar hand om barn.
Läs mer: Barns hälsa.
Rådgivningsbyråernas kontaktuppgifterfinska _ engelska
Skolhälsovårdfinska _ svenska _ engelska
Hälsostationerna enligt stadsdelfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
Jourpolikliniken vid Barnklinikenfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
När ett barn insjuknar - råd till föräldrarnasvenska _ engelska
Tandvård
Offentlig tandvård
Tidsbeställningsnumret till tandvården i Helsingfors är (09) 310 51400.
Du kan ringa tidsbeställningen mån–fre kl. 7–15.
Om du är i akut behov av vård, ring tidsbeställningen direkt på morgonen.
Om du behöver akut hjälp av tandläkaren på kvällen eller veckoslutet, ring jouren på tfn 09 471 71110.
Information om tandvårdenfinska _ svenska _ engelska
Information om tandvårdsjourenfinska _ svenska _ engelska
Film om munhälsovårdfinska _ engelska _ somaliska _ arabiska
Privat tandvård
I Helsingfors finns det också många privata tandläkare.
Du kan besöka en privat tandläkare även om du inte har rätt att anlita tjänster inom den offentliga hälso- och sjukvården.
Privat tandvård är dyrare än offentlig tandvård.
Läs mer: Tandvård.
Mental hälsa
Om du behöver psykiatrisk vård kan du kontakta din hälsocentral.
Vid behov skriver läkaren en remiss till den psykiatriska polikliniken för dig.
Föreningen för mental hälsa i Finland (Suomen Mielenterveysseura) har en krismottagning för invandrare som bor i Helsingforsregionen.
Vid krismottagningen får du hjälp och stöd i svåra situationer.
Du kan ringa och boka tid.
Krismottagningen betjänar på finska, svenska och engelska samt på andra språk med hjälp av tolk.
Boka tid per telefon på nummer (09) 413 50 510.
Läs mer: Mental hälsa.
Mentalvårdstjänsterfinska _ svenska _ engelska
Filmklipp om tjänster inom mental hälsafinska _ engelska _ somaliska _ arabiska
linkkiFöreningen för mental hälsa i Finland:
Krismottagningfinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Sexuell hälsa och prevention
Om du behöver ett recept för preventivmedel eller om du överväger abort, ta kontakt med din hälsostation (terveysasema).
Om du är under 16 år och behöver preventivmedel, ta kontakt med hälsovårdaren vid din läroinrättning.
Om du misstänker att du har en könssjukdom, men har inga symtom, ska du kontakta din hälsostation.
Om du har symtom kan du utan remiss besöka Helsingfors poliklinik för könssjukdomar mån–fre kl. 8–12.
Adressen är Mejlansvägen 2.
Läs mer: Sexuell hälsa och prevention.
Preventivrådgivningfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Polikliniken för könssjukdomarfinska _ svenska _ engelska
Graviditet och förlossning
På rådgivningen (äitiysneuvola) följer man moderns, barnets och hela familjens välmående under graviditeten.
Kontakta rådgivningsbyrån i ditt område genast när du upptäcker att du väntar barn.
Förlossningssjukhusen i Helsingforsregionen är Kvinnokliniken (Helsingfors) och Jorv sjukhus (Esbo).
Du hittar kontaktuppgifterna på HNS webbplats.
Läs mer: Graviditet och förlossning och När ett barn föds i Finland.
Rådgivningsbyråernas kontaktuppgifterfinska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Förlossningfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Patientens rättigheter
Om du upplever att du behandlats fel inom hälsovårdstjänsterna ska du först reda ut situationen vid din egen vårdenhet.
Om situationen inte löser sig, kontakta överläkaren eller överskötaren vid vårdenheten.
Därefter kan du vid behov kontakta patientombudsmannen (potilasasiamies).
Patientombudsmannens verksamhetfinska _ svenska _ engelska
Handikappade personer
Helsingfors stad ordnar tjänster för personer med funktionsnedsättning, till exempel hjälpmedel, färdtjänst och dagverksamhet.
Även barn med funktionsnedsättning kan få tjänster för personer med funktionsnedsättning.
Om du har en funktionsnedsättning, ta då först kontakt med hälsostationen (terveysasema).
På hälsostationen bedöms din situation.
Närmare information om tjänster för personer med funktionsnedsättning i Helsingfors får du av socialarbetarna vid stadens tjänster för personer med funktionsnedsättning.
Läs mer: Handikappade personer.
Läs mer: Ett handikappat barn.
Tjänster för handikappadefinska
Verksamhetsställen för handikappservicefinska _ engelska
Hälsotjänsterna i Helsingfors
Barns hälsa
Tandvård
Mental hälsa
Sexuell hälsa och prevention
Graviditet och förlossning
Patientens rättigheter
Handikappade personer
I brådskande nödsituationer ska du ringa nödnumret 112.
Ring nödnumret till exempel vid allvarliga olyckor eller om någon får en sjukdomsattack.
Ring inte nödnumret om det inte är fråga om en nödsituation.
Om du har hemkommun i Helsingfors, kan du använda de offentliga hälsotjänsterna.
Offentliga hälsotjänster tillhandahålls vid hälsostationer, tandkliniker, rådgivningsbyråer och sjukhus.
Om du inte har rätt att använda de offentliga hälsotjänsterna kan du söka hjälp på en privat läkarstation.
På en privat läkarstation måste du betala samtliga kostnader själv.
Om du behöver information om hälsotjänsterna, kan du ringa hälsorådgivningen: (09) 310 100 23.
Via tjänsten kan du också fråga om anvisningar för vård av sjukdomar.
Du kan tala finska, svenska eller engelska.
Läs mer: Hälsovårdstjänster i Finland.
Hälsotjänsterna i Helsingfors
När du kontaktar hälsostationen (terveysasema), bedömer en sjukskötare först din situation.
Utgående från bedömningen kan du få en tid hos läkare, hälsovårdare eller sjukskötare.
Hälsostationerna har öppet mån–fre kl. 8.00–16.00.
Om du behöver vård under samma dag ska du kontakta hälsostationen direkt på morgonen när den öppnar.
På Helsingfors stads hälsovårdscentrals webbplats hittar du kontaktuppgifterna till hälsostationerna.
linkkiHälsorådgivning:
Information om hälsorådgivningfinska _ svenska _ engelska
Hälsostationerna enligt stadsdelfinska _ svenska _ engelska
Patientavgifterfinska _ svenska _ engelska
Privata hälsovårdstjänster
Du kan gå till en privat läkarstation även om du inte har rätt att använda den offentliga hälso- och sjukvården i Finland.
På en privat läkarstation måste du betala samtliga kostnader själv.
Privat läkarstationfinska _ svenska _ engelska
Privat läkarstationfinska _ svenska _ engelska
Läkemedel
Du får information om hur du köper läkemedel på InfoFinlands sida Läkemedel.
Hälsovård för papperslösa
Med papperslösa avses invandrare som inte har uppehållstillstånd eller invandrare som inte har sjukförsäkring.
I Helsingfors har papperslösa invandrare rätt att få brådskande och nödvändig vård inom de offentliga hälsovårdstjänsterna.
Personer under 18 år och gravida har rätt att få alla de hälsovårdstjänster som övriga helsingforsare får.
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärhälsovård.
Tjänsterna vid Global Clinic är avgiftsfria för kunderna.
Global Clinic anmäler inte sina kunder till polisen eller andra myndigheter.
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
Telefonnumret till Global Clinic i Helsingfors är 044 977 4547.
Samtalet besvaras av en sjukskötare eller en läkare.
E-postadressen är globalclinic.finland(snabel-a)gmail.com.
Kontaktuppgifterfinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Under kvällar och helger är hälsostationerna stängda.
Om du behöver brådskande vård på kvällen eller veckoslutet, kontakta då jourmottagningen (päivystys).
Ring den kostnadsfria Jourhjälpen på tfn 116 117 innan du kommer till jourmottagningen.
Jourhjälpen (Päivystysapu) betjänar dygnet runt.
Om du bor i östra Helsingfors, sydöstra Helsingfors, nordöstra Helsingfors eller norra Helsingfors hittar du hälsovårdscentraljouren vid Malms sjukhus.
Malms sjukhus
Talvelavägen 6, J-trappan
Tfn (09) 310 6611 / 116 117
Om du bor i södra, mellersta eller västra Helsingfors finns hälsocentralsjouren vid Haartmanska sjukhuset.
Haartmanska sjukhuset
Haartmansgatan 4
Byggnad 12
Tfn (09) 310 5018 / 116 117
Hälsocentralsjourenfinska _ svenska _ engelska
Barns hälsa
På rådgivningsbyrån (neuvola) följs hälsa och uppväxt bland barn under skolåldern.
I Helsingfors kan du bli kund hos rådgivningen om du har ett FPA-kort.
Du kan boka tid på rådgivningsbyrån via din hälsostation.
Skolhälsovårdaren tar hand om skolbarns hälsa.
Du får mer information i skolan.
Om ditt barn plötsligt blir sjukt, ta kontakt med din hälsostation.
Ring hälsostationen direkt på morgonen när den öppnar.
Hälsostationerna har öppet mån–fre kl. 8.00–16.00.
När hälsostationen är stängd, kontakta jourmottagningen på Barnsjukhuset.
På jourmottagningen vårdas endast barn som är i akut behov av hjälp.
Nya barnsjukhuset (Uusi lastensairaala)
Stenbäcksgatan 9
Tfn (09) 87 100 23
Du kan även föra barnet till en privat läkarstation.
I Helsingfors finns många privata läkarstationer som även tar hand om barn.
Läs mer: Barns hälsa.
Rådgivningsbyråernas kontaktuppgifterfinska _ engelska
Skolhälsovårdfinska _ svenska _ engelska
Hälsostationerna enligt stadsdelfinska _ svenska _ engelska
linkkiHUS (Helsingfors och Nylands sjukvårdsdistrikt):
Barnjour i Helsingforsfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
När ett barn insjuknar - råd till föräldrarnafinska _ svenska _ engelska
Tandvård
Offentlig tandvård
Tidsbeställningsnumret till tandvården i Helsingfors är (09) 310 51400.
Du kan ringa tidsbeställningen mån–fre kl. 7–15.
Om du är i akut behov av vård, ring tidsbeställningen direkt på morgonen.
Om du behöver akut hjälp av tandläkaren på kvällen eller veckoslutet, ring jouren på tfn 09 471 71110.
Information om tandvårdenfinska _ svenska _ engelska
Information om tandvårdsjourenfinska _ svenska _ engelska
Film om munhälsovårdfinska _ engelska _ somaliska _ arabiska
Privat tandvård
I Helsingfors finns det också många privata tandläkare.
Du kan besöka en privat tandläkare även om du inte har rätt att anlita tjänster inom den offentliga hälso- och sjukvården.
Privat tandvård är dyrare än offentlig tandvård.
Läs mer: Tandvård.
Mental hälsa
Om du behöver psykiatrisk vård kan du kontakta din hälsocentral.
Vid behov skriver läkaren en remiss till den psykiatriska polikliniken för dig.
Föreningen för mental hälsa i Finland (Suomen Mielenterveysseura) har en krismottagning för invandrare som bor i Helsingforsregionen.
Vid krismottagningen får du hjälp och stöd i svåra situationer.
Du kan ringa och boka tid.
Krismottagningen betjänar på finska, svenska och engelska samt på andra språk med hjälp av tolk.
Boka tid per telefon på nummer (09) 413 50 510.
Läs mer: Mental hälsa.
Mentalvårdstjänsterfinska _ svenska _ engelska
Filmklipp om tjänster inom mental hälsafinska _ engelska _ somaliska _ arabiska
linkkiMIELI Psykisk Hälsa Finland rf:
Krismottagningfinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Sexuell hälsa och prevention
Om du behöver ett recept för preventivmedel eller om du överväger abort, ta kontakt med din hälsostation (terveysasema).
Om du är under 16 år och behöver preventivmedel, ta kontakt med hälsovårdaren vid din läroinrättning.
Om du misstänker att du har en könssjukdom, men har inga symtom, ska du kontakta din hälsostation.
Om du har symtom kan du utan remiss besöka Helsingfors poliklinik för könssjukdomar mån–fre kl. 8–12.
Adressen är Mejlansvägen 2.
Läs mer: Sexuell hälsa och prevention.
Preventivrådgivningfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Polikliniken för könssjukdomarfinska _ svenska _ engelska
Graviditet och förlossning
På rådgivningen (äitiysneuvola) följer man moderns, barnets och hela familjens välmående under graviditeten.
Kontakta rådgivningsbyrån i ditt område genast när du upptäcker att du väntar barn.
Förlossningssjukhusen i Helsingforsregionen är Kvinnokliniken (Helsingfors) och Jorv sjukhus (Esbo).
Du hittar kontaktuppgifterna på HNS webbplats.
Läs mer: Graviditet och förlossning och När ett barn föds i Finland.
Rådgivningsbyråernas kontaktuppgifterfinska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Förlossningfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Patientens rättigheter
Om du upplever att du behandlats fel inom hälsovårdstjänsterna ska du först reda ut situationen vid din egen vårdenhet.
Om situationen inte löser sig, kontakta överläkaren eller överskötaren vid vårdenheten.
Därefter kan du vid behov kontakta patientombudsmannen (potilasasiamies).
Patientombudsmannens verksamhetfinska _ svenska _ engelska
Handikappade personer
Helsingfors stad ordnar tjänster för personer med funktionsnedsättning, till exempel hjälpmedel, färdtjänst och dagverksamhet.
Även barn med funktionsnedsättning kan få tjänster för personer med funktionsnedsättning.
Om du har en funktionsnedsättning, ta då först kontakt med hälsostationen (terveysasema).
På hälsostationen bedöms din situation.
Närmare information om tjänster för personer med funktionsnedsättning i Helsingfors får du av socialarbetarna vid stadens tjänster för personer med funktionsnedsättning.
Läs mer: Handikappade personer.
Läs mer: Ett handikappat barn.
Tjänster för handikappadefinska _ svenska _ engelska
Verksamhetsställen för handikappservicefinska _ svenska _ engelska
Dagvård
Förskoleundervisning
Grundläggande undervisning
Eftermiddagsverksamhet för skolbarn
Modersmålsundervisning för invandrare
Yrkesubildning
Gymnasium
Stöd och handledning för unga
Högskoleutbildning
Andra studiemöjligheter
Dagvård
I Helsingfors finns det flera daghem som drivs av staden och privata daghem.
Stadens daghem är finsk- eller svenskspråkiga.
De flesta är finskspråkiga.
Om du ansöker om en dagvårdsplats i stadens daghem, ska du skicka in din ansökan minst fyra månader före dagvårdsstart.
Du kan ansöka om dagvårdsplats vid staden om familjen har sin adress i Helsingfors.
Ansök om dagvårdsplats på Internet.
När du använder den elektroniska blanketten behöver du finländska nätbankkoder.
Dessutom ska ditt barn ha en finländsk personbeteckning.
Om du inte kan använda den elektroniska blanketten kan du skriva ut ansökningsblanketten på stadens webbplats.
Lämna eller posta blanketten till den dagvårdsenhet där du i första hand söker plats.
Du hittar kontaktuppgifterna till daghemmen på stadens webbplats.
Om du har frågor kring dagvården eller om ansökning av dagvårdsplats, kan du ringa rådgivningstelefonen vid stadens tjänster inom småbarnspedagogiken:
Tfn 09 310 44986 (betjänar även på engelska)
I Helsingfors finns även privata daghem vars verksamhetsspråk är engelska, ryska, tyska, franska eller spanska.
I Helsingfors finns även ett muslimskt daghem vars verksamhetsspråk är arabiska.
Om du ansöker om en plats i ett privat daghem, kontakta direkt det daghem som är föremål för platsansökan.
Läs mer: Dagvård.
Dagvård i Helsingforsfinska _ svenska _ engelska
Daghem med vård på främmande språkfinska _ svenska _ engelska
Ansökan om dagvårdsplatsfinska _ svenska _ engelska
Dagvårdsavgifterfinska _ svenska _ engelska
Förskoleundervisning
I Helsingfors ordnas förskoleundervisning (esiopetus) i många daghem och skolor.
På Helsingfors stads webbplats hittar du en lista över de daghem och skolor som ger förskoleundervisning.
Man ansöker till förskoleundervisningen med en elektronisk blankett.
När du använder den elektroniska blanketten behöver du finländska nätbankkoder.
Dessutom ska ditt barn ha en finländsk personbeteckning.
Om du inte kan använda den elektroniska blanketten ska du skriva ut ansökningsblanketten från stadens webbplats eller hämta den vid ett av stadens daghem.
Lämna eller posta blanketten till den dagvårdsenhet där du i första hand söker plats.
Du hittar mer information om förskoleundervisningen på stadens webbplats.
Du kan även fråga om mer information av daghemsföreståndarna.
Förskoleundervisningen börjar i augusti och ansökningstiden är i januari.
Läs mer: Förskoleundervisning.
Daghem som ger förskoleundervisningfinska _ svenska _ engelska
Ansökan till förskoleundervisningfinska _ svenska _ engelska
Förskoleundervisning i Helsingforsfinska _ svenska _ engelska
Grundläggande undervisning
I Helsingfors finns flera grundskolor (peruskoulu).
Utöver stadens egna skolor finns det privata skolor och statliga skolor i Helsingfors.
Studier vid en privat skola kan vara avgiftsbelagda.
I stadens skolor är undervisningsspråket finska eller svenska.
I Helsingfors finns det också privata skolor med undervisning på t.ex. engelska, tyska, franska eller ryska.
Anmälan till grundskolan sker i början av året.
Du kan anmäla ditt barn till skolan via Internet eller genom att besöka skolan på anmälningsdagen.
Helsingfors stads webbsidor ger dig information om anmälningsdagen.
Om barnet inte har tillräckligt bra kunskaper för att klara grundskolan kan han eller hon få förberedande undervisning.
Den förberedande undervisningen förbereder barnet inför grundskolan.
I den förberedande undervisningen ges undervisning i finska och i grundskolans ämnen.
Du kan fråga om den grundläggande utbildningen och om skolorna i Helsingfors vid rådgivningen och kundtjänsten vid sektorn för fostran och utbildning.
Kontaktuppgifter:
Töysägatan 2D
Tfn (09) 310 86400
Vid Helsingfors vuxengymnasium finns en linje avsedd för invandrare över 17 år, där du kan avlägga hela eller en del av den grundläggande utbildningen.
Mer information finns på Helsingfors vuxengymnasiums webbplats.
Också andra vuxengymnasier ger grundläggande utbildning för vuxna.
Kontaktuppgifterna till vuxengymnasierna finns på Helsingfors stads webbplats.
Grundläggande utbildning.
Broschyren Information om den finska grundskolanengelska _ ryska _ franska _ somaliska _ arabiska
Skolornas kontaktuppgifterfinska _ svenska _ engelska
Mer information om anmälanfinska _ svenska _ engelska
Internationella skolor i huvudstadsregionenfinska
linkkiExpatFinland.fi:
Internationella skolor i huvudstadsregionenengelska
linkkiHelsingfors Vuxengymnasium:
Grundläggande utbildning för vuxna invandrarefinska
Grundläggande utbildning för vuxna invandrarefinska _ engelska
Eftermiddagsverksamhet för skolbarn
Helsingfors stad ordnar eftermiddagsverksamhet för barn i årskurs 1 och 2 i skolor och lekparker efter skoldagen.
Eftermiddagsverksamhet ordnas under läsåret på vardagar högst fram till klockan 17.00.
Verksamheten i lekparkerna är avgiftsfri och öppen för alla.
Du kan anmäla ditt barn till lekparkernas eftermiddagsverksamhet med en anmälningsblankett.
Lämna blanketten till den lekpark som anmälan i första hand gäller.
Lekparks- och eftermiddagsverksamhet för skolbarnfinska _ ryska _ somaliska _ arabiska
Anvisningar om eftermiddagsverksamhetens klientavgiftfinska _ ryska _ somaliska _ arabiska
Modersmålsundervisning för invandrare
Barn som har ett annat modersmål än finska eller svenska kan få modersmålsundervisning.
I Helsingfors ges modersmålsundervisning för invandrare på fler än 40 språk.
Du får information om modersmålsundervisningen vid rådgivningen och kundtjänsten vid sektorn för fostran och utbildning.
rådgivningen och kundtjänsten vid sektorn för fostran och utbildning:
Töysägatan 2D
Tfn (09) 310 86400
Yrkesutbildning
Stadin ammattiopisto är Finlands största yrkesläroanstalt där man kan utbilda sig inom många olika branscher.
I Helsingfors finns även andra yrkesläroanstalter.
Man söker till yrkesutbildning i den gemensamma ansökan.
Vid Stadin ammattiopisto ordnas förberedande utbildning inför yrkesutbildning för invandrare.
Den förberedande utbildningen är avsedd för ungdomar och vuxna som är intresserade av yrkesutbildning och vill förbättra sina kunskaper i finska.
Den förberedande undervisningen pågår i en termin eller ett läsår.
Information om den förberedande utbildningen får du vid rådgivningen och kundtjänsten vid sektorn för fostran och utbildning eller vid Stadin ammattiopisto.
rådgivningen och kundtjänsten vid sektorn för fostran och utbildning:
Töysägatan 2D
Tfn (09) 310 86400
Läs mer: Yrkesutbildning, Förberedande utbildning före yrkesutbildning.
Yrkesinriktad utbildningfinska
Yrkesläroanstalterfinska _ svenska _ engelska
För yrkesutbildning förberedande undervisningfinska _ svenska _ engelska
Gymnasium
I Helsingfors finns många gymnasieskolor.
I Helsingfors finns även några sådana gymnasieskolor där undervisningsspråket är något annat än finska eller svenska.
Utöver dagsgymnasierna som är avsedda för ungdomar finns det tre vuxengymnasier (aikuislukio) i Helsingfors.
I Helsingfors arrangeras förberedande utbildning för gymnasiet för invandrare.
Den förberedande utbildningen tar ett läsår och ger beredskap för gymnasiestudier.
Den förberedande utbildningen är avsedd för unga och vuxna som vill studera vid gymnasium men saknar tillräckliga språkkunskaper för gymnasiestudier.
Information om den förberedande utbildningen får du vid rådgivningen och kundtjänsten vid sektorn för fostran och utbildning.
rådgivningen och kundtjänsten vid sektorn för fostran och utbildning:
Töysägatan 2D
Tfn (09) 310 86400
Läs mer: Gymnasium
Gymnasier i Helsingforsfinska _ svenska _ engelska
Gymnasieansökanfinska _ svenska _ engelska
För gymnasium förberedande undervisningfinska _ engelska
Stöd och handledning för unga
Om du är under 30 år gammal kan du få råd och handledning via Ohjaamo-tjänsten.
Ohjaamos personal hjälper dig om du inte har ett arbete eller en studieplats.
Du kan även fråga om andra saker, som till exempel boende eller ekonomiska frågor.
Kontaktuppgifter:
Fredrikinkatu 48
Tfn: 040 70 46 818
Rådgivning för ungafinska
Högskoleutbildning
I Helsingfors kan du avlägga högskolestudier i många branscher.
I Helsingfors finns såväl universitet som yrkeshögskolor.
Största delen av undervisningen på högskolorna ges på finska.
I nästan alla högskolor erbjuds dock även undervisning på engelska.
I Helsingfors finns ett svenskspråkigt universitet och en svenskspråkig yrkeshögskola.
Kontaktuppgifterna till högskolorna finns på Helsingfors stads webbplats.
Anvisningar om ansökning och närmare information om utbildningsprogrammen finns på högskolornas egna webbplatser.
Läs mer: Universitet och Yrkeshögskolor.
Yrkeshögskolorfinska _ svenska _ engelska
Universitetfinska _ svenska _ engelska
Andra studiemöjligheter
I Helsingfors finns många studiemöjligheter som är öppna för alla.
Dessa studier är vanligtvis avgiftsbelagda.
Det är möjligt att avlägga högskolestudier vid öppna universitet och öppna yrkeshögskolor.
Vem som helst kan studera vid dessa.
Det öppna universitetet och de öppna yrkeshögskolorna har ett brett utbud av kurser också på engelska.
Helsingfors stad har ett finskspråkigt arbetarinstitut och ett svenskspråkigt arbetarinstitut.
Vid arbetarinstituten kan du studera t.ex. språk, handarbete och musik.
Studieutbudet är väldigt mångsidigt.
Största delen av arbetarinstitutens kurser går på finska eller svenska.
Arbetarinstituten ordnar kurser också på engelska och ryska.
Läs mer: Studier som hobby.
Finska arbetarinstitutetfinska
Kurser för invandrareengelska _ ryska
Information om öppna universitetetfinska _ svenska
Information om öppna yrkeshögskolanfinska _ svenska
Dagvård
Förskoleundervisning
Grundläggande undervisning
Eftermiddagsverksamhet för skolbarn
Modersmålsundervisning för invandrare
Yrkesubildning
Gymnasium
Stöd och handledning för unga
Högskoleutbildning
Andra studiemöjligheter
Dagvård
I Helsingfors finns det flera daghem som drivs av staden och privata daghem.
Stadens daghem är finsk- eller svenskspråkiga.
De flesta är finskspråkiga.
Om du ansöker om en dagvårdsplats i stadens daghem, ska du skicka in din ansökan minst fyra månader före dagvårdsstart.
Du kan ansöka om dagvårdsplats vid staden om familjen har sin adress i Helsingfors.
Ansök om dagvårdsplats på Internet.
När du använder den elektroniska blanketten behöver du finländska nätbankkoder.
Dessutom ska ditt barn ha en finländsk personbeteckning.
Om du inte kan använda den elektroniska blanketten kan du skriva ut ansökningsblanketten på stadens webbplats.
Lämna eller posta blanketten till den dagvårdsenhet där du i första hand söker plats.
Du hittar kontaktuppgifterna till daghemmen på stadens webbplats.
Om du har frågor kring dagvården eller om ansökning av dagvårdsplats, kan du ringa rådgivningstelefonen vid stadens tjänster inom småbarnspedagogiken:
Tfn 09 310 44986 (betjänar även på engelska)
I Helsingfors finns även privata daghem vars verksamhetsspråk är engelska, ryska, tyska, franska eller spanska.
I Helsingfors finns även ett muslimskt daghem vars verksamhetsspråk är arabiska.
Om du ansöker om en plats i ett privat daghem, kontakta direkt det daghem som är föremål för platsansökan.
Läs mer: Dagvård.
Dagvård i Helsingforsfinska _ svenska _ engelska
Daghem med vård på främmande språkfinska _ svenska _ engelska
Ansökan om dagvårdsplatsfinska _ svenska _ engelska
Dagvårdsavgifterfinska _ svenska _ engelska
Förskoleundervisning
I Helsingfors ordnas förskoleundervisning (esiopetus) i många daghem och skolor.
På Helsingfors stads webbplats hittar du en lista över de daghem och skolor som ger förskoleundervisning.
Man ansöker till förskoleundervisningen med en elektronisk blankett.
När du använder den elektroniska blanketten behöver du finländska nätbankkoder.
Dessutom ska ditt barn ha en finländsk personbeteckning.
Om du inte kan använda den elektroniska blanketten ska du skriva ut ansökningsblanketten från stadens webbplats eller hämta den vid ett av stadens daghem.
Lämna eller posta blanketten till den dagvårdsenhet där du i första hand söker plats.
Du hittar mer information om förskoleundervisningen på stadens webbplats.
Du kan även fråga om mer information av daghemsföreståndarna.
Förskoleundervisningen börjar i augusti och ansökningstiden är i januari.
Läs mer: Förskoleundervisning.
Daghem som ger förskoleundervisningfinska _ svenska _ engelska
Ansökan till förskoleundervisningfinska _ svenska _ engelska
Förskoleundervisning i Helsingforsfinska _ svenska _ engelska
Grundläggande undervisning
I Helsingfors finns flera grundskolor (peruskoulu).
Utöver stadens egna skolor finns det privata skolor och statliga skolor i Helsingfors.
Studier vid en privat skola kan vara avgiftsbelagda.
I stadens skolor är undervisningsspråket finska eller svenska.
I Helsingfors finns det också privata skolor med undervisning på t.ex. engelska, tyska, franska eller ryska.
Anmälan till grundskolan sker i början av året.
Du kan anmäla ditt barn till skolan via Internet eller genom att besöka skolan på anmälningsdagen.
Helsingfors stads webbsidor ger dig information om anmälningsdagen.
Om barnet inte har tillräckligt bra kunskaper för att klara grundskolan kan han eller hon få förberedande undervisning.
Den förberedande undervisningen förbereder barnet inför grundskolan.
I den förberedande undervisningen ges undervisning i finska och i grundskolans ämnen.
Du kan fråga om den grundläggande utbildningen och om skolorna i Helsingfors vid rådgivningen och kundtjänsten vid sektorn för fostran och utbildning.
Kontaktuppgifter:
Töysägatan 2D
Tfn (09) 310 86400
Vid Helsingfors vuxengymnasium finns en linje avsedd för invandrare över 17 år, där du kan avlägga hela eller en del av den grundläggande utbildningen.
Mer information finns på Helsingfors vuxengymnasiums webbplats.
Också andra vuxengymnasier ger grundläggande utbildning för vuxna.
Kontaktuppgifterna till vuxengymnasierna finns på Helsingfors stads webbplats.
Grundläggande utbildning.
Broschyren Information om den finska grundskolanengelska _ ryska _ franska _ somaliska _ arabiska
Skolornas kontaktuppgifterfinska _ svenska _ engelska
Mer information om anmälanfinska _ svenska _ engelska
Internationella skolor i huvudstadsregionenfinska
linkkiExpatFinland.fi:
Internationella skolor i huvudstadsregionenengelska
linkkiHelsingfors Vuxengymnasium:
Grundläggande utbildning för vuxna invandrarefinska
Grundläggande utbildning för vuxna invandrarefinska _ engelska
Eftermiddagsverksamhet för skolbarn
Helsingfors stad ordnar eftermiddagsverksamhet för barn i årskurs 1 och 2 i skolor och lekparker efter skoldagen.
Eftermiddagsverksamhet ordnas under läsåret på vardagar högst fram till klockan 17.00.
Verksamheten i lekparkerna är avgiftsfri och öppen för alla.
Du kan anmäla ditt barn till lekparkernas eftermiddagsverksamhet med en anmälningsblankett.
Lämna blanketten till den lekpark som anmälan i första hand gäller.
Lekparks- och eftermiddagsverksamhet för skolbarnfinska _ ryska _ somaliska _ arabiska
Anvisningar om eftermiddagsverksamhetens klientavgiftfinska _ ryska _ somaliska _ arabiska
Modersmålsundervisning för invandrare
Barn som har ett annat modersmål än finska eller svenska kan få modersmålsundervisning.
I Helsingfors ges modersmålsundervisning för invandrare på fler än 40 språk.
Du får information om modersmålsundervisningen vid rådgivningen och kundtjänsten vid sektorn för fostran och utbildning.
rådgivningen och kundtjänsten vid sektorn för fostran och utbildning:
Töysägatan 2D
Tfn (09) 310 86400
Yrkesutbildning
Stadin ammatti- ja aikuisopisto är Finlands största yrkesläroanstalt där man kan utbilda sig inom många olika branscher.
I Helsingfors finns även andra yrkesläroanstalter.
Man söker till yrkesutbildning i den gemensamma ansökan.
Vid Stadin ammatti- ja aikuisopisto ordnas förberedande utbildning inför yrkesutbildning för invandrare.
Den förberedande utbildningen är avsedd för ungdomar och vuxna som är intresserade av yrkesutbildning och vill förbättra sina kunskaper i finska.
Den förberedande undervisningen pågår i en termin eller ett läsår.
Information om den förberedande utbildningen får du vid rådgivningen och kundtjänsten vid Stadin ammatti- ja aikuisopisto.
Kontaktuppgifter:
Hattulavägen 2
Tfn (09) 310 8415
Läs mer: Yrkesutbildning, Förberedande utbildning före yrkesutbildning.
Yrkesinriktad utbildningfinska
Yrkesläroanstalterfinska _ svenska _ engelska
För yrkesutbildning förberedande undervisningfinska _ svenska _ engelska
Gymnasium
I Helsingfors finns många gymnasieskolor.
I Helsingfors finns även några sådana gymnasieskolor där undervisningsspråket är något annat än finska eller svenska.
Utöver dagsgymnasierna som är avsedda för ungdomar finns det tre vuxengymnasier (aikuislukio) i Helsingfors.
I Helsingfors arrangeras förberedande utbildning för gymnasiet för invandrare.
Den förberedande utbildningen tar ett läsår och ger beredskap för gymnasiestudier.
Den förberedande utbildningen är avsedd för unga och vuxna som vill studera vid gymnasium men saknar tillräckliga språkkunskaper för gymnasiestudier.
Information om den förberedande utbildningen får du vid rådgivningen och kundtjänsten vid sektorn för fostran och utbildning.
rådgivningen och kundtjänsten vid sektorn för fostran och utbildning:
Töysägatan 2D
Tfn (09) 310 86400
Läs mer: Gymnasium
Gymnasier i Helsingforsfinska _ svenska _ engelska
Gymnasieansökanfinska _ svenska _ engelska
För gymnasium förberedande undervisningfinska _ engelska
Stöd och handledning för unga
Om du är under 30 år gammal kan du få råd och handledning via Ohjaamo-tjänsten.
Ohjaamos personal hjälper dig om du inte har ett arbete eller en studieplats.
Du kan även fråga om andra saker, som till exempel boende eller ekonomiska frågor.
Kontaktuppgifter:
Fredrikinkatu 48
Tfn: 040 70 46 818
Rådgivning för ungafinska
Högskoleutbildning
I Helsingfors kan du avlägga högskolestudier i många branscher.
I Helsingfors finns såväl universitet som yrkeshögskolor.
Största delen av undervisningen på högskolorna ges på finska.
I nästan alla högskolor erbjuds dock även undervisning på engelska.
I Helsingfors finns ett svenskspråkigt universitet och en svenskspråkig yrkeshögskola.
Kontaktuppgifterna till högskolorna finns på Helsingfors stads webbplats.
Anvisningar om ansökning och närmare information om utbildningsprogrammen finns på högskolornas egna webbplatser.
Läs mer: Universitet och Yrkeshögskolor.
Yrkeshögskolorfinska _ svenska _ engelska
Universitetfinska _ svenska _ engelska
Andra studiemöjligheter
I Helsingfors finns många studiemöjligheter som är öppna för alla.
Dessa studier är vanligtvis avgiftsbelagda.
Det är möjligt att avlägga högskolestudier vid öppna universitet och öppna yrkeshögskolor.
Vem som helst kan studera vid dessa.
Det öppna universitetet och de öppna yrkeshögskolorna har ett brett utbud av kurser också på engelska.
Helsingfors stad har ett finskspråkigt arbetarinstitut och ett svenskspråkigt arbetarinstitut.
Vid arbetarinstituten kan du studera t.ex. språk, handarbete och musik.
Studieutbudet är väldigt mångsidigt.
Största delen av arbetarinstitutens kurser går på finska eller svenska.
Arbetarinstituten ordnar kurser också på engelska och ryska.
Läs mer: Studier som hobby.
Finska arbetarinstitutetfinska
Svenskspråkiga arbetarinstitutet Arbisfinska _ svenska _ engelska _ ryska
Kurser för invandrarefinska _ engelska _ ryska
Information om öppna universitetetfinska _ svenska
Information om öppna yrkeshögskolanfinska _ svenska
Dagvård
Förskoleundervisning
Grundläggande undervisning
Eftermiddagsverksamhet för skolbarn
Modersmålsundervisning för invandrare
Yrkesubildning
Gymnasium
Stöd och handledning för unga
Högskoleutbildning
Andra studiemöjligheter
Dagvård
I Helsingfors finns det flera daghem som drivs av staden och privata daghem.
Stadens daghem är finsk- eller svenskspråkiga.
De flesta är finskspråkiga.
Om du ansöker om en dagvårdsplats i stadens daghem, ska du skicka in din ansökan minst fyra månader före dagvårdsstart.
Du kan ansöka om dagvårdsplats vid staden om familjen har sin adress i Helsingfors.
Ansök om dagvårdsplats på Internet.
När du använder den elektroniska blanketten behöver du finländska nätbankkoder.
Dessutom ska ditt barn ha en finländsk personbeteckning.
Om du inte kan använda den elektroniska blanketten kan du skriva ut ansökningsblanketten på stadens webbplats.
Lämna eller posta blanketten till den dagvårdsenhet där du i första hand söker plats.
Du hittar kontaktuppgifterna till daghemmen på stadens webbplats.
Om du har frågor kring dagvården eller om ansökning av dagvårdsplats, kan du ringa rådgivningstelefonen vid stadens tjänster inom småbarnspedagogiken:
Tfn 09 310 44986 (betjänar även på engelska)
I Helsingfors finns även privata daghem vars verksamhetsspråk är engelska, ryska, tyska, franska eller spanska.
I Helsingfors finns även ett muslimskt daghem vars verksamhetsspråk är arabiska.
Om du ansöker om en plats i ett privat daghem, kontakta direkt det daghem som är föremål för platsansökan.
Läs mer: Dagvård.
Dagvård i Helsingforsfinska _ svenska _ engelska
Daghem med vård på främmande språkfinska _ svenska _ engelska
Ansökan om dagvårdsplatsfinska _ svenska _ engelska
Dagvårdsavgifterfinska _ svenska _ engelska
Förskoleundervisning
I Helsingfors ordnas förskoleundervisning (esiopetus) i många daghem och skolor.
På Helsingfors stads webbplats hittar du en lista över de daghem och skolor som ger förskoleundervisning.
Man ansöker till förskoleundervisningen med en elektronisk blankett.
När du använder den elektroniska blanketten behöver du finländska nätbankkoder.
Dessutom ska ditt barn ha en finländsk personbeteckning.
Om du inte kan använda den elektroniska blanketten ska du skriva ut ansökningsblanketten från stadens webbplats eller hämta den vid ett av stadens daghem.
Lämna eller posta blanketten till den dagvårdsenhet där du i första hand söker plats.
Du hittar mer information om förskoleundervisningen på stadens webbplats.
Du kan även fråga om mer information av daghemsföreståndarna.
Förskoleundervisningen börjar i augusti och ansökningstiden är i januari.
Läs mer: Förskoleundervisning.
Daghem som ger förskoleundervisningfinska _ svenska _ engelska
Ansökan till förskoleundervisningfinska _ svenska _ engelska
Förskoleundervisning i Helsingforsfinska _ svenska _ engelska
Grundläggande undervisning
I Helsingfors finns flera grundskolor (peruskoulu).
Utöver stadens egna skolor finns det privata skolor och statliga skolor i Helsingfors.
Studier vid en privat skola kan vara avgiftsbelagda.
I stadens skolor är undervisningsspråket finska eller svenska.
I Helsingfors finns det också privata skolor med undervisning på t.ex. engelska, tyska, franska eller ryska.
Anmälan till grundskolan sker i början av året.
Du kan anmäla ditt barn till skolan via Internet eller genom att besöka skolan på anmälningsdagen.
Helsingfors stads webbsidor ger dig information om anmälningsdagen.
Om barnet inte har tillräckligt bra kunskaper för att klara grundskolan kan han eller hon få förberedande undervisning.
Den förberedande undervisningen förbereder barnet inför grundskolan.
I den förberedande undervisningen ges undervisning i finska och i grundskolans ämnen.
Du kan fråga om den grundläggande utbildningen och om skolorna i Helsingfors vid rådgivningen och kundtjänsten vid sektorn för fostran och utbildning.
Kontaktuppgifter:
Töysägatan 2D
Tfn (09) 310 86400
Vid Helsingfors vuxengymnasium finns en linje avsedd för invandrare över 17 år, där du kan avlägga hela eller en del av den grundläggande utbildningen.
Mer information finns på Helsingfors vuxengymnasiums webbplats.
Också andra vuxengymnasier ger grundläggande utbildning för vuxna.
Kontaktuppgifterna till vuxengymnasierna finns på Helsingfors stads webbplats.
Grundläggande utbildning.
Broschyren Information om den finska grundskolanengelska _ ryska _ franska _ somaliska _ arabiska
Skolornas kontaktuppgifterfinska _ svenska _ engelska
Mer information om anmälanfinska _ svenska _ engelska
Internationella skolor i huvudstadsregionenfinska
linkkiExpatFinland.fi:
Internationella skolor i huvudstadsregionenengelska
linkkiHelsingfors Vuxengymnasium:
Grundläggande utbildning för vuxna invandrarefinska
Grundläggande utbildning för vuxna invandrarefinska _ engelska
Eftermiddagsverksamhet för skolbarn
Helsingfors stad ordnar eftermiddagsverksamhet för barn i årskurs 1 och 2 i skolor och lekparker efter skoldagen.
Eftermiddagsverksamhet ordnas under läsåret på vardagar högst fram till klockan 17.00.
Verksamheten i lekparkerna är avgiftsfri och öppen för alla.
Du kan anmäla ditt barn till lekparkernas eftermiddagsverksamhet med en anmälningsblankett.
Lämna blanketten till den lekpark som anmälan i första hand gäller.
Lekparks- och eftermiddagsverksamhet för skolbarnfinska _ engelska _ ryska _ somaliska _ arabiska
Anvisningar om eftermiddagsverksamhetens klientavgiftfinska _ engelska _ ryska _ somaliska _ arabiska
Modersmålsundervisning för invandrare
Barn som har ett annat modersmål än finska eller svenska kan få modersmålsundervisning.
I Helsingfors ges modersmålsundervisning för invandrare på fler än 40 språk.
Du får information om modersmålsundervisningen vid rådgivningen och kundtjänsten vid sektorn för fostran och utbildning.
rådgivningen och kundtjänsten vid sektorn för fostran och utbildning:
Töysägatan 2D
Tfn (09) 310 86400
Yrkesutbildning
Stadin ammatti- ja aikuisopisto är Finlands största yrkesläroanstalt där man kan utbilda sig inom många olika branscher.
I Helsingfors finns även andra yrkesläroanstalter.
Man söker till yrkesutbildning i den gemensamma ansökan.
Vid Stadin ammatti- ja aikuisopisto ordnas förberedande utbildning inför yrkesutbildning för invandrare.
Den förberedande utbildningen är avsedd för ungdomar och vuxna som är intresserade av yrkesutbildning och vill förbättra sina kunskaper i finska.
Den förberedande undervisningen pågår i en termin eller ett läsår.
Information om den förberedande utbildningen får du vid rådgivningen och kundtjänsten vid Stadin ammatti- ja aikuisopisto.
Kontaktuppgifter:
Hattulavägen 2
Tfn (09) 310 8415
Läs mer: Yrkesutbildning, Förberedande utbildning före yrkesutbildning.
Yrkesinriktad utbildningfinska
Yrkesläroanstalterfinska _ svenska _ engelska
För yrkesutbildning förberedande undervisningfinska _ svenska _ engelska
Gymnasium
I Helsingfors finns många gymnasieskolor.
I Helsingfors finns även några sådana gymnasieskolor där undervisningsspråket är något annat än finska eller svenska.
Utöver dagsgymnasierna som är avsedda för ungdomar finns det tre vuxengymnasier (aikuislukio) i Helsingfors.
I Helsingfors arrangeras förberedande utbildning för gymnasiet för invandrare.
Den förberedande utbildningen tar ett läsår och ger beredskap för gymnasiestudier.
Den förberedande utbildningen är avsedd för unga och vuxna som vill studera vid gymnasium men saknar tillräckliga språkkunskaper för gymnasiestudier.
Information om den förberedande utbildningen får du vid rådgivningen och kundtjänsten vid sektorn för fostran och utbildning.
rådgivningen och kundtjänsten vid sektorn för fostran och utbildning:
Töysägatan 2D
Tfn (09) 310 86400
Läs mer: Gymnasium
Gymnasier i Helsingforsfinska _ svenska _ engelska
Gymnasieansökanfinska _ svenska _ engelska
För gymnasium förberedande undervisningfinska _ engelska
Stöd och handledning för unga
Om du är under 30 år gammal kan du få råd och handledning via Ohjaamo-tjänsten.
Ohjaamos personal hjälper dig om du inte har ett arbete eller en studieplats.
Du kan även fråga om andra saker, som till exempel boende eller ekonomiska frågor.
Kontaktuppgifter:
Fredrikinkatu 48
Tfn: 040 70 46 818
Rådgivning för ungafinska
Högskoleutbildning
I Helsingfors kan du avlägga högskolestudier i många branscher.
I Helsingfors finns såväl universitet som yrkeshögskolor.
Största delen av undervisningen på högskolorna ges på finska.
I nästan alla högskolor erbjuds dock även undervisning på engelska.
I Helsingfors finns ett svenskspråkigt universitet och en svenskspråkig yrkeshögskola.
Kontaktuppgifterna till högskolorna finns på Helsingfors stads webbplats.
Anvisningar om ansökning och närmare information om utbildningsprogrammen finns på högskolornas egna webbplatser.
Läs mer: Universitet och Yrkeshögskolor.
Yrkeshögskolorfinska _ svenska _ engelska
Universitetfinska _ svenska _ engelska
Andra studiemöjligheter
I Helsingfors finns många studiemöjligheter som är öppna för alla.
Dessa studier är vanligtvis avgiftsbelagda.
Det är möjligt att avlägga högskolestudier vid öppna universitet och öppna yrkeshögskolor.
Vem som helst kan studera vid dessa.
Det öppna universitetet och de öppna yrkeshögskolorna har ett brett utbud av kurser också på engelska.
Helsingfors stad har ett finskspråkigt arbetarinstitut och ett svenskspråkigt arbetarinstitut.
Vid arbetarinstituten kan du studera t.ex. språk, handarbete och musik.
Studieutbudet är väldigt mångsidigt.
Största delen av arbetarinstitutens kurser går på finska eller svenska.
Arbetarinstituten ordnar kurser också på engelska och ryska.
Läs mer: Studier som hobby.
Finska arbetarinstitutetfinska _ engelska _ ryska
Svenskspråkiga arbetarinstitutet Arbisfinska _ svenska _ engelska _ ryska
Kurser för invandrarefinska _ engelska _ ryska
Information om öppna universitetetfinska _ svenska
Information om öppna yrkeshögskolanfinska _ svenska
Hyresbostad
Köpa bostad
Bostadsrättsbostad
Boende i en krissituation
Bostadslöshet
Stöd- och serviceboende
Avfallshantering och återvinning
Hyresbostad
Hyresnivån är hög i Helsingfors.
Förbered dig på att det kan ta lång tid att hitta en bostad.
Du kan hyra en bostad av privata hyresvärdar eller ansöka om en av Helsingfors stads hyresbostäder.
Du är själv ansvarig för att skaffa en bostad åt dig.
Varken staden eller andra hyresvärdar är skyldiga att erbjuda dig en bostad.
Det lönar sig att söka efter en bostad på ett stort område.
Då har du bättre chanser att hitta en bostad.
Hyrorna för bostäder i Helsingfors grannkommuner (till exempel i Vanda, Esbo eller Kervo) är lite förmånligare än i Helsingfors.
Privata hyresbostäder
I Helsingfors finns många privata hyresvärdar som du kan söka bostad hos.
Till exempel Sato, Vvo och Avara äger hyresbostäder i Helsingfors.
Även försäkringsbolag, banker och många privatpersoner hyr ut bostäder.
Hos en privat hyresvärd kan du få en bostad snabbt.
Om du är studerande kan du söka hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS.
Sökning av hyresbostäderfinska
Sökning av hyresbostäderfinska _ engelska
linkkiHOAS:
Hyresbostäder för studerandefinska _ svenska _ engelska
Stadens hyresbostäder
Hyrorna för Helsingfors stads hyresbostäder är lägre än de för privata hyresbostäder.
Det finns emellertid många sökanden till stadens bostäder och bara en liten del av alla sökanden får en bostad.
För att du ska kunna söka en hyresbostad hos staden, ska du ha uppehållstillstånd för minst ett år.
Om du har en finländsk personbeteckning kan du söka hyresbostad hos Helsingfors stad via internettjänsten stadinasunnot.fi.
Du kan också lämna in en ansökan vid ett serviceställe.
Medarbetaren vid servicestället kan hjälpa dig att fylla i ansökningen.
Du kan få betjäning på finska och engelska.
Serviceställets kontaktuppgifter:
Stadin asunnot
Adress: Östersjögatan 3
Tfn (09) 310 13030
En bostadsansökan är giltig i tre månader.
Därefter ska en ny ansökning göras.
Läs mer:
Hyresbostad och Hyresavtal.
Stadin asunnotfinska _ svenska _ engelska
Köpa bostad
I Helsingfors är bostäderna i allmänhet dyra, men priserna varierar mycket mellan olika områden.
Du hittar bostäder till försäljning på sidor för bostadssökande på internet.
Du får information om hur du köper en bostad på InfoFinlands sida Köpa bostad.
Bostadsrättsbostad
Du kan ansöka om bostadsrättsbostad (asumisoikeusasunto), om du inte har en ägarbostad, och inte heller råd att skaffa en sådan.
Om du vill ansöka om ägarbostad i Helsingfors, Esbo eller Vanda, ska du först skaffa ett könummer.
Du kan skaffa könumret via internet.
Du kan också skriva ut en ansökningsblankett och fylla i den för hand.
När du har fått ett könummer, kan du höra dig för om lediga bostäder hos ägare och byggherrar.
Kontaktuppgifter finns på webbplatsen för Helsingfors stad.
Du kan söka bostad samtidigt på många olika områden.
Läs mer: Bostadsrättsbostad.
Bostadsrättsbostäderfinska _ svenska _ engelska
Ansökan om ordningsnummerfinska
Byggherrarnas kontaktuppgifterfinska
Boende i en krissituation
Om din bostad har skadats, till exempel till följd av brand eller vattenskada, kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
Kontakta ditt försäkringsbolag direkt när skadan har inträffat.
Om en familjemedlem är våldsam eller hotar med våld, ta kontakt med ett skyddshem (turvakoti).
Skyddshemmet Mona är avsett för invandrarkvinnor och deras barn.
Tfn 045 639 6274 (24h)
Du kan också vända dig till Huvudstadens Skyddshem (Pääkaupungin Turvakoti).
Adress: Steniusvägen 20
Tfn (09) 4777 180 (24h)
Unga i åldern 12–19 år kan kontakta Röda Korsets De ungas skyddshus (Nuorten turvatalo).
Öppet varje dag kl. 17–10.
Tfn (09) 622 4322.
Du kan ringa skyddshuset under alla tider på dygnet.
E-postadress: turvatalo.helsinki(snabel-a)redcross.fi
Information för bostadslösafinska _ svenska _ engelska
Servicepunkt för socialarbete och socialhandledningfinska
Hjälp till offer för familjevåldfinska
linkkiFinlands Röda Kors:
De ungas skyddshus i Helsingforsfinska _ svenska
Bostadslöshet
Om du blir bostadslös, ta då kontakt med servicestället för socialarbete på ditt område.
En socialarbetare kan hjälpa dig att hitta bostad.
De bostadslösas servicecenter på Sanduddsgatan har öppet dygnet runt varje dag.
Där kan du vid behov övernatta.
Servicecentret erbjuder nattlogi åt helsingforsare med missbruksproblem, om de inte har något annat ställe att övernatta.
Sanduddsgatan 5 B
Tfn (09) 310 466 28
Vailla vakinaista asuntoa ry. är en förening som hjälper bostadslösa.
Vailla vakinaista asuntoa ry har ett nattcenter, Kalkkers, som erbjuder varmt nattlogi för bostadslösa från höst till vår.
Kalkkers håller öppet kl. 22–6.
Till Kalkkers kan du även komma utan uppehållstillstånd.
Adress: Vasagatan 5
Tfn 050 443 1068
Läs mer: Bostadslöshet.
Information för bostadslösafinska _ svenska _ engelska
Servicepunkt för socialarbete och socialhandledningfinska
Föreningen för bostadslösafinska
Serviceguide för bostadslösa i Helsingforsfinska _ engelska _ ryska _ somaliska _ persiska _ arabiska _ bulgariska
Stöd- och serviceboende
Vissa personer, till exempel äldre eller personer med funktionsnedsättning, har svårt att klara av de dagliga sysslorna utan hjälp.
Staden ordnar tjänster för dem, så att de kan bo självständigt.
Äldre eller personer med funktionsnedsättning som inte kan bo självständigt kan bo i ett servicehus eller på en anstalt.
Du kan fråga mer om tjänsterna vid enheten för socialarbete i ditt bostadsområde.
Läs mer: Stöd- och serviceboende
Enheterna för socialt arbete och närarbetefinska _ svenska _ engelska
Serviceboendefinska _ svenska _ engelska
Boendetjänster för handikappadefinska _ svenska _ engelska
Avfallshantering och återvinning
På InfoFinlands sida Avfallshantering och återvinning hittar du information om sortering av avfall.
Information om avfallshanteringfinska _ svenska _ engelska
linkkiHelsingforsregionens miljötjänster:
Sopsorteringsanvisningarfinska _ svenska _ engelska
linkkiHelsingforsregionens miljötjänster:
Återvinningsstationerfinska _ svenska _ engelska
Avfallsinsamlingsstationerfinska
Hyresbostad
Köpa bostad
Bostadsrättsbostad
Boende i en krissituation
Bostadslöshet
Stöd- och serviceboende
Avfallshantering och återvinning
Hyresbostad
Hyresnivån är hög i Helsingfors.
Förbered dig på att det kan ta lång tid att hitta en bostad.
Du kan hyra en bostad av privata hyresvärdar eller ansöka om en av Helsingfors stads hyresbostäder.
Du är själv ansvarig för att skaffa en bostad åt dig.
Varken staden eller andra hyresvärdar är skyldiga att erbjuda dig en bostad.
Det lönar sig att söka efter en bostad på ett stort område.
Då har du bättre chanser att hitta en bostad.
Hyrorna för bostäder i Helsingfors grannkommuner (till exempel i Vanda, Esbo eller Kervo) är lite förmånligare än i Helsingfors.
Privata hyresbostäder
I Helsingfors finns många privata hyresvärdar som du kan söka bostad hos.
Till exempel Sato, Vvo och Avara äger hyresbostäder i Helsingfors.
Även försäkringsbolag, banker och många privatpersoner hyr ut bostäder.
Hos en privat hyresvärd kan du få en bostad snabbt.
Om du är studerande kan du söka hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS.
Sökning av hyresbostäderfinska
Sökning av hyresbostäderfinska _ engelska
linkkiHOAS:
Hyresbostäder för studerandefinska _ svenska _ engelska
Stadens hyresbostäder
Hyrorna för Helsingfors stads hyresbostäder är lägre än de för privata hyresbostäder.
Det finns emellertid många sökanden till stadens bostäder och bara en liten del av alla sökanden får en bostad.
För att du ska kunna söka en hyresbostad hos staden, ska du ha uppehållstillstånd för minst ett år.
Om du har en finländsk personbeteckning kan du söka hyresbostad hos Helsingfors stad via internettjänsten stadinasunnot.fi.
Du kan också lämna in en ansökan vid ett serviceställe.
Medarbetaren vid servicestället kan hjälpa dig att fylla i ansökningen.
Du kan få betjäning på finska och engelska.
Serviceställets kontaktuppgifter:
Stadin asunnot
Adress: Östersjögatan 3
Tfn (09) 310 13030
En bostadsansökan är giltig i tre månader.
Därefter ska en ny ansökning göras.
Läs mer:
Hyresbostad och Hyresavtal.
Stadin asunnotfinska _ svenska _ engelska
Köpa bostad
I Helsingfors är bostäderna i allmänhet dyra, men priserna varierar mycket mellan olika områden.
Du hittar bostäder till försäljning på sidor för bostadssökande på internet.
Du får information om hur du köper en bostad på InfoFinlands sida Köpa bostad.
Bostadsrättsbostad
Du kan ansöka om bostadsrättsbostad (asumisoikeusasunto), om du inte har en ägarbostad, och inte heller råd att skaffa en sådan.
Om du vill ansöka om ägarbostad i Helsingfors, Esbo eller Vanda, ska du först skaffa ett könummer.
Du kan skaffa könumret via internet.
Du kan också skriva ut en ansökningsblankett och fylla i den för hand.
När du har fått ett könummer, kan du höra dig för om lediga bostäder hos ägare och byggherrar.
Kontaktuppgifter finns på webbplatsen för Helsingfors stad.
Du kan söka bostad samtidigt på många olika områden.
Läs mer: Bostadsrättsbostad.
Bostadsrättsbostäderfinska _ svenska _ engelska
Ansökan om ordningsnummerfinska
Byggherrarnas kontaktuppgifterfinska
Boende i en krissituation
Om din bostad har skadats, till exempel till följd av brand eller vattenskada, kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
Kontakta ditt försäkringsbolag direkt när skadan har inträffat.
Om en familjemedlem är våldsam eller hotar med våld, ta kontakt med ett skyddshem (turvakoti).
Skyddshemmet Mona är avsett för invandrarkvinnor och deras barn.
Tfn 045 639 6274 (24h)
Du kan också vända dig till Huvudstadens Skyddshem (Pääkaupungin Turvakoti).
Adress: Steniusvägen 20
Tfn (09) 4777 180 (24h)
Unga i åldern 12–19 år kan kontakta Röda Korsets De ungas skyddshus (Nuorten turvatalo).
Öppet varje dag kl. 17–10.
Tfn (09) 622 4322.
Du kan ringa skyddshuset under alla tider på dygnet.
E-postadress: turvatalo.helsinki(snabel-a)redcross.fi
Information för bostadslösafinska _ svenska _ engelska
Servicepunkt för socialarbete och socialhandledningfinska
Hjälp till offer för familjevåldfinska
linkkiFinlands Röda Kors:
De ungas skyddshus i Helsingforsfinska _ svenska
Bostadslöshet
Om du blir bostadslös, ta då kontakt med servicestället för socialarbete på ditt område.
En socialarbetare kan hjälpa dig att hitta bostad.
De bostadslösas servicecenter på Sanduddsgatan har öppet dygnet runt varje dag.
Där kan du vid behov övernatta.
Servicecentret erbjuder nattlogi åt helsingforsare med missbruksproblem, om de inte har något annat ställe att övernatta.
Sanduddsgatan 5 B
Tfn (09) 310 466 28
Vailla vakinaista asuntoa ry. är en förening som hjälper bostadslösa.
Vailla vakinaista asuntoa ry har ett nattcenter, Kalkkers, som erbjuder varmt nattlogi för bostadslösa från höst till vår.
Kalkkers håller öppet kl. 22–6.
Till Kalkkers kan du även komma utan uppehållstillstånd.
Adress: Vasagatan 5
Tfn 050 443 1068
Läs mer: Bostadslöshet.
Information för bostadslösafinska _ svenska _ engelska
Servicepunkt för socialarbete och socialhandledningfinska
Föreningen för bostadslösafinska
Serviceguide för bostadslösa i Helsingforsfinska _ engelska _ ryska _ somaliska _ persiska _ arabiska _ bulgariska
Stöd- och serviceboende
Vissa personer, till exempel äldre eller personer med funktionsnedsättning, har svårt att klara av de dagliga sysslorna utan hjälp.
Staden ordnar tjänster för dem, så att de kan bo självständigt.
Äldre eller personer med funktionsnedsättning som inte kan bo självständigt kan bo i ett servicehus eller på en anstalt.
Du kan fråga mer om tjänsterna vid enheten för socialarbete i ditt bostadsområde.
Läs mer: Stöd- och serviceboende
Enheterna för socialt arbete och närarbetefinska _ svenska _ engelska
Serviceboendefinska _ svenska _ engelska
Boendetjänster för handikappadefinska _ svenska _ engelska
Avfallshantering och återvinning
På InfoFinlands sida Avfallshantering och återvinning hittar du information om sortering av avfall.
Information om avfallshanteringfinska _ svenska _ engelska
linkkiHelsingforsregionens miljötjänster:
Sopsorteringsanvisningarfinska _ svenska _ engelska
linkkiHelsingforsregionens miljötjänster:
Återvinningsstationerfinska _ svenska _ engelska
Avfallsinsamlingsstationerfinska
Hyresbostad
Köpa bostad
Bostadsrättsbostad
Boende i en krissituation
Bostadslöshet
Stöd- och serviceboende
Avfallshantering och återvinning
Hyresbostad
Hyresnivån är hög i Helsingfors.
Förbered dig på att det kan ta lång tid att hitta en bostad.
Du kan hyra en bostad av privata hyresvärdar eller ansöka om en av Helsingfors stads hyresbostäder.
Du är själv ansvarig för att skaffa en bostad åt dig.
Varken staden eller andra hyresvärdar är skyldiga att erbjuda dig en bostad.
Det lönar sig att söka efter en bostad på ett stort område.
Då har du bättre chanser att hitta en bostad.
Hyrorna för bostäder i Helsingfors grannkommuner (till exempel i Vanda, Esbo eller Kervo) är lite förmånligare än i Helsingfors.
Privata hyresbostäder
I Helsingfors finns många privata hyresvärdar som du kan söka bostad hos.
Till exempel Sato, Vvo och Avara äger hyresbostäder i Helsingfors.
Även försäkringsbolag, banker och många privatpersoner hyr ut bostäder.
Hos en privat hyresvärd kan du få en bostad snabbt.
Om du är studerande kan du söka hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS.
Sökning av hyresbostäderfinska
Sökning av hyresbostäderfinska _ engelska
linkkiHOAS:
Hyresbostäder för studerandefinska _ svenska _ engelska
Stadens hyresbostäder
Hyrorna för Helsingfors stads hyresbostäder är lägre än de för privata hyresbostäder.
Det finns emellertid många sökanden till stadens bostäder och bara en liten del av alla sökanden får en bostad.
För att du ska kunna söka en hyresbostad hos staden, ska du ha uppehållstillstånd för minst ett år.
Om du har en finländsk personbeteckning kan du söka hyresbostad hos Helsingfors stad via internettjänsten stadinasunnot.fi.
Du kan också lämna in en ansökan vid ett serviceställe.
Medarbetaren vid servicestället kan hjälpa dig att fylla i ansökningen.
Du kan få betjäning på finska och engelska.
Serviceställets kontaktuppgifter:
Stadin asunnot
Adress: Sörnäsgatan 1
Tfn (09) 310 13030
En bostadsansökan är giltig i tre månader.
Därefter ska en ny ansökning göras.
Läs mer:
Hyresbostad och Hyresavtal.
Stadin asunnotfinska _ svenska _ engelska
Köpa bostad
I Helsingfors är bostäderna i allmänhet dyra, men priserna varierar mycket mellan olika områden.
Du hittar bostäder till försäljning på sidor för bostadssökande på internet.
Du får information om hur du köper en bostad på InfoFinlands sida Köpa bostad.
Bostadsrättsbostad
Du kan ansöka om bostadsrättsbostad (asumisoikeusasunto), om du inte har en ägarbostad, och inte heller råd att skaffa en sådan.
Om du vill ansöka om ägarbostad i Helsingfors, Esbo eller Vanda, ska du först skaffa ett könummer.
Du kan skaffa könumret via internet.
Du kan också skriva ut en ansökningsblankett och fylla i den för hand.
När du har fått ett könummer, kan du höra dig för om lediga bostäder hos ägare och byggherrar.
Kontaktuppgifter finns på webbplatsen för Helsingfors stad.
Du kan söka bostad samtidigt på många olika områden.
Läs mer: Bostadsrättsbostad.
Bostadsrättsbostäderfinska _ svenska _ engelska
Ansökan om ordningsnummerfinska _ svenska _ engelska
Byggherrarnas kontaktuppgifterfinska _ svenska _ engelska
Boende i en krissituation
Om din bostad har skadats, till exempel till följd av brand eller vattenskada, kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
Kontakta ditt försäkringsbolag direkt när skadan har inträffat.
Om en familjemedlem är våldsam eller hotar med våld, ta kontakt med ett skyddshem (turvakoti).
Skyddshemmet Mona är avsett för invandrarkvinnor och deras barn.
Tfn 045 639 6274 (24h)
Du kan också vända dig till Huvudstadens Skyddshem (Pääkaupungin Turvakoti).
Adress: Steniusvägen 20, 00320 Helsingfors
Tfn (09) 4777 180 (24h)
Tfn 050 5650 636 (24h)
Unga i åldern 12–19 år kan kontakta Röda Korsets De ungas skyddshus (Nuorten turvatalo).
Öppet varje dag kl. 17–10.
Tfn (09) 622 4322.
Du kan ringa skyddshuset under alla tider på dygnet.
E-postadress: turvatalo.helsinki(snabel-a)redcross.fi
Information för bostadslösafinska _ svenska _ engelska
Servicepunkt för socialarbete och socialhandledningfinska _ svenska _ engelska
Hjälp till offer för familjevåldfinska
linkkiFinlands Röda Kors:
De ungas skyddshus i Helsingforsfinska _ svenska
Bostadslöshet
Om du blir bostadslös, ta då kontakt med servicestället för socialarbete på ditt område.
En socialarbetare kan hjälpa dig att hitta bostad.
De bostadslösas servicecenter på Sanduddsgatan har öppet dygnet runt varje dag.
Där kan du vid behov övernatta.
Servicecentret erbjuder nattlogi åt helsingforsare med missbruksproblem, om de inte har något annat ställe att övernatta.
Sanduddsgatan 5 B
Tfn (09) 310 466 28
Vailla vakinaista asuntoa ry. är en förening som hjälper bostadslösa.
Vailla vakinaista asuntoa ry har ett nattcenter, Kalkkers, som erbjuder varmt nattlogi för bostadslösa från höst till vår.
Kalkkers håller öppet kl. 22–6.
Till Kalkkers kan du även komma utan uppehållstillstånd.
Adress: Vasagatan 5
Tfn 050 443 1068
Läs mer: Bostadslöshet.
Information för bostadslösafinska _ svenska _ engelska
Servicepunkt för socialarbete och socialhandledningfinska _ svenska _ engelska
Föreningen för bostadslösafinska _ engelska
Serviceguide för bostadslösa i Helsingfors(pdf, 3,7 MB)finska _ engelska _ ryska _ somaliska _ persiska _ arabiska _ bulgariska
Stöd- och serviceboende
Vissa personer, till exempel äldre eller personer med funktionsnedsättning, har svårt att klara av de dagliga sysslorna utan hjälp.
Staden ordnar tjänster för dem, så att de kan bo självständigt.
Äldre eller personer med funktionsnedsättning som inte kan bo självständigt kan bo i ett servicehus eller på en anstalt.
Du kan fråga mer om tjänsterna vid enheten för socialarbete i ditt bostadsområde.
Läs mer: Stöd- och serviceboende
Enheterna för socialt arbete och närarbetefinska _ svenska _ engelska
Serviceboendefinska _ svenska _ engelska
Boendetjänster för handikappadefinska _ svenska _ engelska
Avfallshantering och återvinning
På InfoFinlands sida Avfallshantering och återvinning hittar du information om sortering av avfall.
Information om avfallshanteringfinska _ svenska _ engelska
linkkiHelsingforsregionens miljötjänster:
Sopsorteringsanvisningarfinska _ svenska _ engelska
linkkiHelsingforsregionens miljötjänster:
Återvinningsstationerfinska _ svenska _ engelska
Avfallsinsamlingsstationerfinska
Studier i finska och svenska
Språkkurser
Med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig finskakurs i Helsingfors, Vanda, Esbo eller Grankulla.
Kurserna i svenska finns under en länk på tjänstens förstasida.
Du kan använda tjänsten på finska, engelska och ryska.
Anmälan till språkkurserna görs vanligtvis ungefär 2–8 veckor före kursstart.
Till en del kurser måste du ansöka.
Till en del kurser kan du anmäla dig på Internet.
Kurser i finska och svenska språketfinska _ engelska _ ryska
Du kan studera finska och svenska till exempel på kurser vid arbetarinstitut och i anslutning till yrkesstudier.
Helsingfors svenskspråkiga arbetarinstitut Arbis erbjuder många kurser i svenska.
På adressen Ilmonet.fi hittar du hela kursutbudet vid arbetar- och medborgarinstitut i huvudstadsregionen.
linkkiIlmonet.fi:
Kurssökningfinska _ svenska _ engelska
linkkiArbis:
Kurser i svenskafinska _ svenska _ engelska
Till arbets- och näringsbyråns (työ- ja elinkeinotoimisto) kurser i finska eller svenska ansöker du via arbets- och näringsbyrån.
Fråga mer vid din egen arbets- och näringsbyrå.
Samtala på finska
På biblioteken i Helsingfors ordnas språkkaféer, där man kan öva sig i att prata finska.
De är avsedda för alla som vill lära sig att prata finska.
På språkkaféerna samtalar man på finska, så det är bra om du redan kan lite finska.
Språkkaféerna är avgiftsfria.
Du kan fråga mer om språkkaféerna på biblioteken.
Språkkaféerfinska _ svenska _ engelska _ ryska
Allmän språkexamen
I Helsingfors kan du avlägga allmän språkexamen (yleinen kielitutkinto) i finska eller svenska.
På utbildningsstyrelsens (opetushallitus) webbplats finns en sökmotor med vilken du kan se var och när du kan avlägga examen.
Läs mer: Officiellt intyg om språkkunskaper.
linkkiUtbildningsstyrelsen:
Examenssökningfinska
Läs mer: Finska och svenska språket.
Studier i finska och svenska
Språkkurser
Med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig finskakurs i Helsingfors, Vanda, Esbo eller Grankulla.
Kurserna i svenska finns under en länk på tjänstens förstasida.
Du kan använda tjänsten på finska, engelska och ryska.
Anmälan till språkkurserna görs vanligtvis ungefär 2–8 veckor före kursstart.
Till en del kurser måste du ansöka.
Till en del kurser kan du anmäla dig på Internet.
Kurser i finska och svenska språketfinska _ engelska _ ryska
Du kan studera finska och svenska till exempel på kurser vid arbetarinstitut och i anslutning till yrkesstudier.
Helsingfors svenskspråkiga arbetarinstitut Arbis erbjuder många kurser i svenska.
På adressen Ilmonet.fi hittar du hela kursutbudet vid arbetar- och medborgarinstitut i huvudstadsregionen.
linkkiIlmonet.fi:
Kurssökningfinska _ svenska _ engelska
linkkiArbis:
Kurser i svenskafinska _ svenska _ engelska
Till arbets- och näringsbyråns (työ- ja elinkeinotoimisto) kurser i finska eller svenska ansöker du via arbets- och näringsbyrån.
Fråga mer vid din egen arbets- och näringsbyrå.
Samtala på finska
På biblioteken i Helsingfors ordnas språkkaféer, där man kan öva sig i att prata finska.
De är avsedda för alla som vill lära sig att prata finska.
På språkkaféerna samtalar man på finska, så det är bra om du redan kan lite finska.
Språkkaféerna är avgiftsfria.
Du kan fråga mer om språkkaféerna på biblioteken.
Språkkaféerfinska _ svenska _ engelska _ ryska
Allmän språkexamen
I Helsingfors kan du avlägga allmän språkexamen (yleinen kielitutkinto) i finska eller svenska.
På utbildningsstyrelsens (opetushallitus) webbplats finns en sökmotor med vilken du kan se var och när du kan avlägga examen.
Läs mer: Officiellt intyg om språkkunskaper.
linkkiUtbildningsstyrelsen:
Examenssökningfinska
Läs mer: Finska och svenska språket.
Studier i finska och svenska
Språkkurser
Med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig finskakurs i Helsingfors, Vanda, Esbo eller Grankulla.
Kurserna i svenska finns under en länk på tjänstens förstasida.
Du kan använda tjänsten på finska, engelska och ryska.
Anmälan till språkkurserna görs vanligtvis ungefär 2–8 veckor före kursstart.
Till en del kurser måste du ansöka.
Till en del kurser kan du anmäla dig på Internet.
Kurser i finska och svenska språketfinska _ engelska _ ryska
Du kan studera finska och svenska till exempel på kurser vid arbetarinstitut och i anslutning till yrkesstudier.
Helsingfors svenskspråkiga arbetarinstitut Arbis erbjuder många kurser i svenska.
På adressen Ilmonet.fi hittar du hela kursutbudet vid arbetar- och medborgarinstitut i huvudstadsregionen.
linkkiIlmonet.fi:
Kurssökningfinska _ svenska _ engelska
linkkiArbis:
Kurser i svenskafinska _ svenska _ engelska
Till arbets- och näringsbyråns (työ- ja elinkeinotoimisto) kurser i finska eller svenska ansöker du via arbets- och näringsbyrån.
Fråga mer vid din egen arbets- och näringsbyrå.
Samtala på finska
På biblioteken i Helsingfors ordnas språkkaféer, där man kan öva sig i att prata finska.
De är avsedda för alla som vill lära sig att prata finska.
På språkkaféerna samtalar man på finska, så det är bra om du redan kan lite finska.
Språkkaféerna är avgiftsfria.
Du kan fråga mer om språkkaféerna på biblioteken.
Språkkaféerfinska _ engelska
Allmän språkexamen
I Helsingfors kan du avlägga allmän språkexamen (yleinen kielitutkinto) i finska eller svenska.
På utbildningsstyrelsens (opetushallitus) webbplats finns en sökmotor med vilken du kan se var och när du kan avlägga examen.
Läs mer: Officiellt intyg om språkkunskaper.
linkkiUtbildningsstyrelsen:
Examenssökningfinska
Läs mer: Finska och svenska språket.
Var hittar jag jobb?
Hjälp med att söka jobb
Att grunda ett företag
Beskattning
Var hittar jag jobb?
TE-byråns tjänster
Du får hjälp med jobbsökningen på arbets- och näringsbyrån (Työ- ja elinkeinotoimisto), d.v.s. TE-byrån.
Om du är arbetslös och söker jobb, anmäl dig som arbetssökande till TE-byrån.
Du kan anmäla dig antingen via webbtjänsten eller personligen på TE-byrån.
Medborgare i ett EU-land, Norge, Island, Lichtenstein och Schweiz kan anmäla sig som arbetssökande via TE-byråns webbtjänst.
Medborgare från övriga länder måste anmäla sig personligen på TE-byrån.
Ta med dig identitetsbevis och uppehållstillstånd.
Du hittar information om TE-byråns tjänster på InfoFinlands sida Om du blir arbetslös.
Information om att söka jobb i Finland hittar du på InfoFinlands sida Var hittar jag jobb?
I Helsingfors finns tre TE-byråer.
Adress:
Kundgatan 3 A, 4:e våningen
Telefon: 0295 025 500
Öppettider: mån–fre kl. 9.00–16.00
Verksamhetsstället i centrum
Adress: Anttigatan 1, 2. våningen
Telefon: 0295 025 500
Öppettider: mån–fre kl. 9.00–16.00
Böle verksamhetsställe
Adress: Bangårdsvägen 7 (ingång via Loktorget)
Telefon: 0295 025 500
Öppettider: mån–fre kl. 9.00–16.00
Arbetslöshetsersättning
Information om att ansöka om arbetslöshetsersättning hittar du på InfoFinlands sida Arbetslöshetsförsäkring.
linkkiArbets- och näringsförvaltningen:
Länkar till jobbsajterfinska _ svenska _ engelska
linkkiArbets- och näringsministeriet:
Lediga jobbfinska _ svenska
linkkiTE-tjänster:
Videoklipp och broschyrer för invandrarefinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska
Hjälp med att söka jobb
Stadens tjänster för arbetslösa
Helsingfors stad hjälper arbetslösa helsingforsare att hitta jobb eller utbildning.
Om du behöver råd eller stöd för att hitta sysselsättning eller utbildning i finska språket, kontakta Helsingfors stads sysselsättningstjänster.
Stadens tjänster för arbetslösafinska _ svenska _ engelska
Integrationscentret Kotoutumiskeskus Monika hjälper arbetslösa invandrarkvinnor att hitta jobb.
Du kan få hjälp med att skriva din CV eller en jobbansökan, studera vardagsfinska och digitala färdigheter.
Luckan integration
Luckan Integration är en rådgivningstjänst som erbjuder invandrare personlig rådgivning, och ordnar bland annat möten och grupper i anslutning till arbetssökande.
Mötesspråket är engelska.
Råd om jobbsökningfinska _ svenska _ engelska _ spanska
Väestöliittos mentorskap i fråga om arbetskarriär är avsett för utbildade invandrare.
Via det kan du få en mentor som stöder dig när du söker arbete eller studieplats eller grundar ett företag.
Verksamheten är finskspråkig.
Mentorskap i fråga om arbetskarriärfinska _ engelska
Om du är under 30 år, kan du fråga råd om jobbsökande på Ohjaamo.
Ohjaamo är en rådgivningstjänst som är avsedd för unga vuxna.
Kompetenscentret Stadin osaamiskeskus (Stadin osaamiskeskus) förbereder invandrare för arbetsmarknaden och hjälper dem att hitta ett jobb eller en praktikplats.
Kompetenscentret erbjuder sina kunder bland annat undervisning i finska och yrkesutbildning.
Du kan bli kund vid Kompetenscentret via TE-byrån eller social -eller hälsovårdsverket.
Tjänsterna är avsedda för invandrare i Helsingfors som fyllt 17 år och har uppehållstillstånd.
Kompetenscenterfinska
Att grunda ett företag
Vid NewCo Helsinki får du råd och hjälp med att starta ett företag.
Du kan få personlig rådgivning om startande av ett företag på finska, svenska, engelska, ryska, arabiska, estniska, tyska och italienska.
NewCo Helsinki ordnar infomöten för invandrare om startande av ett företag.
Infomöten ordnas på finska, engelska, ryska, arabiska och estniska.
Infomötena är avgiftsfria.
Mer information och anmälan finns på NewCo Helsinkis webbplats.
NewCo Helsinki ordnar företagarutbildning på finska, engelska och ryska.
En del av kurserna är avsedda för personer som vill grunda ett företag, och en del för dem som redan har ett eget företag.
Kurser hålls på finska, engelska och ryska.
Mer information och anmälan finns på NewCo Helsinkis webbplats.
NewCo Helsinki ordnar också möten för nätverkande för nya företagare.
Från NewCo Helsinki får du också hjälp med att utveckla uppstartsföretag.
Om du har ett företag i Helsingfors kan du bli medlem i Helsingfors företagare (Helsingin Yrittäjät).
Helsingfors företagare är företagarnas intressebevakningsorganisation som erbjuder sina medlemmar till exempel utbildning, nätverk och rådgivning.
Mer information hittar du på organisationens webbplats.
Läs mer: Att grunda ett företag.
Som företagare till Finland:
Vilka tillstånd behöver du?(pdf, 384 kt)finska _ engelska
Guiden Bli företagare i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ turkiska _ kinesiska _ arabiska _ kurdiska
linkkiHelsingfors Företagare:
Företagarnas intressebevakningsorganisationfinska
Beskattning
Skattebyrån (verotoimisto) har ett serviceställe i centrala Helsingfors.
Kontaktuppgifter till skattebyråns andra serviceställen och telefonrådgivning hittar du på Skatteförvaltningens (verohallinto) webbplats.
Invandrare kan även sköta ärenden vid servicestället International House Helsinki.
På servicestället hjälper FPA:s och Skatteförvaltningens experter invandrare som kommer till Finland för att arbeta i frågor som rör beskattning och social trygghet.
Kontaktuppgifter till skattebyrån:
Alexandersgatan 9, 4:e våningen (Köpcentret Kluuvi)
Kontaktuppgifter till servicestället International House Helsinki:
Albertsgatan 25
Läs mer: Beskattning.
linkkiSkatteförvaltningen:
Kontaktuppgifter till skattebyråerfinska _ svenska _ engelska
IHH – serviceställe för dig som flyttar till Finland engelska
Var hittar jag jobb?
Hjälp med att söka jobb
Att grunda ett företag
Beskattning
Var hittar jag jobb?
TE-byråns tjänster
Du får hjälp med jobbsökningen på arbets- och näringsbyrån (Työ- ja elinkeinotoimisto), d.v.s. TE-byrån.
Om du är arbetslös och söker jobb, anmäl dig som arbetssökande till TE-byrån.
Du kan anmäla dig antingen via webbtjänsten eller personligen på TE-byrån.
Medborgare i ett EU-land, Norge, Island, Lichtenstein och Schweiz kan anmäla sig som arbetssökande via TE-byråns webbtjänst.
Medborgare från övriga länder måste anmäla sig personligen på TE-byrån.
Ta med dig identitetsbevis och uppehållstillstånd.
Du hittar information om TE-byråns tjänster på InfoFinlands sida Om du blir arbetslös.
Information om att söka jobb i Finland hittar du på InfoFinlands sida Var hittar jag jobb?
I Helsingfors finns tre TE-byråer.
Adress:
Kundgatan 3 A, 4:e våningen
Telefon: 0295 025 500
Öppettider: mån–fre kl. 9.00–16.00
Verksamhetsstället i centrum
Adress: Anttigatan 1, 2. våningen
Telefon: 0295 025 500
Öppettider: mån–fre kl. 9.00–16.00
Böle verksamhetsställe
Adress: Bangårdsvägen 7 (ingång via Loktorget)
Telefon: 0295 025 500
Öppettider: mån–fre kl. 9.00–16.00
Arbetslöshetsersättning
Information om att ansöka om arbetslöshetsersättning hittar du på InfoFinlands sida Arbetslöshetsförsäkring.
linkkiArbets- och näringsförvaltningen:
Länkar till jobbsajterfinska _ svenska _ engelska
linkkiArbets- och näringsministeriet:
Lediga jobbfinska _ svenska
linkkiTE-tjänster:
Videoklipp och broschyrer för invandrarefinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska
Hjälp med att söka jobb
Stadens tjänster för arbetslösa
Helsingfors stad hjälper arbetslösa helsingforsare att hitta jobb eller utbildning.
Om du behöver råd eller stöd för att hitta sysselsättning eller utbildning i finska språket, kontakta Helsingfors stads sysselsättningstjänster.
Stadens tjänster för arbetslösafinska _ svenska _ engelska
Integrationscentret Kotoutumiskeskus Monika hjälper arbetslösa invandrarkvinnor att hitta jobb.
Du kan få hjälp med att skriva din CV eller en jobbansökan, studera vardagsfinska och digitala färdigheter.
Luckan integration
Luckan Integration är en rådgivningstjänst som erbjuder invandrare personlig rådgivning, och ordnar bland annat möten och grupper i anslutning till arbetssökande.
Mötesspråket är engelska.
Råd om jobbsökningfinska _ svenska _ engelska _ spanska
Väestöliittos mentorskap i fråga om arbetskarriär är avsett för utbildade invandrare.
Via det kan du få en mentor som stöder dig när du söker arbete eller studieplats eller grundar ett företag.
Verksamheten är finskspråkig.
Mentorskap i fråga om arbetskarriärfinska _ engelska
Om du är under 30 år, kan du fråga råd om jobbsökande på Ohjaamo.
Ohjaamo är en rådgivningstjänst som är avsedd för unga vuxna.
Kompetenscentret Stadin osaamiskeskus (Stadin osaamiskeskus) förbereder invandrare för arbetsmarknaden och hjälper dem att hitta ett jobb eller en praktikplats.
Kompetenscentret erbjuder sina kunder bland annat undervisning i finska och yrkesutbildning.
Du kan bli kund vid Kompetenscentret via TE-byrån eller social -eller hälsovårdsverket.
Tjänsterna är avsedda för invandrare i Helsingfors som fyllt 17 år och har uppehållstillstånd.
Kompetenscenterfinska
Att grunda ett företag
Vid NewCo Helsinki får du råd och hjälp med att starta ett företag.
Du kan få personlig rådgivning om startande av ett företag på finska, svenska, engelska, ryska, arabiska, estniska, tyska och italienska.
NewCo Helsinki ordnar infomöten för invandrare om startande av ett företag.
Infomöten ordnas på finska, engelska, ryska, arabiska och estniska.
Infomötena är avgiftsfria.
Mer information och anmälan finns på NewCo Helsinkis webbplats.
NewCo Helsinki ordnar företagarutbildning på finska, engelska och ryska.
En del av kurserna är avsedda för personer som vill grunda ett företag, och en del för dem som redan har ett eget företag.
Kurser hålls på finska, engelska och ryska.
Mer information och anmälan finns på NewCo Helsinkis webbplats.
NewCo Helsinki ordnar också möten för nätverkande för nya företagare.
Från NewCo Helsinki får du också hjälp med att utveckla uppstartsföretag.
Om du har ett företag i Helsingfors kan du bli medlem i Helsingfors företagare (Helsingin Yrittäjät).
Helsingfors företagare är företagarnas intressebevakningsorganisation som erbjuder sina medlemmar till exempel utbildning, nätverk och rådgivning.
Mer information hittar du på organisationens webbplats.
Läs mer: Att grunda ett företag i Finland.
Som företagare till Finland:
Vilka tillstånd behöver du?(pdf, 384 kt)finska _ engelska
Guiden Bli företagare i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ turkiska _ kinesiska _ arabiska _ kurdiska
linkkiHelsingfors Företagare:
Företagarnas intressebevakningsorganisationfinska
Beskattning
Skattebyrån (verotoimisto) har ett serviceställe i centrala Helsingfors.
Kontaktuppgifter till skattebyråns andra serviceställen och telefonrådgivning hittar du på Skatteförvaltningens (verohallinto) webbplats.
Invandrare kan även sköta ärenden vid servicestället International House Helsinki.
På servicestället hjälper FPA:s och Skatteförvaltningens experter invandrare som kommer till Finland för att arbeta i frågor som rör beskattning och social trygghet.
Kontaktuppgifter till skattebyrån:
Alexandersgatan 9, 4:e våningen (Köpcentret Kluuvi)
Kontaktuppgifter till servicestället International House Helsinki:
Läs mer: Beskattning.
linkkiSkatteförvaltningen:
Kontaktuppgifter till skattebyråerfinska _ svenska _ engelska
IHH – serviceställe för dig som flyttar till Finland engelska
Var hittar jag jobb?
Hjälp med att söka jobb
Att grunda ett företag
Beskattning
Var hittar jag jobb?
TE-byråns tjänster
Du får hjälp med jobbsökningen på arbets- och näringsbyrån (Työ- ja elinkeinotoimisto), d.v.s. TE-byrån.
Om du är arbetslös och söker jobb, anmäl dig som arbetssökande till TE-byrån.
Du kan anmäla dig antingen via webbtjänsten eller personligen på TE-byrån.
Medborgare i ett EU-land, Norge, Island, Lichtenstein och Schweiz kan anmäla sig som arbetssökande via TE-byråns webbtjänst.
Medborgare från övriga länder måste anmäla sig personligen på TE-byrån.
Ta med dig identitetsbevis och uppehållstillstånd.
Du hittar information om TE-byråns tjänster på InfoFinlands sida Om du blir arbetslös.
Information om att söka jobb i Finland hittar du på InfoFinlands sida Var hittar jag jobb?
I Helsingfors finns tre TE-byråer.
Adress:
Kundgatan 3 A, 4:e våningen
Telefon: 0295 025 500
Öppettider: mån–fre kl. 9.00–16.00
Verksamhetsstället i centrum
Adress: Anttigatan 1, 2. våningen
Telefon: 0295 025 500
Öppettider: mån–fre kl. 9.00–16.00
Böle verksamhetsställe
Adress: Bangårdsvägen 7 (ingång via Loktorget)
Telefon: 0295 025 500
Öppettider: mån–fre kl. 9.00–16.00
Seure (Seure) är ett bemanningsbolag som erbjuder kortvariga jobb vid Helsingfors, Vanda, Esbo och Grankulla städer.
Jobben finns till exempel på skolor, daghem och sjukhus.
Arbetsplatser i kommunernafinska _ svenska _ engelska
Arbetslöshetsersättning
Information om att ansöka om arbetslöshetsersättning hittar du på InfoFinlands sida Arbetslöshetsförsäkring.
linkkiArbets- och näringsförvaltningen:
Länkar till jobbsajterfinska _ svenska _ engelska
linkkiArbets- och näringsministeriet:
Lediga jobbfinska _ svenska
linkkiTE-tjänster:
Videoklipp och broschyrer för invandrarefinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska
Hjälp med att söka jobb
Stadens tjänster för arbetslösa
Helsingfors stad hjälper arbetslösa helsingforsare att hitta jobb eller utbildning.
Om du behöver råd eller stöd för att hitta sysselsättning eller utbildning i finska språket, kontakta Helsingfors stads sysselsättningstjänster.
Stadens tjänster för arbetslösafinska _ svenska _ engelska
Integrationscentret Kotoutumiskeskus Monika hjälper arbetslösa invandrarkvinnor att hitta jobb.
Du kan få hjälp med att skriva din CV eller en jobbansökan, studera vardagsfinska och digitala färdigheter.
Luckan integration
Luckan Integration är en rådgivningstjänst som erbjuder invandrare personlig rådgivning, och ordnar bland annat möten och grupper i anslutning till arbetssökande.
Mötesspråket är engelska.
Råd om jobbsökningfinska _ svenska _ engelska _ spanska
Väestöliittos mentorskap i fråga om arbetskarriär är avsett för utbildade invandrare.
Via det kan du få en mentor som stöder dig när du söker arbete eller studieplats eller grundar ett företag.
Verksamheten är finskspråkig.
Mentorskap i fråga om arbetskarriärfinska _ engelska
Om du är under 30 år, kan du fråga råd om jobbsökande på Ohjaamo.
Ohjaamo är en rådgivningstjänst som är avsedd för unga vuxna.
Kompetenscentret Stadin osaamiskeskus (Stadin osaamiskeskus) förbereder invandrare för arbetsmarknaden och hjälper dem att hitta ett jobb eller en praktikplats.
Kompetenscentret erbjuder sina kunder bland annat undervisning i finska och yrkesutbildning.
Du kan bli kund vid Kompetenscentret via TE-byrån eller social -eller hälsovårdsverket.
Tjänsterna är avsedda för invandrare i Helsingfors som fyllt 17 år och har uppehållstillstånd.
Kompetenscenterfinska
Att grunda ett företag
Vid NewCo Helsinki får du råd och hjälp med att starta ett företag.
Du kan få personlig rådgivning om startande av ett företag på finska, svenska, engelska, ryska, arabiska, estniska, tyska och italienska.
NewCo Helsinki ordnar infomöten för invandrare om startande av ett företag.
Infomöten ordnas på finska, engelska, ryska, arabiska och estniska.
Infomötena är avgiftsfria.
Mer information och anmälan finns på NewCo Helsinkis webbplats.
NewCo Helsinki ordnar företagarutbildning på finska, engelska och ryska.
En del av kurserna är avsedda för personer som vill grunda ett företag, och en del för dem som redan har ett eget företag.
Kurser hålls på finska, engelska och ryska.
Mer information och anmälan finns på NewCo Helsinkis webbplats.
NewCo Helsinki ordnar också möten för nätverkande för nya företagare.
Från NewCo Helsinki får du också hjälp med att utveckla uppstartsföretag.
Om du har ett företag i Helsingfors kan du bli medlem i Helsingfors företagare (Helsingin Yrittäjät).
Helsingfors företagare är företagarnas intressebevakningsorganisation som erbjuder sina medlemmar till exempel utbildning, nätverk och rådgivning.
Mer information hittar du på organisationens webbplats.
Läs mer: Att grunda ett företag i Finland.
Som företagare till Finland:
Vilka tillstånd behöver du?(pdf, 384 kt)finska _ engelska
Guiden Bli företagare i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ turkiska _ kinesiska _ arabiska _ kurdiska
linkkiHelsingfors Företagare:
Företagarnas intressebevakningsorganisationfinska
Beskattning
Skattebyrån (verotoimisto) har ett serviceställe i centrala Helsingfors.
Kontaktuppgifter till skattebyråns andra serviceställen och telefonrådgivning hittar du på Skatteförvaltningens (verohallinto) webbplats.
Invandrare kan även sköta ärenden vid servicestället International House Helsinki.
På servicestället hjälper FPA:s och Skatteförvaltningens experter invandrare som kommer till Finland för att arbeta i frågor som rör beskattning och social trygghet.
Kontaktuppgifter till skattebyrån:
Alexandersgatan 9, 4:e våningen (Köpcentret Kluuvi)
Kontaktuppgifter till servicestället International House Helsinki:
Läs mer: Beskattning.
linkkiSkatteförvaltningen:
Kontaktuppgifter till skattebyråerfinska _ svenska _ engelska
IHH – serviceställe för dig som flyttar till Finland engelska
Rådgivning för och integration av invandrare
Inledande kartläggning och integrationsplan
Behöver du en tolk?
Rådgivning för och integration av invandrare
Helsingfors-info är ett rådgivningsställe där du kan fråga om aktuell information om Helsingfors, stadens tjänster, boendemöjligheter, arbete och studier.
Du kan även be om hjälp om du inte vet vilken myndighet du ska kontakta.
Helsinki-info erbjuder även digital rådgivning och hjälper dig med alla frågor kring invandring.
Helsinki-info betjänar på många olika språk per telefon, ansikte mot ansikte och elektroniskt.
Telefon: 09 310 11111, mån.–tors. kl. 9–16, fre. kl. 10–15
Tjänsteställen:
Centrumbiblioteket Oodi, adress: Tölöviksgatan 1
Elektroniskt:
Rådgivning på chattenfinska _ svenska _ engelska
Skicka en fråga eller ge oss responsfinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
Du kan få:
kostnadsfri rådgivning och information kring att flytta på flera olika språk
en finländsk personbeteckning, registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1-intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
I tjänsten medverkar Helsingfors-info, magistraten i Nyland, Skatteförvaltningen, FPA, NTM-centralen i Nyland, Pensionsskyddscentralen och Helsingforsregionens handelskammare.
Albertsgatan 25
IHH – serviceställe för dig som flyttar till Finland engelska
Webbappen IHH Service Advisor App engelska
Inledande kartläggning och integrationsplan
En anställd vid arbets- och näringsbyrån (työ- ja elinkeinotoimisto) upprättar en inledande kartläggning (alkukartoitus) och en integrationsplan (kotoutumissuunnitelma) tillsammans med dig när du registrerar dig som arbetssökande.
TE-byråerna i Östra centrum och Böle gör inledande kartläggningar.
För att få en inledande kartläggning gjord, ska du anmäla dig som arbetssökande via Internet på adressen te-palvelut.fi.
Du kan anmäla dig via Internet om du har finländska webbankkoder.
Du kan också anmäla dig till den inledande kartläggningen vid TE-byrån.
Adress:
Kundgatan 3 A, 4:e våningen
Telefonnummer: 0295 025 500
Öppettider: mån–fre kl. 9.00–16.00
Böle verksamhetsställe
Adress: Bangårdsvägen 7 (ingång via Loktorget)
Telefonnummer: 0295 025 500
Öppettider: mån–fre kl. 9.00–16.00
linkkiTE-tjänster:
Videoklipp och broschyrer för invandrarefinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska
Invandrarenheten
Invandrarenheten vid Helsingfors stads social- och hälsovårdstjänster hjälper invandrare bosatta i staden att integrera sig.
Invandrarenhetens tjänster är till exempel vägledning, rådgivning och inledande kartläggning.
Invandrarenheten hjälper också personer som fallit offer för människohandel.
Om du inte söker jobb men vill få den inledande kartläggningen och en integrationsplan upprättade, ska du kontakta invandrarenheten vid Helsingfors stads social- och hälsovårdstjänster.
Kontaktuppgifter till invandrarenheten:
Rådgivningsnumret för socialarbete (09) 310 37 577 mån–fre kl. 8.15–16
Invandrarenhetenfinska _ svenska _ engelska
Behöver du en tolk?
Om du inte kan finska eller svenska kan du anlita en tolk när du sköter ärenden med myndigheter.
I vissa fall får du en tolk via myndigheten.
Då är tolkningen kostnadsfri för dig.
Du kan i förväg fråga om tolkningen hos ifrågavarande myndighet eller få råd vid Helsingfors stads invandrarrådgivning.
Till exempel FPA och migrationsverket (Maahanmuuttovirasto) beställer i vissa fall en tolk för kunden.
Du kan anlita en tolk när som helst om du bokar tolken och betalar kostnaderna själv.
Också många företag erbjuder tolktjänster.
Du kan söka dessa företag till exempel med sökmotorer på Internet.
På webbplatsen för Finlands översättar- och tolkförbund finns en sökmotor med vilken du kan söka en tolk eller en översättare.
Tjänsterna vid Helsingforsregionens kontakttolkcentral är främst avsedda för myndigheter som arbetar med invandrare.
Läs mer: Behöver du en tolk?
linkkiFinlands översättar- och tolkförbund:
Sök tolk eller översättarefinska _ svenska _ engelska
linkkiHelsingforsnejdens kontakttolkcentral:
Tolkningfinska
Rådgivning för och integration av invandrare
Inledande kartläggning och integrationsplan
Behöver du en tolk?
Rådgivning för och integration av invandrare
Helsingfors-info är ett rådgivningsställe där du kan fråga om aktuell information om Helsingfors, stadens tjänster, boendemöjligheter, arbete och studier.
Du kan även be om hjälp om du inte vet vilken myndighet du ska kontakta.
Helsinki-info erbjuder även digital rådgivning och hjälper dig med alla frågor kring invandring.
Helsinki-info betjänar på många olika språk per telefon, ansikte mot ansikte och elektroniskt.
Telefon: 09 310 11111, mån.–tors. kl. 9–16, fre. kl. 10–15
Tjänsteställen:
Centrumbiblioteket Oodi, adress: Tölöviksgatan 1
Elektroniskt:
Rådgivning på chattenfinska _ svenska _ engelska
Skicka en fråga eller ge oss responsfinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
Du kan få:
kostnadsfri rådgivning och information kring att flytta på flera olika språk
registrering av uppehållsrätten om du är EU-medborgare
en finländsk personbeteckning, registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1-intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
I tjänsten medverkar Helsingfors-info, Esbo stad, magistraten i Nyland, Migrationsverket, Skatteförvaltningen, FPA, NTM-centralen i Nyland, Pensionsskyddscentralen, Helsingforsregionens handelskammare och Finlands Fackförbunds Centralorganisation FFC.
IHH – serviceställe för dig som flyttar till Finland engelska
Webbappen IHH Service Advisor App engelska
Inledande kartläggning och integrationsplan
En anställd vid arbets- och näringsbyrån (työ- ja elinkeinotoimisto) upprättar en inledande kartläggning (alkukartoitus) och en integrationsplan (kotoutumissuunnitelma) tillsammans med dig när du registrerar dig som arbetssökande.
TE-byråerna i Östra centrum och Böle gör inledande kartläggningar.
För att få en inledande kartläggning gjord, ska du anmäla dig som arbetssökande via Internet på adressen te-palvelut.fi.
Du kan anmäla dig via Internet om du har finländska webbankkoder.
Du kan också anmäla dig till den inledande kartläggningen vid TE-byrån.
Adress:
Kundgatan 3 A, 4:e våningen
Telefonnummer: 0295 025 500
Öppettider: mån–fre kl. 9.00–16.00
Böle verksamhetsställe
Adress: Bangårdsvägen 7 (ingång via Loktorget)
Telefonnummer: 0295 025 500
Öppettider: mån–fre kl. 9.00–16.00
linkkiTE-tjänster:
Videoklipp och broschyrer för invandrarefinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska
Invandrarenheten
Invandrarenheten vid Helsingfors stads social- och hälsovårdstjänster hjälper invandrare bosatta i staden att integrera sig.
Invandrarenhetens tjänster är till exempel vägledning, rådgivning och inledande kartläggning.
Invandrarenheten hjälper också personer som fallit offer för människohandel.
Om du inte söker jobb men vill få den inledande kartläggningen och en integrationsplan upprättade, ska du kontakta invandrarenheten vid Helsingfors stads social- och hälsovårdstjänster.
Kontaktuppgifter till invandrarenheten:
Rådgivningsnumret för socialarbete (09) 310 37 577 mån–fre kl. 8.15–16
Invandrarenhetenfinska _ svenska _ engelska
Behöver du en tolk?
Om du inte kan finska eller svenska kan du anlita en tolk när du sköter ärenden med myndigheter.
I vissa fall får du en tolk via myndigheten.
Då är tolkningen kostnadsfri för dig.
Du kan i förväg fråga om tolkningen hos ifrågavarande myndighet eller få råd vid Helsingfors stads invandrarrådgivning.
Till exempel FPA och migrationsverket (Maahanmuuttovirasto) beställer i vissa fall en tolk för kunden.
Du kan anlita en tolk när som helst om du bokar tolken och betalar kostnaderna själv.
Också många företag erbjuder tolktjänster.
Du kan söka dessa företag till exempel med sökmotorer på Internet.
På webbplatsen för Finlands översättar- och tolkförbund finns en sökmotor med vilken du kan söka en tolk eller en översättare.
Tjänsterna vid Helsingforsregionens kontakttolkcentral är främst avsedda för myndigheter som arbetar med invandrare.
Läs mer: Behöver du en tolk?
linkkiFinlands översättar- och tolkförbund:
Sök tolk eller översättarefinska _ svenska _ engelska
linkkiHelsingforsnejdens kontakttolkcentral:
Tolkningfinska
Rådgivning för och integration av invandrare
Inledande kartläggning och integrationsplan
Behöver du en tolk?
Rådgivning för och integration av invandrare
Helsingfors-info är ett rådgivningsställe där du kan fråga om aktuell information om Helsingfors, stadens tjänster, boendemöjligheter, arbete och studier.
Du kan även be om hjälp om du inte vet vilken myndighet du ska kontakta.
Helsinki-info erbjuder även digital rådgivning och hjälper dig med alla frågor kring invandring.
Helsinki-info betjänar på många olika språk per telefon, ansikte mot ansikte och elektroniskt.
Telefon: 09 310 11111, mån.–tors. kl. 9–16, fre. kl. 10–15
Tjänsteställen:
Centrumbiblioteket Oodi, adress: Tölöviksgatan 4
Elektroniskt:
Rådgivning på chattenfinska _ svenska _ engelska
Skicka en fråga eller ge oss responsfinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
Du kan få:
kostnadsfri rådgivning och information kring att flytta på flera olika språk
registrering av uppehållsrätten om du är EU-medborgare
en finländsk personbeteckning, registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1-intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
I tjänsten medverkar Helsingfors-info, Esbo stad, magistraten i Nyland, Migrationsverket, Skatteförvaltningen, FPA, NTM-centralen i Nyland, Pensionsskyddscentralen, Helsingforsregionens handelskammare och Finlands Fackförbunds Centralorganisation FFC.
IHH – serviceställe för dig som flyttar till Finland engelska
Webbappen IHH Service Advisor App engelska
Inledande kartläggning och integrationsplan
En anställd vid arbets- och näringsbyrån (työ- ja elinkeinotoimisto) upprättar en inledande kartläggning (alkukartoitus) och en integrationsplan (kotoutumissuunnitelma) tillsammans med dig när du registrerar dig som arbetssökande.
TE-byråerna i Östra centrum och Böle gör inledande kartläggningar.
För att få en inledande kartläggning gjord, ska du anmäla dig som arbetssökande via Internet på adressen te-palvelut.fi.
Du kan anmäla dig via Internet om du har finländska webbankkoder.
Du kan också anmäla dig till den inledande kartläggningen vid TE-byrån.
Adress:
Kundgatan 3 A, 4:e våningen
Telefonnummer: 0295 025 500
Öppettider: mån–fre kl. 9.00–16.00
Böle verksamhetsställe
Adress: Bangårdsvägen 7 (ingång via Loktorget)
Telefonnummer: 0295 025 500
Öppettider: mån–fre kl. 9.00–16.00
linkkiTE-tjänster:
Videoklipp och broschyrer för invandrarefinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska
Invandrarenheten
Invandrarenheten vid Helsingfors stads social- och hälsovårdstjänster hjälper invandrare bosatta i staden att integrera sig.
Invandrarenhetens tjänster är till exempel vägledning, rådgivning och inledande kartläggning.
Invandrarenheten hjälper också personer som fallit offer för människohandel.
Om du inte söker jobb men vill få den inledande kartläggningen och en integrationsplan upprättade, ska du kontakta invandrarenheten vid Helsingfors stads social- och hälsovårdstjänster.
Kontaktuppgifter till invandrarenheten:
Rådgivningsnumret för socialarbete (09) 310 37 577 mån–fre kl. 8.15–16
Invandrarenhetenfinska _ svenska _ engelska
Behöver du en tolk?
Om du inte kan finska eller svenska kan du anlita en tolk när du sköter ärenden med myndigheter.
Till exempel FPA (Kela) och Migrationsverket (Maahanmuuttovirasto) bokar i vissa situationer en tolk för klienten.
Då behöver du inte betala för tolken.
Fråga alltid i förväg om tolk hos den aktuella myndigheten eller be om råd vid Helsinki-info.
Om du själv bokar tolken och betalar kostnaderna kan du anlita en tolk när som helst.
I Helsingfors erbjuds tolktjänster av flera företag.
Du kan söka dessa företag på till exempel internet.
Till exempel A-tulkkaus förmedlar i Helsingforsregionen kontakttolkar för tillfällen där du uträttar ärenden hos myndigheter.
Du kan söka en tolk eller översättare med hjälp av sökfunktionen på Finlands översättar- och tolkförbunds webbplats.
Läs mer: Behöver du en tolk?
linkkiFinlands översättar- och tolkförbund:
Sök tolk eller översättarefinska _ svenska _ engelska
Tolkningfinska
Tillståndsärenden
På Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU-medborgarens uppehållsrätt.
Migrationsverkets tjänsteställe i Helsingfors :
Göksgränd 3A
Du kan också ansöka om många slags uppehållstillstånd och EU-registrering på internet i tjänsten Enter Finland.
Om du inte är van vid att använda en dator, fyll i en ansökan på papper och lämna in den på Migrationsverkets tjänsteställe.
Dät är alltid bra att boka en tid i förväg på tjänstestället.
Du kan boka en tid på Migrationsverkets tidsbokningstjänst.
Observera att tjänstestället inte kan ge rådgivning om tillståndsärenden.
Läs mer: Flytta till Finland.
Elektronisk tidsbokningfinska _ svenska _ engelska
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Registrering som invånare
När du flyttar ditt stadigvarande boende till Helsingfors, ska du registrera dig som invånare i kommunen.
Du kan registrera dig vid Helsingfors magistrat.
Kontaktuppgifter till magistraten i Helsingfors:
Magistraten i Nyland, servicestället i Helsingfors
Albertsgatan 25
Tfn 029 55 39391
När du besöker magistraten ska du ta med dig
legitimation (till exempel pass)
uppehållstillstånd och uppehållskort (om du behöver uppehållstillstånd i Finland)
registreringsintyg över uppehållsrätten (oleskeluoikeuden rekisteröintitodistus) (om du är medborgare i ett EU-land)
äktenskapsintyg
dina barns födelseattester.
Observera att utländska handlingar ska vara legaliserade.
På magistratens webbplats finns mer information om registreringen av utlänningar.
Läs mer: Registrering som invånare.
Registrering av utlänningarfinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
Du kan få:
kostnadsfri rådgivning och information kring att flytta på flera olika språk
en finländsk personbeteckning, registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1-intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
I tjänsten medverkar Helsingfors-info, magistraten i Nyland, Skatteförvaltningen, FPA, NTM-centralen i Nyland, Pensionsskyddscentralen och Helsingforsregionens handelskammare.
Adress
Albertsgatan 25
IHH – serviceställe för dig som flyttar till Finland engelska
Webbappen IHH Service Advisor App engelska
Tjänster för invandrarefinska _ svenska _ engelska
Tillståndsärenden
På Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU-medborgarens uppehållsrätt.
Migrationsverkets tjänsteställe i Helsingfors :
Göksgränd 3A
Du kan också ansöka om många slags uppehållstillstånd och EU-registrering på internet i tjänsten Enter Finland.
Om du inte är van vid att använda en dator, fyll i en ansökan på papper och lämna in den på Migrationsverkets tjänsteställe.
Dät är alltid bra att boka en tid i förväg på tjänstestället.
Du kan boka en tid på Migrationsverkets tidsbokningstjänst.
Observera att tjänstestället inte kan ge rådgivning om tillståndsärenden.
Läs mer: Flytta till Finland.
Elektronisk tidsbokningfinska _ svenska _ engelska
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Registrering som invånare
När du flyttar ditt stadigvarande boende till Helsingfors, ska du registrera dig som invånare i kommunen.
Du kan registrera dig vid Helsingfors magistrat.
Kontaktuppgifter till magistraten i Helsingfors:
Magistraten i Nyland, servicestället i Helsingfors
Tfn 029 55 39391
När du besöker magistraten ska du ta med dig
legitimation (till exempel pass)
uppehållstillstånd och uppehållskort (om du behöver uppehållstillstånd i Finland)
registreringsintyg över uppehållsrätten (oleskeluoikeuden rekisteröintitodistus) (om du är medborgare i ett EU-land)
äktenskapsintyg
dina barns födelseattester.
Observera att utländska handlingar ska vara legaliserade.
På magistratens webbplats finns mer information om registreringen av utlänningar.
Läs mer: Registrering som invånare.
Registrering av utlänningarfinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
Du kan få:
kostnadsfri rådgivning och information kring att flytta på flera olika språk
registrering av uppehållsrätten om du är EU-medborgare
en finländsk personbeteckning, registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1-intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
I tjänsten medverkar Helsingfors-info, Esbo stad, magistraten i Nyland, Migrationsverket, Skatteförvaltningen, FPA, NTM-centralen i Nyland, Pensionsskyddscentralen, Helsingforsregionens handelskammare och Finlands Fackförbunds Centralorganisation FFC.
Adress
IHH – serviceställe för dig som flyttar till Finland engelska
Webbappen IHH Service Advisor App engelska
Tjänster för invandrarefinska _ svenska _ engelska
Tillståndsärenden
På Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU-medborgarens uppehållsrätt.
Migrationsverkets tjänsteställe i Helsingfors :
Göksgränd 3A
Du kan också ansöka om många slags uppehållstillstånd och EU-registrering på internet i tjänsten Enter Finland.
Om du inte är van vid att använda en dator, fyll i en ansökan på papper och lämna in den på Migrationsverkets tjänsteställe.
Dät är alltid bra att boka en tid i förväg på tjänstestället.
Du kan boka en tid på Migrationsverkets tidsbokningstjänst.
Observera att tjänstestället inte kan ge rådgivning om tillståndsärenden.
Läs mer: Flytta till Finland.
Elektronisk tidsbokningfinska _ svenska _ engelska
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Registrering som invånare
När du flyttar ditt stadigvarande boende till Helsingfors, ska du registrera dig som invånare i kommunen.
Du kan registrera dig vid Helsingfors magistrat.
Kontaktuppgifter till magistraten i Helsingfors:
Magistraten i Nyland, servicestället i Helsingfors
Tfn 029 55 39391
När du besöker magistraten ska du ta med dig
legitimation (till exempel pass)
uppehållstillstånd och uppehållskort (om du behöver uppehållstillstånd i Finland)
registreringsintyg över uppehållsrätten (oleskeluoikeuden rekisteröintitodistus) (om du är medborgare i ett EU-land)
äktenskapsintyg
dina barns födelseattester.
Observera att utländska handlingar ska vara legaliserade.
På magistratens webbplats finns mer information om registreringen av utlänningar.
Läs mer: Registrering som invånare.
Registrering av utlänningarfinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
Du kan få:
kostnadsfri rådgivning och information kring att flytta på flera olika språk
registrering av uppehållsrätten om du är EU-medborgare
en finländsk personbeteckning, registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1-intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
I tjänsten medverkar Helsingfors-info, Esbo stad, magistraten i Nyland, Migrationsverket, Skatteförvaltningen, FPA, NTM-centralen i Nyland, Pensionsskyddscentralen, Helsingforsregionens handelskammare och Finlands Fackförbunds Centralorganisation FFC.
Adress
IHH – serviceställe för dig som flyttar till Finland engelska
Webbappen IHH Service Advisor App engelska
Tjänster för invandrarefinska _ svenska _ engelska
Var ligger närmaste magistrat, hälsostation eller bibliotek?
På InfoFinlands sida Städer hittar du information om de lokala tjänsterna i InfoFinlands medlemskommuner.
Var ligger närmaste magistrat, hälsostation eller bibliotek?
På InfoFinlands sida Städer hittar du information om de lokala tjänsterna i InfoFinlands medlemskommuner.
Var ligger närmaste magistrat, hälsostation eller bibliotek?
På InfoFinlands sida Städer hittar du information om de lokala tjänsterna i InfoFinlands medlemskommuner.
Dessa telefontjänster upprätthålls av olika myndigheter och organisationer.
InfoFinland-tjänsten ger dock ingen rådgivning och du kan inte ringa InfoFinland.
Information om offentliga tjänster
Information om den sociala tryggheten i Finland
Juridisk rådgivning
Tjänster för arbetstagare och företagare
Stöd vid ekonomiska problem
Diskriminering och rasism
Stöd för familjer
Rådgivning i frågor om hälsa
Hjälp med att få slut på våld
Hjälp till offer för människohandel
Information om offentliga tjänster
Behöver du information om offentliga tjänster eller hjälp med dem?
Statskontorets tjänsten Medborgarrådgivning hjälper medborgarna att snabbt och smidigt hitta rätt myndighet eller elektronisk myndighetstjänst.
Medborgarrådgivningen guidar dig till den rätta tjänsten, hjälper med digital ärendehantering och besvarar allmänna frågor om de offentliga tjänsterna.
Du kan inte anhängiggöra myndighetsärenden hos Medborgarrådgivningen – däremot så styr vi dig till rätta myndighet.
Tjänsten ger service på finska, svenska och engelska.
Ring 0295 000
Mån–fre 8–21
lör 9–15
Information om den sociala tryggheten i Finland
FPA:s telefontjänst
Ärenden rörande den sociala tryggheten när du flyttar till Finland eller utomlands:
020 634 0200 (på finska och på engelska)
FPA ger rådgivning på telefon även på ryska och arabiska.
Tjänsten är avsedd för personer som har bristfälliga kunskaper i finska, svenska eller engelska.
Rysktalande klienter: 020 634 4901
Arabisktalande klienter: 020 634 4902
Om det är kö till kundtjänsten, kan du även lämna ett meddelande och bli uppringd.
Du kan även boka en telefontid vid FPA.
Du kan boka tiden via telefontjänsten eller på FPA:s webbplats.
När du har bokat en telefontid, ringer FPA:s servicerådgivare upp dig vid överenskommen tidpunkt.
Om du behöver en tolk, ska du uppge detta när du bokar tiden.
Om du behöver en tolk, ska du boka din telefontid minst en vecka i förväg.
Vanligtvis går det inte att få tag på en tolk snabbare än så.
FPA beställer tolken.
Juridisk rådgivning
Flyktingrådgivningen r.f.
Flyktingrådgivningen ger juridisk hjälp och rådgivning för asylsökande, flyktingar och andra utlänningar.
Rådgivning ges på finska och engelska.
09 2313 9325 (mån.–fre. ll. 10–12)
Rådgivning för papperslösa utlänningar: 045 2377 104 (måndagar kl. 14–16).
Brottsofferjouren
Hjälptelefon 116 006
Telefonrådgivning av en jurist 0800 161 177
Brottsofferjouren (RIKU) har till uppgift att främja brottsoffrets ställning samt ställningen för deras närstående och brottsmålsvittnen.
Du kan ringa brottsofferjouren om du eller en närstående har blivit utsatt för ett brott eller om du har bevittnat ett brott.
Du behöver inte uppge ditt namn när du ringer.
På hjälptelefonen får du stöd och vid behov råd om var du kan få hjälp.
På juristernas telefonrådgivning får du information om dina juridiska rättigheter.
Tjänster för arbetstagare och företagare
Anställningsrådgivning för invandrare
Om du har frågor om eller problem med din anställning, kan du kontakta anställningsrådgivningen för invandrare.
Rådgivningen ges av Finlands Fackförbunds Centralorganisation FFC.
Du kan få rådgivning även om du inte är medlem i fackförbundet.
En jurist svarar på dina frågor till exempel om arbetsavtal, lön eller arbetstider.
Den kostnadsfria rådgivningen ges på finska och engelska.
Anställningsrådgivningen har öppet måndag–torsdag klockan 9–11 och 12–15.
Telefon: 0800 414 004
Arbets- och näringstjänsten
Rådgivning på finska : 0295 025 500
Rådgivning på svenska: 0295 025 510
Rådgivning på engelska: 0295 020 713
I telefontjänsten får du rådgivning om tjänsterna vid arbets- och näringsbyrån.
Du får även handledning om hur du sköter ärenden och rådgivning om uppehållstillstånd för arbetstagare.
FöretagsFinland
Telefontjänst: 0295 020 500
På FöretagsFinlands telefontjänst får du information, handledning och rådgivning kring start av företagsverksamhet och de offentliga företagstjänsterna.
Skatteförvaltningen
Rådgivning på engelska om beskattningen i Finland: 029 497 050
Tjänsten Internationell personbeskattning tillhandahåller information om beskattningen av inkomster från utlandet och beskattningen av arbete utomlands samt hur en flytt utomlands påverkar beskattningen.
Tjänsten ger även råd om beskattningen för personer som kommer från utlandet till Finland för att arbeta och skyldigheterna för dem som betalar skatter i internationella sammanhang.
Stöd vid ekonomiska problem
Skuldlinjen
Telefonrådgivning: 0800 9 8009
Du kan ringa skuldlinjen kostnadsfritt från hela Finland och diskutera anonymt dina egna eller en närstående persons ekonomiska bekymmer.
Svårigheterna kan vara stora eller små.
Under samtalet får den som ringer hjälp med att kartlägga sin situation, råd och vid behov vägledning till något ställe där man kan få hjälp.
Diskriminering och rasism
Diskrimineringsombudsmannen
Du kan kontakta diskrimineringsombudsmannen byrå om du har råkat ut för diskriminering eller upplever att du har bemötts rasistiskt eller osakligt på grund av ditt etniska ursprung eller för att du är utlänning.
På telefonen ger den jourhavande överinspektören råd om hur du kan utreda saken och kommer överens om eventuella fortsatta åtgärder för att föra saken vidare.
På telefon kan vi betjäna dig på finska, svenska och engelska.
Jämställdhetsombudsmannen
Telefonrådgivning: 0295 666 842
Om du misstänker att en arbetsgivare, en läroanstalt eller någon annan instans har diskriminerat dig på grund av ditt kön och brutit mot lagen om jämställdhet mellan kvinnor och män, kan du be jämställdhetsombudsmannen om råd och anvisningar samt hjälp med att utreda ärendet.
Jämställdhetsombudsmannen ger dig även övrig information om lagen om jämställdhet mellan kvinnor och män.
Stöd för familjer
Kostnadsfri rådgivning för invandrare i frågor som rör familjens välbefinnande eller fostran av barn.
Rådgivning på olika språk:
Ryska och engelska: 050 325 7173
Rådgivning i frågor om hälsa
Föreningen för mental hälsa i Finland
Riksomfattande kristelefon: 010 195 202
Kristelefon för arabisktalande: 040 195 8202.
Du kan även ringa och prata på engelska.
Föreningen för mental hälsa i Finlands kristelefon erbjuder omedelbar samtalshjälp för människor i kris och deras närstående.
Samtalen besvaras av krisarbetare och utbildade frivilliga stödpersoner.
Du behöver inte uppge ditt namn när du ringer.
På kristelefonen kan du prata om en oväntad händelse eller en svår livssituation i en tillåtande och stödande atmosfär.
Stödcentret Hilma för handikappade invandrare
Du får handledning och råd om att ansöka om socialtjänster och förmåner avsedda för handikappade samt med att fylla i blanketter.
Du kan också fråga om möjligheterna till rehabilitering, studier, arbete och hobbyer.
Telefonen betjänar på finska, svenska, engelska och tyska.
Förgiftningar, vård och förebyggande: (09) 471 977
Vid Giftinformationscentralen kan du fråga om förebyggande och vård av akuta förgiftningar.
Hjälp med att få slut på våld
Nollalinja
Tfn 080 005 005
Öppet: varje dag
Nollalinja är en hjälptelefon som du kan ringa om du har blivit utsatt för våld i familjen, sexuellt våld eller hot om våld.
Du kan ringa när som helst.
Medarbetarna pratar finska, svenska och engelska.
Samtal till Nollalinja är kostnadsfria och de syns inte i telefonräkningen.
Du behöver inte uppge ditt namn när du ringer.
Nollalinja är avsedd för både kvinnor och män.
Manslinjen
Hjälptelefon: (09) 276 62 899
Manslinjen är en tjänst som hjälper invandrarmän som har utövat våld eller är oroliga för att de kommer att utöva våld mot en närstående människa eller någon i familjen.
Vi ger stöd och råd åt invandrarkvinnor som blivit utsatt för våld eller lever under hot om våld.
Du behöver inte uppge ditt namn när du ringer.
Maria Akademi
Öppna linjen: 09 7562 2260
Stöd och hjälp för kvinnor som utövar våld eller är oroliga för att de kommer att göra det.
Samtalen är konfidentiella.
Den öppna linjen betjänar på finska, svenska och engelska.
Hjälp till offer för människohandel
Nationellt hjälpsystem till offer för människohandel i Finland
Hjälptelefon: 02954 63177
Ta kontakt med hjälpsystemet till offer för människohandel om du upplever att du blivit offer för utnyttjande.
Du får hjälp även om du
vistas i landet illegalt
inte har identitetsbevis eller pass
blir utsatt för hot, eller om en närstående till dig blir utsatt för hot
endast talar ditt modersmål
står i skuld till någon
Dessa telefontjänster upprätthålls av olika myndigheter och organisationer.
InfoFinland-tjänsten ger dock ingen rådgivning och du kan inte ringa InfoFinland.
Information om offentliga tjänster
Information om den sociala tryggheten i Finland
Juridisk rådgivning
Tjänster för arbetstagare och företagare
Stöd vid ekonomiska problem
Diskriminering och rasism
Stöd för familjer
Rådgivning i frågor om hälsa
Hjälp med att få slut på våld
Hjälp till offer för människohandel
Information om offentliga tjänster
Behöver du information om offentliga tjänster eller hjälp med dem?
Statskontorets tjänsten Medborgarrådgivning hjälper medborgarna att snabbt och smidigt hitta rätt myndighet eller elektronisk myndighetstjänst.
Medborgarrådgivningen guidar dig till den rätta tjänsten, hjälper med digital ärendehantering och besvarar allmänna frågor om de offentliga tjänsterna.
Du kan inte anhängiggöra myndighetsärenden hos Medborgarrådgivningen – däremot så styr vi dig till rätta myndighet.
Tjänsten ger service på finska, svenska och engelska.
Ring 0295 000
Mån–fre 8–21
lör 9–15
Information om den sociala tryggheten i Finland
FPA:s telefontjänst
Ärenden rörande den sociala tryggheten när du flyttar till Finland eller utomlands:
020 634 0200 (på finska och på engelska)
FPA ger rådgivning på telefon även på ryska och arabiska.
Tjänsten är avsedd för personer som har bristfälliga kunskaper i finska, svenska eller engelska.
Rysktalande klienter: 020 634 4901
Arabisktalande klienter: 020 634 4902
Om det är kö till kundtjänsten, kan du även lämna ett meddelande och bli uppringd.
Du kan även boka en telefontid vid FPA.
Du kan boka tiden via telefontjänsten eller på FPA:s webbplats.
När du har bokat en telefontid, ringer FPA:s servicerådgivare upp dig vid överenskommen tidpunkt.
Om du behöver en tolk, ska du uppge detta när du bokar tiden.
Om du behöver en tolk, ska du boka din telefontid minst en vecka i förväg.
Vanligtvis går det inte att få tag på en tolk snabbare än så.
FPA beställer tolken.
Juridisk rådgivning
Flyktingrådgivningen r.f.
Flyktingrådgivningen ger juridisk hjälp och rådgivning för asylsökande, flyktingar och andra utlänningar.
Rådgivning ges på finska och engelska.
09 2313 9325 (mån.–fre. ll. 10–12)
Rådgivning för papperslösa utlänningar: 045 2377 104 (måndagar kl. 14–16).
Brottsofferjouren
Hjälptelefon 116 006
Telefonrådgivning av en jurist 0800 161 177
Brottsofferjouren (RIKU) har till uppgift att främja brottsoffrets ställning samt ställningen för deras närstående och brottsmålsvittnen.
Du kan ringa brottsofferjouren om du eller en närstående har blivit utsatt för ett brott eller om du har bevittnat ett brott.
Du behöver inte uppge ditt namn när du ringer.
På hjälptelefonen får du stöd och vid behov råd om var du kan få hjälp.
På juristernas telefonrådgivning får du information om dina juridiska rättigheter.
Tjänster för arbetstagare och företagare
Anställningsrådgivning för invandrare
Om du har frågor om eller problem med din anställning, kan du kontakta anställningsrådgivningen för invandrare.
Rådgivningen ges av Finlands Fackförbunds Centralorganisation FFC.
Du kan få rådgivning även om du inte är medlem i fackförbundet.
En jurist svarar på dina frågor till exempel om arbetsavtal, lön eller arbetstider.
Den kostnadsfria rådgivningen ges på finska och engelska.
Anställningsrådgivningen har öppet måndag–torsdag klockan 9–11 och 12–15.
Telefon: 0800 414 004
Arbets- och näringstjänsten
Rådgivning på finska : 0295 025 500
Rådgivning på svenska: 0295 025 510
Rådgivning på engelska: 0295 020 713
I telefontjänsten får du rådgivning om tjänsterna vid arbets- och näringsbyrån.
Du får även handledning om hur du sköter ärenden och rådgivning om uppehållstillstånd för arbetstagare.
FöretagsFinland
Telefontjänst: 0295 020 500
På FöretagsFinlands telefontjänst får du information, handledning och rådgivning kring start av företagsverksamhet och de offentliga företagstjänsterna.
Skatteförvaltningen
Rådgivning på engelska om beskattningen i Finland: 029 497 050
Tjänsten Internationell personbeskattning tillhandahåller information om beskattningen av inkomster från utlandet och beskattningen av arbete utomlands samt hur en flytt utomlands påverkar beskattningen.
Tjänsten ger även råd om beskattningen för personer som kommer från utlandet till Finland för att arbeta och skyldigheterna för dem som betalar skatter i internationella sammanhang.
Stöd vid ekonomiska problem
Skuldlinjen
Telefonrådgivning: 0800 9 8009
Du kan ringa skuldlinjen kostnadsfritt från hela Finland och diskutera anonymt dina egna eller en närstående persons ekonomiska bekymmer.
Svårigheterna kan vara stora eller små.
Under samtalet får den som ringer hjälp med att kartlägga sin situation, råd och vid behov vägledning till något ställe där man kan få hjälp.
Diskriminering och rasism
Diskrimineringsombudsmannen
Du kan kontakta diskrimineringsombudsmannen byrå om du har råkat ut för diskriminering eller upplever att du har bemötts rasistiskt eller osakligt på grund av ditt etniska ursprung eller för att du är utlänning.
På telefonen ger den jourhavande överinspektören råd om hur du kan utreda saken och kommer överens om eventuella fortsatta åtgärder för att föra saken vidare.
På telefon kan vi betjäna dig på finska, svenska och engelska.
Jämställdhetsombudsmannen
Telefonrådgivning: 0295 666 842
Om du misstänker att en arbetsgivare, en läroanstalt eller någon annan instans har diskriminerat dig på grund av ditt kön och brutit mot lagen om jämställdhet mellan kvinnor och män, kan du be jämställdhetsombudsmannen om råd och anvisningar samt hjälp med att utreda ärendet.
Jämställdhetsombudsmannen ger dig även övrig information om lagen om jämställdhet mellan kvinnor och män.
Stöd för familjer
Kostnadsfri rådgivning för invandrare i frågor som rör familjens välbefinnande eller fostran av barn.
Rådgivning på olika språk:
Ryska och engelska: 050 325 7173
Rådgivning i frågor om hälsa
Föreningen för mental hälsa i Finland
Riksomfattande kristelefon: 010 195 202
Kristelefon för arabisktalande: 040 195 8202.
Du kan även ringa och prata på engelska.
Föreningen för mental hälsa i Finlands kristelefon erbjuder omedelbar samtalshjälp för människor i kris och deras närstående.
Samtalen besvaras av krisarbetare och utbildade frivilliga stödpersoner.
Du behöver inte uppge ditt namn när du ringer.
På kristelefonen kan du prata om en oväntad händelse eller en svår livssituation i en tillåtande och stödande atmosfär.
Stödcentret Hilma för handikappade invandrare
Du får handledning och råd om att ansöka om socialtjänster och förmåner avsedda för handikappade samt med att fylla i blanketter.
Du kan också fråga om möjligheterna till rehabilitering, studier, arbete och hobbyer.
Telefonen betjänar på finska, svenska, engelska och tyska.
Förgiftningar, vård och förebyggande: (09) 471 977
Vid Giftinformationscentralen kan du fråga om förebyggande och vård av akuta förgiftningar.
Hjälp med att få slut på våld
Nollalinja
Tfn 080 005 005
Öppet: varje dag
Nollalinja är en hjälptelefon som du kan ringa om du har blivit utsatt för våld i familjen, sexuellt våld eller hot om våld.
Du kan ringa när som helst.
Medarbetarna pratar finska, svenska och engelska.
Samtal till Nollalinja är kostnadsfria och de syns inte i telefonräkningen.
Du behöver inte uppge ditt namn när du ringer.
Nollalinja är avsedd för både kvinnor och män.
Manslinjen
Hjälptelefon: (09) 276 62 899
Manslinjen är en tjänst som hjälper invandrarmän som har utövat våld eller är oroliga för att de kommer att utöva våld mot en närstående människa eller någon i familjen.
Vi ger stöd och råd åt invandrarkvinnor som blivit utsatt för våld eller lever under hot om våld.
Du behöver inte uppge ditt namn när du ringer.
Maria Akademi
Öppna linjen: 09 7562 2260
Stöd och hjälp för kvinnor som utövar våld eller är oroliga för att de kommer att göra det.
Samtalen är konfidentiella.
Den öppna linjen betjänar på finska, svenska och engelska.
Hjälp till offer för människohandel
Nationellt hjälpsystem till offer för människohandel i Finland
Hjälptelefon: 02954 63177
Ta kontakt med hjälpsystemet till offer för människohandel om du upplever att du blivit offer för utnyttjande.
Du får hjälp även om du
vistas i landet illegalt
inte har identitetsbevis eller pass
blir utsatt för hot, eller om en närstående till dig blir utsatt för hot
endast talar ditt modersmål
står i skuld till någon
Dessa telefontjänster upprätthålls av olika myndigheter och organisationer.
InfoFinland-tjänsten ger dock ingen rådgivning och du kan inte ringa InfoFinland.
Information om offentliga tjänster
Information om den sociala tryggheten i Finland
Juridisk rådgivning
Tjänster för arbetstagare och företagare
Stöd vid ekonomiska problem
Diskriminering och rasism
Stöd för familjer
Rådgivning i frågor om hälsa
Hjälp med att få slut på våld
Hjälp till offer för människohandel
Information om offentliga tjänster
Behöver du information om offentliga tjänster eller hjälp med dem?
Statskontorets tjänsten Medborgarrådgivning hjälper medborgarna att snabbt och smidigt hitta rätt myndighet eller elektronisk myndighetstjänst.
Medborgarrådgivningen guidar dig till den rätta tjänsten, hjälper med digital ärendehantering och besvarar allmänna frågor om de offentliga tjänsterna.
Du kan inte anhängiggöra myndighetsärenden hos Medborgarrådgivningen – däremot så styr vi dig till rätta myndighet.
Tjänsten ger service på finska, svenska och engelska.
Ring 0295 000
Mån–fre 8–21
lör 9–15
Information om den sociala tryggheten i Finland
FPA:s telefontjänst
Ärenden rörande den sociala tryggheten när du flyttar till Finland eller utomlands:
020 634 0200 (på finska och på engelska)
FPA:s telefontjänst är öppen måndag till fredag klockan 9–16.
FPA ger rådgivning på telefon även på ryska, arabiska och somaliska.
Tjänsten är avsedd för personer som har bristfälliga kunskaper i finska, svenska eller engelska.
Rysktalande klienter: 020 634 4901 (mån.–fre. kl. 10–12 och 13–15)
Arabisktalande klienter: 020 634 4902 (tis.–tors. kl. 10–12 och 13–15)
Somalisktalande klienter 020 634 4905 (mån. och fre. 10–12 och 13–15)
Du kan även boka en telefontid vid FPA.
Du kan boka tiden via telefontjänsten eller på FPA:s webbplats.
När du har bokat en telefontid, ringer FPA:s servicerådgivare upp dig vid överenskommen tidpunkt.
Om du behöver en tolk, ska du uppge detta när du bokar tiden.
Om du behöver en tolk, ska du boka din telefontid minst en vecka i förväg.
Vanligtvis går det inte att få tag på en tolk snabbare än så.
FPA beställer tolken.
Juridisk rådgivning
Flyktingrådgivningen r.f.
Flyktingrådgivningen ger juridisk hjälp och rådgivning för asylsökande, flyktingar och andra utlänningar.
Rådgivning ges på finska och engelska.
09 2313 9325 (mån.–fre. ll. 10–12)
Rådgivning för papperslösa utlänningar: 045 2377 104 (måndagar kl. 14–16).
Brottsofferjouren
Hjälptelefon 116 006
Telefonrådgivning av en jurist 0800 161 177
Brottsofferjouren (RIKU) har till uppgift att främja brottsoffrets ställning samt ställningen för deras närstående och brottsmålsvittnen.
Du kan ringa brottsofferjouren om du eller en närstående har blivit utsatt för ett brott eller om du har bevittnat ett brott.
Du behöver inte uppge ditt namn när du ringer.
På hjälptelefonen får du stöd och vid behov råd om var du kan få hjälp.
På juristernas telefonrådgivning får du information om dina juridiska rättigheter.
Tjänster för arbetstagare och företagare
Anställningsrådgivning för invandrare
Om du har frågor om eller problem med din anställning, kan du kontakta anställningsrådgivningen för invandrare.
Rådgivningen ges av Finlands Fackförbunds Centralorganisation FFC.
Du kan få rådgivning även om du inte är medlem i fackförbundet.
En jurist svarar på dina frågor till exempel om arbetsavtal, lön eller arbetstider.
Den kostnadsfria rådgivningen ges på finska och engelska.
Anställningsrådgivningen har öppet måndag–torsdag klockan 9–11 och 12–15.
Telefon: 0800 414 004
Arbets- och näringstjänsten
Rådgivning på finska : 0295 025 500
Rådgivning på svenska: 0295 025 510
Rådgivning på engelska: 0295 020 713
I telefontjänsten får du rådgivning om tjänsterna vid arbets- och näringsbyrån.
Du får även handledning om hur du sköter ärenden och rådgivning om uppehållstillstånd för arbetstagare.
FöretagsFinland
Telefontjänst: 0295 020 500
På FöretagsFinlands telefontjänst får du information, handledning och rådgivning kring start av företagsverksamhet och de offentliga företagstjänsterna.
Skatteförvaltningen
Rådgivning på engelska om beskattningen i Finland: 029 497 050
Tjänsten Internationell personbeskattning tillhandahåller information om beskattningen av inkomster från utlandet och beskattningen av arbete utomlands samt hur en flytt utomlands påverkar beskattningen.
Tjänsten ger även råd om beskattningen för personer som kommer från utlandet till Finland för att arbeta och skyldigheterna för dem som betalar skatter i internationella sammanhang.
Stöd vid ekonomiska problem
Skuldlinjen
Telefonrådgivning: 0800 9 8009
Du kan ringa skuldlinjen kostnadsfritt från hela Finland och diskutera anonymt dina egna eller en närstående persons ekonomiska bekymmer.
Svårigheterna kan vara stora eller små.
Under samtalet får den som ringer hjälp med att kartlägga sin situation, råd och vid behov vägledning till något ställe där man kan få hjälp.
Diskriminering och rasism
Diskrimineringsombudsmannen
Du kan kontakta diskrimineringsombudsmannen byrå om du har råkat ut för diskriminering eller upplever att du har bemötts rasistiskt eller osakligt på grund av ditt etniska ursprung eller för att du är utlänning.
På telefonen ger den jourhavande överinspektören råd om hur du kan utreda saken och kommer överens om eventuella fortsatta åtgärder för att föra saken vidare.
På telefon kan vi betjäna dig på finska, svenska och engelska.
Jämställdhetsombudsmannen
Telefonrådgivning: 0295 666 842
Om du misstänker att en arbetsgivare, en läroanstalt eller någon annan instans har diskriminerat dig på grund av ditt kön och brutit mot lagen om jämställdhet mellan kvinnor och män, kan du be jämställdhetsombudsmannen om råd och anvisningar samt hjälp med att utreda ärendet.
Jämställdhetsombudsmannen ger dig även övrig information om lagen om jämställdhet mellan kvinnor och män.
Stöd för familjer
Kostnadsfri rådgivning för invandrare i frågor som rör familjens välbefinnande eller fostran av barn.
Rådgivning på olika språk:
Ryska och engelska: 050 325 7173
Rådgivning i frågor om hälsa
MIELI Psykisk Hälsa Finland rf
Kristelefon på finska: 09 2525 0111
Kristelefon för arabisktalande: 09 2525 0113.
Du kan även ringa och prata på engelska.
MIELI rf:s kristelefon erbjuder omedelbar samtalshjälp för människor i kris och deras närstående.
Samtalen besvaras av krisarbetare och utbildade frivilliga stödpersoner.
Du behöver inte uppge ditt namn när du ringer.
På kristelefonen kan du prata om en oväntad händelse eller en svår livssituation i en tillåtande och stödande atmosfär.
Stödcentret Hilma för handikappade invandrare
Du får handledning och råd om att ansöka om socialtjänster och förmåner avsedda för handikappade samt med att fylla i blanketter.
Du kan också fråga om möjligheterna till rehabilitering, studier, arbete och hobbyer.
Telefonen betjänar på finska, svenska, engelska och tyska.
Förgiftningar, vård och förebyggande: (09) 471 977
Vid Giftinformationscentralen kan du fråga om förebyggande och vård av akuta förgiftningar.
Hjälp med att få slut på våld
Nollalinja
Tfn 080 005 005
Öppet: varje dag
Nollalinja är en hjälptelefon som du kan ringa om du har blivit utsatt för våld i familjen, sexuellt våld eller hot om våld.
Du kan ringa när som helst.
Medarbetarna pratar finska, svenska och engelska.
Samtal till Nollalinja är kostnadsfria och de syns inte i telefonräkningen.
Du behöver inte uppge ditt namn när du ringer.
Nollalinja är avsedd för både kvinnor och män.
Manslinjen
Hjälptelefon: (09) 276 62 899
Manslinjen är en tjänst som hjälper invandrarmän som har utövat våld eller är oroliga för att de kommer att utöva våld mot en närstående människa eller någon i familjen.
Vi ger stöd och råd åt invandrarkvinnor som blivit utsatt för våld eller lever under hot om våld.
Du behöver inte uppge ditt namn när du ringer.
Maria Akademi
Öppna linjen: 09 7562 2260
Stöd och hjälp för kvinnor som utövar våld eller är oroliga för att de kommer att göra det.
Samtalen är konfidentiella.
Den öppna linjen betjänar på finska, svenska och engelska.
Hjälp till offer för människohandel
Nationellt hjälpsystem till offer för människohandel i Finland
Hjälptelefon: 02954 63177
Ta kontakt med hjälpsystemet till offer för människohandel om du upplever att du blivit offer för utnyttjande.
Du får hjälp även om du
vistas i landet illegalt
inte har identitetsbevis eller pass
blir utsatt för hot, eller om en närstående till dig blir utsatt för hot
endast talar ditt modersmål
står i skuld till någon
Basfakta
Trafiken
Religion
Beslutsfattande och påverkan
Basfakta
Staden Rovaniemi är belägen mellan två stora älvar, Ounasälv och Kemi älv, och har blivit ett framstegsvänligt och internationellt centrum för handel, administration och utbildning.
Rovaniemi har alltid haft rollen som porten till Lappland och staden har varit det administrativa centret för Lapplands län ända sedan år 1938.
Staden och landskommunen slogs samman till nya Rovaniemi stad år 2006.
Naturen är som bäst en källa till kraft och inspiration.
Att bo i Rovaniemi betyder att man har tillgång till både en livfull urban miljö och den positiva lappländska atmosfären.
Skogarna, kärren, ängarna, åkrarna, älvarna och de små insjöarna skapar en bild av Lappland och Rovaniemi, vars uttryck och stämning ändras och förnyas i takt med årstiderna.
Rovaniemis färger bär ett budskap för övriga Finland och Europa om de anpassningsbara nordliga breddgraderna, den arktiska kulturen och människorna.
Vid Rovaniemi Turistinformation får du den senaste informationen om aktiviteter och evenemang i Rovaniemi.
På turistbyrån finns bland annat broschyrer om Rovaniemi, kartor, tidtabeller och information om evenemang.
Tfn 016 346 270 eller 040 829 0676
Läs mer:
Trafiken
Läs mer:
InfoFinlands
Trafiken i Finland
Bussar
Tidtabeller, biljettpriser och linjekartor hittar du enklast på Matkahuoltos webbplats på finska, svenska och engelska.
Läs mer:
Ruttsökning
Taxi
Rovaniemi regiontaxi erbjuder taxitjänster i Rovaniemiområdet dygnet runt.
Du kan ringa efter en taxi eller ta en vid en taxistolpe där lediga taxibilar väntar på passagerare.
Du kan betala för taxin med kontanter eller med bank- eller kreditkort.
Läs mer:
Att köra bil och parkera
I centrum är parkeringsplatserna i regel avgiftsbelagda.
Parkeringsavgiften är 1,40 € per timme på alla avgiftsbelagda platser.
Det finns 73 parkeringsautomater och du betalar parkeringsavgiften i en parkeringsautomat.
Automaten skriver ut en parkeringsbiljett som du placerar innanför bilens vindruta så att hela parkeringsbiljetten kan läsas från utsidan.
Med parkeringsbiljetter köpta i parkeringsautomater kan man parkera på alla avgiftsbelagda parkeringsplatser i centrum (på mätarplatser längs gator, på torg och parkeringar) om det finns parkeringstid kvar på biljetten.
Läs mer:
Parkering
Cykling
Att cykla är ett fint och smidigt sätt att röra sig i Rovaniemi.
I staden finns flera cykelleder och vägar som lämpar sig för cykling.
En av de mest populära cykelrutterna bland stadsborna är turen som går över de tre broarna.
Läs mer:
Rovaniemi karttjänstfinska _ svenska _ engelska
Trafiklänkar
Flera av Matkahuoltos bussar i lokal- och regiontrafiken avgår från Rovaniemi busstation.
Från Rovaniemi järnvägsstation finns flera förbindelser med VR till övriga Finland.
Från Rovaniemi flygplats finns flera flyg till Helsingfors, andra städer i landet och utrikes resmål.
Läs mer:
Religion
Läs mer:
InfoFinlands
Kulturer och religioner i Finland
Beslutsfattande och påverkan
Beslutsfattande
Stadsfullmäktige är det högsta beslutsorganet i staden.
Stadsfullmäktige styr stadens utveckling på ett konkret sätt genom att utöva den ekonomiska makten.
Fullmäktige beslutar om grunderna för ekonomin och finansieringen, skattesatsen och de allmänna avgiftsgrunderna, samt ställer upp kvalitets- och verksamhetsmål för förvaltningarna.
Rovaniemi stadsstyrelse svarar för stadens administration och ekonomi, förbereder ärenden som beslutas av stadsfullmäktige samt ser till att fullmäktiges beslut verkställs och är lagliga.
Stadsstyrelsen representerar kommunen: den använder stadens yttranderätt och vidtar olika juridiska åtgärder för staden.
De högsta tjänstemännen i Rovaniemi stad är stadsdirektören och två biträdande stadsdirektörer.
Läs mer:
Beslutsfattande
Påverkan
Kommuninvånarna kan delta i och påverka stadens ärenden vid kommunalvalet som hålls vart fjärde år.
Kommuninvånarna kan dessutom väcka initiativ, svara på förfrågningar, delta i diskussionen och ge feedback till tjänstemännen.
Läs mer:
Delaktighet
Basfakta
Trafiken
Religion
Beslutsfattande och påverkan
Basfakta
Staden Rovaniemi är belägen mellan två stora älvar, Ounasälv och Kemi älv, och har blivit ett framstegsvänligt och internationellt centrum för handel, administration och utbildning.
Rovaniemi har alltid haft rollen som porten till Lappland och staden har varit det administrativa centret för Lapplands län ända sedan år 1938.
Staden och landskommunen slogs samman till nya Rovaniemi stad år 2006.
Naturen är som bäst en källa till kraft och inspiration.
Att bo i Rovaniemi betyder att man har tillgång till både en livfull urban miljö och den positiva lappländska atmosfären.
Skogarna, kärren, ängarna, åkrarna, älvarna och de små insjöarna skapar en bild av Lappland och Rovaniemi, vars uttryck och stämning ändras och förnyas i takt med årstiderna.
Rovaniemis färger bär ett budskap för övriga Finland och Europa om de anpassningsbara nordliga breddgraderna, den arktiska kulturen och människorna.
Vid Rovaniemi Turistinformation får du den senaste informationen om aktiviteter och evenemang i Rovaniemi.
På turistbyrån finns bland annat broschyrer om Rovaniemi, kartor, tidtabeller och information om evenemang.
Tfn 016 346 270 eller 040 829 0676
Läs mer:
Trafiken
Läs mer:
InfoFinlands
Trafiken i Finland
Bussar
Tidtabeller, biljettpriser och linjekartor hittar du enklast på Matkahuoltos webbplats på finska, svenska och engelska.
Läs mer:
Ruttsökning
Taxi
Rovaniemi regiontaxi erbjuder taxitjänster i Rovaniemiområdet dygnet runt.
Du kan ringa efter en taxi eller ta en vid en taxistolpe där lediga taxibilar väntar på passagerare.
Du kan betala för taxin med kontanter eller med bank- eller kreditkort.
Läs mer:
Att köra bil och parkera
I centrum är parkeringsplatserna i regel avgiftsbelagda.
Parkeringsavgiften är 1,40 € per timme på alla avgiftsbelagda platser.
Det finns 73 parkeringsautomater och du betalar parkeringsavgiften i en parkeringsautomat.
Automaten skriver ut en parkeringsbiljett som du placerar innanför bilens vindruta så att hela parkeringsbiljetten kan läsas från utsidan.
Med parkeringsbiljetter köpta i parkeringsautomater kan man parkera på alla avgiftsbelagda parkeringsplatser i centrum (på mätarplatser längs gator, på torg och parkeringar) om det finns parkeringstid kvar på biljetten.
Läs mer:
Parkering
Cykling
Att cykla är ett fint och smidigt sätt att röra sig i Rovaniemi.
I staden finns flera cykelleder och vägar som lämpar sig för cykling.
En av de mest populära cykelrutterna bland stadsborna är turen som går över de tre broarna.
Läs mer:
Rovaniemi karttjänstfinska _ svenska _ engelska
Trafiklänkar
Flera av Matkahuoltos bussar i lokal- och regiontrafiken avgår från Rovaniemi busstation.
Från Rovaniemi järnvägsstation finns flera förbindelser med VR till övriga Finland.
Från Rovaniemi flygplats finns flera flyg till Helsingfors, andra städer i landet och utrikes resmål.
Läs mer:
Religion
Läs mer:
InfoFinlands
Kulturer och religioner i Finland
Beslutsfattande och påverkan
Beslutsfattande
Stadsfullmäktige är det högsta beslutsorganet i staden.
Stadsfullmäktige styr stadens utveckling på ett konkret sätt genom att utöva den ekonomiska makten.
Fullmäktige beslutar om grunderna för ekonomin och finansieringen, skattesatsen och de allmänna avgiftsgrunderna, samt ställer upp kvalitets- och verksamhetsmål för förvaltningarna.
Rovaniemi stadsstyrelse svarar för stadens administration och ekonomi, förbereder ärenden som beslutas av stadsfullmäktige samt ser till att fullmäktiges beslut verkställs och är lagliga.
Stadsstyrelsen representerar kommunen: den använder stadens yttranderätt och vidtar olika juridiska åtgärder för staden.
De högsta tjänstemännen i Rovaniemi stad är stadsdirektören och två biträdande stadsdirektörer.
Läs mer:
Beslutsfattande
Påverkan
Kommuninvånarna kan delta i och påverka stadens ärenden vid kommunalvalet som hålls vart fjärde år.
Kommuninvånarna kan dessutom väcka initiativ, svara på förfrågningar, delta i diskussionen och ge feedback till tjänstemännen.
Läs mer:
Delaktighet
Basfakta
Trafiken
Religion
Beslutsfattande och påverkan
Basfakta
Staden Rovaniemi är belägen mellan två stora älvar, Ounasälv och Kemi älv, och har blivit ett framstegsvänligt och internationellt centrum för handel, administration och utbildning.
Rovaniemi har alltid haft rollen som porten till Lappland och staden har varit det administrativa centret för Lapplands län ända sedan år 1938.
Staden och landskommunen slogs samman till nya Rovaniemi stad år 2006.
Naturen är som bäst en källa till kraft och inspiration.
Att bo i Rovaniemi betyder att man har tillgång till både en livfull urban miljö och den positiva lappländska atmosfären.
Skogarna, kärren, ängarna, åkrarna, älvarna och de små insjöarna skapar en bild av Lappland och Rovaniemi, vars uttryck och stämning ändras och förnyas i takt med årstiderna.
Rovaniemis färger bär ett budskap för övriga Finland och Europa om de anpassningsbara nordliga breddgraderna, den arktiska kulturen och människorna.
Vid Rovaniemi Turistinformation får du den senaste informationen om aktiviteter och evenemang i Rovaniemi.
På turistbyrån finns bland annat broschyrer om Rovaniemi, kartor, tidtabeller och information om evenemang.
Tfn 016 346 270 eller 040 829 0676
Läs mer:
Trafiken
Läs mer:
InfoFinlands
Trafiken i Finland
Bussar
Tidtabeller, biljettpriser och linjekartor hittar du enklast på Matkahuoltos webbplats på finska, svenska och engelska.
Läs mer:
Ruttsökning
Taxi
Rovaniemi regiontaxi erbjuder taxitjänster i Rovaniemiområdet dygnet runt.
Du kan ringa efter en taxi eller ta en vid en taxistolpe där lediga taxibilar väntar på passagerare.
Du kan betala för taxin med kontanter eller med bank- eller kreditkort.
Läs mer:
Att köra bil och parkera
I centrum är parkeringsplatserna i regel avgiftsbelagda.
Parkeringsavgiften är 1,40 € per timme på alla avgiftsbelagda platser.
Det finns 73 parkeringsautomater och du betalar parkeringsavgiften i en parkeringsautomat.
Automaten skriver ut en parkeringsbiljett som du placerar innanför bilens vindruta så att hela parkeringsbiljetten kan läsas från utsidan.
Med parkeringsbiljetter köpta i parkeringsautomater kan man parkera på alla avgiftsbelagda parkeringsplatser i centrum (på mätarplatser längs gator, på torg och parkeringar) om det finns parkeringstid kvar på biljetten.
Läs mer:
Parkering
Cykling
Att cykla är ett fint och smidigt sätt att röra sig i Rovaniemi.
I staden finns flera cykelleder och vägar som lämpar sig för cykling.
En av de mest populära cykelrutterna bland stadsborna är turen som går över de tre broarna.
Läs mer:
Rovaniemi karttjänstfinska _ svenska _ engelska
Trafiklänkar
Flera av Matkahuoltos bussar i lokal- och regiontrafiken avgår från Rovaniemi busstation.
Från Rovaniemi järnvägsstation finns flera förbindelser med VR till övriga Finland.
Från Rovaniemi flygplats finns flera flyg till Helsingfors, andra städer i landet och utrikes resmål.
Läs mer:
Religion
Läs mer:
InfoFinlands
Kulturer och religioner i Finland
Beslutsfattande och påverkan
Beslutsfattande
Stadsfullmäktige är det högsta beslutsorganet i staden.
Stadsfullmäktige styr stadens utveckling på ett konkret sätt genom att utöva den ekonomiska makten.
Fullmäktige beslutar om grunderna för ekonomin och finansieringen, skattesatsen och de allmänna avgiftsgrunderna, samt ställer upp kvalitets- och verksamhetsmål för förvaltningarna.
Rovaniemi stadsstyrelse svarar för stadens administration och ekonomi, förbereder ärenden som beslutas av stadsfullmäktige samt ser till att fullmäktiges beslut verkställs och är lagliga.
Stadsstyrelsen representerar kommunen: den använder stadens yttranderätt och vidtar olika juridiska åtgärder för staden.
De högsta tjänstemännen i Rovaniemi stad är stadsdirektören och två biträdande stadsdirektörer.
Läs mer:
Beslutsfattande
Påverkan
Kommuninvånarna kan delta i och påverka stadens ärenden vid kommunalvalet som hålls vart fjärde år.
Kommuninvånarna kan dessutom väcka initiativ, svara på förfrågningar, delta i diskussionen och ge feedback till tjänstemännen.
Läs mer:
Delaktighet
Polisen
FPA
Arbets- och näringsbyrån
Socialbyrån
Skattebyrån
Migrationsverket
Ambassader och konsulat
Diskrimineringsombudsmannen
Polisen
Polisens uppgifter i Finland
Polisens uppgifter omfattar tryggande av ordning och säkerhet i samhället samt förebyggande och utredning av brott.
Broschyren Information om polisen i Finlandfinska _ svenska _ engelska
Brottsutredning
I Finland har polisen ansvaret för att reda ut brott och lämna dem till åtalsprövning.
Brott kan anmälas per telefon eller fax, på polisens webbplats eller genom personligt besök till polisstationen.
Polisen inleder utredningen om det finns skäl att misstänka ett brott.
Mer information om brottsanmälan hittar du på InfoFinlands sida Brott.
Information om brottfinska _ svenska _ engelska
Pass
Polisen utfärdar pass för finska medborgare.
Pass ansöks på polisstationen.
Du kan lämna in din passansökan på vilken av polisens tillståndsenheter som helst.
Att ansöka om finskt passfinska _ svenska _ engelska
Identitetskort
Polisen utfärdar identitetskort.
Identitetskort ansöks på polisstationen.
Du kan lämna in din ansökan om identitetskort på vilken av polisens tillståndsenheter som helst.
Identitetskort för utlänningar
Polisen kan utfärda identitetskort för en utlänning som
bor stadigvarande i Finland
är införd i befolkningsdatasystemet
kan på ett pålitligt sätt styrka sin identitet
Identitetskortet för utlänningar kan användas som identitetsbevis i Finland, men inte som resedokument när man reser utomlands.
ID-kortfinska _ svenska _ engelska
Tidsbeställning
När du ska sköta ärenden vid polisens tillståndsenhet, kan du boka tid på förhand på polisens webbplats.
På så sätt undviker du köandet.
Observera att tidsbokningen är obligatorisk på vissa polisstationer.
Tidsbeställning till tillståndstjänstenfinska _ svenska _ engelska _ samiska
FPA
Folkpensionsanstalten, det vill säga FPA, betalar ut ekonomiskt stöd under olika livsskeden.
Vanligtvis kan man få FPA:s bidrag då de övriga inkomsterna är låga.
FPA:s stöd är till exempel
utkomststöd
folkpensionen, garantipensionen och andra bidrag för pensionärer
bostadsbidraget
stöd, som man kan få när man är sjuk
grundtryggheten för arbetslösa
stöd för studerande
stöd avsedda för barnfamiljer.
På InfoFinlands sida Den sociala tryggheten i Finland hittar du information om vem som kan få FPA:s stöd.
Information om FPAfinska _ svenska _ engelska
Arbets- och näringsbyrån
Arbets- och näringsbyråerna tillhandahåller till exempel följande tjänster:
arbetsförmedling
arbetskraftsutbildning
tjänster för företagare
yrkesvägledning
Arbets- och näringsbyråeran upprättar även integrationsplaner för invandrare som är klienter vid arbets- och näringsbyrån.
Via arbets- och näringsbyråerna kan man till exempel söka till kurser i det finska språket.
På arbets- och näringsbyrån får man information om lediga jobb.
Arbets- och näringsbyråns klienter kan ansöka om arbetslöshetspenning vid FPA.
Information om arbets- och näringsbyråernas tjänster hittar du på InfoFinlands sida Tjänsterna vid arbets- och näringsbyrån.
linkkiArbets- och näringsministeriet:
Arbets- och näringsbyråerfinska _ svenska
Socialbyrån
Socialbyråerna betjänar kommuninvånarna till exempel i följande ärenden:
tjänster för äldre
tjänster för handikappade
barnskydd
stöd för närståendevården
missbrukarvård
skuldrådgivning
Kontaktuppgifterna till närmaste socialbyrå hittar du på din hemkommuns webbplats.
Socialbyrån kan ha olika namn i olika kommuner.
linkkiSocial- och hälsovårdsministeriet:
Information om socialtjänsterfinska _ svenska _ engelska
Skattebyrån
På skattebyrån (verotoimisto) kan du sköta ärenden rörande skatter.
På skattebyrån kan du till exempel få skattekort, ändra din skatteprocent eller fråga om sådant som rör beskattningen.
I webbtjänsten MinSkatt kan du sköta många skatterelaterade ärenden elektroniskt.
Du kan till exempel beställa ett nytt skattekort om du ha nätbankskoder eller ett mobilcertifikat.
På skatteförvaltningens webbplats finns mycket information om beskattningen i Finland.
linkkiSkatteförvaltningen:
Information om skatteförvaltningenfinska _ svenska _ engelska
Migrationsverket
När du flyttar till Finland måste du ansöka om uppehållstillstånd hos Migrationsverket eller registrera din uppehållsrätt.
Huruvida du behöver ett uppehållstillstånd beror på i vilket land du är medborgare, varför du kommer till Finland och hur länge du ska stanna.
Migrationsverket (Maahanmuuttovirasto) behandlar även asylansökningarna och ansökningarna om medborgarskap.
Information om Migrationsverketfinska _ svenska _ engelska
Magistraterna (maistraatti) är lokala statliga förvaltningsmyndigheter.
Magistraterna lagrar information om invånarna i sitt område i befolkningsregistret.
I befolkningsregistret registreras alla personer som bor i Finland.
Man ska göra en anmälan till magistraten när man flyttar till Finland.
Anmälan ska även göras då man flyttar inom eller bort från Finland.
Magistraten har även många andra uppgifter.
förrättar civilvigslar och registrerar parförhållanden,
utfärdar personbeteckningar för personer bosatta i Finland,
utfärdar hemortsintyg med vilket man kan bevisa var man bor.
Information om magistraternafinska _ svenska _ engelska
Ambassader och konsulat
Ambassader och konsulat är statliga beskickningar i en annan stat.
Finlands beskickningar utomlands
Finlands beskickningar utomlands
tar emot ansökan om uppehållstillstånd i Finland
utfärdar visum för Finland
betjänar utomlands bosatta finländare när de behöver sköta ärenden med finska myndigheter, till exempel ansöka om nytt pass
hjälper finska medborgare som råkat ut för en nödsituation utomlands
På utrikesministeriets sida finns en lista över Finlands beskickningar utomlands.
Utländska beskickningar i Finland
Information om utländska beskickningar i Finland och deras tjänster hittar du på InfoFinlands sida Ambassader i Finland.
Finlands beskickningar utomlandsfinska _ svenska _ engelska
Inresetillstånd för utlänningarfinska _ svenska _ engelska
Andra länders beskickningar i Finlandfinska _ svenska _ engelska
Information om konsultjänsternafinska _ svenska _ engelska
Diskrimineringsombudsmannen
Diskrimineringsombudsmannen är en myndighet vars uppgift är att främja likabehandling och ingripa i diskriminering.
Du kan vända dig till diskrimineringsombudsmannen till exempel om du själv har råkat ut för etnisk diskriminering eller observerat att en annan person diskrimineras.
Diskrimineringsombudsmannen kan ge anvisningar, råd och rekommendationer samt hjälpa parterna att åstadkomma förlikning i diskrimineringsfall.
Du får kontakt med diskrimineringsombudsmannens byrå:
Per telefon får du betjäning på finska, svenska och engelska.
Möten måste avtalas på förhand.
Byråns tjänster är avgiftsfria.
Om du inte kan finska, svenska eller engelska kan du skriva e-post eller brev även på andra språk.
Hjälp till diskrimineringsofferfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ thai _ vietnamesiska _ portugisiska _ tagalog _ polska
Polisen
FPA
Arbets- och näringsbyrån
Socialbyrån
Skattebyrån
Migrationsverket
Ambassader och konsulat
Diskrimineringsombudsmannen
Polisen
Polisens uppgifter i Finland
Polisens uppgifter omfattar tryggande av ordning och säkerhet i samhället samt förebyggande och utredning av brott.
Broschyren Information om polisen i Finlandfinska _ svenska _ engelska
Brottsutredning
I Finland har polisen ansvaret för att reda ut brott och lämna dem till åtalsprövning.
Brott kan anmälas per telefon eller fax, på polisens webbplats eller genom personligt besök till polisstationen.
Polisen inleder utredningen om det finns skäl att misstänka ett brott.
Mer information om brottsanmälan hittar du på InfoFinlands sida Brott.
Information om brottfinska _ svenska _ engelska
Pass
Polisen utfärdar pass för finska medborgare.
Pass ansöks på polisstationen.
Du kan lämna in din passansökan på vilken av polisens tillståndsenheter som helst.
Att ansöka om finskt passfinska _ svenska _ engelska
Identitetskort
Polisen utfärdar identitetskort.
Identitetskort ansöks på polisstationen.
Du kan lämna in din ansökan om identitetskort på vilken av polisens tillståndsenheter som helst.
Identitetskort för utlänningar
Polisen kan utfärda identitetskort för en utlänning som
bor stadigvarande i Finland
är införd i befolkningsdatasystemet
kan på ett pålitligt sätt styrka sin identitet
Identitetskortet för utlänningar kan användas som identitetsbevis i Finland, men inte som resedokument när man reser utomlands.
ID-kortfinska _ svenska _ engelska
Tidsbeställning
När du ska sköta ärenden vid polisens tillståndsenhet, kan du boka tid på förhand på polisens webbplats.
På så sätt undviker du köandet.
Observera att tidsbokningen är obligatorisk på vissa polisstationer.
Tidsbeställning till tillståndstjänstenfinska _ svenska _ engelska _ samiska
FPA
Folkpensionsanstalten, det vill säga FPA, betalar ut ekonomiskt stöd under olika livsskeden.
Vanligtvis kan man få FPA:s bidrag då de övriga inkomsterna är låga.
FPA:s stöd är till exempel
utkomststöd
folkpensionen, garantipensionen och andra bidrag för pensionärer
bostadsbidraget
stöd, som man kan få när man är sjuk
grundtryggheten för arbetslösa
stöd för studerande
stöd avsedda för barnfamiljer.
På InfoFinlands sida Den sociala tryggheten i Finland hittar du information om vem som kan få FPA:s stöd.
Information om FPAfinska _ svenska _ engelska
Arbets- och näringsbyrån
Arbets- och näringsbyråerna tillhandahåller till exempel följande tjänster:
arbetsförmedling
arbetskraftsutbildning
tjänster för företagare
yrkesvägledning
Arbets- och näringsbyråeran upprättar även integrationsplaner för invandrare som är klienter vid arbets- och näringsbyrån.
Via arbets- och näringsbyråerna kan man till exempel söka till kurser i det finska språket.
På arbets- och näringsbyrån får man information om lediga jobb.
Arbets- och näringsbyråns klienter kan ansöka om arbetslöshetspenning vid FPA.
Information om arbets- och näringsbyråernas tjänster hittar du på InfoFinlands sida Tjänsterna vid arbets- och näringsbyrån.
linkkiArbets- och näringsministeriet:
Arbets- och näringsbyråerfinska _ svenska
Socialbyrån
Socialbyråerna betjänar kommuninvånarna till exempel i följande ärenden:
tjänster för äldre
tjänster för handikappade
barnskydd
stöd för närståendevården
missbrukarvård
skuldrådgivning
Kontaktuppgifterna till närmaste socialbyrå hittar du på din hemkommuns webbplats.
Socialbyrån kan ha olika namn i olika kommuner.
linkkiSocial- och hälsovårdsministeriet:
Information om socialtjänsterfinska _ svenska _ engelska
Skattebyrån
På skattebyrån (verotoimisto) kan du sköta ärenden rörande skatter.
På skattebyrån kan du till exempel få skattekort, ändra din skatteprocent eller fråga om sådant som rör beskattningen.
I webbtjänsten MinSkatt kan du sköta många skatterelaterade ärenden elektroniskt.
Du kan till exempel beställa ett nytt skattekort om du ha nätbankskoder eller ett mobilcertifikat.
På skatteförvaltningens webbplats finns mycket information om beskattningen i Finland.
linkkiSkatteförvaltningen:
Information om skatteförvaltningenfinska _ svenska _ engelska
Migrationsverket
När du flyttar till Finland måste du ansöka om uppehållstillstånd hos Migrationsverket eller registrera din uppehållsrätt.
Huruvida du behöver ett uppehållstillstånd beror på i vilket land du är medborgare, varför du kommer till Finland och hur länge du ska stanna.
Migrationsverket (Maahanmuuttovirasto) behandlar även asylansökningarna och ansökningarna om medborgarskap.
Information om Migrationsverketfinska _ svenska _ engelska
Magistraterna (maistraatti) är lokala statliga förvaltningsmyndigheter.
Magistraterna lagrar information om invånarna i sitt område i befolkningsregistret.
I befolkningsregistret registreras alla personer som bor i Finland.
Man ska göra en anmälan till magistraten när man flyttar till Finland.
Anmälan ska även göras då man flyttar inom eller bort från Finland.
Magistraten har även många andra uppgifter.
förrättar civilvigslar och registrerar parförhållanden,
utfärdar personbeteckningar för personer bosatta i Finland,
utfärdar hemortsintyg med vilket man kan bevisa var man bor.
Information om magistraternafinska _ svenska _ engelska
Ambassader och konsulat
Ambassader och konsulat är statliga beskickningar i en annan stat.
Finlands beskickningar utomlands
Finlands beskickningar utomlands
tar emot ansökan om uppehållstillstånd i Finland
utfärdar visum för Finland
betjänar utomlands bosatta finländare när de behöver sköta ärenden med finska myndigheter, till exempel ansöka om nytt pass
hjälper finska medborgare som råkat ut för en nödsituation utomlands
På utrikesministeriets sida finns en lista över Finlands beskickningar utomlands.
Utländska beskickningar i Finland
Information om utländska beskickningar i Finland och deras tjänster hittar du på InfoFinlands sida Ambassader i Finland.
Finlands beskickningar utomlandsfinska _ svenska _ engelska
Inresetillstånd för utlänningarfinska _ svenska _ engelska
Andra länders beskickningar i Finlandfinska _ svenska _ engelska
Information om konsultjänsternafinska _ svenska _ engelska
Diskrimineringsombudsmannen
Diskrimineringsombudsmannen är en myndighet vars uppgift är att främja likabehandling och ingripa i diskriminering.
Du kan vända dig till diskrimineringsombudsmannen till exempel om du själv har råkat ut för etnisk diskriminering eller observerat att en annan person diskrimineras.
Diskrimineringsombudsmannen kan ge anvisningar, råd och rekommendationer samt hjälpa parterna att åstadkomma förlikning i diskrimineringsfall.
Du får kontakt med diskrimineringsombudsmannens byrå:
Per telefon får du betjäning på finska, svenska och engelska.
Möten måste avtalas på förhand.
Byråns tjänster är avgiftsfria.
Om du inte kan finska, svenska eller engelska kan du skriva e-post eller brev även på andra språk.
Hjälp till diskrimineringsofferfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ thai _ vietnamesiska _ portugisiska _ tagalog _ polska
Polisen
FPA
Arbets- och näringsbyrån
Socialbyrån
Skattebyrån
Migrationsverket
Ambassader och konsulat
Diskrimineringsombudsmannen
Polisen
Polisens uppgifter i Finland
Polisens uppgifter omfattar tryggande av ordning och säkerhet i samhället samt förebyggande och utredning av brott.
Broschyren Information om polisen i Finlandfinska _ svenska _ engelska
Brottsutredning
I Finland har polisen ansvaret för att reda ut brott och lämna dem till åtalsprövning.
Brott kan anmälas per telefon eller fax, på polisens webbplats eller genom personligt besök till polisstationen.
Polisen inleder utredningen om det finns skäl att misstänka ett brott.
Mer information om brottsanmälan hittar du på InfoFinlands sida Brott.
Information om brottfinska _ svenska _ engelska
Pass
Polisen utfärdar pass för finska medborgare.
Pass ansöks på polisstationen.
Du kan lämna in din passansökan på vilken av polisens tillståndsenheter som helst.
Att ansöka om finskt passfinska _ svenska _ engelska
Identitetskort
Polisen utfärdar identitetskort.
Identitetskort ansöks på polisstationen.
Du kan lämna in din ansökan om identitetskort på vilken av polisens tillståndsenheter som helst.
Identitetskort för utlänningar
Polisen kan utfärda identitetskort för en utlänning som
bor stadigvarande i Finland
är införd i befolkningsdatasystemet
kan på ett pålitligt sätt styrka sin identitet
Identitetskortet för utlänningar kan användas som identitetsbevis i Finland, men inte som resedokument när man reser utomlands.
ID-kortfinska _ svenska _ engelska
Tidsbeställning
När du ska sköta ärenden vid polisens tillståndsenhet, kan du boka tid på förhand på polisens webbplats.
På så sätt undviker du köandet.
Observera att tidsbokningen är obligatorisk på vissa polisstationer.
Tidsbeställning till tillståndstjänstenfinska _ svenska _ engelska _ samiska
FPA
Folkpensionsanstalten, det vill säga FPA, betalar ut ekonomiskt stöd under olika livsskeden.
Vanligtvis kan man få FPA:s bidrag då de övriga inkomsterna är låga.
FPA:s stöd är till exempel
utkomststöd
folkpensionen, garantipensionen och andra bidrag för pensionärer
bostadsbidraget
stöd, som man kan få när man är sjuk
grundtryggheten för arbetslösa
stöd för studerande
stöd avsedda för barnfamiljer.
På InfoFinlands sida Den sociala tryggheten i Finland hittar du information om vem som kan få FPA:s stöd.
Information om FPAfinska _ svenska _ engelska
Arbets- och näringsbyrån
Arbets- och näringsbyråerna tillhandahåller till exempel följande tjänster:
arbetsförmedling
arbetskraftsutbildning
tjänster för företagare
yrkesvägledning
Arbets- och näringsbyråeran upprättar även integrationsplaner för invandrare som är klienter vid arbets- och näringsbyrån.
Via arbets- och näringsbyråerna kan man till exempel söka till kurser i det finska språket.
På arbets- och näringsbyrån får man information om lediga jobb.
Arbets- och näringsbyråns klienter kan ansöka om arbetslöshetspenning vid FPA.
linkkiArbets- och näringsministeriet:
Arbets- och näringsbyråerfinska _ svenska
Socialbyrån
Socialbyråerna betjänar kommuninvånarna till exempel i följande ärenden:
tjänster för äldre
tjänster för handikappade
barnskydd
stöd för närståendevården
missbrukarvård
skuldrådgivning
Kontaktuppgifterna till närmaste socialbyrå hittar du på din hemkommuns webbplats.
Socialbyrån kan ha olika namn i olika kommuner.
linkkiSocial- och hälsovårdsministeriet:
Information om socialtjänsterfinska _ svenska _ engelska
Skattebyrån
På skattebyrån (verotoimisto) kan du sköta ärenden rörande skatter.
På skattebyrån kan du till exempel få skattekort, ändra din skatteprocent eller fråga om sådant som rör beskattningen.
I webbtjänsten MinSkatt kan du sköta många skatterelaterade ärenden elektroniskt.
Du kan till exempel beställa ett nytt skattekort om du ha nätbankskoder eller ett mobilcertifikat.
På skatteförvaltningens webbplats finns mycket information om beskattningen i Finland.
linkkiSkatteförvaltningen:
Information om skatteförvaltningenfinska _ svenska _ engelska
Migrationsverket
När du flyttar till Finland måste du ansöka om uppehållstillstånd hos Migrationsverket eller registrera din uppehållsrätt.
Huruvida du behöver ett uppehållstillstånd beror på i vilket land du är medborgare, varför du kommer till Finland och hur länge du ska stanna.
Migrationsverket (Maahanmuuttovirasto) behandlar även asylansökningarna och ansökningarna om medborgarskap.
Information om Migrationsverketfinska _ svenska _ engelska
Magistraterna (maistraatti) är lokala statliga förvaltningsmyndigheter.
Magistraterna lagrar information om invånarna i sitt område i befolkningsregistret.
I befolkningsregistret registreras alla personer som bor i Finland.
Man ska göra en anmälan till magistraten när man flyttar till Finland.
Anmälan ska även göras då man flyttar inom eller bort från Finland.
Magistraten har även många andra uppgifter.
förrättar civilvigslar och registrerar parförhållanden,
utfärdar personbeteckningar för personer bosatta i Finland,
utfärdar hemortsintyg med vilket man kan bevisa var man bor.
Information om magistraternafinska _ svenska _ engelska
Ambassader och konsulat
Ambassader och konsulat är statliga beskickningar i en annan stat.
Finlands beskickningar utomlands
Finlands beskickningar utomlands
tar emot ansökan om uppehållstillstånd i Finland
utfärdar visum för Finland
betjänar utomlands bosatta finländare när de behöver sköta ärenden med finska myndigheter, till exempel ansöka om nytt pass
hjälper finska medborgare som råkat ut för en nödsituation utomlands
På utrikesministeriets sida finns en lista över Finlands beskickningar utomlands.
Utländska beskickningar i Finland
Information om utländska beskickningar i Finland och deras tjänster hittar du på InfoFinlands sida Ambassader i Finland.
Finlands beskickningar utomlandsfinska _ svenska _ engelska
Inresetillstånd för utlänningarfinska _ svenska _ engelska
Andra länders beskickningar i Finlandfinska _ svenska _ engelska
Information om konsultjänsternafinska _ svenska _ engelska
Diskrimineringsombudsmannen
Diskrimineringsombudsmannen är en myndighet vars uppgift är att främja likabehandling och ingripa i diskriminering.
Du kan vända dig till diskrimineringsombudsmannen till exempel om du själv har råkat ut för etnisk diskriminering eller observerat att en annan person diskrimineras.
Diskrimineringsombudsmannen kan ge anvisningar, råd och rekommendationer samt hjälpa parterna att åstadkomma förlikning i diskrimineringsfall.
Du får kontakt med diskrimineringsombudsmannens byrå:
Per telefon får du betjäning på finska, svenska och engelska.
Möten måste avtalas på förhand.
Byråns tjänster är avgiftsfria.
Om du inte kan finska, svenska eller engelska kan du skriva e-post eller brev även på andra språk.
Hjälp till diskrimineringsofferfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ thai _ vietnamesiska _ portugisiska _ tagalog _ polska
Jämställdhet mellan män och kvinnor
Enligt Finlands lag har män och kvinnor samma rättigheter.
Även gifta kvinnor har samma rättigheter som män.
I Finland är det vanligt att också kvinnor arbetar, trots att de har barn.
Ansvaret för skötseln av barnen och hemmet hör till både kvinnan och mannen.
En kvinna behöver inte sin makes eller sina föräldrars tillåtelse för att arbeta eller studera.
Kvinnor och män kan själva besluta om vem de gifter sig med.
Att tvinga någon till äktenskap är ett brott i Finland.
Exempelvis föräldrarna har inte rätt att tvinga eller utöva påtryckning på sitt barn att gifta sig.
Både kvinnan och mannen har rätt att söka skilsmässa.
Man kan också söka skilsmässa utan makens eller makans samtycke.
Våld är alltid ett brott i Finland.
Även våld i familjen och parförhållandet, till exempel slag och sexuellt våld är alltid ett brott.
Läs mer på InfoFinlands sida Våld och Hedersrelaterat våld.
Jämställdhet i arbetslivet
I arbetslivet ska kvinnor och män behandlas lika.
Diskriminering på grund av kön är förbjudet.
Detta innebär till exempel att man inte får betala högre lön till en man än till en kvinna på grund av kön eller säga upp en anställd på grund av att hon är gravid.
Jämställdhetslagen förbjuder diskriminering på grund av kön.
Jämställdhetsombudsmannen är en myndighet, som övervakar att jämställdhetslagen följs.
Om du misstänker att du har blivit diskriminerad i arbetslivet på grund av ditt kön, kan du kontakta jämställdhetsombudsmannen (tasa-arvovaltuutettu) eller ditt fackförbund.
Läs mer på InfoFinlands sida Jämlikhet och jämställdhet i arbetslivet.
linkkiJämställdhetsombudsman:
Information om jämställdhetfinska _ svenska _ engelska
Likabehandling
Enligt Finlands lag ska alla människor behandlas likvärdigt.
Diskriminering är ett brott.
På InfoFinlands sida Diskriminering och rasism finns information om var du kan få hjälp om du har upplevt diskriminering eller blivit offer för ett rasistiskt brott.
Sexuella minoriteter och könsminoriteters rättigheter
Enligt Finlands lag får en människa inte diskrimineras på grund av sin sexuella läggning.
Lagen förbjuder även diskriminering på grund av könsidentitet eller uttryck för kön.
Den som har blivit förföljd på grund av sin sexuella läggning eller könsidentitet någon annanstans kan söka asyl i Finland.
Det är dock inte givet att man får asyl, utan varje fall utreds separat.
I utredningen klarläggs situationen för den sökande och landet där denna kommer ifrån så noga som möjligt.
I Finland finns flera organisationer för sexuella minoriteter och könsminoriteter.
De strävar efter att förbättra dessa minoriteters ställning i samhället.
Många organisationer erbjuder även utbildning, rådgivning och olika stödtjänster.
Transsexuella personer, transvestiter, intersexuella personer och andra människor med mångfacetterad könsidentitet kan få hjälp av jämställdhetsombudsmannen om de upplever diskriminering.
I Finland kan också två män eller två kvinnor gifta sig med varandra.
Läs mer på InfoFinlands sida Äktenskap.
På InfoFinlands sida Vad är en familj?
finns information om familjer som bildas av samkönade par.
linkkiSeta:
Information om sexuellt likaberättigandefinska _ svenska _ engelska _ ryska
linkkiTrasek ry.:
Information för könsminoriteterfinska _ svenska _ engelska
linkkiDreamwearclub ry.:
Information för könsminoriteterfinska
Information för könsminoriteterfinska _ svenska _ engelska
Barns rättigheter
I Finland har barn rätt till särskilt skydd och särskild omsorg.
Barn har även rätt att uttrycka sina egna åsikter.
Barn har rätt till att deras åsikt tas i beaktande när man fattar beslut om sådant som rör dem.
Enligt Finlands lag är kroppsaga mot barn förbjudet och den kan ha straffpåföljd.
Mer information om barns rättigheter i Finland hittar du också på InfoFinlands sidor Barn.
linkkiBarnombudsmannen:
Broschyren Barnets rättigheterfinska _ svenska _ engelska _ ryska
Handikappades rättigheter
Enligt lag få handikappade personer inte diskrimineras.
En handikappad har rätt att leva ett vanligt liv, till exempel studera, arbeta och bilda familj.
Enligt lagen om likabehandling måste arbetsgivare och utbildningsanordnare förbättra handikappade personers möjligheter att få arbete och utbildning.
Till exempel kan arbetsmiljön modifieras så att den handikappade lättare kan röra sig där.
Information om tjänster för handikappade hittar du på InfoFinlands sida Handikappade.
Jämställdhet mellan män och kvinnor
Enligt Finlands lag har män och kvinnor samma rättigheter.
Även gifta kvinnor har samma rättigheter som män.
I Finland är det vanligt att också kvinnor arbetar, trots att de har barn.
Ansvaret för skötseln av barnen och hemmet hör till både kvinnan och mannen.
En kvinna behöver inte sin makes eller sina föräldrars tillåtelse för att arbeta eller studera.
Kvinnor och män kan själva besluta om vem de gifter sig med.
Att tvinga någon till äktenskap är ett brott i Finland.
Exempelvis föräldrarna har inte rätt att tvinga eller utöva påtryckning på sitt barn att gifta sig.
Både kvinnan och mannen har rätt att söka skilsmässa.
Man kan också söka skilsmässa utan makens eller makans samtycke.
Våld är alltid ett brott i Finland.
Även våld i familjen och parförhållandet, till exempel slag och sexuellt våld är alltid ett brott.
Läs mer på InfoFinlands sida Våld och Hedersrelaterat våld.
Jämställdhet i arbetslivet
I arbetslivet ska kvinnor och män behandlas lika.
Diskriminering på grund av kön är förbjudet.
Detta innebär till exempel att man inte får betala högre lön till en man än till en kvinna på grund av kön eller säga upp en anställd på grund av att hon är gravid.
Jämställdhetslagen förbjuder diskriminering på grund av kön.
Jämställdhetsombudsmannen är en myndighet, som övervakar att jämställdhetslagen följs.
Om du misstänker att du har blivit diskriminerad i arbetslivet på grund av ditt kön, kan du kontakta jämställdhetsombudsmannen (tasa-arvovaltuutettu) eller ditt fackförbund.
Läs mer på InfoFinlands sida Jämlikhet och jämställdhet i arbetslivet.
linkkiJämställdhetsombudsman:
Information om jämställdhetfinska _ svenska _ engelska
Likabehandling
Enligt Finlands lag ska alla människor behandlas likvärdigt.
Diskriminering är ett brott.
På InfoFinlands sida Diskriminering och rasism finns information om var du kan få hjälp om du har upplevt diskriminering eller blivit offer för ett rasistiskt brott.
Sexuella minoriteter och könsminoriteters rättigheter
Enligt Finlands lag får en människa inte diskrimineras på grund av sin sexuella läggning.
Lagen förbjuder även diskriminering på grund av könsidentitet eller uttryck för kön.
Den som har blivit förföljd på grund av sin sexuella läggning eller könsidentitet någon annanstans kan söka asyl i Finland.
Det är dock inte givet att man får asyl, utan varje fall utreds separat.
I utredningen klarläggs situationen för den sökande och landet där denna kommer ifrån så noga som möjligt.
I Finland finns flera organisationer för sexuella minoriteter och könsminoriteter.
De strävar efter att förbättra dessa minoriteters ställning i samhället.
Många organisationer erbjuder även utbildning, rådgivning och olika stödtjänster.
Transsexuella personer, transvestiter, intersexuella personer och andra människor med mångfacetterad könsidentitet kan få hjälp av jämställdhetsombudsmannen om de upplever diskriminering.
I Finland kan också två män eller två kvinnor gifta sig med varandra.
Läs mer på InfoFinlands sida Äktenskap.
På InfoFinlands sida Vad är en familj?
finns information om familjer som bildas av samkönade par.
linkkiSeta:
Information om sexuellt likaberättigandefinska _ svenska _ engelska _ ryska
linkkiTrasek ry.:
Information för könsminoriteterfinska _ svenska _ engelska
linkkiDreamwearclub ry.:
Information för könsminoriteterfinska
Information för könsminoriteterfinska _ svenska _ engelska
Barns rättigheter
I Finland har barn rätt till särskilt skydd och särskild omsorg.
Barn har även rätt att uttrycka sina egna åsikter.
Barn har rätt till att deras åsikt tas i beaktande när man fattar beslut om sådant som rör dem.
Enligt Finlands lag är kroppsaga mot barn förbjudet och den kan ha straffpåföljd.
Mer information om barns rättigheter i Finland hittar du också på InfoFinlands sidor Barn.
linkkiBarnombudsmannen:
Broschyren Barnets rättigheterfinska _ svenska _ engelska _ ryska
Handikappades rättigheter
Enligt lag få handikappade personer inte diskrimineras.
En handikappad har rätt att leva ett vanligt liv, till exempel studera, arbeta och bilda familj.
Enligt lagen om likabehandling måste arbetsgivare och utbildningsanordnare förbättra handikappade personers möjligheter att få arbete och utbildning.
Till exempel kan arbetsmiljön modifieras så att den handikappade lättare kan röra sig där.
Information om tjänster för handikappade hittar du på InfoFinlands sida Handikappade.
Jämställdhet mellan män och kvinnor
Enligt Finlands lag har män och kvinnor samma rättigheter.
Även gifta kvinnor har samma rättigheter som män.
I Finland är det vanligt att också kvinnor arbetar, trots att de har barn.
Ansvaret för skötseln av barnen och hemmet hör till både kvinnan och mannen.
En kvinna behöver inte sin makes eller sina föräldrars tillåtelse för att arbeta eller studera.
Kvinnor och män kan själva besluta om vem de gifter sig med.
Att tvinga någon till äktenskap är ett brott i Finland.
Exempelvis föräldrarna har inte rätt att tvinga eller utöva påtryckning på sitt barn att gifta sig.
Både kvinnan och mannen har rätt att söka skilsmässa.
Man kan också söka skilsmässa utan makens eller makans samtycke.
Våld är alltid ett brott i Finland.
Även våld i familjen och parförhållandet, till exempel slag och sexuellt våld är alltid ett brott.
Läs mer på InfoFinlands sida Våld och Hedersrelaterat våld.
Jämställdhet i arbetslivet
I arbetslivet ska kvinnor och män behandlas lika.
Diskriminering på grund av kön är förbjudet.
Detta innebär till exempel att man inte får betala högre lön till en man än till en kvinna på grund av kön eller säga upp en anställd på grund av att hon är gravid.
Jämställdhetslagen förbjuder diskriminering på grund av kön.
Jämställdhetsombudsmannen är en myndighet, som övervakar att jämställdhetslagen följs.
Om du misstänker att du har blivit diskriminerad i arbetslivet på grund av ditt kön, kan du kontakta jämställdhetsombudsmannen (tasa-arvovaltuutettu) eller ditt fackförbund.
Läs mer på InfoFinlands sida Jämlikhet och jämställdhet i arbetslivet.
linkkiJämställdhetsombudsman:
Information om jämställdhetfinska _ svenska _ engelska
Likabehandling
Enligt Finlands lag ska alla människor behandlas likvärdigt.
Diskriminering är ett brott.
På InfoFinlands sida Diskriminering och rasism finns information om var du kan få hjälp om du har upplevt diskriminering eller blivit offer för ett rasistiskt brott.
Sexuella minoriteter och könsminoriteters rättigheter
Enligt Finlands lag får en människa inte diskrimineras på grund av sin sexuella läggning.
Lagen förbjuder även diskriminering på grund av könsidentitet eller uttryck för kön.
Den som har blivit förföljd på grund av sin sexuella läggning eller könsidentitet någon annanstans kan söka asyl i Finland.
Det är dock inte givet att man får asyl, utan varje fall utreds separat.
I utredningen klarläggs situationen för den sökande och landet där denna kommer ifrån så noga som möjligt.
I Finland finns flera organisationer för sexuella minoriteter och könsminoriteter.
De strävar efter att förbättra dessa minoriteters ställning i samhället.
Många organisationer erbjuder även utbildning, rådgivning och olika stödtjänster.
Transsexuella personer, transvestiter, intersexuella personer och andra människor med mångfacetterad könsidentitet kan få hjälp av jämställdhetsombudsmannen om de upplever diskriminering.
I Finland kan också två män eller två kvinnor gifta sig med varandra.
Läs mer på InfoFinlands sida Äktenskap.
På InfoFinlands sida Vad är en familj?
finns information om familjer som bildas av samkönade par.
linkkiSeta:
Information om sexuellt likaberättigandefinska _ svenska _ engelska _ ryska
linkkiTrasek ry.:
Information för könsminoriteterfinska _ svenska _ engelska
linkkiDreamwearclub ry.:
Information för könsminoriteterfinska
Information för könsminoriteterfinska _ svenska _ engelska
Barns rättigheter
I Finland har barn rätt till särskilt skydd och särskild omsorg.
Barn har även rätt att uttrycka sina egna åsikter.
Barn har rätt till att deras åsikt tas i beaktande när man fattar beslut om sådant som rör dem.
Enligt Finlands lag är kroppsaga mot barn förbjudet och den kan ha straffpåföljd.
Mer information om barns rättigheter i Finland hittar du också på InfoFinlands sidor Barn.
linkkiBarnombudsmannen:
Broschyren Barnets rättigheterfinska _ svenska _ engelska _ ryska
Handikappades rättigheter
Enligt lag få handikappade personer inte diskrimineras.
En handikappad har rätt att leva ett vanligt liv, till exempel studera, arbeta och bilda familj.
Enligt lagen om likabehandling måste arbetsgivare och utbildningsanordnare förbättra handikappade personers möjligheter att få arbete och utbildning.
Till exempel kan arbetsmiljön modifieras så att den handikappade lättare kan röra sig där.
Information om tjänster för handikappade hittar du på InfoFinlands sida Handikappade.
Grundläggande rättigheter
Alla som är bosatta i Finland har rättigheter och skyldigheter enligt lag.
Utlänningar som är bosatta i Finland har nästan samma rättigheter och skyldigheter som finska medborgare.
Följande rättigheter och skyldigheter gäller även utlänningar bosatta i Finland.
Rättigheter
Alla har rätt att bli jämlikt bemötta.
Ingen får behandlas annorlunda till exempel på grund av kön, ålder, religion eller handikapp.
Var och en får fritt yttra sina åsikter i tal och skrift.
Människor får ordna sammankomster och demonstrationer samt delta i dem.
En demonstration ska anmälas till polisen på förhand.
Ingen får dömas till döden eller torteras.
Alla kan själv välja var de vill bo och fritt röra sig i Finland.
Alla har rätt till integritetsskydd.
Ett brev som tillhör en annan person får inte läsas och en annan persons telefonsamtal får inte avlyssnas.
Var och en får själv välja sin religion.
Om man inte vill, måste man inte välja någon religion alls.
Utlänningar som bor stadigvarande i Finland och som har fyllt 18 år har rätt att rösta i kommunalval.
Utlänningar som har rösträtt i kommunalval har även rätt att ställa upp som kandidat i kommunalval.
EU-medborgare som har sin hemkommun i Finland kan rösta i val till Europaparlamentet i Finland om de har anmält sig till rösträttsregistret.
EU-medborgare som är i det finska rösträttsregistret kan också ställa upp som kandidat i Finlands Europaparlamentsval.
Läs mer om utlänningarnas rösträtt på InfoFinlands sida Val och röstning i Finland.
Skyldigheter
Alla som bor eller vistas i Finland måste följa Finlands lag.
Barn i åldern 7–17 år har läroplikt, det vill säga skyldighet att avlägga grundskolans lärokurs.
Ofta måste de som arbetar i Finland betala skatt på sin lön till Finland.
Alla har skyldighet att vittna inför domstol om de blir kallade.
Föräldrar är skyldiga att ta hand om sina barn.
Alla har skyldighet att hjälpa vid en olycka.
Läs mer om beskattningen i Finland på InfoFinlands sida Beskattning.
Finska medborgares rättigheter och skyldigheter
Finska medborgare har utöver det ovan nämnda också några ytterligare rättigheter och skyldigheter som utlänningar bosatta i Finland inte har.
Läs mer om finska medborgares rättigheter och skyldigheter på InfoFinlands sida Finskt medborgarskap.
Det finländska samhället och dess verksamhet styrs av lagar.
Den viktigaste lagen är grundlagen( perustuslaki).
Alla som bor i Finland måste följa Finlands lag.
Också myndigheterna måste följa lagen.
Lagarna stiftas av riksdagen.
Vem som helst kan framföra ett klagomål till justitiekanslern (oikeuskansleri) eller till riksdagens justitieombudsman (eduskunnan oikeusasiamies) om man misstänker att en myndighet har brutit mot lagen.
Finland och alla som är bosatta i Finland måste dessutom följa Europeiska unionens lagar.
Finlands lagarfinska _ svenska _ engelska
Några lagar
Grundlagen
Med grundlagen stadgas till exempel de grundläggande rättigheterna för alla som är bosatta i Finland samt regler för hur den finska staten fungerar.
Information om grundlagenfinska _ svenska _ engelska _ ryska
Enligt lagen om likabehandling (Yhdenvertaisuuslaki) får ingen diskrimineras på grund av ålder, etniskt eller nationellt ursprung, nationalitet, språk, religion, övertygelse, åsikt, hälsotillstånd, funktionshinder, sexuell läggning eller av någon annan orsak som gäller hans eller hennes person.
Mer information om likabehandling hittar du på InfoFinlands sida Jämställdhet och likabehandling.
Lag om jämställdhet mellan kvinnor och män
Lagen om jämställdhet mellan kvinnor och män (Tasa-arvolaki) förbjuder diskriminering på grund av kön.
Enligt lagen om jämställdhet ska myndigheter, arbetsgivare och läroanstalter främja jämställdheten mellan kvinnor och män.
Mer information om jämställdhet hittar du på InfoFinlands sida Jämställdhet och likabehandling.
linkkiJämställdhetsombudsman:
Information om jämställdhetfinska _ svenska _ engelska
Barnskyddslag
Barnskyddslagen (Lastensuojelulaki) säger att alla barn bosatta i Finland har rätt till omsorg och en trygg uppväxtmiljö.
Mer information om barns rättigheter i Finland hittar du på InfoFinlands sida Barn.
Information om barnskyddslagenfinska _ svenska _ engelska _ ryska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
Konsumentens rättigheter
Alla som köper varor och tjänster är konsumenter.
Konsumentskyddslagen (Kuluttajansuojalaki) tryggar konsumentens rättigheter i Finland.
Du har rätt till gottgörelse till exempel då varan som du köpt har fel som inte du har orsakat.
Du kan till exempel ersättas med en felfri vara eller få dina pengar tillbaka.
Om en vara som du köpt har brister ska du först kontakt säljaren.
Om du inte kan komma överens om saken med säljaren, ta då kontakt med konsumentrådgivningen.
linkkiKonkurrens- och konsumentverket:
Konsumentrådgivningfinska _ svenska _ engelska
Information om konsumenträttigheterfinska _ svenska _ engelska
Grundläggande rättigheter
Alla som är bosatta i Finland har rättigheter och skyldigheter enligt lag.
Utlänningar som är bosatta i Finland har nästan samma rättigheter och skyldigheter som finska medborgare.
Följande rättigheter och skyldigheter gäller även utlänningar bosatta i Finland.
Rättigheter
Alla har rätt att bli jämlikt bemötta.
Ingen får behandlas annorlunda till exempel på grund av kön, ålder, religion eller handikapp.
Var och en får fritt yttra sina åsikter i tal och skrift.
Människor får ordna sammankomster och demonstrationer samt delta i dem.
En demonstration ska anmälas till polisen på förhand.
Ingen får dömas till döden eller torteras.
Alla kan själv välja var de vill bo och fritt röra sig i Finland.
Alla har rätt till integritetsskydd.
Ett brev som tillhör en annan person får inte läsas och en annan persons telefonsamtal får inte avlyssnas.
Var och en får själv välja sin religion.
Om man inte vill, måste man inte välja någon religion alls.
Utlänningar som bor stadigvarande i Finland och som har fyllt 18 år har rätt att rösta i kommunalval.
Utlänningar som har rösträtt i kommunalval har även rätt att ställa upp som kandidat i kommunalval.
EU-medborgare som har sin hemkommun i Finland kan rösta i val till Europaparlamentet i Finland om de har anmält sig till rösträttsregistret.
EU-medborgare som är i det finska rösträttsregistret kan också ställa upp som kandidat i Finlands Europaparlamentsval.
Läs mer om utlänningarnas rösträtt på InfoFinlands sida Val och röstning i Finland.
Skyldigheter
Alla som bor eller vistas i Finland måste följa Finlands lag.
Barn i åldern 7–17 år har läroplikt, det vill säga skyldighet att avlägga grundskolans lärokurs.
Ofta måste de som arbetar i Finland betala skatt på sin lön till Finland.
Alla har skyldighet att vittna inför domstol om de blir kallade.
Föräldrar är skyldiga att ta hand om sina barn.
Alla har skyldighet att hjälpa vid en olycka.
Läs mer om beskattningen i Finland på InfoFinlands sida Beskattning.
Finska medborgares rättigheter och skyldigheter
Finska medborgare har utöver det ovan nämnda också några ytterligare rättigheter och skyldigheter som utlänningar bosatta i Finland inte har.
Läs mer om finska medborgares rättigheter och skyldigheter på InfoFinlands sida Finskt medborgarskap.
Det finländska samhället och dess verksamhet styrs av lagar.
Den viktigaste lagen är grundlagen( perustuslaki).
Alla som bor i Finland måste följa Finlands lag.
Också myndigheterna måste följa lagen.
Lagarna stiftas av riksdagen.
Vem som helst kan framföra ett klagomål till justitiekanslern (oikeuskansleri) eller till riksdagens justitieombudsman (eduskunnan oikeusasiamies) om man misstänker att en myndighet har brutit mot lagen.
Finland och alla som är bosatta i Finland måste dessutom följa Europeiska unionens lagar.
Finlands lagarfinska _ svenska _ engelska
Några lagar
Grundlagen
Med grundlagen stadgas till exempel de grundläggande rättigheterna för alla som är bosatta i Finland samt regler för hur den finska staten fungerar.
Information om grundlagenfinska _ svenska _ engelska _ ryska
Enligt lagen om likabehandling (Yhdenvertaisuuslaki) får ingen diskrimineras på grund av ålder, etniskt eller nationellt ursprung, nationalitet, språk, religion, övertygelse, åsikt, hälsotillstånd, funktionshinder, sexuell läggning eller av någon annan orsak som gäller hans eller hennes person.
Mer information om likabehandling hittar du på InfoFinlands sida Jämställdhet och likabehandling.
Lag om jämställdhet mellan kvinnor och män
Lagen om jämställdhet mellan kvinnor och män (Tasa-arvolaki) förbjuder diskriminering på grund av kön.
Enligt lagen om jämställdhet ska myndigheter, arbetsgivare och läroanstalter främja jämställdheten mellan kvinnor och män.
Mer information om jämställdhet hittar du på InfoFinlands sida Jämställdhet och likabehandling.
linkkiJämställdhetsombudsman:
Information om jämställdhetfinska _ svenska _ engelska
Barnskyddslag
Barnskyddslagen (Lastensuojelulaki) säger att alla barn bosatta i Finland har rätt till omsorg och en trygg uppväxtmiljö.
Mer information om barns rättigheter i Finland hittar du på InfoFinlands sida Barn.
Information om barnskyddslagenfinska _ svenska _ engelska _ ryska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
Konsumentens rättigheter
Alla som köper varor och tjänster är konsumenter.
Konsumentskyddslagen (Kuluttajansuojalaki) tryggar konsumentens rättigheter i Finland.
Du har rätt till gottgörelse till exempel då varan som du köpt har fel som inte du har orsakat.
Du kan till exempel ersättas med en felfri vara eller få dina pengar tillbaka.
Om en vara som du köpt har brister ska du först kontakt säljaren.
Om du inte kan komma överens om saken med säljaren, ta då kontakt med konsumentrådgivningen.
linkkiKonkurrens- och konsumentverket:
Konsumentrådgivningfinska _ svenska _ engelska
Information om konsumenträttigheterfinska _ svenska _ engelska
Grundläggande rättigheter
Alla som är bosatta i Finland har rättigheter och skyldigheter enligt lag.
Utlänningar som är bosatta i Finland har nästan samma rättigheter och skyldigheter som finska medborgare.
Följande rättigheter och skyldigheter gäller även utlänningar bosatta i Finland.
Rättigheter
Alla har rätt att bli jämlikt bemötta.
Ingen får behandlas annorlunda till exempel på grund av kön, ålder, religion eller handikapp.
Var och en får fritt yttra sina åsikter i tal och skrift.
Människor får ordna sammankomster och demonstrationer samt delta i dem.
En demonstration ska anmälas till polisen på förhand.
Ingen får dömas till döden eller torteras.
Alla kan själv välja var de vill bo och fritt röra sig i Finland.
Alla har rätt till integritetsskydd.
Ett brev som tillhör en annan person får inte läsas och en annan persons telefonsamtal får inte avlyssnas.
Var och en får själv välja sin religion.
Om man inte vill, måste man inte välja någon religion alls.
Utlänningar som bor stadigvarande i Finland och som har fyllt 18 år har rätt att rösta i kommunalval.
Utlänningar som har rösträtt i kommunalval har även rätt att ställa upp som kandidat i kommunalval.
EU-medborgare som har sin hemkommun i Finland kan rösta i val till Europaparlamentet i Finland om de har anmält sig till rösträttsregistret.
EU-medborgare som är i det finska rösträttsregistret kan också ställa upp som kandidat i Finlands Europaparlamentsval.
Läs mer om utlänningarnas rösträtt på InfoFinlands sida Val och röstning i Finland.
Skyldigheter
Alla som bor eller vistas i Finland måste följa Finlands lag.
Barn i åldern 7–17 år har läroplikt, det vill säga skyldighet att avlägga grundskolans lärokurs.
Ofta måste de som arbetar i Finland betala skatt på sin lön till Finland.
Alla har skyldighet att vittna inför domstol om de blir kallade.
Föräldrar är skyldiga att ta hand om sina barn.
Alla har skyldighet att hjälpa vid en olycka.
Läs mer om beskattningen i Finland på InfoFinlands sida Beskattning.
Finska medborgares rättigheter och skyldigheter
Finska medborgare har utöver det ovan nämnda också några ytterligare rättigheter och skyldigheter som utlänningar bosatta i Finland inte har.
Läs mer om finska medborgares rättigheter och skyldigheter på InfoFinlands sida Finskt medborgarskap.
Det finländska samhället och dess verksamhet styrs av lagar.
Den viktigaste lagen är grundlagen( perustuslaki).
Alla som bor i Finland måste följa Finlands lag.
Också myndigheterna måste följa lagen.
Lagarna stiftas av riksdagen.
Vem som helst kan framföra ett klagomål till justitiekanslern (oikeuskansleri) eller till riksdagens justitieombudsman (eduskunnan oikeusasiamies) om man misstänker att en myndighet har brutit mot lagen.
Finland och alla som är bosatta i Finland måste dessutom följa Europeiska unionens lagar.
Finlands lagarfinska _ svenska _ engelska
Några lagar
Grundlagen
Med grundlagen stadgas till exempel de grundläggande rättigheterna för alla som är bosatta i Finland samt regler för hur den finska staten fungerar.
Information om grundlagenfinska _ svenska _ engelska _ ryska
Enligt lagen om likabehandling (Yhdenvertaisuuslaki) får ingen diskrimineras på grund av ålder, etniskt eller nationellt ursprung, nationalitet, språk, religion, övertygelse, åsikt, hälsotillstånd, funktionshinder, sexuell läggning eller av någon annan orsak som gäller hans eller hennes person.
Mer information om likabehandling hittar du på InfoFinlands sida Jämställdhet och likabehandling.
Lag om jämställdhet mellan kvinnor och män
Lagen om jämställdhet mellan kvinnor och män (Tasa-arvolaki) förbjuder diskriminering på grund av kön.
Enligt lagen om jämställdhet ska myndigheter, arbetsgivare och läroanstalter främja jämställdheten mellan kvinnor och män.
Mer information om jämställdhet hittar du på InfoFinlands sida Jämställdhet och likabehandling.
linkkiJämställdhetsombudsman:
Information om jämställdhetfinska _ svenska _ engelska
Barnskyddslag
Barnskyddslagen (Lastensuojelulaki) säger att alla barn bosatta i Finland har rätt till omsorg och en trygg uppväxtmiljö.
Mer information om barns rättigheter i Finland hittar du på InfoFinlands sida Barn.
Information om barnskyddslagenfinska _ svenska _ engelska _ ryska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
Konsumentens rättigheter
Alla som köper varor och tjänster är konsumenter.
Konsumentskyddslagen (Kuluttajansuojalaki) tryggar konsumentens rättigheter i Finland.
Du har rätt till gottgörelse till exempel då varan som du köpt har fel som inte du har orsakat.
Du kan till exempel ersättas med en felfri vara eller få dina pengar tillbaka.
Om en vara som du köpt har brister ska du först kontakt säljaren.
Om du inte kan komma överens om saken med säljaren, ta då kontakt med konsumentrådgivningen.
linkkiKonkurrens- och konsumentverket:
Konsumentrådgivningfinska _ svenska _ engelska
Information om konsumenträttigheterfinska _ svenska _ engelska
Röstning
I regel har alla finska medborgare som fyllt 18 år rätt att rösta vid val.
Vid kommunalval och Europaparlamentsval har dock också andra länders medborgare som bor i Finland rösträtt.
Också andra EU-länders medborgare som registrerat sig till rösträttsregistret i Finland har rösträtt vid Europaparlamentsval.
Medborgare i alla länder, vilka haft en hemkommun i Finland i minst två år, har rösträtt vid kommunalval.
Meddelandet om rösträtt vid ett val skickas hem till dig per post cirka en månad före valdagen.
Ditt röstningsställe har antecknats på meddelandekortet.
Om du röstar på valdagen, kan du rösta endast på det ställe som anges på kortet.
I alla val är det möjligt att rösta också före valdagen, under förhandsröstningstiden.
Om du röstar på förhand kan du rösta vid vilket allmänt förhandsröstningsställe som helst i Finland eller utomlands.
Kontakta magistraten på din hemort om meddelandet om rösträtt inte skickas hem till dig.
Du måste ha med ett ID-kort när du röstar.
Det lönar sig också att ta med meddelandet om rösträtt.
Kommunalval
Beslut i viktiga kommunala ärenden fattas av kommunfullmäktige (kunnanvaltuusto).
Ledamöterna i kommunfullmäktige, eller bara kommunfullmäktige, utses i kommunalval.
Kommunalval förrättas vart fjärde år.
Antalet kommunfullmäktige beror på kommunens invånarantal.
Vem kan rösta?
Du kan rösta i kommunalvalet om:
du är medborgare i Finland, ett annat EU-land, Norge eller Island och fyller 18 år senast på valdagen.
Dessutom ska den ifrågavarande kommunen vara din hemkommun senast den 51:a dagen före valdagen.
du är medborgare i vilket annat land som helst och fyller 18 år senast på valdagen.
Dessutom ska den ifrågavarande kommunen vara din hemkommun den 51:a dagen före valdagen.
Dessutom krävs det att du har haft din hemkommun i Finland i minst två år i rad.
Vem kan ställa upp som kandidat?
Kandidater kan nomineras av
partier som finns i partiregistret och
röstberättigade personer som har grundat en valmansförening.
Valmansföreningen ska ha minst tio medlemmar.
Kandidaten ska vara en person
som har rösträtt i kommunalval,
som har ifrågavarande kommun som hemkommun och
som inte står under förmyndarskap.
Information om kommunvalfinska _ svenska _ engelska
Riksdagsval
Riksdagen (eduskunta) är finska statens viktigaste organ för beslutsfattande.
Riksdagsledamöterna väljs i riksdagsval.
Riksdagsval förrättas vart fjärde år.
I riksdagsval är landet indelat i valkretsar.
Från varje valkrets väljs ett visst antal ledamöter.
Antalet ledamöter beror på invånarantalet i valkretsen.
Sammanlagt väljer man 200 riksdagsledamöter.
Vem kan rösta?
Du kan rösta i riksdagsval om du är finsk medborgare och fyller 18 år senast på valdagen.
Även utomlands bosatta finska medborgare har rösträtt.
Vem kan ställa upp som kandidat?
Kandidater kan nomineras av
partier som finns i partiregistret och
röstberättigade personer som har grundat en valmansförening.
Valmansföreningen ska ha minst 100 medlemmar.
Kandidaten ska vara en person
som har rösträtt i riksdagsval och
som inte står under förmyndarskap
Information om riksdagsvalfinska _ svenska _ engelska
linkkiRiksdagen:
Information om riksdagsvalfinska _ svenska _ engelska
Presidentval
Presidenten är Finlands statsöverhuvud.
Presidenten väljs i presidentval.
Presidentval förrättas vart sjätte år.
Samma person kan väljas till president högst två gånger.
Presidentvalet har vanligen två steg.
Om ingen av kandidaterna får mer än hälften av de givna rösterna vid första valomgången, förrättas en andra valomgång.
I den andra valomgången kandiderar de två kandidater som fick flest röster vid första valomgången.
Den person som får flest röster vid andra valomgången väljs till president.
Vem kan rösta?
Du kan rösta i presidentval om du är finsk medborgare och fyller 18 år senast på valdagen.
Även utomlands bosatta finska medborgare har rösträtt.
Vem kan ställa upp som kandidat?
Presidentkandidater kan nomineras av
de partier som har minst en riksdagsledamot,
röstberättigade personer som har grundat en valmansförening.
Valmansföreningen ska ha minst 20 000 medlemmar.
Kandidaten ska vara en person
som är infödd finsk medborgare,
som har rösträtt i presidentval och
som inte står under förmyndarskap.
Information om presidentvalfinska _ svenska _ engelska
Val till Europaparlamentet
I Europeiska unionens råd är regeringarna för medlemsländerna representerade.
Parlamentet har 754 ledamöter och tretton av dem har valts i Finland.
Parlamentsledamöterna utses genom val.
Valet förrättas vart femte år.
Vem kan rösta?
Du kan rösta i valet till Europaparlamentet om
du är finsk medborgare och fyller 18 år senast på valdagen,
du är medborgare i ett annat EU-land och fyller 18 år senast på valdagen.
Dessutom ska du ha hemkommun i Finland den 51:a dagen före valdagen.
Du måste också anmäla dig till rösträttsregistret i Finland.
Anmälningen ska göras till magistraten senast den 80:e dagen före valdagen.
I samma val kan du rösta i endast ett EU-land.
Vem kan ställa upp som kandidat?
Kandidater kan nomineras av
partier som finns i partiregistret och
röstberättigade personer som har grundat en valmansförening.
Valmansföreningen ska ha minst 2 000 medlemmar.
Kandidaten ska vara en person
som har rösträtt i val till Europaparlamentet och
som inte står under förmyndarskap
Information om Europaparlamentsvalfinska _ svenska _ engelska
Röstning
I regel har alla finska medborgare som fyllt 18 år rätt att rösta vid val.
Vid kommunalval och Europaparlamentsval har dock också andra länders medborgare som bor i Finland rösträtt.
Också andra EU-länders medborgare som registrerat sig till rösträttsregistret i Finland har rösträtt vid Europaparlamentsval.
Medborgare i alla länder, vilka haft en hemkommun i Finland i minst två år, har rösträtt vid kommunalval.
Meddelandet om rösträtt vid ett val skickas hem till dig per post cirka en månad före valdagen.
Ditt röstningsställe har antecknats på meddelandekortet.
Om du röstar på valdagen, kan du rösta endast på det ställe som anges på kortet.
I alla val är det möjligt att rösta också före valdagen, under förhandsröstningstiden.
Om du röstar på förhand kan du rösta vid vilket allmänt förhandsröstningsställe som helst i Finland eller utomlands.
Kontakta magistraten på din hemort om meddelandet om rösträtt inte skickas hem till dig.
Du måste ha med ett ID-kort när du röstar.
Det lönar sig också att ta med meddelandet om rösträtt.
Kommunalval
Beslut i viktiga kommunala ärenden fattas av kommunfullmäktige (kunnanvaltuusto).
Ledamöterna i kommunfullmäktige, eller bara kommunfullmäktige, utses i kommunalval.
Kommunalval förrättas vart fjärde år.
Antalet kommunfullmäktige beror på kommunens invånarantal.
Vem kan rösta?
Du kan rösta i kommunalvalet om:
du är medborgare i Finland, ett annat EU-land, Norge eller Island och fyller 18 år senast på valdagen.
Dessutom ska den ifrågavarande kommunen vara din hemkommun senast den 51:a dagen före valdagen.
du är medborgare i vilket annat land som helst och fyller 18 år senast på valdagen.
Dessutom ska den ifrågavarande kommunen vara din hemkommun den 51:a dagen före valdagen.
Dessutom krävs det att du har haft din hemkommun i Finland i minst två år i rad.
Vem kan ställa upp som kandidat?
Kandidater kan nomineras av
partier som finns i partiregistret och
röstberättigade personer som har grundat en valmansförening.
Valmansföreningen ska ha minst tio medlemmar.
Kandidaten ska vara en person
som har rösträtt i kommunalval,
som har ifrågavarande kommun som hemkommun och
som inte står under förmyndarskap.
Information om kommunvalfinska _ svenska _ engelska
Riksdagsval
Riksdagen (eduskunta) är finska statens viktigaste organ för beslutsfattande.
Riksdagsledamöterna väljs i riksdagsval.
Riksdagsval förrättas vart fjärde år.
I riksdagsval är landet indelat i valkretsar.
Från varje valkrets väljs ett visst antal ledamöter.
Antalet ledamöter beror på invånarantalet i valkretsen.
Sammanlagt väljer man 200 riksdagsledamöter.
Vem kan rösta?
Du kan rösta i riksdagsval om du är finsk medborgare och fyller 18 år senast på valdagen.
Även utomlands bosatta finska medborgare har rösträtt.
Vem kan ställa upp som kandidat?
Kandidater kan nomineras av
partier som finns i partiregistret och
röstberättigade personer som har grundat en valmansförening.
Valmansföreningen ska ha minst 100 medlemmar.
Kandidaten ska vara en person
som har rösträtt i riksdagsval och
som inte står under förmyndarskap
Information om riksdagsvalfinska _ svenska _ engelska
linkkiRiksdagen:
Information om riksdagsvalfinska _ svenska _ engelska
Presidentval
Presidenten är Finlands statsöverhuvud.
Presidenten väljs i presidentval.
Presidentval förrättas vart sjätte år.
Samma person kan väljas till president högst två gånger.
Presidentvalet har vanligen två steg.
Om ingen av kandidaterna får mer än hälften av de givna rösterna vid första valomgången, förrättas en andra valomgång.
I den andra valomgången kandiderar de två kandidater som fick flest röster vid första valomgången.
Den person som får flest röster vid andra valomgången väljs till president.
Vem kan rösta?
Du kan rösta i presidentval om du är finsk medborgare och fyller 18 år senast på valdagen.
Även utomlands bosatta finska medborgare har rösträtt.
Vem kan ställa upp som kandidat?
Presidentkandidater kan nomineras av
de partier som har minst en riksdagsledamot,
röstberättigade personer som har grundat en valmansförening.
Valmansföreningen ska ha minst 20 000 medlemmar.
Kandidaten ska vara en person
som är infödd finsk medborgare,
som har rösträtt i presidentval och
som inte står under förmyndarskap.
Information om presidentvalfinska _ svenska _ engelska
Val till Europaparlamentet
I Europeiska unionens råd är regeringarna för medlemsländerna representerade.
Parlamentet har 754 ledamöter och tretton av dem har valts i Finland.
Parlamentsledamöterna utses genom val.
Valet förrättas vart femte år.
Vem kan rösta?
Du kan rösta i valet till Europaparlamentet om
du är finsk medborgare och fyller 18 år senast på valdagen,
du är medborgare i ett annat EU-land och fyller 18 år senast på valdagen.
Dessutom ska du ha hemkommun i Finland den 51:a dagen före valdagen.
Du måste också anmäla dig till rösträttsregistret i Finland.
Anmälningen ska göras till magistraten senast den 80:e dagen före valdagen.
I samma val kan du rösta i endast ett EU-land.
Vem kan ställa upp som kandidat?
Kandidater kan nomineras av
partier som finns i partiregistret och
röstberättigade personer som har grundat en valmansförening.
Valmansföreningen ska ha minst 2 000 medlemmar.
Kandidaten ska vara en person
som har rösträtt i val till Europaparlamentet och
som inte står under förmyndarskap
Information om Europaparlamentsvalfinska _ svenska _ engelska
Instruktionsfilmer om att rösta
Röstning
I regel har alla finska medborgare som fyllt 18 år rätt att rösta vid val.
Vid kommunalval och Europaparlamentsval har dock också andra länders medborgare som bor i Finland rösträtt.
Också andra EU-länders medborgare som registrerat sig till rösträttsregistret i Finland har rösträtt vid Europaparlamentsval.
Medborgare i alla länder, vilka haft en hemkommun i Finland i minst två år, har rösträtt vid kommunalval.
Meddelandet om rösträtt vid ett val skickas hem till dig per post cirka en månad före valdagen.
Ditt röstningsställe har antecknats på meddelandekortet.
Om du röstar på valdagen, kan du rösta endast på det ställe som anges på kortet.
I alla val är det möjligt att rösta också före valdagen, under förhandsröstningstiden.
Om du röstar på förhand kan du rösta vid vilket allmänt förhandsröstningsställe som helst i Finland eller utomlands.
Kontakta magistraten på din hemort om meddelandet om rösträtt inte skickas hem till dig.
Du måste ha med ett ID-kort när du röstar.
Det lönar sig också att ta med meddelandet om rösträtt.
Kommunalval
Beslut i viktiga kommunala ärenden fattas av kommunfullmäktige (kunnanvaltuusto).
Ledamöterna i kommunfullmäktige, eller bara kommunfullmäktige, utses i kommunalval.
Kommunalval förrättas vart fjärde år.
Antalet kommunfullmäktige beror på kommunens invånarantal.
Vem kan rösta?
Du kan rösta i kommunalvalet om:
du är medborgare i Finland, ett annat EU-land, Norge eller Island och fyller 18 år senast på valdagen.
Dessutom ska den ifrågavarande kommunen vara din hemkommun senast den 51:a dagen före valdagen.
du är medborgare i vilket annat land som helst och fyller 18 år senast på valdagen.
Dessutom ska den ifrågavarande kommunen vara din hemkommun den 51:a dagen före valdagen.
Dessutom krävs det att du har haft din hemkommun i Finland i minst två år i rad.
Vem kan ställa upp som kandidat?
Kandidater kan nomineras av
partier som finns i partiregistret och
röstberättigade personer som har grundat en valmansförening.
Valmansföreningen ska ha minst tio medlemmar.
Kandidaten ska vara en person
som har rösträtt i kommunalval,
som har ifrågavarande kommun som hemkommun och
som inte står under förmyndarskap.
Information om kommunvalfinska _ svenska _ engelska
Riksdagsval
Riksdagen (eduskunta) är finska statens viktigaste organ för beslutsfattande.
Riksdagsledamöterna väljs i riksdagsval.
Riksdagsval förrättas vart fjärde år.
I riksdagsval är landet indelat i valkretsar.
Från varje valkrets väljs ett visst antal ledamöter.
Antalet ledamöter beror på invånarantalet i valkretsen.
Sammanlagt väljer man 200 riksdagsledamöter.
Vem kan rösta?
Du kan rösta i riksdagsval om du är finsk medborgare och fyller 18 år senast på valdagen.
Även utomlands bosatta finska medborgare har rösträtt.
Vem kan ställa upp som kandidat?
Kandidater kan nomineras av
partier som finns i partiregistret och
röstberättigade personer som har grundat en valmansförening.
Valmansföreningen ska ha minst 100 medlemmar.
Kandidaten ska vara en person
som har rösträtt i riksdagsval och
som inte står under förmyndarskap
Information om riksdagsvalfinska _ svenska _ engelska
linkkiRiksdagen:
Information om riksdagsvalfinska _ svenska _ engelska
Presidentval
Presidenten är Finlands statsöverhuvud.
Presidenten väljs i presidentval.
Presidentval förrättas vart sjätte år.
Samma person kan väljas till president högst två gånger.
Presidentvalet har vanligen två steg.
Om ingen av kandidaterna får mer än hälften av de givna rösterna vid första valomgången, förrättas en andra valomgång.
I den andra valomgången kandiderar de två kandidater som fick flest röster vid första valomgången.
Den person som får flest röster vid andra valomgången väljs till president.
Vem kan rösta?
Du kan rösta i presidentval om du är finsk medborgare och fyller 18 år senast på valdagen.
Även utomlands bosatta finska medborgare har rösträtt.
Vem kan ställa upp som kandidat?
Presidentkandidater kan nomineras av
de partier som har minst en riksdagsledamot,
röstberättigade personer som har grundat en valmansförening.
Valmansföreningen ska ha minst 20 000 medlemmar.
Kandidaten ska vara en person
som är infödd finsk medborgare,
som har rösträtt i presidentval och
som inte står under förmyndarskap.
Information om presidentvalfinska _ svenska _ engelska
Val till Europaparlamentet
I Europeiska unionens råd är regeringarna för medlemsländerna representerade.
Parlamentet har 754 ledamöter och tretton av dem har valts i Finland.
Parlamentsledamöterna utses genom val.
Valet förrättas vart femte år.
Vem kan rösta?
Du kan rösta i valet till Europaparlamentet om
du är finsk medborgare och fyller 18 år senast på valdagen,
du är medborgare i ett annat EU-land och fyller 18 år senast på valdagen.
Dessutom ska du ha hemkommun i Finland den 51:a dagen före valdagen.
Du måste också anmäla dig till rösträttsregistret i Finland.
Anmälningen ska göras till magistraten senast den 80:e dagen före valdagen.
I samma val kan du rösta i endast ett EU-land.
Vem kan ställa upp som kandidat?
Kandidater kan nomineras av
partier som finns i partiregistret och
röstberättigade personer som har grundat en valmansförening.
Valmansföreningen ska ha minst 2 000 medlemmar.
Kandidaten ska vara en person
som har rösträtt i val till Europaparlamentet och
som inte står under förmyndarskap
Information om Europaparlamentsvalfinska _ svenska _ engelska
Instruktionsfilmer om att rösta
Statsförvaltningen
Finland är en republik.
De högsta statliga organen är riksdagen, presidenten och statsrådet, det vill säga regeringen.
Riksdagen
Riksdagen (eduskunta) stiftar lagarna i Finland och beslutar om statens budget.
Dessutom övervakar riksdagen regeringens verksamhet.
I riksdagen sitter 200 riksdagsledamöter.
Riksdagsledamöterna utses genom val för fyra år i taget.
På InfoFinlands sida Val och röstning i Finland finns information om vem som kan rösta i riksdagsvalet.
Finlands statsöverhuvud är republikens president (tasavallan presidentti).
Presidenten utses genom val.
Presidentens mandat är sex år.
Samma person kan väljas till president för högst två mandatperioder efter varandra, det vill säga för tolv år.
stadfäster lagarna,
utnämner högsta tjänstemän, leder
Finlands utrikespolitik i samverkan med statsrådet och
är överbefälhavare för Finlands försvarsmakt.
På InfoFinlands sida Val och röstning i Finland finns information om vem som kan rösta i presidentvalet.
Regeringen (hallitus) består av statsministern och de andra ministrarna.
Riksdagen utser statsministern och republikens president tillsätter honom eller henne.
De övriga ministrarna utnämner presidenten i enlighet med förslag av statsministern.
Regeringen bereder och verkställer riksdagens beslut.
Regeringen svarar för sin verksamhet inför riksdagen, vilket betyder att ministrarna ska ha riksdagens förtroende.
Ministerierna bereder de ärenden som regeringen fattar beslut om.
Ministrarna leder arbetet för ministeriernas tjänstemän.
Under ministerierna verkar flera ämbetsverk och inrättningar.
Till exempel är Migrationsverket ett ämbetsverk som lyder under inrikesministeriet.
Information om förvaltningen i Finlandfinska _ svenska _ engelska
linkkiRiksdagen:
Information om riksdagenfinska _ svenska _ engelska
Regeringens verksamhetfinska _ svenska _ engelska
Den nuvarande regeringenfinska _ svenska _ engelska
Information om presidentens uppgifterfinska _ svenska _ engelska
Statens lokalförvaltning
Med statens lokalförvaltning avses de myndigheter som sköter statliga ärenden i en viss region.
Följande myndigheter hör till statens lokalförvaltning:
polisen,
åklagarväsendet,
utsökningen,
arbets- och näringsbyråerna,
skattebyråerna,
tullen,
rättshjälpsbyråerna.
Mer information om myndigheterna och deras uppgifter hittar du på InfoFinlands sida Viktiga myndigheter.
Regionförvaltningen
Regionförvaltningen sköts av regionförvaltningsverken (aluehallintovirasto) och ELY-centralerna, det vill säga närings-, trafik- och miljöcentralerna (elinkeino- liikenne- ja ympäristökeskus).
I Finland finns sex regionförvaltningsverk.
Regionförvaltningsverken sköter om verkställighets- och tillsynsuppgifter rörande Finlands lag i sina egna regioner.
Regionförvaltningsverken sköter följande:
grundläggande service, rättsskydd och tillstånd
räddningsväsendet och beredskap
polisen
arbetarskydd
miljötillstånd
I Finland finns femton ELY-centraler.
I deras uppgifter ingår till exempel
företagsrådgivning
miljöskydd
främjande av trafiksäkerhet
främjande av invandrares integration
linkkiFinansministeriet:
Statens lokalförvaltningfinska _ svenska
linkkiFinansministeriet:
Regionförvaltningenfinska _ svenska
linkkiRegionförvaltningsverket:
Regionförvaltningsverkenfinska _ svenska _ engelska
ELY-centralernafinska _ svenska _ engelska
Kommuner
Finland är indelat i kommuner.
Kommunerna har självstyre, vilket betyder att de själva kan besluta om ärenden i kommunen.
Kommunerna har beskattningsrätt, det vill säga rätt att uppbära kommunalskatt av sina invånare.
Kommunerna är skyldiga att ordna många olika tjänster för sina invånare.
Sådana tjänster är till exempel hälsovård, barndagvård och undervisning.
De kan dessutom tillhandahålla andra tjänster.
Mer information hittar du på InfoFinlands sida Hemkommun i Finland.
Beslut i kommunens ärenden fattas av kommunfullmäktige.
Ledamöterna till kommunfullmäktige utses i kommunalval som förrättas vart fjärde år.
Fullmäktige väljer ledamöterna till kommunstyrelsen, som har som uppgift att bereda och verkställa fullmäktiges beslut.
På InfoFinlands sida Val och röstning i Finland finns information om vem som kan rösta i kommunaval.
Kommunförvaltningenfinska _ svenska _ engelska
linkkiKommunförbundet:
Kommunernas verksamhetfinska _ svenska
Statsförvaltningen
Finland är en republik.
De högsta statliga organen är riksdagen, presidenten och statsrådet, det vill säga regeringen.
Riksdagen
Riksdagen (eduskunta) stiftar lagarna i Finland och beslutar om statens budget.
Dessutom övervakar riksdagen regeringens verksamhet.
I riksdagen sitter 200 riksdagsledamöter.
Riksdagsledamöterna utses genom val för fyra år i taget.
På InfoFinlands sida Val och röstning i Finland finns information om vem som kan rösta i riksdagsvalet.
Finlands statsöverhuvud är republikens president (tasavallan presidentti).
Presidenten utses genom val.
Presidentens mandat är sex år.
Samma person kan väljas till president för högst två mandatperioder efter varandra, det vill säga för tolv år.
stadfäster lagarna,
utnämner högsta tjänstemän, leder
Finlands utrikespolitik i samverkan med statsrådet och
är överbefälhavare för Finlands försvarsmakt.
På InfoFinlands sida Val och röstning i Finland finns information om vem som kan rösta i presidentvalet.
Regeringen (hallitus) består av statsministern och de andra ministrarna.
Riksdagen utser statsministern och republikens president tillsätter honom eller henne.
De övriga ministrarna utnämner presidenten i enlighet med förslag av statsministern.
Regeringen bereder och verkställer riksdagens beslut.
Regeringen svarar för sin verksamhet inför riksdagen, vilket betyder att ministrarna ska ha riksdagens förtroende.
Ministerierna bereder de ärenden som regeringen fattar beslut om.
Ministrarna leder arbetet för ministeriernas tjänstemän.
Under ministerierna verkar flera ämbetsverk och inrättningar.
Till exempel är Migrationsverket ett ämbetsverk som lyder under inrikesministeriet.
Information om förvaltningen i Finlandfinska _ svenska _ engelska
linkkiRiksdagen:
Information om riksdagenfinska _ svenska _ engelska
Regeringens verksamhetfinska _ svenska _ engelska
Den nuvarande regeringenfinska _ svenska _ engelska
Information om presidentens uppgifterfinska _ svenska _ engelska
Statens lokalförvaltning
Med statens lokalförvaltning avses de myndigheter som sköter statliga ärenden i en viss region.
Följande myndigheter hör till statens lokalförvaltning:
polisen,
åklagarväsendet,
utsökningen,
arbets- och näringsbyråerna,
skattebyråerna,
tullen,
rättshjälpsbyråerna.
Mer information om myndigheterna och deras uppgifter hittar du på InfoFinlands sida Viktiga myndigheter.
Regionförvaltningen
Regionförvaltningen sköts av regionförvaltningsverken (aluehallintovirasto) och ELY-centralerna, det vill säga närings-, trafik- och miljöcentralerna (elinkeino- liikenne- ja ympäristökeskus).
I Finland finns sex regionförvaltningsverk.
Regionförvaltningsverken sköter om verkställighets- och tillsynsuppgifter rörande Finlands lag i sina egna regioner.
Regionförvaltningsverken sköter följande:
grundläggande service, rättsskydd och tillstånd
räddningsväsendet och beredskap
polisen
arbetarskydd
miljötillstånd
I Finland finns femton ELY-centraler.
I deras uppgifter ingår till exempel
företagsrådgivning
miljöskydd
främjande av trafiksäkerhet
främjande av invandrares integration
linkkiFinansministeriet:
Statens lokalförvaltningfinska _ svenska
linkkiFinansministeriet:
Regionförvaltningenfinska _ svenska
linkkiRegionförvaltningsverket:
Regionförvaltningsverkenfinska _ svenska _ engelska
ELY-centralernafinska _ svenska _ engelska
Kommuner
Finland är indelat i kommuner.
Kommunerna har självstyre, vilket betyder att de själva kan besluta om ärenden i kommunen.
Kommunerna har beskattningsrätt, det vill säga rätt att uppbära kommunalskatt av sina invånare.
Kommunerna är skyldiga att ordna många olika tjänster för sina invånare.
Sådana tjänster är till exempel hälsovård, barndagvård och undervisning.
De kan dessutom tillhandahålla andra tjänster.
Mer information hittar du på InfoFinlands sida Hemkommun i Finland.
Beslut i kommunens ärenden fattas av kommunfullmäktige.
Ledamöterna till kommunfullmäktige utses i kommunalval som förrättas vart fjärde år.
Fullmäktige väljer ledamöterna till kommunstyrelsen, som har som uppgift att bereda och verkställa fullmäktiges beslut.
På InfoFinlands sida Val och röstning i Finland finns information om vem som kan rösta i kommunaval.
Kommunförvaltningenfinska _ svenska _ engelska
linkkiKommunförbundet:
Kommunernas verksamhetfinska _ svenska
Statsförvaltningen
Finland är en republik.
De högsta statliga organen är riksdagen, presidenten och statsrådet, det vill säga regeringen.
Riksdagen
Riksdagen (eduskunta) stiftar lagarna i Finland och beslutar om statens budget.
Dessutom övervakar riksdagen regeringens verksamhet.
I riksdagen sitter 200 riksdagsledamöter.
Riksdagsledamöterna utses genom val för fyra år i taget.
På InfoFinlands sida Val och röstning i Finland finns information om vem som kan rösta i riksdagsvalet.
Finlands statsöverhuvud är republikens president (tasavallan presidentti).
Presidenten utses genom val.
Presidentens mandat är sex år.
Samma person kan väljas till president för högst två mandatperioder efter varandra, det vill säga för tolv år.
stadfäster lagarna,
utnämner högsta tjänstemän, leder
Finlands utrikespolitik i samverkan med statsrådet och
är överbefälhavare för Finlands försvarsmakt.
På InfoFinlands sida Val och röstning i Finland finns information om vem som kan rösta i presidentvalet.
Regeringen (hallitus) består av statsministern och de andra ministrarna.
Riksdagen utser statsministern och republikens president tillsätter honom eller henne.
De övriga ministrarna utnämner presidenten i enlighet med förslag av statsministern.
Regeringen bereder och verkställer riksdagens beslut.
Regeringen svarar för sin verksamhet inför riksdagen, vilket betyder att ministrarna ska ha riksdagens förtroende.
Ministerierna bereder de ärenden som regeringen fattar beslut om.
Ministrarna leder arbetet för ministeriernas tjänstemän.
Under ministerierna verkar flera ämbetsverk och inrättningar.
Till exempel är Migrationsverket ett ämbetsverk som lyder under inrikesministeriet.
Information om förvaltningen i Finlandfinska _ svenska _ engelska
linkkiRiksdagen:
Information om riksdagenfinska _ svenska _ engelska
Regeringens verksamhetfinska _ svenska _ engelska
Den nuvarande regeringenfinska _ svenska _ engelska
Information om presidentens uppgifterfinska _ svenska _ engelska
Statens lokalförvaltning
Med statens lokalförvaltning avses de myndigheter som sköter statliga ärenden i en viss region.
Följande myndigheter hör till statens lokalförvaltning:
polisen,
åklagarväsendet,
utsökningen,
arbets- och näringsbyråerna,
skattebyråerna,
tullen,
rättshjälpsbyråerna.
Mer information om myndigheterna och deras uppgifter hittar du på InfoFinlands sida Viktiga myndigheter.
Regionförvaltningen
Regionförvaltningen sköts av regionförvaltningsverken (aluehallintovirasto) och ELY-centralerna, det vill säga närings-, trafik- och miljöcentralerna (elinkeino- liikenne- ja ympäristökeskus).
I Finland finns sex regionförvaltningsverk.
Regionförvaltningsverken sköter om verkställighets- och tillsynsuppgifter rörande Finlands lag i sina egna regioner.
Regionförvaltningsverken sköter följande:
grundläggande service, rättsskydd och tillstånd
räddningsväsendet och beredskap
polisen
arbetarskydd
miljötillstånd
I Finland finns femton ELY-centraler.
I deras uppgifter ingår till exempel
företagsrådgivning
miljöskydd
främjande av trafiksäkerhet
främjande av invandrares integration
linkkiFinansministeriet:
Statens lokalförvaltningfinska _ svenska
linkkiFinansministeriet:
Regionförvaltningenfinska _ svenska
linkkiRegionförvaltningsverket:
Regionförvaltningsverkenfinska _ svenska _ engelska
ELY-centralernafinska _ svenska _ engelska
Kommuner
Finland är indelat i kommuner.
Kommunerna har självstyre, vilket betyder att de själva kan besluta om ärenden i kommunen.
Kommunerna har beskattningsrätt, det vill säga rätt att uppbära kommunalskatt av sina invånare.
Kommunerna är skyldiga att ordna många olika tjänster för sina invånare.
Sådana tjänster är till exempel hälsovård, barndagvård och undervisning.
De kan dessutom tillhandahålla andra tjänster.
Mer information hittar du på InfoFinlands sida Hemkommun i Finland.
Beslut i kommunens ärenden fattas av kommunfullmäktige.
Ledamöterna till kommunfullmäktige utses i kommunalval som förrättas vart fjärde år.
Fullmäktige väljer ledamöterna till kommunstyrelsen, som har som uppgift att bereda och verkställa fullmäktiges beslut.
På InfoFinlands sida Val och röstning i Finland finns information om vem som kan rösta i kommunaval.
Kommunförvaltningenfinska _ svenska _ engelska
linkkiKommunförbundet:
Kommunernas verksamhetfinska _ svenska
På den här sidan har vi samlat länkar till andra webbplatser på språk som inte finns bland InfoFinlands urval av språk.
InfoFinland är en webbtjänst på 12 språk där alla språkversioner är identiska.
Du hittar urvalet av språk i tjänsten i menyn uppe på sidan.
Tyska
Thai
Kurdiska
Polska
Portugisiska
Rumänska
Tyska
Flytta till Finland
linkkiEuropa.eu:
EU-länderfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Rådgivning för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropa.eu:
Information för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
Arbete och entreprenörskap
linkkiArbetshälsoinstitutet:
Handboken Jobba i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ kurdiska _ tyska _ thai _ vietnamesiska
linkkiEuropass.eu:
Information om CVfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropass.eu:
CV-mallarfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiWebbtjänsten Suomi.fi:
Arbetsavtalsmallar på olika språkfinska _ svenska _ engelska _ ryska _ estniska _ franska _ tyska
linkkiEuropeiska unionen:
Information om att arbeta och driva ett företag i den europeiska unionenfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEures-portalen:
information om arbetsplatser i Europafinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropeiska arbetsmiljöbyrån:
Information om arbetarskyddfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Ta med dig dina arbetslöshetsförmånerfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Finska och svenska språket
linkkiEuropass.eu:
Utvärdera nivån på din språkkunskapfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Nybörjarkurs i finska, Tavataan taasengelska _ franska _ tyska _ bulgariska
linkkiWordDive:
Nybörjarkurs i finskafinska _ svenska _ engelska _ ryska _ kinesiska _ tyska
Webbkurs med många hjälpspråksvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ portugisiska
linkkiWordDive:
Finskans grammatikfinska _ svenska _ engelska _ ryska _ spanska _ tyska _ japanska
Boende
Heminkvarteringengelska _ franska _ spanska _ kinesiska _ tyska _ portugisiska _ italienska
Utbildning
linkkiUtbildningsstyrelsen:
Eget språk, eget sinnefinska _ engelska _ ryska _ estniska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ burmesiska _ bosniska
linkkiStudentexamensnämnden:
Information om studentexamenfinska _ svenska _ engelska _ franska _ tyska
Hälsa
linkkiNödcentralsverket:
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
linkkiEuropeiska kommissionen:
Europeiska sjukvårdskortetfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Privat psykoterapitjänst på Internetfinska _ svenska _ engelska _ ryska _ franska _ spanska _ turkiska _ kinesiska _ tyska _ portugisiska _ norska
_ holländska _ japanska _ italienska
_ danska
Hjälp till diskrimineringsofferfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ thai _ vietnamesiska _ portugisiska _ tagalog _ polska
linkkiBrottsofferjouren:
Hjälp för brottsofferfinska _ svenska _ engelska
linkkiBortförda barn rf:
Stöd och information för offer för barnkidnappningfinska _ svenska _ engelska _ turkiska _ arabiska _ tyska _ italienska
_ danska
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Information om Finland
Information om Finlandengelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ portugisiska
linkkiVisitFinland.com:
Information om Finland till turistersvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ japanska _ italienska
Information om finländska sederengelska _ spanska _ kinesiska _ tyska _ portugisiska
Information om Finlands historiaengelska _ ryska _ franska _ spanska _ tyska _ portugisiska
linkkiSkype:
Förmånliga utlandssamtalfinska _ svenska _ engelska _ ryska _ estniska _ franska _ spanska _ turkiska _ kinesiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ ungerska _ japanska
Länder som är anslutna till Apostilleavtaletengelska _ franska _ spanska _ tyska _ portugisiska
Thai
Arbete och entreprenörskap
linkkiArbetshälsoinstitutet:
Handboken Jobba i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ kurdiska _ tyska _ thai _ vietnamesiska
Guide för arbets- och näringsbyråns invandrarkunder(pdf, 5,1 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska _ kurdiska _ thai _ vietnamesiska
linkkiTE-tjänster:
Videoklipp och broschyrer för invandrarefinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska
Utbildning
linkkiKervo stad:
Så här använder du Wilma(pdf, 239 kt)finska _ engelska _ ryska _ estniska _ turkiska _ kurdiska _ thai _ vietnamesiska
Hälsä
linkkiStödcentralen Hilma för handikappade invandrare:
Serviceguide för handikappade invandrare(pdf, 797,26)finska _ svenska _ engelska _ ryska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ thai _ burmesiska
linkkiHivpoint:
Broschyren Information om sexuellt överförda sjukdomar(pdf, 1500kt)finska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Rådgivning för personer som säljer sexuella tjänsterfinska _ engelska
Anvisning för identifiering av bröstcancer(pdf, 440kt)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ kinesiska _ thai _ rumänska _ samiska
Familij
Handbok för familjer med två kulturer (pdf, 4,74 Mt)finska _ engelska _ ryska _ franska _ spanska _ thai
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Hjälp till diskrimineringsofferfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ thai _ vietnamesiska _ portugisiska _ tagalog _ polska
linkkiBrottsofferjouren:
Hjälp för brottsofferfinska _ svenska _ engelska
Hjälp till offer för människohandelfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska _ polska _ rumänska _ bulgariska
Fritid
linkkiFinlands Simundervisnings- och Livräddningsförbund rf:
Kom till simhallen!(pdf, 2 MB)finska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ arabiska _ kurdiska _ thai
Medborgarinstitut i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Information om Finland
linkkiArbets- och näringsministeriet:
Guiden Välkommen till Finland(pdf, 3,40 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
Kurdiska
Flytta till Finland
Information för flyktingarfinska _ engelska _ franska _ persiska _ arabiska _ kurdiska
Broschyren Information till asylsökandefinska _ svenska _ engelska _ ryska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
Arbete och entreprenörskap
linkkiArbetshälsoinstitutet:
Handboken Jobba i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ kurdiska _ tyska _ thai _ vietnamesiska
Guiden Bli företagare i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ turkiska _ kinesiska _ arabiska _ kurdiska
Guide om att grunda ett företagfinska _ engelska _ kinesiska
Guide för arbets- och näringsbyråns invandrarkunder(pdf, 5,1 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska _ kurdiska _ thai _ vietnamesiska
linkkiTE-tjänster:
Videoklipp och broschyrer för invandrarefinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska
linkkiKervo stad:
Så här använder du Wilma(pdf, 239 kt)finska _ engelska _ ryska _ estniska _ turkiska _ kurdiska _ thai _ vietnamesiska
linkki4V:
Tips för boende(pdf, 1,5 Mt)finska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Utbildning
linkkiKervo stad:
Så här använder du Wilma(pdf, 239 kt)finska _ engelska _ ryska _ estniska _ turkiska _ kurdiska _ thai _ vietnamesiska
Hälsä
linkkiNödcentralsverket:
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
linkkiStödcentralen Hilma för funktionshindrade invandrare :
Handbok med ordlista i hälso- och sjukvård på finska(pdf, 341,02 kt)finska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska
linkkiFöreningen för Mental Hälsa i Finland:
Information om mental hälsafinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
linkkiTuberkuloosi.fi:
Information om tuberkulosfinska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
linkkiStödcentralen Hilma för handikappade invandrare:
Stöd och hjälp för handikappade invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ persiska _ arabiska _ kurdiska
linkkiStödcentralen Hilma för handikappade invandrare:
Serviceguide för handikappade invandrare(pdf, 797,26)finska _ svenska _ engelska _ ryska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ thai _ burmesiska
linkkiSäg nej till droger -projektet:
Information om droger och faror som anknyter till dem särskilt för ungafinska _ somaliska _ arabiska _ kurdiska _ albanska
Familij
Uppfostring av barn i Finland(pdf, 8,08 Mt)finska _ engelska _ ryska _ somaliska _ kurdiska _ albanska _ burmesiska
Information om barnskyddslagenfinska _ svenska _ engelska _ ryska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
linkkiUtbildningsstyrelsen:
Eget språk, eget sinnefinska _ engelska _ ryska _ estniska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ burmesiska _ bosniska
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Hjälp till diskrimineringsofferfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ thai _ vietnamesiska _ portugisiska _ tagalog _ polska
Depression(pdf, 110,37 kt)finska _ engelska _ ryska _ franska _ somaliska _ turkiska _ persiska _ arabiska _ kurdiska _ albanska _ vietnamesiska _ burmesiska _ bosniska _ serbiska _ swahili
Information om posttraumatiskt stressyndromfinska _ engelska _ ryska _ franska _ somaliska _ turkiska _ persiska _ arabiska _ kurdiska _ albanska _ vietnamesiska _ burmesiska _ bosniska _ serbiska _ swahili
linkkiBrottsofferjouren:
Hjälp för brottsofferfinska _ svenska _ engelska
linkkiAndra ämbetsverk:
Broschyr om besöksförbud(pdf, 418,92 kt)finska _ svenska _ engelska
Diskrimineringsombudsmannenfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ persiska _ arabiska _ kurdiska
Hjälp till offer för människohandelfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska _ polska _ rumänska _ bulgariska
Information om krissituationer och sorgfinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Fritid
linkkiFinlands Simundervisnings- och Livräddningsförbund rf:
Kom till simhallen!(pdf, 2 MB)finska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ arabiska _ kurdiska _ thai
Medborgarinstitut i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Polska
Flytta till Finland
linkkiEuropa.eu:
EU-länderfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Rådgivning för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropa.eu:
Information för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
Arbete och entreprenörskap
linkkiArbets- och näringsbyrån:
Broschyren Jobba i Finland(pdf, 5,51 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ polska
linkkiEures-portalen:
information om arbetsplatser i Europafinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropass.eu:
Information om CVfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropass.eu:
CV-mallarfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropeiska arbetsmiljöbyrån:
Information om arbetarskyddfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Ta med dig dina arbetslöshetsförmånerfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Finska och svenska språket
linkkiEuropass.eu:
Utvärdera nivån på din språkkunskapfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Hälsä
linkkiEuropeiska kommissionen:
Europeiska sjukvårdskortetfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Hjälp till diskrimineringsofferfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ thai _ vietnamesiska _ portugisiska _ tagalog _ polska
linkkiBrottsofferjouren:
Hjälp för brottsofferfinska _ svenska _ engelska
Hjälp till offer för människohandelfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska _ polska _ rumänska _ bulgariska
Portugisiska
Flytta till Finland
linkkiEuropa.eu:
EU-länderfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Rådgivning för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropa.eu:
Information för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
Arbete och entreprenörskap
linkkiEures-portalen:
information om arbetsplatser i Europafinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropass.eu:
Information om CVfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropass.eu:
CV-mallarfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropeiska arbetsmiljöbyrån:
Information om arbetarskyddfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Ta med dig dina arbetslöshetsförmånerfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Finska och svenska språket
linkkiEuropass.eu:
Utvärdera nivån på din språkkunskapfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Webbkurs med många hjälpspråksvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ portugisiska
Hälsä
linkkiEuropeiska kommissionen:
Europeiska sjukvårdskortetfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Privat psykoterapitjänst på Internetfinska _ svenska _ engelska _ ryska _ franska _ spanska _ turkiska _ kinesiska _ tyska _ portugisiska _ norska
_ holländska _ japanska _ italienska
_ danska
Hjälp till diskrimineringsofferfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ thai _ vietnamesiska _ portugisiska _ tagalog _ polska
Information om Finland
Information om Finlandengelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ portugisiska
Information om Finlands historiaengelska _ ryska _ franska _ spanska _ tyska _ portugisiska
Länder som är anslutna till Apostilleavtaletengelska _ franska _ spanska _ tyska _ portugisiska
Rumänska
Flytta till Finland
linkkiEuropa.eu:
EU-länderfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Rådgivning för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropa.eu:
Information för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
Arbete och entreprenörskap
linkkiEures-portalen:
information om arbetsplatser i Europafinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropass.eu:
Information om CVfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropass.eu:
CV-mallarfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropeiska arbetsmiljöbyrån:
Information om arbetarskyddfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Ta med dig dina arbetslöshetsförmånerfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Hälsa
linkkiEuropeiska kommissionen:
Europeiska sjukvårdskortetfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Anvisning för identifiering av bröstcancer(pdf, 440kt)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ kinesiska _ thai _ rumänska _ samiska
Hjälp till offer för människohandelfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska _ polska _ rumänska _ bulgariska
På den här sidan har vi samlat länkar till andra webbplatser på språk som inte finns bland InfoFinlands urval av språk.
InfoFinland är en webbtjänst på 12 språk där alla språkversioner är identiska.
Du hittar urvalet av språk i tjänsten i menyn uppe på sidan.
Tyska
Thai
Kurdiska
Polska
Portugisiska
Rumänska
Tyska
Flytta till Finland
linkkiEuropa.eu:
EU-länderfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Rådgivning för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropa.eu:
Information för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
Arbete och entreprenörskap
linkkiArbetshälsoinstitutet:
Handboken Jobba i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ kurdiska _ tyska _ thai _ vietnamesiska
linkkiEuropass.eu:
Information om CVfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropass.eu:
CV-mallarfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiWebbtjänsten Suomi.fi:
Arbetsavtalsmallar på olika språkfinska _ svenska _ engelska _ ryska _ estniska _ franska _ tyska
linkkiEuropeiska unionen:
Information om att arbeta och driva ett företag i den europeiska unionenfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEures-portalen:
information om arbetsplatser i Europafinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropeiska arbetsmiljöbyrån:
Information om arbetarskyddfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Ta med dig dina arbetslöshetsförmånerfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Finska och svenska språket
linkkiEuropass.eu:
Utvärdera nivån på din språkkunskapfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Nybörjarkurs i finska, Tavataan taasengelska _ franska _ tyska _ bulgariska
linkkiWordDive:
Nybörjarkurs i finskafinska _ svenska _ engelska _ ryska _ kinesiska _ tyska
Webbkurs med många hjälpspråksvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ portugisiska
linkkiWordDive:
Finskans grammatikfinska _ svenska _ engelska _ ryska _ spanska _ tyska _ japanska
Boende
Heminkvarteringengelska _ franska _ spanska _ kinesiska _ tyska _ portugisiska _ italienska
Utbildning
linkkiUtbildningsstyrelsen:
Eget språk, eget sinnefinska _ engelska _ ryska _ estniska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ burmesiska _ bosniska
linkkiStudentexamensnämnden:
Information om studentexamenfinska _ svenska _ engelska _ franska _ tyska
Hälsa
linkkiNödcentralsverket:
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
linkkiEuropeiska kommissionen:
Europeiska sjukvårdskortetfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Privat psykoterapitjänst på Internetfinska _ svenska _ engelska _ ryska _ franska _ spanska _ turkiska _ kinesiska _ tyska _ portugisiska _ norska
_ holländska _ japanska _ italienska
_ danska
Hjälp till diskrimineringsofferfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ thai _ vietnamesiska _ portugisiska _ tagalog _ polska
linkkiBrottsofferjouren:
Hjälp för brottsofferfinska _ svenska _ engelska
linkkiBortförda barn rf:
Stöd och information för offer för barnkidnappningfinska _ svenska _ engelska _ turkiska _ arabiska _ tyska _ italienska
_ danska
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Information om Finland
Information om Finlandengelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ portugisiska
linkkiVisitFinland.com:
Information om Finland till turistersvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ japanska _ italienska
Information om finländska sederengelska _ spanska _ kinesiska _ tyska _ portugisiska
Information om Finlands historiaengelska _ ryska _ franska _ spanska _ tyska _ portugisiska
linkkiSkype:
Förmånliga utlandssamtalfinska _ svenska _ engelska _ ryska _ estniska _ franska _ spanska _ turkiska _ kinesiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ ungerska _ japanska
Länder som är anslutna till Apostilleavtaletengelska _ franska _ spanska _ tyska _ portugisiska
Thai
Arbete och entreprenörskap
linkkiArbetshälsoinstitutet:
Handboken Jobba i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ kurdiska _ tyska _ thai _ vietnamesiska
Guide för arbets- och näringsbyråns invandrarkunder(pdf, 5,1 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska _ kurdiska _ thai _ vietnamesiska
linkkiTE-tjänster:
Videoklipp och broschyrer för invandrarefinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska
Utbildning
linkkiKervo stad:
Så här använder du Wilma(pdf, 239 kt)finska _ engelska _ ryska _ estniska _ turkiska _ kurdiska _ thai _ vietnamesiska
Hälsä
linkkiStödcentralen Hilma för handikappade invandrare:
Serviceguide för handikappade invandrare(pdf, 797,26)finska _ svenska _ engelska _ ryska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ thai _ burmesiska
linkkiHivpoint:
Broschyren Information om sexuellt överförda sjukdomar(pdf, 1500kt)finska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Rådgivning för personer som säljer sexuella tjänsterfinska _ engelska
Anvisning för identifiering av bröstcancer(pdf, 440kt)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ kinesiska _ thai _ rumänska _ samiska
Familij
Handbok för familjer med två kulturer (pdf, 4,74 Mt)finska _ engelska _ ryska _ franska _ spanska _ thai
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Hjälp till diskrimineringsofferfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ thai _ vietnamesiska _ portugisiska _ tagalog _ polska
linkkiBrottsofferjouren:
Hjälp för brottsofferfinska _ svenska _ engelska
Hjälp till offer för människohandelfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska _ polska _ rumänska _ bulgariska
Fritid
linkkiFinlands Simundervisnings- och Livräddningsförbund rf:
Kom till simhallen!(pdf, 2 MB)finska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ arabiska _ kurdiska _ thai
Medborgarinstitut i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Information om Finland
linkkiArbets- och näringsministeriet:
Guiden Välkommen till Finland(pdf, 3,40 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
Kurdiska
Flytta till Finland
Information för flyktingarfinska _ engelska _ franska _ persiska _ arabiska _ kurdiska
Broschyren Information till asylsökandefinska _ svenska _ engelska _ ryska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
Arbete och entreprenörskap
linkkiArbetshälsoinstitutet:
Handboken Jobba i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ kurdiska _ tyska _ thai _ vietnamesiska
Guiden Bli företagare i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ turkiska _ kinesiska _ arabiska _ kurdiska
Guide om att grunda ett företagfinska _ engelska _ kinesiska
Guide för arbets- och näringsbyråns invandrarkunder(pdf, 5,1 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska _ kurdiska _ thai _ vietnamesiska
linkkiTE-tjänster:
Videoklipp och broschyrer för invandrarefinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska
linkkiKervo stad:
Så här använder du Wilma(pdf, 239 kt)finska _ engelska _ ryska _ estniska _ turkiska _ kurdiska _ thai _ vietnamesiska
linkki4V:
Tips för boende(pdf, 1,5 Mt)finska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Utbildning
linkkiKervo stad:
Så här använder du Wilma(pdf, 239 kt)finska _ engelska _ ryska _ estniska _ turkiska _ kurdiska _ thai _ vietnamesiska
Hälsä
linkkiNödcentralsverket:
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
linkkiStödcentralen Hilma för funktionshindrade invandrare :
Handbok med ordlista i hälso- och sjukvård på finska(pdf, 341,02 kt)finska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska
linkkiFöreningen för Mental Hälsa i Finland:
Information om mental hälsafinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
linkkiTuberkuloosi.fi:
Information om tuberkulosfinska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
linkkiStödcentralen Hilma för handikappade invandrare:
Stöd och hjälp för handikappade invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ persiska _ arabiska _ kurdiska
linkkiStödcentralen Hilma för handikappade invandrare:
Serviceguide för handikappade invandrare(pdf, 797,26)finska _ svenska _ engelska _ ryska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ thai _ burmesiska
linkkiSäg nej till droger -projektet:
Information om droger och faror som anknyter till dem särskilt för ungafinska _ somaliska _ arabiska _ kurdiska _ albanska
Familij
Uppfostring av barn i Finland(pdf, 8,08 Mt)finska _ engelska _ ryska _ somaliska _ kurdiska _ albanska _ burmesiska
Information om barnskyddslagenfinska _ svenska _ engelska _ ryska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
linkkiUtbildningsstyrelsen:
Eget språk, eget sinnefinska _ engelska _ ryska _ estniska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ burmesiska _ bosniska
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Hjälp till diskrimineringsofferfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ thai _ vietnamesiska _ portugisiska _ tagalog _ polska
Depression(pdf, 110,37 kt)finska _ engelska _ ryska _ franska _ somaliska _ turkiska _ persiska _ arabiska _ kurdiska _ albanska _ vietnamesiska _ burmesiska _ bosniska _ serbiska _ swahili
Information om posttraumatiskt stressyndromfinska _ engelska _ ryska _ franska _ somaliska _ turkiska _ persiska _ arabiska _ kurdiska _ albanska _ vietnamesiska _ burmesiska _ bosniska _ serbiska _ swahili
linkkiBrottsofferjouren:
Hjälp för brottsofferfinska _ svenska _ engelska
linkkiAndra ämbetsverk:
Broschyr om besöksförbud(pdf, 418,92 kt)finska _ svenska _ engelska
Diskrimineringsombudsmannenfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ persiska _ arabiska _ kurdiska
Hjälp till offer för människohandelfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska _ polska _ rumänska _ bulgariska
Information om krissituationer och sorgfinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Fritid
linkkiFinlands Simundervisnings- och Livräddningsförbund rf:
Kom till simhallen!(pdf, 2 MB)finska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ arabiska _ kurdiska _ thai
Medborgarinstitut i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Polska
Flytta till Finland
linkkiEuropa.eu:
EU-länderfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Rådgivning för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropa.eu:
Information för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
Arbete och entreprenörskap
linkkiArbets- och näringsbyrån:
Broschyren Jobba i Finland(pdf, 5,51 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ polska
linkkiEures-portalen:
information om arbetsplatser i Europafinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropass.eu:
Information om CVfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropass.eu:
CV-mallarfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropeiska arbetsmiljöbyrån:
Information om arbetarskyddfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Ta med dig dina arbetslöshetsförmånerfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Finska och svenska språket
linkkiEuropass.eu:
Utvärdera nivån på din språkkunskapfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Hälsä
linkkiEuropeiska kommissionen:
Europeiska sjukvårdskortetfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Hjälp till diskrimineringsofferfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ thai _ vietnamesiska _ portugisiska _ tagalog _ polska
linkkiBrottsofferjouren:
Hjälp för brottsofferfinska _ svenska _ engelska
Hjälp till offer för människohandelfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska _ polska _ rumänska _ bulgariska
Portugisiska
Flytta till Finland
linkkiEuropa.eu:
EU-länderfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Rådgivning för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropa.eu:
Information för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
Arbete och entreprenörskap
linkkiEures-portalen:
information om arbetsplatser i Europafinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropass.eu:
Information om CVfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropass.eu:
CV-mallarfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropeiska arbetsmiljöbyrån:
Information om arbetarskyddfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Ta med dig dina arbetslöshetsförmånerfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Finska och svenska språket
linkkiEuropass.eu:
Utvärdera nivån på din språkkunskapfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Webbkurs med många hjälpspråksvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ portugisiska
Hälsä
linkkiEuropeiska kommissionen:
Europeiska sjukvårdskortetfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Privat psykoterapitjänst på Internetfinska _ svenska _ engelska _ ryska _ franska _ spanska _ turkiska _ kinesiska _ tyska _ portugisiska _ norska
_ holländska _ japanska _ italienska
_ danska
Hjälp till diskrimineringsofferfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ thai _ vietnamesiska _ portugisiska _ tagalog _ polska
Information om Finland
Information om Finlandengelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ portugisiska
Information om Finlands historiaengelska _ ryska _ franska _ spanska _ tyska _ portugisiska
Länder som är anslutna till Apostilleavtaletengelska _ franska _ spanska _ tyska _ portugisiska
Rumänska
Flytta till Finland
linkkiEuropa.eu:
EU-länderfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Rådgivning för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropa.eu:
Information för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
Arbete och entreprenörskap
linkkiEures-portalen:
information om arbetsplatser i Europafinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropass.eu:
Information om CVfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropass.eu:
CV-mallarfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropeiska arbetsmiljöbyrån:
Information om arbetarskyddfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Ta med dig dina arbetslöshetsförmånerfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Hälsa
linkkiEuropeiska kommissionen:
Europeiska sjukvårdskortetfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Anvisning för identifiering av bröstcancer(pdf, 440kt)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ kinesiska _ thai _ rumänska _ samiska
Hjälp till offer för människohandelfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska _ polska _ rumänska _ bulgariska
På den här sidan har vi samlat länkar till andra webbplatser på språk som inte finns bland InfoFinlands urval av språk.
InfoFinland är en webbtjänst på 12 språk där alla språkversioner är identiska.
Du hittar urvalet av språk i tjänsten i menyn uppe på sidan.
Tyska
Thai
Kurdiska
Polska
Portugisiska
Rumänska
Tyska
Flytta till Finland
linkkiEuropa.eu:
EU-länderfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Rådgivning för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropa.eu:
Information för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
Arbete och entreprenörskap
linkkiArbetshälsoinstitutet:
Handboken Jobba i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ kurdiska _ tyska _ thai _ vietnamesiska
linkkiEuropass.eu:
Information om CVfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropass.eu:
CV-mallarfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiWebbtjänsten Suomi.fi:
Arbetsavtalsmallar på olika språkfinska _ svenska _ engelska _ ryska _ estniska _ franska _ tyska
linkkiEuropeiska unionen:
Information om att arbeta och driva ett företag i den europeiska unionenfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEures-portalen:
information om arbetsplatser i Europafinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropeiska arbetsmiljöbyrån:
Information om arbetarskyddfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Ta med dig dina arbetslöshetsförmånerfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Finska och svenska språket
linkkiEuropass.eu:
Utvärdera nivån på din språkkunskapfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Nybörjarkurs i finska, Tavataan taasengelska _ franska _ tyska _ bulgariska
linkkiWordDive:
Nybörjarkurs i finskafinska _ svenska _ engelska _ ryska _ kinesiska _ tyska
Webbkurs med många hjälpspråksvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ portugisiska
linkkiWordDive:
Finskans grammatikfinska _ svenska _ engelska _ ryska _ spanska _ tyska _ japanska
Boende
Heminkvarteringengelska _ franska _ spanska _ kinesiska _ tyska _ portugisiska _ italienska
Utbildning
linkkiUtbildningsstyrelsen:
Eget språk, eget sinnefinska _ engelska _ ryska _ estniska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ burmesiska _ bosniska
linkkiStudentexamensnämnden:
Information om studentexamenfinska _ svenska _ engelska _ franska _ tyska
Hälsa
linkkiNödcentralsverket:
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
linkkiEuropeiska kommissionen:
Europeiska sjukvårdskortetfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Privat psykoterapitjänst på Internetfinska _ svenska _ engelska _ ryska _ franska _ spanska _ turkiska _ kinesiska _ tyska _ portugisiska _ norska
_ holländska _ japanska _ italienska
_ danska
Hjälp till diskrimineringsofferfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ thai _ vietnamesiska _ portugisiska _ tagalog _ polska
linkkiBrottsofferjouren:
Hjälp för brottsofferfinska _ svenska _ engelska
linkkiBortförda barn rf:
Stöd och information för offer för barnkidnappningfinska _ svenska _ engelska _ turkiska _ arabiska _ tyska _ italienska
_ danska
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Information om Finland
Information om Finlandengelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ portugisiska
linkkiVisitFinland.com:
Information om Finland till turistersvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ japanska _ italienska
Information om finländska sederengelska _ spanska _ kinesiska _ tyska _ portugisiska
Information om Finlands historiaengelska _ ryska _ franska _ spanska _ tyska _ portugisiska
linkkiSkype:
Förmånliga utlandssamtalfinska _ svenska _ engelska _ ryska _ estniska _ franska _ spanska _ turkiska _ kinesiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ japanska _ italienska
_ danska
_ bulgariska
_ grekiska
_ tjeckiska
Länder som är anslutna till Apostilleavtaletengelska _ franska _ spanska _ tyska _ portugisiska
Thai
Arbete och entreprenörskap
linkkiArbetshälsoinstitutet:
Handboken Jobba i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ kurdiska _ tyska _ thai _ vietnamesiska
Guide för arbets- och näringsbyråns invandrarkunder(pdf, 5,1 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska _ kurdiska _ thai _ vietnamesiska
linkkiTE-tjänster:
Videoklipp och broschyrer för invandrarefinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska
Utbildning
linkkiKervo stad:
Så här använder du Wilma(pdf, 239 kt)finska _ engelska _ ryska _ estniska _ turkiska _ kurdiska _ thai _ vietnamesiska
Hälsä
linkkiStödcentralen Hilma för handikappade invandrare:
Serviceguide för handikappade invandrare(pdf, 797,26)finska _ engelska _ ryska _ arabiska
linkkiHivpoint:
Broschyren Information om sexuellt överförda sjukdomar(pdf, 1500kt)finska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Rådgivning för personer som säljer sexuella tjänsterfinska _ engelska
Anvisning för identifiering av bröstcancer(pdf, 440kt)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ kinesiska _ thai _ rumänska _ samiska
Familij
Handbok för familjer med två kulturer (pdf, 4,74 Mt)finska _ engelska _ ryska _ franska _ spanska _ thai
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Hjälp till diskrimineringsofferfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ thai _ vietnamesiska _ portugisiska _ tagalog _ polska
linkkiBrottsofferjouren:
Hjälp för brottsofferfinska _ svenska _ engelska
Hjälp till offer för människohandelfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska _ polska _ rumänska _ bulgariska
Fritid
linkkiFinlands Simundervisnings- och Livräddningsförbund rf:
Kom till simhallen!(pdf, 2 MB)finska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ arabiska _ kurdiska _ thai
Medborgarinstitut i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Information om Finland
linkkiArbets- och näringsministeriet:
Guiden Välkommen till Finland(pdf, 3,40 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
Kurdiska
Flytta till Finland
Information för flyktingarfinska _ engelska _ franska _ persiska _ arabiska _ kurdiska
Broschyren Information till asylsökandefinska _ svenska _ engelska _ ryska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
Arbete och entreprenörskap
linkkiArbetshälsoinstitutet:
Handboken Jobba i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ kurdiska _ tyska _ thai _ vietnamesiska
Guiden Bli företagare i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ turkiska _ kinesiska _ arabiska _ kurdiska
Guide om att grunda ett företagfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ turkiska _ kinesiska _ arabiska
Guide för arbets- och näringsbyråns invandrarkunder(pdf, 5,1 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska _ kurdiska _ thai _ vietnamesiska
linkkiTE-tjänster:
Videoklipp och broschyrer för invandrarefinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska
linkkiKervo stad:
Så här använder du Wilma(pdf, 239 kt)finska _ engelska _ ryska _ estniska _ turkiska _ kurdiska _ thai _ vietnamesiska
linkki4V:
Tips för boende(pdf, 1,5 Mt)finska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Utbildning
linkkiKervo stad:
Så här använder du Wilma(pdf, 239 kt)finska _ engelska _ ryska _ estniska _ turkiska _ kurdiska _ thai _ vietnamesiska
Hälsä
linkkiNödcentralsverket:
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
linkkiStödcentralen Hilma för funktionshindrade invandrare :
Handbok med ordlista i hälso- och sjukvård på finska(pdf, 341,02 kt)finska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska
linkkiFöreningen för Mental Hälsa i Finland:
Information om mental hälsafinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
linkkiTuberkuloosi.fi:
Information om tuberkulosfinska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska _ portugisiska _ tagalog _ polska _ bosniska _ rumänska _ swahili
_ lettiska
_ litauiska
linkkiStödcentralen Hilma för handikappade invandrare:
Stöd och hjälp för handikappade invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ persiska _ arabiska _ kurdiska
linkkiStödcentralen Hilma för handikappade invandrare:
Serviceguide för handikappade invandrare(pdf, 797,26)finska _ engelska _ ryska _ arabiska
linkkiSäg nej till droger -projektet:
Information om droger och faror som anknyter till dem särskilt för ungafinska _ somaliska _ arabiska _ kurdiska _ albanska
Familij
Uppfostring av barn i Finland(pdf, 8,08 Mt)finska _ engelska _ ryska _ somaliska _ kurdiska _ albanska _ burmesiska
Information om barnskyddslagenfinska _ svenska _ engelska _ ryska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
linkkiUtbildningsstyrelsen:
Eget språk, eget sinnefinska _ engelska _ ryska _ estniska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ burmesiska _ bosniska
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Hjälp till diskrimineringsofferfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ thai _ vietnamesiska _ portugisiska _ tagalog _ polska
Depression(pdf, 110,37 kt)finska _ engelska _ ryska _ franska _ somaliska _ turkiska _ persiska _ arabiska _ kurdiska _ albanska _ vietnamesiska _ burmesiska _ bosniska _ serbiska _ swahili
Information om posttraumatiskt stressyndromfinska _ engelska _ ryska _ franska _ somaliska _ turkiska _ persiska _ arabiska _ kurdiska _ albanska _ vietnamesiska _ burmesiska _ bosniska _ serbiska _ swahili
linkkiBrottsofferjouren:
Hjälp för brottsofferfinska _ svenska _ engelska
linkkiAndra ämbetsverk:
Broschyr om besöksförbud(pdf, 418,92 kt)finska _ svenska _ engelska
Diskrimineringsombudsmannenfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ persiska _ arabiska _ kurdiska
Hjälp till offer för människohandelfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska _ polska _ rumänska _ bulgariska
Information om krissituationer och sorgfinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Fritid
linkkiFinlands Simundervisnings- och Livräddningsförbund rf:
Kom till simhallen!(pdf, 2 MB)finska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ arabiska _ kurdiska _ thai
Medborgarinstitut i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Polska
Flytta till Finland
linkkiEuropa.eu:
EU-länderfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Rådgivning för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropa.eu:
Information för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
Arbete och entreprenörskap
linkkiArbets- och näringsbyrån:
Broschyren Jobba i Finland(pdf, 5,51 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ polska
linkkiEures-portalen:
information om arbetsplatser i Europafinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropass.eu:
Information om CVfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropass.eu:
CV-mallarfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropeiska arbetsmiljöbyrån:
Information om arbetarskyddfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Ta med dig dina arbetslöshetsförmånerfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Finska och svenska språket
linkkiEuropass.eu:
Utvärdera nivån på din språkkunskapfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Hälsä
linkkiEuropeiska kommissionen:
Europeiska sjukvårdskortetfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Hjälp till diskrimineringsofferfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ thai _ vietnamesiska _ portugisiska _ tagalog _ polska
linkkiBrottsofferjouren:
Hjälp för brottsofferfinska _ svenska _ engelska
Hjälp till offer för människohandelfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska _ polska _ rumänska _ bulgariska
Portugisiska
Flytta till Finland
linkkiEuropa.eu:
EU-länderfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Rådgivning för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropa.eu:
Information för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
Arbete och entreprenörskap
linkkiEures-portalen:
information om arbetsplatser i Europafinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropass.eu:
Information om CVfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropass.eu:
CV-mallarfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropeiska arbetsmiljöbyrån:
Information om arbetarskyddfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Ta med dig dina arbetslöshetsförmånerfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Finska och svenska språket
linkkiEuropass.eu:
Utvärdera nivån på din språkkunskapfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Webbkurs med många hjälpspråksvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ portugisiska
Hälsä
linkkiEuropeiska kommissionen:
Europeiska sjukvårdskortetfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Privat psykoterapitjänst på Internetfinska _ svenska _ engelska _ ryska _ franska _ spanska _ turkiska _ kinesiska _ tyska _ portugisiska _ norska
_ holländska _ japanska _ italienska
_ danska
Hjälp till diskrimineringsofferfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ thai _ vietnamesiska _ portugisiska _ tagalog _ polska
Information om Finland
Information om Finlandengelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ portugisiska
Information om Finlands historiaengelska _ ryska _ franska _ spanska _ tyska _ portugisiska
Länder som är anslutna till Apostilleavtaletengelska _ franska _ spanska _ tyska _ portugisiska
Rumänska
Flytta till Finland
linkkiEuropa.eu:
EU-länderfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Rådgivning för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropa.eu:
Information för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
Arbete och entreprenörskap
linkkiEures-portalen:
information om arbetsplatser i Europafinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropass.eu:
Information om CVfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropass.eu:
CV-mallarfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropeiska arbetsmiljöbyrån:
Information om arbetarskyddfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Ta med dig dina arbetslöshetsförmånerfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Hälsa
linkkiEuropeiska kommissionen:
Europeiska sjukvårdskortetfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Anvisning för identifiering av bröstcancer(pdf, 440kt)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ kinesiska _ thai _ rumänska _ samiska
Hjälp till offer för människohandelfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska _ polska _ rumänska _ bulgariska
I Finland har många helgdagar rötterna i kristendomen.
En del av helgdagarna, till exempel jul och påsk, är allmänna lediga dagar.
Då är också många butiker och ämbetsverk stängda.
Ett sätt att fira en helgdag är att hissa flaggan.
I Finland flaggar man på bestämda dagar som är intagna i kalendern.
Både myndigheter och vanliga människor deltar i flaggdagarna.
I Finland är flaggan något högtidligt.
På den här sidan finns kortfattad information om några finländska helgdagar.
Om flaggdagarna hittar du mer information på webbplatsen för Helsingfors universitets almanacksbyrå.
Om kristna fester kan du läsa mer på webbplatsen för evangelisk-lutherska kyrkan i Finland.
linkkiUniversitetets almanacksbyrå:
Högtidsdagarna i den finska kalendernfinska _ svenska _ engelska
linkkiEvangelisk-lutherska kyrkan i Finland:
Nyår
Nyårsaftonen den 31 december är årets sista dag.
Då ordnas fyrverkerier.
Fyrverkeripjäser kan köpas i affären.
För fyrverkerierna har man satt exakta tidsgränser.
Trettondagen
Trettondagen den 6 januari är julens sista dag.
Då minns man de tre vise männen som kom med gåvor till Jesusbarnet.
Runebergsdagen
Johan Ludvig Runeberg (1804–1877) är en viktig finländsk skald.
På Runebergsdagen den 5 februari äter man Runebergstårtor.
Vändagen
På vändagen den 14 februari kan man minnas sina vänner till exempel med blommor eller ett kort.
I Finland firas vändagen inte med lika mycket pompa och ståt som till exempel i USA.
Fastlagen
Fastlagen inleder förberedelserna för påsken.
På fastlagen åker man i Finland backe och äter fastlagsbullar som har bland annat grädde som fyllning.
Påsk
Påsken är en kristen fest.
Tidpunkten varierar men oftast firas påsk i mars eller april.
Före påsken firas palmsöndagen.
Då klär barn sig ut till häxor och går runt i grannskapet för att dela ut videkvistar som de dekorerat.
Barnen får oftast en liten present, till exempel lite godis.
På långfredagen minns man Jesu död.
Söndagen är påskdagen och då minns man Jesu uppståndelse.
Påskfirandet fortsätter ännu på måndagen som är annandag påsk.
På påsken äter man ofta lamm, chokladägg och memma.
Kristi himmelsfärdsdag
Kristi himmelsfärdsdag har sina rötter i kristendomen.
Då minns man Jesu himmelsfärd.
Valborgsmässoafton och första maj
Första maj är vårens och arbetarnas fest.
I Finland firas Valborgsmässoafton och första maj på många olika sätt.
Människorna samlas på picknick.
På första maj äter man munkar och dricker mjöd, som liknar läsk.
Många firar också med mousserande vin.
Studenterna tar på sig sina vita studentmössor.
Arbetarna ordnar Valborgsmarscher.
Morsdag
I Finland firas morsdag den andra söndagen i maj.
Mammorna firas till exempel med presenter och blommor.
Midsommar
Midsommar firas i slutet av juni.
Midsommar är en högtid som firas nära sommarsolståndet.
Många finländare åker gärna till stugan på midsommaren.
Stora midsommareldar hör till de finländska midsommartraditionerna.
I södra Finland reser man ibland också midsommarstången.
Alla helgons dag
Alla helgons dag firas i början av november.
Då minns man sina avlidna.
Människorna tänder ljus på sina anhörigas gravar.
Samtidigt firas också Halloween.
Alla helgons dag är emellertid inte en karneval som Halloween, utan en högtidlig och stilla fest.
Farsdag
Farsdag firas i Finland den andra söndagen i november.
Självständighetsdagen
Finland blev självständigt 1917.
Det firas på självständighetsdagen den 6 december.
Då tittar många finländare på självständighetsdagens mottagning med presidenten som värd på TV.
Julen
Julen är den viktigaste kristna festen i Finland.
Då minns man Jesu födelse.
Den egentliga dagen för firandet är julafton den 24 december.
Många skaffar sig en julgran som pyntas.
Julklapparna delas oftast ut på julafton.
Till den finländska julen hör många slags festmat, såsom julskinka, rosoll som är en rödbetssallad, olika slags lådor, julstjärnor och pepparkakor.
På julen sjunger man julsånger och umgås med familjen och andra nära och kära.
I Finland har många helgdagar rötterna i kristendomen.
En del av helgdagarna, till exempel jul och påsk, är allmänna lediga dagar.
Då är också många butiker och ämbetsverk stängda.
Ett sätt att fira en helgdag är att hissa flaggan.
I Finland flaggar man på bestämda dagar som är intagna i kalendern.
Både myndigheter och vanliga människor deltar i flaggdagarna.
I Finland är flaggan något högtidligt.
På den här sidan finns kortfattad information om några finländska helgdagar.
Om flaggdagarna hittar du mer information på webbplatsen för Helsingfors universitets almanacksbyrå.
Om kristna fester kan du läsa mer på webbplatsen för evangelisk-lutherska kyrkan i Finland.
linkkiUniversitetets almanacksbyrå:
Högtidsdagarna i den finska kalendernfinska _ svenska _ engelska
linkkiEvangelisk-lutherska kyrkan i Finland:
Nyår
Nyårsaftonen den 31 december är årets sista dag.
Då ordnas fyrverkerier.
Fyrverkeripjäser kan köpas i affären.
För fyrverkerierna har man satt exakta tidsgränser.
Trettondagen
Trettondagen den 6 januari är julens sista dag.
Då minns man de tre vise männen som kom med gåvor till Jesusbarnet.
Runebergsdagen
Johan Ludvig Runeberg (1804–1877) är en viktig finländsk skald.
På Runebergsdagen den 5 februari äter man Runebergstårtor.
Vändagen
På vändagen den 14 februari kan man minnas sina vänner till exempel med blommor eller ett kort.
I Finland firas vändagen inte med lika mycket pompa och ståt som till exempel i USA.
Fastlagen
Fastlagen inleder förberedelserna för påsken.
På fastlagen åker man i Finland backe och äter fastlagsbullar som har bland annat grädde som fyllning.
Påsk
Påsken är en kristen fest.
Tidpunkten varierar men oftast firas påsk i mars eller april.
Före påsken firas palmsöndagen.
Då klär barn sig ut till häxor och går runt i grannskapet för att dela ut videkvistar som de dekorerat.
Barnen får oftast en liten present, till exempel lite godis.
På långfredagen minns man Jesu död.
Söndagen är påskdagen och då minns man Jesu uppståndelse.
Påskfirandet fortsätter ännu på måndagen som är annandag påsk.
På påsken äter man ofta lamm, chokladägg och memma.
Kristi himmelsfärdsdag
Kristi himmelsfärdsdag har sina rötter i kristendomen.
Då minns man Jesu himmelsfärd.
Valborgsmässoafton och första maj
Första maj är vårens och arbetarnas fest.
I Finland firas Valborgsmässoafton och första maj på många olika sätt.
Människorna samlas på picknick.
På första maj äter man munkar och dricker mjöd, som liknar läsk.
Många firar också med mousserande vin.
Studenterna tar på sig sina vita studentmössor.
Arbetarna ordnar Valborgsmarscher.
Morsdag
I Finland firas morsdag den andra söndagen i maj.
Mammorna firas till exempel med presenter och blommor.
Midsommar
Midsommar firas i slutet av juni.
Midsommar är en högtid som firas nära sommarsolståndet.
Många finländare åker gärna till stugan på midsommaren.
Stora midsommareldar hör till de finländska midsommartraditionerna.
I södra Finland reser man ibland också midsommarstången.
Alla helgons dag
Alla helgons dag firas i början av november.
Då minns man sina avlidna.
Människorna tänder ljus på sina anhörigas gravar.
Samtidigt firas också Halloween.
Alla helgons dag är emellertid inte en karneval som Halloween, utan en högtidlig och stilla fest.
Farsdag
Farsdag firas i Finland den andra söndagen i november.
Självständighetsdagen
Finland blev självständigt 1917.
Det firas på självständighetsdagen den 6 december.
Då tittar många finländare på självständighetsdagens mottagning med presidenten som värd på TV.
Julen
Julen är den viktigaste kristna festen i Finland.
Då minns man Jesu födelse.
Den egentliga dagen för firandet är julafton den 24 december.
Många skaffar sig en julgran som pyntas.
Julklapparna delas oftast ut på julafton.
Till den finländska julen hör många slags festmat, såsom julskinka, rosoll som är en rödbetssallad, olika slags lådor, julstjärnor och pepparkakor.
På julen sjunger man julsånger och umgås med familjen och andra nära och kära.
I Finland har många helgdagar rötterna i kristendomen.
En del av helgdagarna, till exempel jul och påsk, är allmänna lediga dagar.
Då är också många butiker och ämbetsverk stängda.
Ett sätt att fira en helgdag är att hissa flaggan.
I Finland flaggar man på bestämda dagar som är intagna i kalendern.
Både myndigheter och vanliga människor deltar i flaggdagarna.
I Finland är flaggan något högtidligt.
På den här sidan finns kortfattad information om några finländska helgdagar.
Om flaggdagarna hittar du mer information på webbplatsen för Helsingfors universitets almanacksbyrå.
Om kristna fester kan du läsa mer på webbplatsen för evangelisk-lutherska kyrkan i Finland.
linkkiUniversitetets almanacksbyrå:
Högtidsdagarna i den finska kalendernfinska _ svenska _ engelska
linkkiEvangelisk-lutherska kyrkan i Finland:
Nyår
Nyårsaftonen den 31 december är årets sista dag.
Då ordnas fyrverkerier.
Fyrverkeripjäser kan köpas i affären.
För fyrverkerierna har man satt exakta tidsgränser.
Trettondagen
Trettondagen den 6 januari är julens sista dag.
Då minns man de tre vise männen som kom med gåvor till Jesusbarnet.
Runebergsdagen
Johan Ludvig Runeberg (1804–1877) är en viktig finländsk skald.
På Runebergsdagen den 5 februari äter man Runebergstårtor.
Vändagen
På vändagen den 14 februari kan man minnas sina vänner till exempel med blommor eller ett kort.
I Finland firas vändagen inte med lika mycket pompa och ståt som till exempel i USA.
Fastlagen
Fastlagen inleder förberedelserna för påsken.
På fastlagen åker man i Finland backe och äter fastlagsbullar som har bland annat grädde som fyllning.
Påsk
Påsken är en kristen fest.
Tidpunkten varierar men oftast firas påsk i mars eller april.
Före påsken firas palmsöndagen.
Då klär barn sig ut till häxor och går runt i grannskapet för att dela ut videkvistar som de dekorerat.
Barnen får oftast en liten present, till exempel lite godis.
På långfredagen minns man Jesu död.
Söndagen är påskdagen och då minns man Jesu uppståndelse.
Påskfirandet fortsätter ännu på måndagen som är annandag påsk.
På påsken äter man ofta lamm, chokladägg och memma.
Kristi himmelsfärdsdag
Kristi himmelsfärdsdag har sina rötter i kristendomen.
Då minns man Jesu himmelsfärd.
Valborgsmässoafton och första maj
Första maj är vårens och arbetarnas fest.
I Finland firas Valborgsmässoafton och första maj på många olika sätt.
Människorna samlas på picknick.
På första maj äter man munkar och dricker mjöd, som liknar läsk.
Många firar också med mousserande vin.
Studenterna tar på sig sina vita studentmössor.
Arbetarna ordnar Valborgsmarscher.
Morsdag
I Finland firas morsdag den andra söndagen i maj.
Mammorna firas till exempel med presenter och blommor.
Midsommar
Midsommar firas i slutet av juni.
Midsommar är en högtid som firas nära sommarsolståndet.
Många finländare åker gärna till stugan på midsommaren.
Stora midsommareldar hör till de finländska midsommartraditionerna.
I södra Finland reser man ibland också midsommarstången.
Alla helgons dag
Alla helgons dag firas i början av november.
Då minns man sina avlidna.
Människorna tänder ljus på sina anhörigas gravar.
Samtidigt firas också Halloween.
Alla helgons dag är emellertid inte en karneval som Halloween, utan en högtidlig och stilla fest.
Farsdag
Farsdag firas i Finland den andra söndagen i november.
Självständighetsdagen
Finland blev självständigt 1917.
Det firas på självständighetsdagen den 6 december.
Då tittar många finländare på självständighetsdagens mottagning med presidenten som värd på TV.
Julen
Julen är den viktigaste kristna festen i Finland.
Då minns man Jesu födelse.
Den egentliga dagen för firandet är julafton den 24 december.
Många skaffar sig en julgran som pyntas.
Julklapparna delas oftast ut på julafton.
Till den finländska julen hör många slags festmat, såsom julskinka, rosoll som är en rödbetssallad, olika slags lådor, julstjärnor och pepparkakor.
På julen sjunger man julsånger och umgås med familjen och andra nära och kära.
På den här sidan finns allmän information om finländska seder.
Du hittar information om den finländska arbetskulturen på InfoFinlands sida Den finländska arbetskulturen.
Den finländska värdegrunden
Jämlikhet och rättvisa är värden som finländarna skattar högt.
I det finländska samhället är alla jämlika och alla ska behandlas rättvist.
Information om jämlikhet och likabehandling hittar du på InfoFinlands sida Jämställdhet och jämlikhet.
Jämställdhet
Enligt finsk lag är kvinnor och män jämställda.
I Finland är det vanligt att kvinnor arbetar, även om de har barn.
Mannen och kvinnan ansvarar båda för att ta hand om barnen och hemmet.
Tillit
Det är vanligt att finländarna litar på andra människor och på myndigheter.
I Finland värdesätts också demokrati och yttrandefrihet.
Varje människa har rätt att delta i samhällslivet.
I Finland råder också yttrandefrihet.
I den finländska kulturen framhävs individualism mer än i många andra kulturer.
Individens frihet syns starkt i den finländska lagstiftningen.
Eget utrymme
Finländarna värdesätter också sin integritet och privatsfär.
Till exempel uppmuntras unga vuxna att bli självständiga och flytta hemifrån.
Ärlighet och punktlighet
I Finland värdesätts ärlighet.
Det är viktigt att hålla sina löften och tala sanning.
Också punktlighet är viktigt för finländarna.
När du har ett möte ska du komma i tid.
Om du till exempel har bokat tid hos en myndighet eller läkaren är det speciellt viktigt att du är på plats i tid.
Om du till exempel har en tid klockan tolv, var på plats strax före tolv.
Om du kommer klockan 12.10 är du försenad.
Anspråkslöshet
Många finländare uppskattar anspråkslöshet.
Människor framhäver sig inte i gruppen; de talar inte högljutt och skryter inte.
I Finland anses det vara välartat att ta hänsyn till och lyssna på andra.
Också arbetsamhet och flit värdesätts högt.
Naturen
Naturen är mycket viktig för finländarna.
Många finländare trivs i naturen, till exempel vandrar eller plockar bär.
I Finland gäller allemansrätten (jokamiehenoikeus).
Enligt allemansrätten får alla röra sig fritt i naturen utan att behöva be om markägarens tillstånd till allt.
Läs mer om allemansrätten på InfoFinlands sida Att röra sig i naturen.
Att hälsa
Att skaka hand är ett vanligt sätt att hälsa på människor i officiella situationer.
Också män och kvinnor skakar hand med varandra.
Nära vänner eller släktingar kan även hälsa på varandra genom att krama om varandra.
Kindpussar är dock ovanliga.
När du pratar med någon, ta ögonkontakt med personen du pratar med.
I Finland uppfattas ögonkontakt som uppriktighet och ärlighet gentemot den andra.
På finska duar man oftast.
Man duar också folk man inte känner, likaså sina kollegor.
Niande hör hemma endast i mycket formella situationer.
Det är också bra att nia äldre människor.
Samtal och växelverkan
Finländare går gärna rakt på sak i samtal.
Det finländska sättet att kommunicera är rakt och okomplicerat.
I Finland förväntar människorna sig att man verkligen menar det man säger.
Det du säger tas på allvar och andra förväntar sig att du står bakom dina ord.
När finländare samtalar, kan det ibland uppstå tysta stunder.
Tystnaden är inte negativ utan upplevs som något naturligt.
De tysta stunderna behöver inte fyllas med prat.
Högljutt prat kan anses vara obekvämt eller hotfullt.
I Finland är det oartigt att avbryta andra när de talar.
Finländare väntar vanligtvis att samtalspartnern har sagt sitt innan de själva tar till ordet.
I Finland är det inte vanligt att visa sina känslor offentligt.
När man talar är det oartigt att höja rösten, speciellt på allmänna platser.
Finländare äter relativt typisk europeisk mat som ofta innehåller kött, fisk, potatis, ris eller pasta.
Vegetarism har blivit allt populärare.
Det är vanligt att man äter två varma måltider om dagen, lunch och middag.
I Finland dricker också vuxna ofta mjölk.
I Finland äter man lunch tidigare än i många andra länder.
På arbetsplatser och i skolor serveras lunch vanligtvis kl. 11–12.
Middag äts ofta vid femtiden på eftermiddagen.
I Finland betonas ofta att maten ska vara hälsosam.
Bland annat rågbröd och olika gröträtter är en viktig del av den finländska matkulturen.
Olika regioner i Finland har olika matkulturer.
Till exempel i Lappland äts mycket renkött, medan man i kustregionerna äter fisk.
Till exempel syns italienska pastarätter och asiatiska matkulturer också i Finland.
Barn och unga serveras mat i daghem och skolor.
Skolmaten är gratis för alla och man behöver inte ta med sig en matsäck till skolan.
I Finland dricker man mycket kaffe.
Till exempel på fester serveras det nästan alltid kaffe.
På möten på arbetsplatsen dricker man ofta kaffe.
Alkoholdrycker är relativt dyra i Finland och köpet av dem begränsas med åldersgränser för unga personer.
I mataffären säljs endast milda alkoholdrycker.
Starka alkoholdrycker köper man i de statligt reglerade Alko-butikerna.
Att köra bil under alkoholpåverkan är förbjudet enligt lag och det kan ge ett hårt straff.
Att äta på restaurang är ofta dyrare i Finland än i andra länder.
Också alkoholdrycker är dyra på restaurang.
Du behöver inte lämna dricks, men du kan göra det om du vill tacka för en speciellt bra service.
linkkiVisitFinland.com:
Den finska matkulturenengelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ japanska _ italienska
Bastu
Bastun är en viktig del av den finländska kulturen.
Bastun är avsedd för att man ska göra sig ren och koppla av och därför förknippas den med tystnad och lugn.
Många finländare badar bastu varje vecka.
Man badar bastu med såväl familjemedlemmar och vänner som med affärspartner.
Män och kvinnor badar bastu olika tider.
Vanligtvis badar man bastu naken.
På bastulaven sitter man oftast på ett litet sittunderlag.
Som gäst i ett finländskt hem
I Finland ska man alltid på förhand komma överens om besök hos andra, även hos goda vänner.
Finländare lägger speciellt stort värde på sitt privatliv och sitt eget lugn.
Finländare använder inte skor inomhus.
Det är artigt att ta av sig skorna när du går in i någons hem.
När du besöker ett finländskt hem, ta av dig skorna eller fråga om du kan ha dem på.
Information om finländska sederengelska _ spanska _ kinesiska _ tyska _ portugisiska
På den här sidan finns allmän information om finländska seder.
Du hittar information om den finländska arbetskulturen på InfoFinlands sida Den finländska arbetskulturen.
Den finländska värdegrunden
Jämlikhet och rättvisa är värden som finländarna skattar högt.
I det finländska samhället är alla jämlika och alla ska behandlas rättvist.
Information om jämlikhet och likabehandling hittar du på InfoFinlands sida Jämställdhet och jämlikhet.
Jämställdhet
Enligt finsk lag är kvinnor och män jämställda.
I Finland är det vanligt att kvinnor arbetar, även om de har barn.
Mannen och kvinnan ansvarar båda för att ta hand om barnen och hemmet.
Tillit
Det är vanligt att finländarna litar på andra människor och på myndigheter.
I Finland värdesätts också demokrati och yttrandefrihet.
Varje människa har rätt att delta i samhällslivet.
I Finland råder också yttrandefrihet.
I den finländska kulturen framhävs individualism mer än i många andra kulturer.
Individens frihet syns starkt i den finländska lagstiftningen.
Eget utrymme
Finländarna värdesätter också sin integritet och privatsfär.
Till exempel uppmuntras unga vuxna att bli självständiga och flytta hemifrån.
Ärlighet och punktlighet
I Finland värdesätts ärlighet.
Det är viktigt att hålla sina löften och tala sanning.
Också punktlighet är viktigt för finländarna.
När du har ett möte ska du komma i tid.
Om du till exempel har bokat tid hos en myndighet eller läkaren är det speciellt viktigt att du är på plats i tid.
Om du till exempel har en tid klockan tolv, var på plats strax före tolv.
Om du kommer klockan 12.10 är du försenad.
Anspråkslöshet
Många finländare uppskattar anspråkslöshet.
Människor framhäver sig inte i gruppen; de talar inte högljutt och skryter inte.
I Finland anses det vara välartat att ta hänsyn till och lyssna på andra.
Också arbetsamhet och flit värdesätts högt.
Naturen
Naturen är mycket viktig för finländarna.
Många finländare trivs i naturen, till exempel vandrar eller plockar bär.
I Finland gäller allemansrätten (jokamiehenoikeus).
Enligt allemansrätten får alla röra sig fritt i naturen utan att behöva be om markägarens tillstånd till allt.
Läs mer om allemansrätten på InfoFinlands sida Att röra sig i naturen.
Att hälsa
Att skaka hand är ett vanligt sätt att hälsa på människor i officiella situationer.
Också män och kvinnor skakar hand med varandra.
Nära vänner eller släktingar kan även hälsa på varandra genom att krama om varandra.
Kindpussar är dock ovanliga.
När du pratar med någon, ta ögonkontakt med personen du pratar med.
I Finland uppfattas ögonkontakt som uppriktighet och ärlighet gentemot den andra.
På finska duar man oftast.
Man duar också folk man inte känner, likaså sina kollegor.
Niande hör hemma endast i mycket formella situationer.
Det är också bra att nia äldre människor.
Samtal och växelverkan
Finländare går gärna rakt på sak i samtal.
Det finländska sättet att kommunicera är rakt och okomplicerat.
I Finland förväntar människorna sig att man verkligen menar det man säger.
Det du säger tas på allvar och andra förväntar sig att du står bakom dina ord.
När finländare samtalar, kan det ibland uppstå tysta stunder.
Tystnaden är inte negativ utan upplevs som något naturligt.
De tysta stunderna behöver inte fyllas med prat.
Högljutt prat kan anses vara obekvämt eller hotfullt.
I Finland är det oartigt att avbryta andra när de talar.
Finländare väntar vanligtvis att samtalspartnern har sagt sitt innan de själva tar till ordet.
I Finland är det inte vanligt att visa sina känslor offentligt.
När man talar är det oartigt att höja rösten, speciellt på allmänna platser.
Finländare äter relativt typisk europeisk mat som ofta innehåller kött, fisk, potatis, ris eller pasta.
Vegetarism har blivit allt populärare.
Det är vanligt att man äter två varma måltider om dagen, lunch och middag.
I Finland dricker också vuxna ofta mjölk.
I Finland äter man lunch tidigare än i många andra länder.
På arbetsplatser och i skolor serveras lunch vanligtvis kl. 11–12.
Middag äts ofta vid femtiden på eftermiddagen.
I Finland betonas ofta att maten ska vara hälsosam.
Bland annat rågbröd och olika gröträtter är en viktig del av den finländska matkulturen.
Olika regioner i Finland har olika matkulturer.
Till exempel i Lappland äts mycket renkött, medan man i kustregionerna äter fisk.
Till exempel syns italienska pastarätter och asiatiska matkulturer också i Finland.
Barn och unga serveras mat i daghem och skolor.
Skolmaten är gratis för alla och man behöver inte ta med sig en matsäck till skolan.
I Finland dricker man mycket kaffe.
Till exempel på fester serveras det nästan alltid kaffe.
På möten på arbetsplatsen dricker man ofta kaffe.
Alkoholdrycker är relativt dyra i Finland och köpet av dem begränsas med åldersgränser för unga personer.
I mataffären säljs endast milda alkoholdrycker.
Starka alkoholdrycker köper man i de statligt reglerade Alko-butikerna.
Att köra bil under alkoholpåverkan är förbjudet enligt lag och det kan ge ett hårt straff.
Att äta på restaurang är ofta dyrare i Finland än i andra länder.
Också alkoholdrycker är dyra på restaurang.
Du behöver inte lämna dricks, men du kan göra det om du vill tacka för en speciellt bra service.
linkkiVisitFinland.com:
Den finska matkulturenengelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ japanska _ italienska
Bastu
Bastun är en viktig del av den finländska kulturen.
Bastun är avsedd för att man ska göra sig ren och koppla av och därför förknippas den med tystnad och lugn.
Många finländare badar bastu varje vecka.
Man badar bastu med såväl familjemedlemmar och vänner som med affärspartner.
Män och kvinnor badar bastu olika tider.
Vanligtvis badar man bastu naken.
På bastulaven sitter man oftast på ett litet sittunderlag.
Som gäst i ett finländskt hem
I Finland ska man alltid på förhand komma överens om besök hos andra, även hos goda vänner.
Finländare lägger speciellt stort värde på sitt privatliv och sitt eget lugn.
Finländare använder inte skor inomhus.
Det är artigt att ta av sig skorna när du går in i någons hem.
När du besöker ett finländskt hem, ta av dig skorna eller fråga om du kan ha dem på.
Information om finländska sederengelska _ spanska _ kinesiska _ tyska _ portugisiska
På den här sidan finns allmän information om finländska seder.
Du hittar information om den finländska arbetskulturen på InfoFinlands sida Den finländska arbetskulturen.
Den finländska värdegrunden
Jämlikhet och rättvisa är värden som finländarna skattar högt.
I det finländska samhället är alla jämlika och alla ska behandlas rättvist.
Information om jämlikhet och likabehandling hittar du på InfoFinlands sida Jämställdhet och jämlikhet.
Jämställdhet
Enligt finsk lag är kvinnor och män jämställda.
I Finland är det vanligt att kvinnor arbetar, även om de har barn.
Mannen och kvinnan ansvarar båda för att ta hand om barnen och hemmet.
Tillit
Det är vanligt att finländarna litar på andra människor och på myndigheter.
I Finland värdesätts också demokrati och yttrandefrihet.
Varje människa har rätt att delta i samhällslivet.
I Finland råder också yttrandefrihet.
I den finländska kulturen framhävs individualism mer än i många andra kulturer.
Individens frihet syns starkt i den finländska lagstiftningen.
Eget utrymme
Finländarna värdesätter också sin integritet och privatsfär.
Till exempel uppmuntras unga vuxna att bli självständiga och flytta hemifrån.
Ärlighet och punktlighet
I Finland värdesätts ärlighet.
Det är viktigt att hålla sina löften och tala sanning.
Också punktlighet är viktigt för finländarna.
När du har ett möte ska du komma i tid.
Om du till exempel har bokat tid hos en myndighet eller läkaren är det speciellt viktigt att du är på plats i tid.
Om du till exempel har en tid klockan tolv, var på plats strax före tolv.
Om du kommer klockan 12.10 är du försenad.
Anspråkslöshet
Många finländare uppskattar anspråkslöshet.
Människor framhäver sig inte i gruppen; de talar inte högljutt och skryter inte.
I Finland anses det vara välartat att ta hänsyn till och lyssna på andra.
Också arbetsamhet och flit värdesätts högt.
Naturen
Naturen är mycket viktig för finländarna.
Många finländare trivs i naturen, till exempel vandrar eller plockar bär.
I Finland gäller allemansrätten (jokamiehenoikeus).
Enligt allemansrätten får alla röra sig fritt i naturen utan att behöva be om markägarens tillstånd till allt.
Läs mer om allemansrätten på InfoFinlands sida Att röra sig i naturen.
Att hälsa
Att skaka hand är ett vanligt sätt att hälsa på människor i officiella situationer.
Också män och kvinnor skakar hand med varandra.
Nära vänner eller släktingar kan även hälsa på varandra genom att krama om varandra.
Kindpussar är dock ovanliga.
När du pratar med någon, ta ögonkontakt med personen du pratar med.
I Finland uppfattas ögonkontakt som uppriktighet och ärlighet gentemot den andra.
På finska duar man oftast.
Man duar också folk man inte känner, likaså sina kollegor.
Niande hör hemma endast i mycket formella situationer.
Det är också bra att nia äldre människor.
Samtal och växelverkan
Finländare går gärna rakt på sak i samtal.
Det finländska sättet att kommunicera är rakt och okomplicerat.
I Finland förväntar människorna sig att man verkligen menar det man säger.
Det du säger tas på allvar och andra förväntar sig att du står bakom dina ord.
När finländare samtalar, kan det ibland uppstå tysta stunder.
Tystnaden är inte negativ utan upplevs som något naturligt.
De tysta stunderna behöver inte fyllas med prat.
Högljutt prat kan anses vara obekvämt eller hotfullt.
I Finland är det oartigt att avbryta andra när de talar.
Finländare väntar vanligtvis att samtalspartnern har sagt sitt innan de själva tar till ordet.
I Finland är det inte vanligt att visa sina känslor offentligt.
När man talar är det oartigt att höja rösten, speciellt på allmänna platser.
Finländare äter relativt typisk europeisk mat som ofta innehåller kött, fisk, potatis, ris eller pasta.
Vegetarism har blivit allt populärare.
Det är vanligt att man äter två varma måltider om dagen, lunch och middag.
I Finland dricker också vuxna ofta mjölk.
I Finland äter man lunch tidigare än i många andra länder.
På arbetsplatser och i skolor serveras lunch vanligtvis kl. 11–12.
Middag äts ofta vid femtiden på eftermiddagen.
I Finland betonas ofta att maten ska vara hälsosam.
Bland annat rågbröd och olika gröträtter är en viktig del av den finländska matkulturen.
Olika regioner i Finland har olika matkulturer.
Till exempel i Lappland äts mycket renkött, medan man i kustregionerna äter fisk.
Till exempel syns italienska pastarätter och asiatiska matkulturer också i Finland.
Barn och unga serveras mat i daghem och skolor.
Skolmaten är gratis för alla och man behöver inte ta med sig en matsäck till skolan.
I Finland dricker man mycket kaffe.
Till exempel på fester serveras det nästan alltid kaffe.
På möten på arbetsplatsen dricker man ofta kaffe.
Alkoholdrycker är relativt dyra i Finland och köpet av dem begränsas med åldersgränser för unga personer.
I mataffären säljs endast milda alkoholdrycker.
Starka alkoholdrycker köper man i de statligt reglerade Alko-butikerna.
Att köra bil under alkoholpåverkan är förbjudet enligt lag och det kan ge ett hårt straff.
Att äta på restaurang är ofta dyrare i Finland än i andra länder.
Också alkoholdrycker är dyra på restaurang.
Du behöver inte lämna dricks, men du kan göra det om du vill tacka för en speciellt bra service.
linkkiVisitFinland.com:
Den finska matkulturenengelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ japanska _ italienska
Bastu
Bastun är en viktig del av den finländska kulturen.
Bastun är avsedd för att man ska göra sig ren och koppla av och därför förknippas den med tystnad och lugn.
Många finländare badar bastu varje vecka.
Man badar bastu med såväl familjemedlemmar och vänner som med affärspartner.
Män och kvinnor badar bastu olika tider.
Vanligtvis badar man bastu naken.
På bastulaven sitter man oftast på ett litet sittunderlag.
Som gäst i ett finländskt hem
I Finland ska man alltid på förhand komma överens om besök hos andra, även hos goda vänner.
Finländare lägger speciellt stort värde på sitt privatliv och sitt eget lugn.
Finländare använder inte skor inomhus.
Det är artigt att ta av sig skorna när du går in i någons hem.
När du besöker ett finländskt hem, ta av dig skorna eller fråga om du kan ha dem på.
Information om finländska sederengelska _ spanska _ kinesiska _ tyska _ portugisiska
Befolkningen i Finland
Finlands folkmängd är cirka 5,5 miljoner människor.
Finland är ett mycket glesbefolkat land.
Befolkningen är framför allt koncentrerad till de stora städerna och tätorterna.
I huvudstadsregionen bor över en miljon människor.
Finlands befolkningfinska _ svenska _ engelska
Finska och svenska är Finlands nationalspråk.
Strax under 4,9 miljoner människor har finska som modersmål, medan strax under 300 000 människor talar svenska.
De största språken efter finska och svenska är ryska, estniska, engelska, somaliska och arabiska.
Till befolkningen i Finland hör olika slags minoriteter som till exempel har ett annat modersmål, en annan kultur eller religion än majoriteten av finländarna.
Traditionella minoriteter i Finland är till exempel finlandssvenskarna, samerna, romerna, judarna och tatarerna.
Dessutom har Finland fått invandrare till exempel från Ryssland, Estland, länderna på Balkan, Somalia och Irak.
Religioner i Finland
De flesta finländarna är kristna.
Det största religiösa samfundet är evangelisk-lutherska kyrkan i Finland, där cirka 70 procent av befolkningen är medlemmar.
Ortodoxa kyrkan i Finland är landets näst största religiösa samfund.
Drygt en procent av befolkningen hör till den ortodoxa kyrkan.
Den evangelisk-lutherska och den ortodoxa kyrkan har en särställning i Finland.
De har till exempel rätt att uppbära skatt.
I Finland bor tiotusentals muslimer.
Av dem hör emellertid endast en del till de islamska samfunden.
I Finland bor även några tusen judar.
I Helsingfors och Åbo finns en synagoga.
Andra religiösa samfund i Finland är till exempel Katolska kyrkan i Finland, Pingstkyrkan i Finland, Frikyrkan i Finland, Adventkyrkan i Finland, mormonkyrkan och Jehovas vittnen.
linkkiUndervisnings- och kulturministeriet:
Religiösa samfundfinska _ svenska _ engelska
Religiösa samfundfinska _ engelska
Religionsfrihet och religionsutövande i Finland
I Finland råder religionsfrihet.
Alla som bor i Finland har rätt att själva välja sin religion och utöva den.
Om man inte vill, måste man inte välja någon religion alls.
Ingen kan heller mot sin vilja tvingas att delta i religionsutövande.
linkkiUndervisnings- och kulturministeriet:
Religionsfrihetfinska _ svenska _ engelska
Minst 20 myndiga personer kan grunda ett religiöst samfund.
Religiösa grupper måste inte registrera sig som samfund, utan de kan även verka utan att ha registrerat sig.
linkkiPatent- och registerstyrelsen:
Registrering av ett religiöst samfundfinska _ svenska _ engelska
Barnets religion
Föräldrarna bestämmer barnets religion.
Om föräldrarna inte är överens, kan modern fatta beslut om religionstillhörigheten för ett barn som inte har fyllt ett år.
Barnet har rätt att få undervisning i sin egen religion i skolan.
Läs mer på InfoFinlands sida Grundläggande utbildning.
En myndig person, alltså en person som har fyllt 18 år, får själv besluta om sin religion.
Befolkningen i Finland
Finlands folkmängd är cirka 5,5 miljoner människor.
Finland är ett mycket glesbefolkat land.
Befolkningen är framför allt koncentrerad till de stora städerna och tätorterna.
I huvudstadsregionen bor över en miljon människor.
Finlands befolkningfinska _ svenska _ engelska
Finska och svenska är Finlands nationalspråk.
Strax under 4,9 miljoner människor har finska som modersmål, medan strax under 300 000 människor talar svenska.
De största språken efter finska och svenska är ryska, estniska, engelska, somaliska och arabiska.
Till befolkningen i Finland hör olika slags minoriteter som till exempel har ett annat modersmål, en annan kultur eller religion än majoriteten av finländarna.
Traditionella minoriteter i Finland är till exempel finlandssvenskarna, samerna, romerna, judarna och tatarerna.
Dessutom har Finland fått invandrare till exempel från Ryssland, Estland, länderna på Balkan, Somalia och Irak.
Religioner i Finland
De flesta finländarna är kristna.
Det största religiösa samfundet är evangelisk-lutherska kyrkan i Finland, där cirka 70 procent av befolkningen är medlemmar.
Ortodoxa kyrkan i Finland är landets näst största religiösa samfund.
Drygt en procent av befolkningen hör till den ortodoxa kyrkan.
Den evangelisk-lutherska och den ortodoxa kyrkan har en särställning i Finland.
De har till exempel rätt att uppbära skatt.
I Finland bor tiotusentals muslimer.
Av dem hör emellertid endast en del till de islamska samfunden.
I Finland bor även några tusen judar.
I Helsingfors och Åbo finns en synagoga.
Andra religiösa samfund i Finland är till exempel Katolska kyrkan i Finland, Pingstkyrkan i Finland, Frikyrkan i Finland, Adventkyrkan i Finland, mormonkyrkan och Jehovas vittnen.
linkkiUndervisnings- och kulturministeriet:
Religiösa samfundfinska _ svenska _ engelska
Religiösa samfundfinska _ engelska
Religionsfrihet och religionsutövande i Finland
I Finland råder religionsfrihet.
Alla som bor i Finland har rätt att själva välja sin religion och utöva den.
Om man inte vill, måste man inte välja någon religion alls.
Ingen kan heller mot sin vilja tvingas att delta i religionsutövande.
linkkiUndervisnings- och kulturministeriet:
Religionsfrihetfinska _ svenska _ engelska
Minst 20 myndiga personer kan grunda ett religiöst samfund.
Religiösa grupper måste inte registrera sig som samfund, utan de kan även verka utan att ha registrerat sig.
linkkiPatent- och registerstyrelsen:
Registrering av ett religiöst samfundfinska _ svenska _ engelska
Barnets religion
Föräldrarna bestämmer barnets religion.
Om föräldrarna inte är överens, kan modern fatta beslut om religionstillhörigheten för ett barn som inte har fyllt ett år.
Barnet har rätt att få undervisning i sin egen religion i skolan.
Läs mer på InfoFinlands sida Grundläggande utbildning.
En myndig person, alltså en person som har fyllt 18 år, får själv besluta om sin religion.
Befolkningen i Finland
Finlands folkmängd är cirka 5,5 miljoner människor.
Finland är ett mycket glesbefolkat land.
Befolkningen är framför allt koncentrerad till de stora städerna och tätorterna.
I huvudstadsregionen bor över en miljon människor.
Finlands befolkningfinska _ svenska _ engelska
Finska och svenska är Finlands nationalspråk.
Strax under 4,9 miljoner människor har finska som modersmål, medan strax under 300 000 människor talar svenska.
De största språken efter finska och svenska är ryska, estniska, engelska, somaliska och arabiska.
Till befolkningen i Finland hör olika slags minoriteter som till exempel har ett annat modersmål, en annan kultur eller religion än majoriteten av finländarna.
Traditionella minoriteter i Finland är till exempel finlandssvenskarna, samerna, romerna, judarna och tatarerna.
Dessutom har Finland fått invandrare till exempel från Ryssland, Estland, länderna på Balkan, Somalia och Irak.
Religioner i Finland
De flesta finländarna är kristna.
Det största religiösa samfundet är evangelisk-lutherska kyrkan i Finland, där cirka 70 procent av befolkningen är medlemmar.
Ortodoxa kyrkan i Finland är landets näst största religiösa samfund.
Drygt en procent av befolkningen hör till den ortodoxa kyrkan.
Den evangelisk-lutherska och den ortodoxa kyrkan har en särställning i Finland.
De har till exempel rätt att uppbära skatt.
I Finland bor tiotusentals muslimer.
Av dem hör emellertid endast en del till de islamska samfunden.
I Finland bor även några tusen judar.
I Helsingfors och Åbo finns en synagoga.
Andra religiösa samfund i Finland är till exempel Katolska kyrkan i Finland, Pingstkyrkan i Finland, Frikyrkan i Finland, Adventkyrkan i Finland, mormonkyrkan och Jehovas vittnen.
linkkiUndervisnings- och kulturministeriet:
Religiösa samfundfinska _ svenska _ engelska
Religiösa samfundfinska _ engelska
Religionsfrihet och religionsutövande i Finland
I Finland råder religionsfrihet.
Alla som bor i Finland har rätt att själva välja sin religion och utöva den.
Om man inte vill, måste man inte välja någon religion alls.
Ingen kan heller mot sin vilja tvingas att delta i religionsutövande.
linkkiUndervisnings- och kulturministeriet:
Religionsfrihetfinska _ svenska _ engelska
Minst 20 myndiga personer kan grunda ett religiöst samfund.
Religiösa grupper måste inte registrera sig som samfund, utan de kan även verka utan att ha registrerat sig.
linkkiPatent- och registerstyrelsen:
Registrering av ett religiöst samfundfinska _ svenska _ engelska
Barnets religion
Föräldrarna bestämmer barnets religion.
Om föräldrarna inte är överens, kan modern fatta beslut om religionstillhörigheten för ett barn som inte har fyllt ett år.
Barnet har rätt att få undervisning i sin egen religion i skolan.
Läs mer på InfoFinlands sida Grundläggande utbildning.
En myndig person, alltså en person som har fyllt 18 år, får själv besluta om sin religion.
Det innebär att staten inte kan bestämma vad som sägs i medier som dagstidningar, television eller internet.
Nyheter och tv-program på internet
linkkiYLE:
linkkiYLE:
Nyheter på ryskaryska
linkkiYLE:
Nyheter på lättläst finskafinska
Nyheter på lättläst finskafinska
Tidningar
I Finland utkommer många tidningar.
Tidningen med den största upplagan är Helsingin Sanomat.
De flesta tidningarna är finskspråkiga.
På vissa orter utkommer även svenskspråkiga tidningar.
I Finland utkommer även den ryskspråkiga tidskriften Spektr.
linkkiTidningarnas föbund:
Tidningar i Finlandfinska
Ryskspråkig tidskriftryska
Television
Om du har en gammal tv, behöver du också en digitalbox för att titta på tv-program.
Nya tv-apparater som säljs i Finland har redan inbyggd digitalbox.
De flesta tv-programmen är finskspråkiga.
I Finland har program på främmande språk text på finska eller svenska, med andra ord kan man också titta på dem på originalspråket (oftast engelska).
Rundradion, det vill säga Yle, äger fyra tv-kanaler som visas i hela landet.
Yle är en offentlig tjänst och dess verksamhet bekostas med skattepengar.
Utöver den finns det flera kommersiella tv-kanaler i Finland, till exempel MTV3 och Nelonen.
Vissa tv-program kan du titta på avgiftsfritt.
Yles kanaler och flera kommersiella kanaler är avgiftsfria.
Du kan också köpa avgiftsbelagda kanaler.
linkkiExpatFinland:
Televisionen i Finlandengelska
linkkitvguido.com:
Programguideengelska
Radio
I Finland finns det flera radiokanaler.
Du kan lyssna på största delen av kanalerna också på webben.
Största delen av kanalerna är finskspråkiga.
Yles radiokanal Mondo erbjuder radioprogram på engelska och många andra språk.
Radio Sputnik är en ryskspråkig radiokanal.
Finest sänder radioprogram på estniska.
Radiokanalerna i Finlandfinska
Det innebär att staten inte kan bestämma vad som sägs i medier som dagstidningar, television eller internet.
Nyheter och tv-program på internet
linkkiYLE:
linkkiYLE:
Nyheter på ryskaryska
linkkiYLE:
Nyheter på lättläst finskafinska
Nyheter på lättläst finskafinska
Tidningar
I Finland utkommer många tidningar.
Tidningen med den största upplagan är Helsingin Sanomat.
De flesta tidningarna är finskspråkiga.
På vissa orter utkommer även svenskspråkiga tidningar.
I Finland utkommer även den ryskspråkiga tidskriften Spektr.
linkkiTidningarnas föbund:
Tidningar i Finlandfinska
Ryskspråkig tidskriftryska
Television
Om du har en gammal tv, behöver du också en digitalbox för att titta på tv-program.
Nya tv-apparater som säljs i Finland har redan inbyggd digitalbox.
De flesta tv-programmen är finskspråkiga.
I Finland har program på främmande språk text på finska eller svenska, med andra ord kan man också titta på dem på originalspråket (oftast engelska).
Rundradion, det vill säga Yle, äger fyra tv-kanaler som visas i hela landet.
Yle är en offentlig tjänst och dess verksamhet bekostas med skattepengar.
Utöver den finns det flera kommersiella tv-kanaler i Finland, till exempel MTV3 och Nelonen.
Vissa tv-program kan du titta på avgiftsfritt.
Yles kanaler och flera kommersiella kanaler är avgiftsfria.
Du kan också köpa avgiftsbelagda kanaler.
linkkiExpatFinland:
Televisionen i Finlandengelska
linkkitvguido.com:
Programguideengelska
Radio
I Finland finns det flera radiokanaler.
Du kan lyssna på största delen av kanalerna också på webben.
Största delen av kanalerna är finskspråkiga.
Yles radiokanal Mondo erbjuder radioprogram på engelska och många andra språk.
Radio Sputnik är en ryskspråkig radiokanal.
Finest sänder radioprogram på estniska.
Radiokanalerna i Finlandfinska
Det innebär att staten inte kan bestämma vad som sägs i medier som dagstidningar, television eller internet.
Nyheter och tv-program på internet
linkkiYLE:
linkkiYLE:
Nyheter på ryskaryska
linkkiYLE:
Nyheter på lättläst finskafinska
Nyheter på lättläst finskafinska
Tidningar
I Finland utkommer många tidningar.
Tidningen med den största upplagan är Helsingin Sanomat.
De flesta tidningarna är finskspråkiga.
På vissa orter utkommer även svenskspråkiga tidningar.
I Finland utkommer även den ryskspråkiga tidskriften Spektr.
linkkiTidningarnas föbund:
Tidningar i Finlandfinska
Ryskspråkig tidskriftryska
Television
Om du har en gammal tv, behöver du också en digitalbox för att titta på tv-program.
Nya tv-apparater som säljs i Finland har redan inbyggd digitalbox.
De flesta tv-programmen är finskspråkiga.
I Finland har program på främmande språk text på finska eller svenska, med andra ord kan man också titta på dem på originalspråket (oftast engelska).
Rundradion, det vill säga Yle, äger fyra tv-kanaler som visas i hela landet.
Yle är en offentlig tjänst och dess verksamhet bekostas med skattepengar.
Utöver den finns det flera kommersiella tv-kanaler i Finland, till exempel MTV3 och Nelonen.
Vissa tv-program kan du titta på avgiftsfritt.
Yles kanaler och flera kommersiella kanaler är avgiftsfria.
Du kan också köpa avgiftsbelagda kanaler.
linkkiExpatFinland:
Televisionen i Finlandengelska
linkkitvguido.com:
Programguideengelska
Radio
I Finland finns det flera radiokanaler.
Du kan lyssna på största delen av kanalerna också på webben.
Största delen av kanalerna är finskspråkiga.
Yles radiokanal Mondo erbjuder radioprogram på engelska och många andra språk.
Radio Sputnik är en ryskspråkig radiokanal.
Finest sänder radioprogram på estniska.
Radiokanalerna i Finlandfinska
På den här sidan finns information om tjänsterna i Rovaniemi.
Motion
I Rovaniemi finns mångsidiga motionsmöjligheter.
Rovaniemi stads idrottstjänster erbjuder personer över 27 år (inte heltidsstuderande) möjlighet till regelbunden motion i hälsomotionsgrupper.
Syftet med verksamheten är att hjälpa nybörjare att komma igång med motion och tillhandahålla motionsformer som passar för nybörjare.
Målet är att med hjälp av motion förbättra både den psykiska hälsan och den fysiska konditionen.
Mer information om Rovaniemi stads idrottstjänster och hälsomotionskalendern hittar du under följande länk:
Rovaniemi stad/idrottstjänster linkkiRovaniemi stad/idrottstjänster:
Hälsomotion för personer i arbetsför ålderfinska
Rovaniemi stad/idrottstjänster linkkiRovaniemi stad/idrottstjänster:
Kontaktuppgifterfinska
Simhallar
Badhuset/simhallen Vesihiisi
Nuortenkatu 11
tfn 016 322 2592
Badhuset/+simhallen Vesihiisifinska
Santa Sport Spa
Hiihtomajantie 2
tfn 020 798 4200
linkkiSanta Sport :
Santa Sport Spafinska
Bibliotek
Lapplands landskapsbibliotek
Lapplands landskapsbibliotek/alla verksamhetsställen linkkiLapplands landskapsbibliotek/alla verksamhetsställen:
Öppettider och kontaktuppgifterfinska
Bybibliotek linkkiBybiblioteken:
Öppettider och kontaktuppgifterfinska
Bokbussarnas rutter och tidtabellerfinska
Tjänster för unga
Rovaniemi stads ungdomstjänster ordnar intressanta aktiviteter och intressant verksamhet för unga.
De viktigaste verksamhetsformerna består av ungdomsgårdarna, stora ungdomsevenemang, utflykter, internationella utbyten för ungdomsgrupper och sommarkollon för barn.
Centralen för ungdomstjänster ordnar verksamhet vanligtvis när ungdomarna är lediga, det vill säga på kvällstid, veckoslut och under lov.
All verksamhet ordnas av utbildade medarbetare.
Byrån för ungdomstjänster
Du hittar byrån för ungdomstjänster vid Salutorget, på övervåningen i Monde ungdomsgård.
Ingången till byrån för ungdomstjänster ligger på torgsidan. Ta trappan upp till andra våningen.
Besöksadress:
LaNuti linkkiLaNuti:
Lapplands rådgivnings- och informationsservice för ungafinska
Ungdomsgårdar
I Rovaniemi finns ungdomsgårdar i åtta olika områden: centrum, Korkalovaara, Nivavaara och Ylikylä samt byarna Muurola, Sinettä, Oikarainen och Vanttauskoski.
Ungdomsgården är centret för ungdomsarbetet i respektive område.
De ordnar verksamhet under 2–5 dagar i veckan med tyngdpunkt på fredagar och lördagar.
Verksamheten är avsedd för alla ungdomar i åldersspannet 13–20 år.
Regionala ungdomstjänsterfinska
Ungdomsgårdarna är ungdomarnas egna lokaler där de tillsammans med ungdomsledarna kan syssla med sådant som är viktigt för dem.
I verksamheten förenas aktiviteter, fostran och social gemenskap i lagom grad.
Den centrala målsättningen är att producera verksamhet som samtidigt är uppfostrande och intressant för de unga, som stöder deras utveckling och uppväxt och som stärker deras samhälleliga delaktighet.
Typiska ledda aktiviteter är olika temadagar och utflykter.
På ungdomsgårdarna har ungdomarna kostnadsfritt tillgång till ett mångsidigt urval av hobbyredskap, så utbudet av aktiviteter är stort.
Teater
Lapplands studentteaters webbplatsfinska _ engelska
Webbplatsen för sommarteatern Konttisen kesäteatterifinska
Bildkonst
Rovaniemi stad/kulturtjänster linkkiRovaniemi stad/kulturtjänster:
Museer
Korundifinska _ engelska
Rovaniemi stad/kulturtjänster linkkiRovaniemi stad/kulturtjänster:
Lapplands landskapsmuseumfinska
Föreningen för Lapplands skogsmuseum rf linkkiFöreningen för Lapplands skogsmuseum rf:
Lapplands skogsmuseumfinska _ engelska
Filmer
Finnkino linkkiFinnkino:
Finnkinos webbplatsfinska _ engelska
MoniNet
MoniNet är ett mångkulturellt center som bedrivs av settlementföreningen Rovalan Setlementti ry.
Vid MoniNet kan du få information om hobbyer, till exempel kurserna vid medborgarinstituten eller föreningsverksamhet.
Etelärinne 32
tfn 040 559 6564
MoniNetfinska _ engelska
På den här sidan finns information om tjänsterna i Rovaniemi.
Motion
I Rovaniemi finns mångsidiga motionsmöjligheter.
Rovaniemi stads idrottstjänster erbjuder personer över 27 år (inte heltidsstuderande) möjlighet till regelbunden motion i hälsomotionsgrupper.
Syftet med verksamheten är att hjälpa nybörjare att komma igång med motion och tillhandahålla motionsformer som passar för nybörjare.
Målet är att med hjälp av motion förbättra både den psykiska hälsan och den fysiska konditionen.
Mer information om Rovaniemi stads idrottstjänster och hälsomotionskalendern hittar du under följande länk:
Rovaniemi stad/idrottstjänster linkkiRovaniemi stad/idrottstjänster:
Hälsomotion för personer i arbetsför ålderfinska
Rovaniemi stad/idrottstjänster linkkiRovaniemi stad/idrottstjänster:
Kontaktuppgifterfinska
Simhallar
Badhuset/simhallen Vesihiisi
Nuortenkatu 11
tfn 016 322 2592
Badhuset/+simhallen Vesihiisifinska
Santa Sport Spa
Hiihtomajantie 2
tfn 020 798 4200
linkkiSanta Sport :
Santa Sport Spafinska _ engelska
Bibliotek
Lapplands landskapsbibliotek
Lapplands landskapsbibliotek/alla verksamhetsställen linkkiLapplands landskapsbibliotek/alla verksamhetsställen:
Öppettider och kontaktuppgifterfinska
Bybibliotek linkkiBybiblioteken:
Öppettider och kontaktuppgifterfinska
Bokbussarnas rutter och tidtabellerfinska
Tjänster för unga
Rovaniemi stads ungdomstjänster ordnar intressanta aktiviteter och intressant verksamhet för unga.
De viktigaste verksamhetsformerna består av ungdomsgårdarna, stora ungdomsevenemang, utflykter, internationella utbyten för ungdomsgrupper och sommarkollon för barn.
Centralen för ungdomstjänster ordnar verksamhet vanligtvis när ungdomarna är lediga, det vill säga på kvällstid, veckoslut och under lov.
All verksamhet ordnas av utbildade medarbetare.
Byrån för ungdomstjänster
Du hittar byrån för ungdomstjänster vid Salutorget, på övervåningen i Monde ungdomsgård.
Ingången till byrån för ungdomstjänster ligger på torgsidan. Ta trappan upp till andra våningen.
Besöksadress:
LaNuti linkkiLaNuti:
Lapplands rådgivnings- och informationsservice för ungafinska
Ungdomsgårdar
I Rovaniemi finns ungdomsgårdar i åtta olika områden: centrum, Korkalovaara, Nivavaara och Ylikylä samt byarna Muurola, Sinettä, Oikarainen och Vanttauskoski.
Ungdomsgården är centret för ungdomsarbetet i respektive område.
De ordnar verksamhet under 2–5 dagar i veckan med tyngdpunkt på fredagar och lördagar.
Verksamheten är avsedd för alla ungdomar i åldersspannet 13–20 år.
Regionala ungdomstjänsterfinska
Ungdomsgårdarna är ungdomarnas egna lokaler där de tillsammans med ungdomsledarna kan syssla med sådant som är viktigt för dem.
I verksamheten förenas aktiviteter, fostran och social gemenskap i lagom grad.
Den centrala målsättningen är att producera verksamhet som samtidigt är uppfostrande och intressant för de unga, som stöder deras utveckling och uppväxt och som stärker deras samhälleliga delaktighet.
Typiska ledda aktiviteter är olika temadagar och utflykter.
På ungdomsgårdarna har ungdomarna kostnadsfritt tillgång till ett mångsidigt urval av hobbyredskap, så utbudet av aktiviteter är stort.
Teater
Lapplands studentteaters webbplatsfinska _ engelska
Webbplatsen för sommarteatern Konttisen kesäteatterifinska
Bildkonst
Rovaniemi stad/kulturtjänster linkkiRovaniemi stad/kulturtjänster:
Museer
Korundifinska _ engelska
Rovaniemi stad/kulturtjänster linkkiRovaniemi stad/kulturtjänster:
Lapplands landskapsmuseumfinska
Föreningen för Lapplands skogsmuseum rf linkkiFöreningen för Lapplands skogsmuseum rf:
Lapplands skogsmuseumfinska _ engelska
MoniNet
MoniNet är ett mångkulturellt center som bedrivs av settlementföreningen Rovalan Setlementti ry.
Vid MoniNet kan du få information om hobbyer, till exempel kurserna vid medborgarinstituten eller föreningsverksamhet.
Etelärinne 32
tfn 040 559 6564
MoniNetfinska _ engelska
På den här sidan finns information om tjänsterna i Rovaniemi.
Motion
I Rovaniemi finns mångsidiga motionsmöjligheter.
Rovaniemi stads idrottstjänster erbjuder personer över 27 år (inte heltidsstuderande) möjlighet till regelbunden motion i hälsomotionsgrupper.
Syftet med verksamheten är att hjälpa nybörjare att komma igång med motion och tillhandahålla motionsformer som passar för nybörjare.
Målet är att med hjälp av motion förbättra både den psykiska hälsan och den fysiska konditionen.
Mer information om Rovaniemi stads idrottstjänster och hälsomotionskalendern hittar du under följande länk:
Rovaniemi stad/idrottstjänster linkkiRovaniemi stad/idrottstjänster:
Hälsomotion för personer i arbetsför ålderfinska
Rovaniemi stad/idrottstjänster linkkiRovaniemi stad/idrottstjänster:
Kontaktuppgifterfinska
Simhallar
Badhuset/simhallen Vesihiisi
Nuortenkatu 11
tfn 016 322 2592
Badhuset/+simhallen Vesihiisifinska
Santa Sport Spa
Hiihtomajantie 2
tfn 020 798 4200
linkkiSanta Sport :
Santa Sport Spafinska _ engelska
Bibliotek
Lapplands landskapsbibliotek
Lapplands landskapsbibliotek/alla verksamhetsställen linkkiLapplands landskapsbibliotek/alla verksamhetsställen:
Öppettider och kontaktuppgifterfinska
Bybibliotek linkkiBybiblioteken:
Öppettider och kontaktuppgifterfinska
Bokbussarnas rutter och tidtabellerfinska
Tjänster för unga
Rovaniemi stads ungdomstjänster ordnar intressanta aktiviteter och intressant verksamhet för unga.
De viktigaste verksamhetsformerna består av ungdomsgårdarna, stora ungdomsevenemang, utflykter, internationella utbyten för ungdomsgrupper och sommarkollon för barn.
Centralen för ungdomstjänster ordnar verksamhet vanligtvis när ungdomarna är lediga, det vill säga på kvällstid, veckoslut och under lov.
All verksamhet ordnas av utbildade medarbetare.
Byrån för ungdomstjänster
Du hittar byrån för ungdomstjänster vid Salutorget, på övervåningen i Monde ungdomsgård.
Ingången till byrån för ungdomstjänster ligger på torgsidan. Ta trappan upp till andra våningen.
Besöksadress:
LaNuti linkkiLaNuti:
Lapplands rådgivnings- och informationsservice för ungafinska
Ungdomsgårdar
I Rovaniemi finns ungdomsgårdar i åtta olika områden: centrum, Korkalovaara, Nivavaara och Ylikylä samt byarna Muurola, Sinettä, Oikarainen och Vanttauskoski.
Ungdomsgården är centret för ungdomsarbetet i respektive område.
De ordnar verksamhet under 2–5 dagar i veckan med tyngdpunkt på fredagar och lördagar.
Verksamheten är avsedd för alla ungdomar i åldersspannet 13–20 år.
Regionala ungdomstjänsterfinska
Ungdomsgårdarna är ungdomarnas egna lokaler där de tillsammans med ungdomsledarna kan syssla med sådant som är viktigt för dem.
I verksamheten förenas aktiviteter, fostran och social gemenskap i lagom grad.
Den centrala målsättningen är att producera verksamhet som samtidigt är uppfostrande och intressant för de unga, som stöder deras utveckling och uppväxt och som stärker deras samhälleliga delaktighet.
Typiska ledda aktiviteter är olika temadagar och utflykter.
På ungdomsgårdarna har ungdomarna kostnadsfritt tillgång till ett mångsidigt urval av hobbyredskap, så utbudet av aktiviteter är stort.
Teater
Lapplands studentteaters webbplatsfinska _ engelska
Webbplatsen för sommarteatern Konttisen kesäteatterifinska
Bildkonst
Rovaniemi stad/kulturtjänster linkkiRovaniemi stad/kulturtjänster:
Museer
Korundifinska _ engelska
Rovaniemi stad/kulturtjänster linkkiRovaniemi stad/kulturtjänster:
Lapplands landskapsmuseumfinska
Föreningen för Lapplands skogsmuseum rf linkkiFöreningen för Lapplands skogsmuseum rf:
Lapplands skogsmuseumfinska _ engelska
MoniNet
MoniNet är ett mångkulturellt center som bedrivs av settlementföreningen Rovalan Setlementti ry.
Vid MoniNet kan du få information om hobbyer, till exempel kurserna vid medborgarinstituten eller föreningsverksamhet.
Etelärinne 32
tfn 040 559 6564
MoniNetfinska _ engelska
Kollektivtrafiken
Kollektivtrafiken fungerar väl i Finland.
Man kan resa nästan över allt i Finland med tåg eller buss.
Man kan också flyga till många städer.
I stora städer och deras näromgivning finns en välfungerande lokaltrafik.
Lokaltrafiken trafikeras vanligtvis med bussar.
Tåg
Tågtrafiken i Finland sköts av bolaget VR.
Du kan köpa tågbiljetter på VR:s webbplats, på järnvägsstationer och ombord på tågen.
Information om tågtidtabellerna hittar du på VR:s webbplats och på järnvägsstationerna.
linkkiVR:
Tågbiljetterfinska _ svenska _ engelska _ ryska
Bussar
Det finns många bussbolag i Finland.
Du kan köpa biljetter på Matkahuoltos verksamhetsställen och webbplats.
Information om busstidtabellerna hittar du på Matkahuoltos webbplats och verksamhetsställen.
Rabatt på bussbiljetter ges åt
barn
studerande
pensionärer
beväringar och civiltjänstgörare
På trafikverkets webbplats finns kollektivtrafikens reseplanerare, matka.fi, där du kan söka den bästa rutten och det bästa resesättet.
Bussbiljetterfinska _ svenska _ engelska
Ruttjänstenfinska _ svenska _ engelska
Flygtrafiken
I Finland finns det 24 flygplatser.
Den största av dem är Helsingfors-Vanda flygplats.
Många flygbolag erbjuder flyg från Finland till utlandet.
De flesta utrikesflygen avgår från Helsingfors-Vanda flygplats.
linkkiFinavia:
Flygplatserna i Finlandfinska _ engelska
Egen bil
Det är relativt dyrt att köpa och använda en bil i Finland.
En välhållen bil kostar flera tusen euro.
Också ägandet och användningen av bilen medför kostnader, till exempel för
bensin
försäkringar
däck
service och reparationer
bilskatter
Om du har en bil måste du teckna en trafikförsäkring (liikennevakuutus).
Trafikförsäkringen tecknar du hos ett försäkringsbolag.
I Finland måste bilen besiktigas och registreras.
Besiktningar görs på besiktningsstationer.
Registreringen kan göras till exempel på besiktningsstationer, vid försäkringsbolag och hos bilhandlare.
Du kan även registrera bilen på Internet.
I Finland är det lag på att bilen ska ha vinterdäck på vintern.
På vintern kan man använda antingen dubbdäck eller friktionsdäck.
En bil med dubbdäck är lättare att manövrera på hala vägar.
Du kan dock inte använda dubbdäcken på sommaren.
I Finland måste du noga iaktta trafikreglerna.
Polisen övervakar att trafikreglerna följs.
Om man bryter mot trafikreglerna kan man få böter.
Att framföra vilket som helst motorfordon i onyktert tillstånd (alkohol eller droger) är ett brott.
linkkiExpatFinland.com:
Bil och körning i Finlandengelska
linkkiTrafiksäkerhetsverket:
Information om registrering av fordonfinska _ svenska _ engelska
linkkiTrafiksäkerhetsverket:
Registrering av fordon på Internetfinska _ svenska _ engelska
linkkiTrafiksäkerhetsverket:
Besiktning av fordonfinska _ svenska
linkkiTrafiksäkerhetsverket:
Information om fordonsbeskattningfinska _ svenska _ engelska
Information om bildäckfinska _ svenska _ engelska
Körkort
För att få köra bil måste du ha körkort.
För att få körkort måste du vara minst 18 år.
Innan du kan få körkort måste du delta i förarutbildning och avlägga förarexamen.
Förarutbildning kan du få i en bilskola.
Också till exempel en släkting eller en bekant som har körkort och erfarenhet av att köra bil kan lära dig.
För detta behövs dock ett undervisningstillstånd från Trafi.
linkkiTrafiksäkerhetsverket Trafi:
Undervisningstillståndfinska _ svenska
För att få köra motorcykel behöver du ett motorcykelkort.
Vilket kort du behöver beror på hurdan motorcykel du vill köra.
För att köra moped behöver du ett mopedkort, om du inte har ett körkort.
Du behöver inget mopedkort om du har fyllt 15 år före den 1 januari 2000.
Du hittar information om körkort på polisens och Trafiksäkerhetsverkets (Liikenteen turvallisuusvirasto) webbplatser.
Utländskt körkort i Finland
Om du har ett körkort som utfärdats i ett av de nordiska länderna eller i ett EU-/EES-land, är det giltigt även i Finland.
Om du bor stadigvarande i Finland kan du byta ut kortet mot ett finländskt körkort.
Om du har ett körkort som utfärdats i ett land som är anslutet till Genève- eller Wien-konventionerna kan du köra med detta kort högst två år i Finland.
Du måste byta ut ditt körkort mot ett finländskt körkort inom två år efter att du flyttat till Finland.
Om du har ett körkort som utfärdats i ett land som inte är anslutet till Genève- eller Wien-konventionerna kan du köra bil med detta kort under ett års tid efter att ha registrerats i befolkningsregistret i Finland.
Du kan byta ut ditt körkort till ett finskt körkort på Ajovarmas serviceställen.
Du kan boka en tid i förväg på Ajovarmas webbplats.
linkkiTrafiksäkerhetsverket:
Information om körkortfinska _ svenska
linkkiTrafiksäkerhetsverket:
Utländskt körkort i Finlandfinska _ svenska _ engelska
Kollektivtrafiken
Kollektivtrafiken fungerar väl i Finland.
Man kan resa nästan över allt i Finland med tåg eller buss.
Man kan också flyga till många städer.
I stora städer och deras näromgivning finns en välfungerande lokaltrafik.
Lokaltrafiken trafikeras vanligtvis med bussar.
Tåg
Tågtrafiken i Finland sköts av bolaget VR.
Du kan köpa tågbiljetter på VR:s webbplats, på järnvägsstationer och ombord på tågen.
Information om tågtidtabellerna hittar du på VR:s webbplats och på järnvägsstationerna.
linkkiVR:
Tågbiljetterfinska _ svenska _ engelska _ ryska
Bussar
Det finns många bussbolag i Finland.
Du kan köpa biljetter på Matkahuoltos verksamhetsställen och webbplats.
Information om busstidtabellerna hittar du på Matkahuoltos webbplats och verksamhetsställen.
Rabatt på bussbiljetter ges åt
barn
studerande
pensionärer
beväringar och civiltjänstgörare
På trafikverkets webbplats finns kollektivtrafikens reseplanerare, matka.fi, där du kan söka den bästa rutten och det bästa resesättet.
Bussbiljetterfinska _ svenska _ engelska
Ruttjänstenfinska _ svenska _ engelska
Flygtrafiken
I Finland finns det 24 flygplatser.
Den största av dem är Helsingfors-Vanda flygplats.
Många flygbolag erbjuder flyg från Finland till utlandet.
De flesta utrikesflygen avgår från Helsingfors-Vanda flygplats.
linkkiFinavia:
Flygplatserna i Finlandfinska _ engelska
Egen bil
Det är relativt dyrt att köpa och använda en bil i Finland.
En välhållen bil kostar flera tusen euro.
Också ägandet och användningen av bilen medför kostnader, till exempel för
bensin
försäkringar
däck
service och reparationer
bilskatter
Om du har en bil måste du teckna en trafikförsäkring (liikennevakuutus).
Trafikförsäkringen tecknar du hos ett försäkringsbolag.
I Finland måste bilen besiktigas och registreras.
Besiktningar görs på besiktningsstationer.
Registreringen kan göras till exempel på besiktningsstationer, vid försäkringsbolag och hos bilhandlare.
Du kan även registrera bilen på Internet.
I Finland är det lag på att bilen ska ha vinterdäck på vintern.
På vintern kan man använda antingen dubbdäck eller friktionsdäck.
En bil med dubbdäck är lättare att manövrera på hala vägar.
Du kan dock inte använda dubbdäcken på sommaren.
I Finland måste du noga iaktta trafikreglerna.
Polisen övervakar att trafikreglerna följs.
Om man bryter mot trafikreglerna kan man få böter.
Att framföra vilket som helst motorfordon i onyktert tillstånd (alkohol eller droger) är ett brott.
linkkiExpatFinland.com:
Bil och körning i Finlandengelska
linkkiTrafiksäkerhetsverket:
Information om registrering av fordonfinska _ svenska _ engelska
linkkiTrafiksäkerhetsverket:
Registrering av fordon på Internetfinska _ svenska _ engelska
linkkiTrafiksäkerhetsverket:
Besiktning av fordonfinska _ svenska
linkkiTrafiksäkerhetsverket:
Information om fordonsbeskattningfinska _ svenska _ engelska
Information om bildäckfinska _ svenska _ engelska
Körkort
För att få köra bil måste du ha körkort.
För att få körkort måste du vara minst 18 år.
Innan du kan få körkort måste du delta i förarutbildning och avlägga förarexamen.
Förarutbildning kan du få i en bilskola.
Också till exempel en släkting eller en bekant som har körkort och erfarenhet av att köra bil kan lära dig.
För detta behövs dock ett undervisningstillstånd från Trafi.
linkkiTrafiksäkerhetsverket Trafi:
Undervisningstillståndfinska _ svenska
För att få köra motorcykel behöver du ett motorcykelkort.
Vilket kort du behöver beror på hurdan motorcykel du vill köra.
För att köra moped behöver du ett mopedkort, om du inte har ett körkort.
Du behöver inget mopedkort om du har fyllt 15 år före den 1 januari 2000.
Du hittar information om körkort på polisens och Trafiksäkerhetsverkets (Liikenteen turvallisuusvirasto) webbplatser.
Utländskt körkort i Finland
Om du har ett körkort som utfärdats i ett av de nordiska länderna eller i ett EU-/EES-land, är det giltigt även i Finland.
Om du bor stadigvarande i Finland kan du byta ut kortet mot ett finländskt körkort.
Om du har ett körkort som utfärdats i ett land som är anslutet till Genève- eller Wien-konventionerna kan du köra med detta kort högst två år i Finland.
Du måste byta ut ditt körkort mot ett finländskt körkort inom två år efter att du flyttat till Finland.
Om du har ett körkort som utfärdats i ett land som inte är anslutet till Genève- eller Wien-konventionerna kan du köra bil med detta kort under ett års tid efter att ha registrerats i befolkningsregistret i Finland.
Du kan byta ut ditt körkort till ett finskt körkort på Ajovarmas serviceställen.
Du kan boka en tid i förväg på Ajovarmas webbplats.
linkkiTrafiksäkerhetsverket:
Information om körkortfinska _ svenska
linkkiTrafiksäkerhetsverket:
Utländskt körkort i Finlandfinska _ svenska _ engelska
Kollektivtrafiken
Kollektivtrafiken fungerar väl i Finland.
Man kan resa nästan över allt i Finland med tåg eller buss.
Man kan också flyga till många städer.
I stora städer och deras näromgivning finns en välfungerande lokaltrafik.
Lokaltrafiken trafikeras vanligtvis med bussar.
Tåg
Tågtrafiken i Finland sköts av bolaget VR.
Du kan köpa tågbiljetter på VR:s webbplats, på järnvägsstationer och ombord på tågen.
Information om tågtidtabellerna hittar du på VR:s webbplats och på järnvägsstationerna.
linkkiVR:
Tågbiljetterfinska _ svenska _ engelska _ ryska
Bussar
Det finns många bussbolag i Finland.
Du kan köpa biljetter på Matkahuoltos verksamhetsställen och webbplats.
Information om busstidtabellerna hittar du på Matkahuoltos webbplats och verksamhetsställen.
Rabatt på bussbiljetter ges åt
barn
studerande
pensionärer
beväringar och civiltjänstgörare
På trafikverkets webbplats finns kollektivtrafikens reseplanerare, matka.fi, där du kan söka den bästa rutten och det bästa resesättet.
Bussbiljetterfinska _ svenska _ engelska
Ruttjänstenfinska _ svenska _ engelska
Flygtrafiken
I Finland finns det 24 flygplatser.
Den största av dem är Helsingfors-Vanda flygplats.
Många flygbolag erbjuder flyg från Finland till utlandet.
De flesta utrikesflygen avgår från Helsingfors-Vanda flygplats.
linkkiFinavia:
Flygplatserna i Finlandfinska _ engelska
Egen bil
Det är relativt dyrt att köpa och använda en bil i Finland.
En välhållen bil kostar flera tusen euro.
Också ägandet och användningen av bilen medför kostnader, till exempel för
bensin
försäkringar
däck
service och reparationer
bilskatter
Om du har en bil måste du teckna en trafikförsäkring (liikennevakuutus).
Trafikförsäkringen tecknar du hos ett försäkringsbolag.
I Finland måste bilen besiktigas och registreras.
Besiktningar görs på besiktningsstationer.
Registreringen kan göras till exempel på besiktningsstationer, vid försäkringsbolag och hos bilhandlare.
Du kan även registrera bilen på Internet.
I Finland är det lag på att bilen ska ha vinterdäck på vintern.
På vintern kan man använda antingen dubbdäck eller friktionsdäck.
En bil med dubbdäck är lättare att manövrera på hala vägar.
Du kan dock inte använda dubbdäcken på sommaren.
I Finland måste du noga iaktta trafikreglerna.
Polisen övervakar att trafikreglerna följs.
Om man bryter mot trafikreglerna kan man få böter.
Att framföra vilket som helst motorfordon i onyktert tillstånd (alkohol eller droger) är ett brott.
linkkiExpatFinland.com:
Bil och körning i Finlandengelska
linkkiTrafiksäkerhetsverket:
Information om registrering av fordonfinska _ svenska _ engelska
linkkiTrafiksäkerhetsverket:
Registrering av fordon på Internetfinska _ svenska _ engelska
linkkiTrafiksäkerhetsverket:
Besiktning av fordonfinska _ svenska
linkkiTrafiksäkerhetsverket:
Information om fordonsbeskattningfinska _ svenska _ engelska
Information om bildäckfinska _ svenska _ engelska
Körkort
För att få köra bil måste du ha körkort.
För att få körkort måste du vara minst 18 år.
Innan du kan få körkort måste du delta i förarutbildning och avlägga förarexamen.
Förarutbildning kan du få i en bilskola.
Också till exempel en släkting eller en bekant som har körkort och erfarenhet av att köra bil kan lära dig.
För detta behövs dock ett undervisningstillstånd från Trafi.
linkkiTrafiksäkerhetsverket Trafi:
Undervisningstillståndfinska _ svenska
För att få köra motorcykel behöver du ett motorcykelkort.
Vilket kort du behöver beror på hurdan motorcykel du vill köra.
För att köra moped behöver du ett mopedkort, om du inte har ett körkort.
Du behöver inget mopedkort om du har fyllt 15 år före den 1 januari 2000.
Du hittar information om körkort på polisens och Trafiksäkerhetsverkets (Liikenteen turvallisuusvirasto) webbplatser.
Utländskt körkort i Finland
Om du har ett körkort som utfärdats i ett av de nordiska länderna eller i ett EU-/EES-land, är det giltigt även i Finland.
Om du bor stadigvarande i Finland kan du byta ut kortet mot ett finländskt körkort.
Om du har ett körkort som utfärdats i ett land som är anslutet till Genève- eller Wien-konventionerna kan du köra med detta kort högst två år i Finland.
Du måste byta ut ditt körkort mot ett finländskt körkort inom två år efter att du flyttat till Finland.
Om du har ett körkort som utfärdats i ett land som inte är anslutet till Genève- eller Wien-konventionerna kan du köra bil med detta kort under ett års tid efter att ha registrerats i befolkningsregistret i Finland.
Du kan byta ut ditt körkort till ett finskt körkort på Ajovarmas serviceställen.
Du kan boka en tid i förväg på Ajovarmas webbplats.
linkkiTrafiksäkerhetsverket:
Information om körkortfinska _ svenska
linkkiTrafiksäkerhetsverket:
Utländskt körkort i Finlandfinska _ svenska _ engelska
Klimatet i Finland är kallare än i många andra länder.
Vädret varierar ändå mycket under olika årstider.
Vinter
På vintern är det kallt och snöar i Finland.
Vanligen stannar snön kvar på marken hela vintern.
Temperaturen är oftast under noll grader celsius.
Temperaturen kan t.ex. dagtid vara -10 Celsiusgrader och ibland till och med -20 grader.
I norra Finland kan temperaturen vara till och med -30 grader.
Om det är snö och is på marken är det också halt.
Det är viktigt att klä sig varmt på vintern.
Det betyder att det är bra att klä på sig åtminstone en täckjacka, ylletröja, mössa, handskar, halsduk och varma vinterskor.
Vid kallt väder lönar det sig att ha på sig flera lager med kläder.
På vintern är det ofta mörkt i Finland, eftersom solen går upp först på förmiddagen och går ner redan på eftermiddagen.
I norra Finland är det mörkare än i södra Finland.
I de nordligaste delarna av Finland går det flera veckor utan att solen går upp överhuvudtaget.
Vintermånaderna är december, januari och februari.
Även i november och mars kan vädret vara kallt och det kan snöa.
Snön smälter vanligen i mars eller april.
Att klä sig på vinternfinska
Vår
Våren börjar i Finlands södra delar i slutet av mars och i de nordligare delarna i slutet av april.
Under våren är vädret ännu svalt, men varmare än på vintern.
Under våren förändras naturen en hel del, när snö och is smälter bort, löven spricker fram på träden och växterna börjar gro.
I södra Finland är medeltemperaturen på sommaren ca 20 grader Celsius, i norr ca 15 grader.
Sommarmånaderna i Finland är juni, juli och augusti.
Den varmaste månaden är juli, då stiger temperaturen dagtid ofta över 20 grader.
På sommaren är det ljust i Finland även på kvällen och natten, eftersom solen går ner sent och går upp tidigt.
I norra Finland är det ljusare än i södra Finland.
Den allra ljusaste månaden är juni.
Då firas i Finland midsommar, som är midnattssolens och högsommarens fest.
I de allra nordligaste delarna av Finland går solen inte alls ner i början av sommaren.
Höst
Hösten börjar vanligen i slutet av augusti eller början av september.
Vädret är svalt och ofta regnar och blåser det också.
På hösten är det också mörkt, eftersom solen går ner tidigare än på sommaren.
Den första snön kommer vanligen i oktober eller november.
Information om klimatet i Finlandfinska _ svenska _ engelska
Klimatet i Finland är kallare än i många andra länder.
Vädret varierar ändå mycket under olika årstider.
Vinter
På vintern är det kallt och snöar i Finland.
Vanligen stannar snön kvar på marken hela vintern.
Temperaturen är oftast under noll grader celsius.
Temperaturen kan t.ex. dagtid vara -10 Celsiusgrader och ibland till och med -20 grader.
I norra Finland kan temperaturen vara till och med -30 grader.
Om det är snö och is på marken är det också halt.
Det är viktigt att klä sig varmt på vintern.
Det betyder att det är bra att klä på sig åtminstone en täckjacka, ylletröja, mössa, handskar, halsduk och varma vinterskor.
Vid kallt väder lönar det sig att ha på sig flera lager med kläder.
På vintern är det ofta mörkt i Finland, eftersom solen går upp först på förmiddagen och går ner redan på eftermiddagen.
I norra Finland är det mörkare än i södra Finland.
I de nordligaste delarna av Finland går det flera veckor utan att solen går upp överhuvudtaget.
Vintermånaderna är december, januari och februari.
Även i november och mars kan vädret vara kallt och det kan snöa.
Snön smälter vanligen i mars eller april.
Att klä sig på vinternfinska
Vår
Våren börjar i Finlands södra delar i slutet av mars och i de nordligare delarna i slutet av april.
Under våren är vädret ännu svalt, men varmare än på vintern.
Under våren förändras naturen en hel del, när snö och is smälter bort, löven spricker fram på träden och växterna börjar gro.
I södra Finland är medeltemperaturen på sommaren ca 20 grader Celsius, i norr ca 15 grader.
Sommarmånaderna i Finland är juni, juli och augusti.
Den varmaste månaden är juli, då stiger temperaturen dagtid ofta över 20 grader.
På sommaren är det ljust i Finland även på kvällen och natten, eftersom solen går ner sent och går upp tidigt.
I norra Finland är det ljusare än i södra Finland.
Den allra ljusaste månaden är juni.
Då firas i Finland midsommar, som är midnattssolens och högsommarens fest.
I de allra nordligaste delarna av Finland går solen inte alls ner i början av sommaren.
Höst
Hösten börjar vanligen i slutet av augusti eller början av september.
Vädret är svalt och ofta regnar och blåser det också.
På hösten är det också mörkt, eftersom solen går ner tidigare än på sommaren.
Den första snön kommer vanligen i oktober eller november.
Information om klimatet i Finlandfinska _ svenska _ engelska
Klimatet i Finland är kallare än i många andra länder.
Vädret varierar ändå mycket under olika årstider.
Vinter
På vintern är det kallt och snöar i Finland.
Vanligen stannar snön kvar på marken hela vintern.
Temperaturen är oftast under noll grader celsius.
Temperaturen kan t.ex. dagtid vara -10 Celsiusgrader och ibland till och med -20 grader.
I norra Finland kan temperaturen vara till och med -30 grader.
Om det är snö och is på marken är det också halt.
Det är viktigt att klä sig varmt på vintern.
Det betyder att det är bra att klä på sig åtminstone en täckjacka, ylletröja, mössa, handskar, halsduk och varma vinterskor.
Vid kallt väder lönar det sig att ha på sig flera lager med kläder.
På vintern är det ofta mörkt i Finland, eftersom solen går upp först på förmiddagen och går ner redan på eftermiddagen.
I norra Finland är det mörkare än i södra Finland.
I de nordligaste delarna av Finland går det flera veckor utan att solen går upp överhuvudtaget.
Vintermånaderna är december, januari och februari.
Även i november och mars kan vädret vara kallt och det kan snöa.
Snön smälter vanligen i mars eller april.
Att klä sig på vinternfinska
Vår
Våren börjar i Finlands södra delar i slutet av mars och i de nordligare delarna i slutet av april.
Under våren är vädret ännu svalt, men varmare än på vintern.
Under våren förändras naturen en hel del, när snö och is smälter bort, löven spricker fram på träden och växterna börjar gro.
I södra Finland är medeltemperaturen på sommaren ca 20 grader Celsius, i norr ca 15 grader.
Sommarmånaderna i Finland är juni, juli och augusti.
Den varmaste månaden är juli, då stiger temperaturen dagtid ofta över 20 grader.
På sommaren är det ljust i Finland även på kvällen och natten, eftersom solen går ner sent och går upp tidigt.
I norra Finland är det ljusare än i södra Finland.
Den allra ljusaste månaden är juni.
Då firas i Finland midsommar, som är midnattssolens och högsommarens fest.
I de allra nordligaste delarna av Finland går solen inte alls ner i början av sommaren.
Höst
Hösten börjar vanligen i slutet av augusti eller början av september.
Vädret är svalt och ofta regnar och blåser det också.
På hösten är det också mörkt, eftersom solen går ner tidigare än på sommaren.
Den första snön kommer vanligen i oktober eller november.
Information om klimatet i Finlandfinska _ svenska _ engelska
Folk flyttar till Finland
Inflyttningen till Finland började för cirka 10 000 år sedan.
Folket kom österifrån från nuvarande Rysslands område och söderifrån via Baltikum.
Finska språket har sina rötter i de mellersta delarna av Ryssland, men har också inslag av baltiska och germanska språk.
Finland har haft svenskspråkig befolkning i över 800 år.
Finland som en del av Sverige och Ryssland
Finland var en del av Sverige i över 600 års tid från medeltiden till 1800-talets början.
Sverige och Ryssland stred under denna tid ett flertal gånger om vem som skulle vara makthavaren över Finland.
Till slut anslöts hela Finland år 1809 till Ryssland, efter att Ryssland besegrat Sverige i krig.
Under den här tiden var Finland autonomt, vilket betyder att finländarna fick själva bestämma om många saker.
Ryska kejsaren var ändå regent i Finland.
Det finska språket och den finländska kulturen och ekonomin utvecklades enormt under Finlands tid som en del av Ryssland.
I början av 1900-talet började dock Ryssland inskränka det finländska självstyret, vilket finländarna inte kunde acceptera.
Finland blir självständigt
Finland ett självständigt land och den 6 december firas än idag som Finlands självständighetsdag.
Våren 1918 befann sig Finland i inbördeskrig som kämpades mellan de röda gardena som representerade arbetarna och de vita skyddskårerna som representerade borgarna och markägarna.
Kriget avslutades i maj 1918 med de vitas seger över de röda.
Det självständiga Finland blev en republik där lagarna stiftas av en folkvald riksdag.
Statsöverhuvud är presidenten, inte en kejsare eller en kung.
Vinterkriget och fortsättningskriget
I slutet av november 1939 anföll sovjetarmén Finland.
Under andra världskriget kämpade Finland två krig mot Sovjetunionen: först vinterkriget åren 1939–1940 och därefter fortsättningskriget åren 1941–1944.
I krigen förlorade Finland områden till Sovjetunionen.
Fler än 400 000 finländare lämnade de förlorade områdena och kom som flyktingar till övriga delar av landet.
För finländarna var det ändå viktigast att ha kunnat bevara landets självständighet.
Efter krigen befarade många finländare att Sovjetunionen skulle försöka göra Finland till ett socialistiskt land, eftersom detta hade hänt Sovjetunionens andra europeiska grannländer.
Finland lyckades dock skapa goda relationer till Sovjetunionen, bibehålla sitt demokratiska system och öka handeln också med västländerna.
I utrikespolitiken tvingades Finland under en lång tid balansera mellan Sovjetunionen och väst.
Finland industrialiserades kunde finländarna sälja allt mer industriprodukter till utlandet.
Finland exporterade speciellt papper och andra produkter från skogsindustrin.
Många saker i det finländska samhället förändrades.
Många människor flyttade från landsbygden till städerna och allt fler kvinnor började arbeta utanför hemmet.
De offentliga tjänsterna började utvecklas och på så sätt skapade man den offentliga hälsovården, sociala tryggheten och grundskolan.
På 1960-talet flyttade tusentals finländare till Sverige, eftersom det fanns mer jobb och betalades högre löner i Sverige än i Finland.
När Sovjetunionen kollapsade i början av 1990-talet, hamnade Finland i ekonomisk lågkonjunktur eftersom handeln med Sovjetunionen upphörde.
Många företag gick i konkurs, vilket fick till följd att många människor förlorade sina jobb.
Efter lågkonjunkturen uppstod det mycket högteknologisk industri och högteknologiska arbetsplatser i Finland.
Allt fler människor jobbade också i olika serviceyrken.
På 1990-talet ökade inflyttningen från andra länder till Finland.
Finland fick flyktingar från många länder och hit flyttade människor med finländskt påbrå från forna Sovjetunionen.
Många flyttade till Finland även för att studera, arbeta eller för att de hade sin familj här.
År 1995 blev Finland medlem i Europeiska unionen (EU).
År 2002 införde Finland bland de första EU-länderna EU:s gemensamma valuta, euro, och gav därmed upp sin egen valuta.
Information om Finlands historiaengelska _ ryska _ franska _ spanska _ tyska _ portugisiska
Folk flyttar till Finland
Inflyttningen till Finland började för cirka 10 000 år sedan.
Folket kom österifrån från nuvarande Rysslands område och söderifrån via Baltikum.
Finska språket har sina rötter i de mellersta delarna av Ryssland, men har också inslag av baltiska och germanska språk.
Finland har haft svenskspråkig befolkning i över 800 år.
Finland som en del av Sverige och Ryssland
Finland var en del av Sverige i över 600 års tid från medeltiden till 1800-talets början.
Sverige och Ryssland stred under denna tid ett flertal gånger om vem som skulle vara makthavaren över Finland.
Till slut anslöts hela Finland år 1809 till Ryssland, efter att Ryssland besegrat Sverige i krig.
Under den här tiden var Finland autonomt, vilket betyder att finländarna fick själva bestämma om många saker.
Ryska kejsaren var ändå regent i Finland.
Det finska språket och den finländska kulturen och ekonomin utvecklades enormt under Finlands tid som en del av Ryssland.
I början av 1900-talet började dock Ryssland inskränka det finländska självstyret, vilket finländarna inte kunde acceptera.
Finland blir självständigt
Finland ett självständigt land och den 6 december firas än idag som Finlands självständighetsdag.
Våren 1918 befann sig Finland i inbördeskrig som kämpades mellan de röda gardena som representerade arbetarna och de vita skyddskårerna som representerade borgarna och markägarna.
Kriget avslutades i maj 1918 med de vitas seger över de röda.
Det självständiga Finland blev en republik där lagarna stiftas av en folkvald riksdag.
Statsöverhuvud är presidenten, inte en kejsare eller en kung.
Vinterkriget och fortsättningskriget
I slutet av november 1939 anföll sovjetarmén Finland.
Under andra världskriget kämpade Finland två krig mot Sovjetunionen: först vinterkriget åren 1939–1940 och därefter fortsättningskriget åren 1941–1944.
I krigen förlorade Finland områden till Sovjetunionen.
Fler än 400 000 finländare lämnade de förlorade områdena och kom som flyktingar till övriga delar av landet.
För finländarna var det ändå viktigast att ha kunnat bevara landets självständighet.
Efter krigen befarade många finländare att Sovjetunionen skulle försöka göra Finland till ett socialistiskt land, eftersom detta hade hänt Sovjetunionens andra europeiska grannländer.
Finland lyckades dock skapa goda relationer till Sovjetunionen, bibehålla sitt demokratiska system och öka handeln också med västländerna.
I utrikespolitiken tvingades Finland under en lång tid balansera mellan Sovjetunionen och väst.
Finland industrialiserades kunde finländarna sälja allt mer industriprodukter till utlandet.
Finland exporterade speciellt papper och andra produkter från skogsindustrin.
Många saker i det finländska samhället förändrades.
Många människor flyttade från landsbygden till städerna och allt fler kvinnor började arbeta utanför hemmet.
De offentliga tjänsterna började utvecklas och på så sätt skapade man den offentliga hälsovården, sociala tryggheten och grundskolan.
På 1960-talet flyttade tusentals finländare till Sverige, eftersom det fanns mer jobb och betalades högre löner i Sverige än i Finland.
När Sovjetunionen kollapsade i början av 1990-talet, hamnade Finland i ekonomisk lågkonjunktur eftersom handeln med Sovjetunionen upphörde.
Många företag gick i konkurs, vilket fick till följd att många människor förlorade sina jobb.
Efter lågkonjunkturen uppstod det mycket högteknologisk industri och högteknologiska arbetsplatser i Finland.
Allt fler människor jobbade också i olika serviceyrken.
På 1990-talet ökade inflyttningen från andra länder till Finland.
Finland fick flyktingar från många länder och hit flyttade människor med finländskt påbrå från forna Sovjetunionen.
Många flyttade till Finland även för att studera, arbeta eller för att de hade sin familj här.
År 1995 blev Finland medlem i Europeiska unionen (EU).
År 2002 införde Finland bland de första EU-länderna EU:s gemensamma valuta, euro, och gav därmed upp sin egen valuta.
Information om Finlands historiaengelska _ ryska _ franska _ spanska _ tyska _ portugisiska
Finland har alltid varit en nordlig och liten plats mellan öst och väst.
Finlands historia är en berättelse om handelsvägar, möten mellan kulturer och livet intill stora grannar.
Finlands förhistoria –1323
Finland har varit bebott sedan istiden, från cirka år 8800 före tideräkningen.
Bosättningen utvecklades först vid vattendrag och det finländska territoriet har alltid använts för livlig handelstrafik.
Namnet på Finlands äldsta stad, Åbo (Turku), betyder handelsplats.
De första skriftliga källorna om Finland är från 1100–1200-talen. Då anslöts
Finlands territorium med hjälp av korståg till påven i Roms maktkrets och det medeltida nätverket av hansaköpmän.
Den katolska kyrkan kom till Finland via Sverige och den ortodoxa kyrkan från Novgorod i öster, nuvarande Rysslands område.
Nöteborgsfreden 1323 avslutade kriget mellan Sverige och Novgorod om herraväldet i området.
Med freden etablerades den katolska tron i Finlands västra delar och den ortodoxa tron i landets östra delar.
Denna gräns mellan religionerna finns fortfarande, men med reformationen byttes den katolska tron till den lutherska.
Sveriges östra del 1323–1809
Efter Nöteborgsfreden 1323 hörde största delen av det finska territoriet till Sverige.
Under cirka 500 år var Finlands historia Sveriges historia.
Finlands område var Sveriges buffert österut och gränserna drogs om flera gånger i samband med olika krig.
Finländarna ser sig själva som västeuropéer, eftersom tiden som en del av det svenska riket knöt finländarna starkt till det västliga kulturarvet.
Till exempel stred finska soldater i Sveriges armé under Trettioåriga kriget i Mellaneuropa.
Samtidigt hade man emellertid även kontakter med handelscentra i öst och den ortodoxa kyrkan.
Viktiga händelser
1523 Gustav Vasa blev kung över Sverige och lösgjorde Sverige från den medeltida nordiska unionen.
Den första finskspråkiga ABC-boken (Aapinen) ges ut i Finland
1550 Helsingfors grundas för att konkurrera med Tallinn om handeln på Östersjön
1640 I Åbo grundas
Finlands första universitet
Finland som en del av Kejsardömet Ryssland 1809–1917
Ryssland erövrade Finlands område från Sverige 1808–1809.
De flesta lagarna från den svenska tiden fortsatte att gälla.
Under Ryssland blev Finland ett speciellt område som utvecklades på kejsarens order.
Till exempel har Helsingfors innerstad byggts under den ryska tiden.
Från 1899 och framåt tog Ryssland ett hårdare grepp om storfurstendömet Finland.
Finland deltog inte i första världskriget, men nationalismen hade inverkan även i det finska området.
Finland fick en egen lantdag 1906 och det första valet ordnades 1907.
Finland förklarade sig självständigt den 6 december 1917 och bolsjevikregeringen som tog makten i samband med oktoberrevolutionen i Ryssland erkände självständigheten den 31 december 1917.
Viktiga händelser
1812 Helsingfors blir huvudstad
Den gamla huvudstaden Åbo förstörs i en brand och Helsingfors får en allt viktigare ställning
1860 Finland inför en egen valuta, mark
1906 Allmän och lika rösträtt, även för kvinnor
Självständighetens tidiga år 1917–1945
Finlands ställning under självständighetens tidiga år var skör.
Snart efter att landet hade blivit självständigt utbröt ett blodigt inbördeskrig i Finland.
Kriget bekämpades mellan den röda arbetarrörelsen och vita regeringsstyrkor.
De vita fick stöd av Tyskland och de röda av Ryssland.
Kriget slutade med de vitas seger.
Finland var starkt knutet till Tysklands inflytandesfär, eftersom Sovjetunionen blev det största hotet mot den nationella säkerheten.
På 1930-talet var många högersinnade och högerextrema rörelser populära i Finland liksom i det övriga Europa.
I augusti 1939 avtalade Nazityskland och Sovjetunionen att Finland hör till Sovjetunionens intressesfär.
Under andra världskriget stred Finland två gånger mot Sovjetunionen på Tysklands sida.
Finland förlorade båda krigen, men Sovjetunionen ockuperade aldrig Finland.
Eftersom Finland lyckades försvara sitt territorium i krigen kort efter att landet hade blivit självständigt har krigen under 1900-talet betraktats som den tid då Finlands självständighet etablerades.
Viktiga händelser
1918 Inbördeskrig mellan röda och vita
1921 Lagen om läroplikt träder i kraft och sexårig folkskola blir obligatorisk för alla
1939–1940 blir Finland inblandat i andra världskriget när vinterkriget mellan Finland och Sovjetunionen utbryter
1941–1944 Andra världskriget fortsätter med fortsättningskriget mellan Finland och Sovjetunionen
Återuppbyggnad, industrialisering och kalla kriget 1945–1991
Finland förlorade kriget och var därför tvunget att betala ett tungt krigsskadestånd till Sovjetunionen i form av varor.
Finland finansierade tillverkningen av varorna med lån och understöd.
I och med produktionen av krigsskadeståndet utvecklades
Finland från ett jordbruksland till ett industriland.
I takt med industrialiseringen började flyttrörelsen från landsbygden till städerna.
Finland och Sovjetunionen ingick 1948 ett avtal om vänskap, samarbete och bistånd, enligt vilket staterna lovade att försvara varandra mot yttre hot.
I praktiken var Finland under hela kalla kriget en del av Sovjetunionens intressesfär och landets utrikes- och inrikespolitik styrdes av rädslan för Sovjetunionen.
Viktiga händelser
1948 VSB-avtalet mellan Finland och Sovjetunionen
1952 OS i Helsingfors
1968 Den finländska grundskoleinstitutionen inrättas
Till följd av Sovjetunionens kollaps och den ekonomiska tillväxten på 1980-talet som baserade sig på lån hamnade Finland i depression på 1990-talet.
Värst var depressionen i början av 1990-talet, då det fanns ett stort antal arbetslösa i Finland, många företag gick i konkurs och staten hade lite pengar.
Efter cirka 1995 började en ekonomisk tillväxt i Finland, varvid det viktigaste företaget var mobiltelefontillverkaren Nokia.
Finland blev medlem i EU 1995 och var ett av de första länderna som införde euro som valuta.
Viktiga händelser
1991 Den hårdaste ekonomiska krisen under
Finlands historia
1995 Finland går med i Europeiska Unionen
2000 Finland placerar sig på första plats i barns läskunnighet i den första PISA-undersökningen
Finland inför euro som kontantvaluta
2007 Nokia säljer 40 procent av alla mobiltelefoner i världen
Staten
Finland är en republik och medlem i Europeiska unionen (EU).
Finlands huvudstad är Helsingfors.
Finland är indelat i kommuner som har självstyre.
Befolkning
Finland har 5,5 miljoner invånare.
Finlands nationalspråk är finska och svenska (cirka fem procent av finländarna har svenska som modersmål).
Många finländare pratar bra engelska.
Klimat och geografi
Finland ligger i Nordeuropa.
Finlands grannländer är Ryssland (i öster), Norge (i norr), Sverige (i väster) och Estland (i söder).
Finlands areal är 338 432 km², vilken omfattar landets markområden och insjöar.
Ekonomi
Valutaenheten i Finland är euro.
Information om Finland på andra ställen på Internet
linkkiArbets- och näringsministeriet:
Guiden Välkommen till Finland(pdf, 3,40 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
Offentliga tjänster på internetfinska _ svenska _ engelska
Information om Finlandengelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ portugisiska
linkkiVisitFinland.com:
Information om Finland till turistersvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ japanska _ italienska
Staten
Finland är en republik och medlem i Europeiska unionen (EU).
Finlands huvudstad är Helsingfors.
Finland är indelat i kommuner som har självstyre.
Befolkning
Finland har 5,5 miljoner invånare.
Finlands nationalspråk är finska och svenska (cirka fem procent av finländarna har svenska som modersmål).
Många finländare pratar bra engelska.
Klimat och geografi
Finland ligger i Nordeuropa.
Finlands grannländer är Ryssland (i öster), Norge (i norr), Sverige (i väster) och Estland (i söder).
Finlands areal är 338 432 km², vilken omfattar landets markområden och insjöar.
Ekonomi
Valutaenheten i Finland är euro.
Information om Finland på andra ställen på Internet
linkkiArbets- och näringsministeriet:
Guiden Välkommen till Finland(pdf, 3,40 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
Offentliga tjänster på internetfinska _ svenska _ engelska
Information om Finlandengelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ portugisiska
linkkiVisitFinland.com:
Information om Finland till turistersvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ japanska _ italienska
Staten
Finland är en republik och medlem i Europeiska unionen (EU).
Finlands huvudstad är Helsingfors.
Finland är indelat i kommuner som har självstyre.
Befolkning
Finland har 5,5 miljoner invånare.
Finlands nationalspråk är finska och svenska (cirka fem procent av finländarna har svenska som modersmål).
Många finländare pratar bra engelska.
Klimat och geografi
Finland ligger i Nordeuropa.
Finlands grannländer är Ryssland (i öster), Norge (i norr), Sverige (i väster) och Estland (i söder).
Finlands areal är 338 432 km², vilken omfattar landets markområden och insjöar.
Ekonomi
Valutaenheten i Finland är euro.
Information om Finland på andra ställen på Internet
linkkiArbets- och näringsministeriet:
Guiden Välkommen till Finland(pdf, 3,40 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
Offentliga tjänster på internetfinska _ svenska _ engelska
Information om Finlandengelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ portugisiska
linkkiVisitFinland.com:
Information om Finland till turistersvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ japanska _ italienska
Frivilligarbete är ett bra sätt att hjälpa, lära känna nya människor och medverka i något som du tycker att är viktigt.
Frivilligarbete är inte samma sak som arbete eller praktik.
Väg in i arbetslivet
Om din arbetserfarenhet i Finland är kort eller om din finska ännu inte är så bra, kan frivilligarbete vara ett bra sätt att få fotfäste i arbetslivet och förbättra språkkunskaperna.
Frivilligarbete är oavlönat arbete, men arbetserfarenheten kan vara nyttig när du söker ett avlönat arbete.
Ta kontakt direkt med den organisation där du vill arbeta som frivillig.
Om du får utkomstskydd för arbetslösa ska du på förhand fråga din TE-byrå huruvida frivilligarbetet påverkar utbetalningen av utkomstskyddet för arbetslösa.
I vissa fall kan frivilligarbete vara en del av din integrationsplan.
En rolig hobby
Frivilligarbete kan dessutom bli en bra hobby.
Du kan själv bestämma när och hur ofta du vill vara med i verksamheten.
I frivilligarbete kan du träffa människor med samma intressen som du själv har och få nya vänner.
Du kan också utnyttja de kontakter som du skapat via frivilligarbetet i arbetslivet.
Volontärarbetefinska
linkkiRöda Korset:
Volontärarbetefinska _ svenska _ engelska
linkkiMedborgararenan:
Volontärarbeteengelska
linkkiGuide till volontärarbete:
Guide till volontärarbetefinska _ engelska
Frivilligarbete är ett bra sätt att hjälpa, lära känna nya människor och medverka i något som du tycker att är viktigt.
Frivilligarbete är inte samma sak som arbete eller praktik.
Väg in i arbetslivet
Om din arbetserfarenhet i Finland är kort eller om din finska ännu inte är så bra, kan frivilligarbete vara ett bra sätt att få fotfäste i arbetslivet och förbättra språkkunskaperna.
Frivilligarbete är oavlönat arbete, men arbetserfarenheten kan vara nyttig när du söker ett avlönat arbete.
Ta kontakt direkt med den organisation där du vill arbeta som frivillig.
Om du får utkomstskydd för arbetslösa ska du på förhand fråga din TE-byrå huruvida frivilligarbetet påverkar utbetalningen av utkomstskyddet för arbetslösa.
I vissa fall kan frivilligarbete vara en del av din integrationsplan.
En rolig hobby
Frivilligarbete kan dessutom bli en bra hobby.
Du kan själv bestämma när och hur ofta du vill vara med i verksamheten.
I frivilligarbete kan du träffa människor med samma intressen som du själv har och få nya vänner.
Du kan också utnyttja de kontakter som du skapat via frivilligarbetet i arbetslivet.
Volontärarbetefinska
linkkiRöda Korset:
Volontärarbetefinska _ svenska _ engelska
linkkiMedborgararenan:
Volontärarbeteengelska
linkkiGuide till volontärarbete:
Guide till volontärarbetefinska _ engelska
Frivilligarbete är ett bra sätt att hjälpa, lära känna nya människor och medverka i något som du tycker att är viktigt.
Frivilligarbete är inte samma sak som arbete eller praktik.
Väg in i arbetslivet
Om din arbetserfarenhet i Finland är kort eller om din finska ännu inte är så bra, kan frivilligarbete vara ett bra sätt att få fotfäste i arbetslivet och förbättra språkkunskaperna.
Frivilligarbete är oavlönat arbete, men arbetserfarenheten kan vara nyttig när du söker ett avlönat arbete.
Ta kontakt direkt med den organisation där du vill arbeta som frivillig.
Om du får utkomstskydd för arbetslösa ska du på förhand fråga din TE-byrå huruvida frivilligarbetet påverkar utbetalningen av utkomstskyddet för arbetslösa.
I vissa fall kan frivilligarbete vara en del av din integrationsplan.
En rolig hobby
Frivilligarbete kan dessutom bli en bra hobby.
Du kan själv bestämma när och hur ofta du vill vara med i verksamheten.
I frivilligarbete kan du träffa människor med samma intressen som du själv har och få nya vänner.
Du kan också utnyttja de kontakter som du skapat via frivilligarbetet i arbetslivet.
Volontärarbetefinska
linkkiRöda Korset:
Volontärarbetefinska _ svenska _ engelska
linkkiMedborgararenan:
Volontärarbeteengelska
linkkiGuide till volontärarbete:
Guide till volontärarbetefinska _ engelska
I Finland finns det många föreningar sett till befolkningens storlek.
Enligt lagen har alla rätt att verka i föreningar.
Föreningsfriheten gäller också utlänningar.
En förening kan till exempel vara ett idrottssällskap, en kulturförening, en vänskapsförening eller en religiös förening.
Registrerade föreningar är ideella föreningar.
En förening bör inte grundas i syfte att idka en näring.
I Finland finns också många föreningar som grundats av invandrare.
En invandrarförening eller det egna landets vänskapsförening kan hjälpa till att bevara och utveckla den egna kulturen i det nya samhället och samarbeta med myndigheter och andra organisationer.
Du kan söka olika föreningar i patent- och registerstyrelsens tjänst Föreningsregistret.
linkkiPatent- och registerstyrelsen:
Föreningsnätetfinska _ svenska _ engelska
linkkiFinlands Flyktinghjälp:
Organisationssmedjanfinska _ svenska _ engelska
Riksomfattande föreningar för invandrare
linkkiMoniheli:
linkkiIESAF:
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
linkkiFaro:
Takorganisation för somaliska föreningarfinska _ engelska _ somaliska
linkkiAFAES:
Motionsföreningfinska _ engelska
linkkiVänskapsföreningarnas samfund:
Vänskapsföreningarfinska
Att grunda en förening
Grundandet av en förening sker i praktiken i tre steg:
beslut om att grunda en förening
upprättande av stadgar
registrering av föreningen.
Registrering av föreningen
Det lönar sig att registrera sin förening.
Då är föreningen en juridisk person vars medlemmar inte personligen bär ansvar för föreningens verksamhet.
En registrerad förening kan ansöka om finansiering och bidrag samt samarbeta med andra föreningar och myndigheter.
Föreningen registreras med anmälan till Patent- och registerstyrelsen.
linkkiPatent- och registerstryrelsen:
Föreningsregisterfinska _ svenska _ engelska
Att grunda en förening när stiftarna är utlänningar
Också utlänningar, d.v.s. personer som inte har finskt medborgarskap, kan grunda en registrerad förening.
I detta fall ska både ordföranden och vice ordföranden ha sin hemort i Finland.
Om ordföranden eller vice ordföranden har sin hemort utomlands kan föreningen ansöka om dispens hos patent- och registerstyrelsen.
Föreningens verksamhet
Föreningar bedriver sin verksamhet vanligen ett år i taget.
De planerar sin verksamhet och sin ekonomi ett år fram i tiden.
Ekonomin och bokföringen ska granskas i slutet av perioden.
I en förening är det medlemmarna som har makten.
De viktigaste besluten fattas på föreningsmöten som är öppna för alla medlemmar.
linkkiUndervisnings- och kulturministeriet:
Bidrag och priserfinska _ svenska _ engelska
Föreningens styrelse
För föreningen väljs en styrelse på föreningsmötet dit alla föreningsmedlemmar sammankallas.
Styrelsen ska bestå av minst ordföranden och två medlemmar.
Styrelsens storlek kan föreskrivas i stadgarna.
Styrelsen har som uppgift att sköta ärenden enligt lagar, föreningens stadgar och föreningens beslut.
Upplösning av föreningen
Föreningen upplöses när merparten av medlemmarna fattar beslut om detta på föreningens möte.
När beslutet om upplösning har fattats och tillgångarna överlåtits görs en anmälan om upplösning av föreningen till registerstyrelsen.
I Finland finns det många föreningar sett till befolkningens storlek.
Enligt lagen har alla rätt att verka i föreningar.
Föreningsfriheten gäller också utlänningar.
En förening kan till exempel vara ett idrottssällskap, en kulturförening, en vänskapsförening eller en religiös förening.
Registrerade föreningar är ideella föreningar.
En förening bör inte grundas i syfte att idka en näring.
I Finland finns också många föreningar som grundats av invandrare.
En invandrarförening eller det egna landets vänskapsförening kan hjälpa till att bevara och utveckla den egna kulturen i det nya samhället och samarbeta med myndigheter och andra organisationer.
Du kan söka olika föreningar i patent- och registerstyrelsens tjänst Föreningsregistret.
linkkiPatent- och registerstyrelsen:
Föreningsnätetfinska _ svenska _ engelska
linkkiFinlands Flyktinghjälp:
Organisationssmedjanfinska _ svenska _ engelska
Riksomfattande föreningar för invandrare
linkkiMoniheli:
linkkiIESAF:
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
linkkiFaro:
Takorganisation för somaliska föreningarfinska _ engelska _ somaliska
linkkiAFAES:
Motionsföreningfinska _ engelska
linkkiVänskapsföreningarnas samfund:
Vänskapsföreningarfinska
Att grunda en förening
Grundandet av en förening sker i praktiken i tre steg:
beslut om att grunda en förening
upprättande av stadgar
registrering av föreningen.
Registrering av föreningen
Det lönar sig att registrera sin förening.
Då är föreningen en juridisk person vars medlemmar inte personligen bär ansvar för föreningens verksamhet.
En registrerad förening kan ansöka om finansiering och bidrag samt samarbeta med andra föreningar och myndigheter.
Föreningen registreras med anmälan till Patent- och registerstyrelsen.
linkkiPatent- och registerstryrelsen:
Föreningsregisterfinska _ svenska _ engelska
Att grunda en förening när stiftarna är utlänningar
Också utlänningar, d.v.s. personer som inte har finskt medborgarskap, kan grunda en registrerad förening.
I detta fall ska både ordföranden och vice ordföranden ha sin hemort i Finland.
Om ordföranden eller vice ordföranden har sin hemort utomlands kan föreningen ansöka om dispens hos patent- och registerstyrelsen.
Föreningens verksamhet
Föreningar bedriver sin verksamhet vanligen ett år i taget.
De planerar sin verksamhet och sin ekonomi ett år fram i tiden.
Ekonomin och bokföringen ska granskas i slutet av perioden.
I en förening är det medlemmarna som har makten.
De viktigaste besluten fattas på föreningsmöten som är öppna för alla medlemmar.
linkkiUndervisnings- och kulturministeriet:
Bidrag och priserfinska _ svenska _ engelska
Föreningens styrelse
För föreningen väljs en styrelse på föreningsmötet dit alla föreningsmedlemmar sammankallas.
Styrelsen ska bestå av minst ordföranden och två medlemmar.
Styrelsens storlek kan föreskrivas i stadgarna.
Styrelsen har som uppgift att sköta ärenden enligt lagar, föreningens stadgar och föreningens beslut.
Upplösning av föreningen
Föreningen upplöses när merparten av medlemmarna fattar beslut om detta på föreningens möte.
När beslutet om upplösning har fattats och tillgångarna överlåtits görs en anmälan om upplösning av föreningen till registerstyrelsen.
I Finland finns det många föreningar sett till befolkningens storlek.
Enligt lagen har alla rätt att verka i föreningar.
Föreningsfriheten gäller också utlänningar.
En förening kan till exempel vara ett idrottssällskap, en kulturförening, en vänskapsförening eller en religiös förening.
Registrerade föreningar är ideella föreningar.
En förening bör inte grundas i syfte att idka en näring.
I Finland finns också många föreningar som grundats av invandrare.
En invandrarförening eller det egna landets vänskapsförening kan hjälpa till att bevara och utveckla den egna kulturen i det nya samhället och samarbeta med myndigheter och andra organisationer.
Du kan söka olika föreningar i patent- och registerstyrelsens tjänst Föreningsregistret.
linkkiPatent- och registerstyrelsen:
Föreningsnätetfinska _ svenska _ engelska
linkkiFinlands Flyktinghjälp:
Riksomfattande föreningar för invandrare
linkkiMoniheli:
linkkiIESAF:
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
linkkiFaro:
Takorganisation för somaliska föreningarfinska _ engelska _ somaliska
linkkiAFAES:
Motionsföreningfinska
linkkiVänskapsföreningarnas samfund:
Vänskapsföreningarfinska
Att grunda en förening
Grundandet av en förening sker i praktiken i tre steg:
beslut om att grunda en förening
upprättande av stadgar
registrering av föreningen.
Registrering av föreningen
Det lönar sig att registrera sin förening.
Då är föreningen en juridisk person vars medlemmar inte personligen bär ansvar för föreningens verksamhet.
En registrerad förening kan ansöka om finansiering och bidrag samt samarbeta med andra föreningar och myndigheter.
Föreningen registreras med anmälan till Patent- och registerstyrelsen.
linkkiPatent- och registerstryrelsen:
Föreningsregisterfinska _ svenska _ engelska
Att grunda en förening när stiftarna är utlänningar
Också utlänningar, d.v.s. personer som inte har finskt medborgarskap, kan grunda en registrerad förening.
I detta fall ska både ordföranden och vice ordföranden ha sin hemort i Finland.
Om ordföranden eller vice ordföranden har sin hemort utomlands kan föreningen ansöka om dispens hos patent- och registerstyrelsen.
Föreningens verksamhet
Föreningar bedriver sin verksamhet vanligen ett år i taget.
De planerar sin verksamhet och sin ekonomi ett år fram i tiden.
Ekonomin och bokföringen ska granskas i slutet av perioden.
I en förening är det medlemmarna som har makten.
De viktigaste besluten fattas på föreningsmöten som är öppna för alla medlemmar.
linkkiUndervisnings- och kulturministeriet:
Bidrag och priserfinska _ svenska _ engelska
Föreningens styrelse
För föreningen väljs en styrelse på föreningsmötet dit alla föreningsmedlemmar sammankallas.
Styrelsen ska bestå av minst ordföranden och två medlemmar.
Styrelsens storlek kan föreskrivas i stadgarna.
Styrelsen har som uppgift att sköta ärenden enligt lagar, föreningens stadgar och föreningens beslut.
Upplösning av föreningen
Föreningen upplöses när merparten av medlemmarna fattar beslut om detta på föreningens möte.
När beslutet om upplösning har fattats och tillgångarna överlåtits görs en anmälan om upplösning av föreningen till registerstyrelsen.
I Finland finns ett rikt hobbyutbud för barn och unga.
Barn och ungdomar kan till exempel ha idrott, dans, musik, bildkonst eller teater som hobby.
En del fritidsaktiviteter är avgiftsbelagda men det finns också tillgång till gratis aktiviteter.
Också kommunerna ordnar aktiviteter för barn och unga.
Barn och motion
Små barn behöver inte nödvändigtvis ledd motion, utan det räcker med vanlig lekverksamhet och utevistelser i olika miljöer.
Det skulle ändå vara bra att se till att små barn får så mångsidig motion som möjligt, eftersom motion utvecklar barnets motoriska färdigheter och är bra för hälsan.
Daghemmet står ofta för en del av motionen eftersom man där ordnar rörelselekar.
Dessutom ordnar även idrottsklubbar motion för små barn.
Daghem och skolor gör sitt för att ordna motion men detta är inte deras huvudsakliga uppgift.
Barn får inte tillräckligt med motion bara genom att delta i gymnastiklektionerna..
Därför skulle det vara bra att barnen hade möjlighet att röra på sig tillräckligt också utanför daghemmet eller skoltiden.
Sport och motion
Mer information om sport som hobby hittar du på InfoFinlands sida Motion.
Bästa stället att fråga om enskilda grenar och var man kan utöva dem är grenförbunden.
Konsthobbyer
Utöver sport har ungdomar också tillgång till många konstaktiviteter, som till exempel bildkonst, musik eller teater.
Dessa finns till exempel på arbetarinstitut, bildkonstskolor, musikskolor och kommunernas ungdomsväsende.
Fråga mer om hobbymöjligheterna, tidtabellerna och priserna direkt hos arrangören.
Ungdomsarbete
Tjänsterna inom kommunernas ungdomsarbete är avsedda för barn och unga vuxna.
De vanligaste tjänsterna är olika klubbar och den öppna verksamheten som pågår på ungdomsgårdarna.
Tjänsterna kan variera något i olika delar av landet.
Mer information om den kommunala ungdomsverksamheten får du hos ungdomsväsendet i din hemkommun.
Många organisationer och församlingar bedriver också ungdomsarbete.
Ungdomsgården är en plats där de unga kan vistas och utöva olika hobbyer.
På ungdomsgårdarna ordnas också ledd verksamhet.
Största delen av verksamheten på ungdomsgårdarna är gratis.
Verksamheten utformas enligt ungdomarnas önskemål och de unga kan själva påverka innehållet i verksamheten.
På ungdomsgården finns alltid någon vuxen, vanligen kommunens ungdomsarbetare eller ungdomsledare.
Åldersgränsen på ungdomsgårdarna varierar.
Ungdomar och påverkan
Ungdomarna har många möjligheter att påverka.
Ett lätt sätt att komma igång är till exempel genom att delta i skolans eller läroanstaltens elevverksamhet.
Deltagande i elev- och föreningsverksamhet är ett bra sätt att bidra till att också de unga får sin röst hör då det fattas beslut om sådant som påverkar deras livsmiljö.
I dag finns det många medborgarorganisationer som specialiserat sig på att främja en viss samhällelig fråga.
Många medborgarorganisationer och föreningar har särskilda ungdomsavdelningar som ordnar verksamhet för unga.
Dessutom finns det speciella organisationer för ungdomar, yngre tonåringar och studerande.
I Finland finns ett rikt hobbyutbud för barn och unga.
Barn och ungdomar kan till exempel ha idrott, dans, musik, bildkonst eller teater som hobby.
En del fritidsaktiviteter är avgiftsbelagda men det finns också tillgång till gratis aktiviteter.
Också kommunerna ordnar aktiviteter för barn och unga.
Barn och motion
Små barn behöver inte nödvändigtvis ledd motion, utan det räcker med vanlig lekverksamhet och utevistelser i olika miljöer.
Det skulle ändå vara bra att se till att små barn får så mångsidig motion som möjligt, eftersom motion utvecklar barnets motoriska färdigheter och är bra för hälsan.
Daghemmet står ofta för en del av motionen eftersom man där ordnar rörelselekar.
Dessutom ordnar även idrottsklubbar motion för små barn.
Daghem och skolor gör sitt för att ordna motion men detta är inte deras huvudsakliga uppgift.
Barn får inte tillräckligt med motion bara genom att delta i gymnastiklektionerna..
Därför skulle det vara bra att barnen hade möjlighet att röra på sig tillräckligt också utanför daghemmet eller skoltiden.
Sport och motion
Mer information om sport som hobby hittar du på InfoFinlands sida Motion.
Bästa stället att fråga om enskilda grenar och var man kan utöva dem är grenförbunden.
Konsthobbyer
Utöver sport har ungdomar också tillgång till många konstaktiviteter, som till exempel bildkonst, musik eller teater.
Dessa finns till exempel på arbetarinstitut, bildkonstskolor, musikskolor och kommunernas ungdomsväsende.
Fråga mer om hobbymöjligheterna, tidtabellerna och priserna direkt hos arrangören.
Ungdomsarbete
Tjänsterna inom kommunernas ungdomsarbete är avsedda för barn och unga vuxna.
De vanligaste tjänsterna är olika klubbar och den öppna verksamheten som pågår på ungdomsgårdarna.
Tjänsterna kan variera något i olika delar av landet.
Mer information om den kommunala ungdomsverksamheten får du hos ungdomsväsendet i din hemkommun.
Många organisationer och församlingar bedriver också ungdomsarbete.
Ungdomsgården är en plats där de unga kan vistas och utöva olika hobbyer.
På ungdomsgårdarna ordnas också ledd verksamhet.
Största delen av verksamheten på ungdomsgårdarna är gratis.
Verksamheten utformas enligt ungdomarnas önskemål och de unga kan själva påverka innehållet i verksamheten.
På ungdomsgården finns alltid någon vuxen, vanligen kommunens ungdomsarbetare eller ungdomsledare.
Åldersgränsen på ungdomsgårdarna varierar.
Ungdomar och påverkan
Ungdomarna har många möjligheter att påverka.
Ett lätt sätt att komma igång är till exempel genom att delta i skolans eller läroanstaltens elevverksamhet.
Deltagande i elev- och föreningsverksamhet är ett bra sätt att bidra till att också de unga får sin röst hör då det fattas beslut om sådant som påverkar deras livsmiljö.
I dag finns det många medborgarorganisationer som specialiserat sig på att främja en viss samhällelig fråga.
Många medborgarorganisationer och föreningar har särskilda ungdomsavdelningar som ordnar verksamhet för unga.
Dessutom finns det speciella organisationer för ungdomar, yngre tonåringar och studerande.
I Finland finns ett rikt hobbyutbud för barn och unga.
Barn och ungdomar kan till exempel ha idrott, dans, musik, bildkonst eller teater som hobby.
En del fritidsaktiviteter är avgiftsbelagda men det finns också tillgång till gratis aktiviteter.
Också kommunerna ordnar aktiviteter för barn och unga.
Barn och motion
Små barn behöver inte nödvändigtvis ledd motion, utan det räcker med vanlig lekverksamhet och utevistelser i olika miljöer.
Det skulle ändå vara bra att se till att små barn får så mångsidig motion som möjligt, eftersom motion utvecklar barnets motoriska färdigheter och är bra för hälsan.
Daghemmet står ofta för en del av motionen eftersom man där ordnar rörelselekar.
Dessutom ordnar även idrottsklubbar motion för små barn.
Daghem och skolor gör sitt för att ordna motion men detta är inte deras huvudsakliga uppgift.
Barn får inte tillräckligt med motion bara genom att delta i gymnastiklektionerna..
Därför skulle det vara bra att barnen hade möjlighet att röra på sig tillräckligt också utanför daghemmet eller skoltiden.
Sport och motion
Mer information om sport som hobby hittar du på InfoFinlands sida Motion.
Bästa stället att fråga om enskilda grenar och var man kan utöva dem är grenförbunden.
Konsthobbyer
Utöver sport har ungdomar också tillgång till många konstaktiviteter, som till exempel bildkonst, musik eller teater.
Dessa finns till exempel på arbetarinstitut, bildkonstskolor, musikskolor och kommunernas ungdomsväsende.
Fråga mer om hobbymöjligheterna, tidtabellerna och priserna direkt hos arrangören.
Ungdomsarbete
Tjänsterna inom kommunernas ungdomsarbete är avsedda för barn och unga vuxna.
De vanligaste tjänsterna är olika klubbar och den öppna verksamheten som pågår på ungdomsgårdarna.
Tjänsterna kan variera något i olika delar av landet.
Mer information om den kommunala ungdomsverksamheten får du hos ungdomsväsendet i din hemkommun.
Många organisationer och församlingar bedriver också ungdomsarbete.
Ungdomsgården är en plats där de unga kan vistas och utöva olika hobbyer.
På ungdomsgårdarna ordnas också ledd verksamhet.
Största delen av verksamheten på ungdomsgårdarna är gratis.
Verksamheten utformas enligt ungdomarnas önskemål och de unga kan själva påverka innehållet i verksamheten.
På ungdomsgården finns alltid någon vuxen, vanligen kommunens ungdomsarbetare eller ungdomsledare.
Åldersgränsen på ungdomsgårdarna varierar.
Ungdomar och påverkan
Ungdomarna har många möjligheter att påverka.
Ett lätt sätt att komma igång är till exempel genom att delta i skolans eller läroanstaltens elevverksamhet.
Deltagande i elev- och föreningsverksamhet är ett bra sätt att bidra till att också de unga får sin röst hör då det fattas beslut om sådant som påverkar deras livsmiljö.
I dag finns det många medborgarorganisationer som specialiserat sig på att främja en viss samhällelig fråga.
Många medborgarorganisationer och föreningar har särskilda ungdomsavdelningar som ordnar verksamhet för unga.
Dessutom finns det speciella organisationer för ungdomar, yngre tonåringar och studerande.
I Finland finns många möjligheter att syssla med musik.
Du kan lära dig att spela ett instrument, sjunga i kör, gå på konserter och festivaler eller till och med sjunga karaoke.
Möjligheter till musikhobbyer finns för såväl vuxna som unga och barn.
På många orter finns medborgarinstitut, som kommunerna upprätthåller.
Medborgarinstituten ordnar förmånlig musikundervisning.
Dessutom erbjuder även privata musikskolor och -institut undervisning.
Medborgarinstitutens musikgrupper är öppna för alla.
Elever antas till undervisningen vanligtvis i anmälningsordning till hösten och våren.
Till musikskolorna ansöker man medelst inträdesprov en gång per år.
Mer information om möjligheter till musikhobby får du via kommunens kulturkontor.
Medborgarinstitut i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Information om körerfinska _ engelska
Konserter och festivaler
Konserter ordnas på olika platser: I konsertsalar, musikhus, kulturcenter, institut, restauranger, på historiska platser och i kyrkor.
En del konserter är avgiftsfria, men vanligtvis har konserter en inträdesavgift.
Mer information om konserter hittar du i lokala tidningar och på internet.
Musikfestivaler är populära, särskilt på sommaren.
Festivalerna ordnas på olika håll i Finland, både i städerna och på landsbygden.
Vanligtvis måste man betala en inträdesavgift till festivaler.
Festivaler i Finlandfinska _ svenska _ engelska _ ryska _ franska _ kinesiska _ tyska _ japanska
linkkiCentralen för främjande av Folkmusik och Folkdans :
Folkmusik och -dans i Finlandfinska _ svenska _ engelska
I Finland finns många möjligheter att syssla med musik.
Du kan lära dig att spela ett instrument, sjunga i kör, gå på konserter och festivaler eller till och med sjunga karaoke.
Möjligheter till musikhobbyer finns för såväl vuxna som unga och barn.
På många orter finns medborgarinstitut, som kommunerna upprätthåller.
Medborgarinstituten ordnar förmånlig musikundervisning.
Dessutom erbjuder även privata musikskolor och -institut undervisning.
Medborgarinstitutens musikgrupper är öppna för alla.
Elever antas till undervisningen vanligtvis i anmälningsordning till hösten och våren.
Till musikskolorna ansöker man medelst inträdesprov en gång per år.
Mer information om möjligheter till musikhobby får du via kommunens kulturkontor.
Medborgarinstitut i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Information om körerfinska _ engelska
Konserter och festivaler
Konserter ordnas på olika platser: I konsertsalar, musikhus, kulturcenter, institut, restauranger, på historiska platser och i kyrkor.
En del konserter är avgiftsfria, men vanligtvis har konserter en inträdesavgift.
Mer information om konserter hittar du i lokala tidningar och på internet.
Musikfestivaler är populära, särskilt på sommaren.
Festivalerna ordnas på olika håll i Finland, både i städerna och på landsbygden.
Vanligtvis måste man betala en inträdesavgift till festivaler.
Festivaler i Finlandfinska _ svenska _ engelska _ ryska _ franska _ kinesiska _ tyska _ japanska
linkkiCentralen för främjande av Folkmusik och Folkdans :
Folkmusik och -dans i Finlandfinska _ svenska _ engelska
I Finland finns många möjligheter att syssla med musik.
Du kan lära dig att spela ett instrument, sjunga i kör, gå på konserter och festivaler eller till och med sjunga karaoke.
Möjligheter till musikhobbyer finns för såväl vuxna som unga och barn.
På många orter finns medborgarinstitut, som kommunerna upprätthåller.
Medborgarinstituten ordnar förmånlig musikundervisning.
Dessutom erbjuder även privata musikskolor och -institut undervisning.
Medborgarinstitutens musikgrupper är öppna för alla.
Elever antas till undervisningen vanligtvis i anmälningsordning till hösten och våren.
Till musikskolorna ansöker man medelst inträdesprov en gång per år.
Mer information om möjligheter till musikhobby får du via kommunens kulturkontor.
Medborgarinstitut i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Information om körerfinska _ engelska
Konserter och festivaler
Konserter ordnas på olika platser: I konsertsalar, musikhus, kulturcenter, institut, restauranger, på historiska platser och i kyrkor.
En del konserter är avgiftsfria, men vanligtvis har konserter en inträdesavgift.
Mer information om konserter hittar du i lokala tidningar och på internet.
Musikfestivaler är populära, särskilt på sommaren.
Festivalerna ordnas på olika håll i Finland, både i städerna och på landsbygden.
Vanligtvis måste man betala en inträdesavgift till festivaler.
Festivaler i Finlandfinska _ svenska _ engelska _ ryska _ franska _ kinesiska _ tyska _ japanska
linkkiCentralen för främjande av Folkmusik och Folkdans :
Folkmusik och -dans i Finlandfinska _ svenska _ engelska
I Finlands finns ungefär ett tusen museer, varav cirka 300 är regelbundet öppna för allmänheten.
De övriga är hembygdsmuseer som vanligen bara har öppet sommartid.
Museerna är avsedda för alla.
De presenterar konst, historia, natur, någon person eller ett specialområde.
Med friluftsmuseum avses ett större museiområde med hela byggnader.
Ett friluftsmuseum kan till exempel vara en traditionell finländsk bondgård eller något annat område som gjorts om till ett museum.
Kända finska friluftsmuseer är till exempel Fölisön i Helsingfors och hantverksmuseet på Klosterbacken i Åbo.
Finsk konst presenteras till exempel i Ateneum som hör till Nationalgalleriet och Esbo moderna konstmuseum (EMMA). Med
Finlands kulturhistoria kan du bekanta dig med bland annat i Finlands nationalmuseum som ligger i Helsingfors.
Utöver detta finns det många museer och museiområden runt omkring i Finland.
Vissa museers samlingar kan du även bekanta dig med på internet.
Mer information om museer och aktuella utställningar får du på webbplatsen museot.fi.
På museerna ordnas ofta också guidade rundvandringar på olika språk.
Museisökningfinska _ svenska _ engelska
Utställningskalenderfinska _ svenska _ engelska
Unescos världsarv
I Finland finns sju Unescos världsarv.
Dessa är Sveaborg, Gamla Raumo, Petäjävesi gamla kyrka, Verla träsliperi och pappfabrik, Sammallahdenmäki fornlämningsområde, Struves kedja och Kvarkens skärgård.
Du hittar mer information om världsarven på Museiverkets webbplats.
Slott
I Finland finns också slott som är öppna för allmänheten, till exempel Olofsborg, Åbo slott och Tavastehus slott.
De är populära turistmål speciellt på sommaren.
I slotten ordnas också guidade rundvandringar där slottets historia och arkitektur presenteras.
Du hittar mer information om slotten och de guidade rundvandringarna på Museiverkets webbplats.
Inträdesavgifter och rabatter
Inträdesavgifterna till museerna varierar.
Inträdet kostar i snitt fem euro för vuxna och två euro för barn.
Många museer ger rabatt på inträdesavgiften till vissa grupper.
Sådana grupper kan till exempel vara besökare under 18 år, studerande, arbetslösa och pensionärer.
Barn kan ha fritt inträde till vissa museer.
Många museer ordnar speciella dagar då alla besökare har fritt inträde.
På museiförbundets sidor hittar du mer information om dagar med fritt inträde.
Många museer har fritt inträde på den internationella museidagen 18.5.
Några museer, som till exempel Helsingfors stadsmuseum, har alltid fritt inträde.
linkkiMuseiverket:
Unescos världsarv i Finlandfinska _ svenska _ engelska
linkkiMuseiverket:
Museer och slottfinska _ svenska _ engelska
I Finlands finns ungefär ett tusen museer, varav cirka 300 är regelbundet öppna för allmänheten.
De övriga är hembygdsmuseer som vanligen bara har öppet sommartid.
Museerna är avsedda för alla.
De presenterar konst, historia, natur, någon person eller ett specialområde.
Med friluftsmuseum avses ett större museiområde med hela byggnader.
Ett friluftsmuseum kan till exempel vara en traditionell finländsk bondgård eller något annat område som gjorts om till ett museum.
Kända finska friluftsmuseer är till exempel Fölisön i Helsingfors och hantverksmuseet på Klosterbacken i Åbo.
Finsk konst presenteras till exempel i Ateneum som hör till Nationalgalleriet och Esbo moderna konstmuseum (EMMA). Med
Finlands kulturhistoria kan du bekanta dig med bland annat i Finlands nationalmuseum som ligger i Helsingfors.
Utöver detta finns det många museer och museiområden runt omkring i Finland.
Vissa museers samlingar kan du även bekanta dig med på internet.
Mer information om museer och aktuella utställningar får du på webbplatsen museot.fi.
På museerna ordnas ofta också guidade rundvandringar på olika språk.
Museisökningfinska _ svenska _ engelska
Utställningskalenderfinska _ svenska _ engelska
Unescos världsarv
I Finland finns sju Unescos världsarv.
Dessa är Sveaborg, Gamla Raumo, Petäjävesi gamla kyrka, Verla träsliperi och pappfabrik, Sammallahdenmäki fornlämningsområde, Struves kedja och Kvarkens skärgård.
Du hittar mer information om världsarven på Museiverkets webbplats.
Slott
I Finland finns också slott som är öppna för allmänheten, till exempel Olofsborg, Åbo slott och Tavastehus slott.
De är populära turistmål speciellt på sommaren.
I slotten ordnas också guidade rundvandringar där slottets historia och arkitektur presenteras.
Du hittar mer information om slotten och de guidade rundvandringarna på Museiverkets webbplats.
Inträdesavgifter och rabatter
Inträdesavgifterna till museerna varierar.
Inträdet kostar i snitt fem euro för vuxna och två euro för barn.
Många museer ger rabatt på inträdesavgiften till vissa grupper.
Sådana grupper kan till exempel vara besökare under 18 år, studerande, arbetslösa och pensionärer.
Barn kan ha fritt inträde till vissa museer.
Många museer ordnar speciella dagar då alla besökare har fritt inträde.
På museiförbundets sidor hittar du mer information om dagar med fritt inträde.
Många museer har fritt inträde på den internationella museidagen 18.5.
Några museer, som till exempel Helsingfors stadsmuseum, har alltid fritt inträde.
linkkiMuseiverket:
Unescos världsarv i Finlandfinska _ svenska _ engelska
linkkiMuseiverket:
Museer och slottfinska _ svenska _ engelska
I Finlands finns ungefär ett tusen museer, varav cirka 300 är regelbundet öppna för allmänheten.
De övriga är hembygdsmuseer som vanligen bara har öppet sommartid.
Museerna är avsedda för alla.
De presenterar konst, historia, natur, någon person eller ett specialområde.
Med friluftsmuseum avses ett större museiområde med hela byggnader.
Ett friluftsmuseum kan till exempel vara en traditionell finländsk bondgård eller något annat område som gjorts om till ett museum.
Kända finska friluftsmuseer är till exempel Fölisön i Helsingfors och hantverksmuseet på Klosterbacken i Åbo.
Finsk konst presenteras till exempel i Ateneum som hör till Nationalgalleriet och Esbo moderna konstmuseum (EMMA). Med
Finlands kulturhistoria kan du bekanta dig med bland annat i Finlands nationalmuseum som ligger i Helsingfors.
Utöver detta finns det många museer och museiområden runt omkring i Finland.
Vissa museers samlingar kan du även bekanta dig med på internet.
Mer information om museer och aktuella utställningar får du på webbplatsen museot.fi.
På museerna ordnas ofta också guidade rundvandringar på olika språk.
Museisökningfinska _ svenska _ engelska
Utställningskalenderfinska _ svenska _ engelska
Unescos världsarv
I Finland finns sju Unescos världsarv.
Dessa är Sveaborg, Gamla Raumo, Petäjävesi gamla kyrka, Verla träsliperi och pappfabrik, Sammallahdenmäki fornlämningsområde, Struves kedja och Kvarkens skärgård.
Du hittar mer information om världsarven på Museiverkets webbplats.
Slott
I Finland finns också slott som är öppna för allmänheten, till exempel Olofsborg, Åbo slott och Tavastehus slott.
De är populära turistmål speciellt på sommaren.
I slotten ordnas också guidade rundvandringar där slottets historia och arkitektur presenteras.
Du hittar mer information om slotten och de guidade rundvandringarna på Museiverkets webbplats.
Inträdesavgifter och rabatter
Inträdesavgifterna till museerna varierar.
Inträdet kostar i snitt fem euro för vuxna och två euro för barn.
Många museer ger rabatt på inträdesavgiften till vissa grupper.
Sådana grupper kan till exempel vara besökare under 18 år, studerande, arbetslösa och pensionärer.
Barn kan ha fritt inträde till vissa museer.
Många museer ordnar speciella dagar då alla besökare har fritt inträde.
På museiförbundets sidor hittar du mer information om dagar med fritt inträde.
Många museer har fritt inträde på den internationella museidagen 18.5.
Några museer, som till exempel Helsingfors stadsmuseum, har alltid fritt inträde.
linkkiMuseiverket:
Unescos världsarv i Finlandfinska _ svenska _ engelska
linkkiMuseiverket:
Museer och slottfinska _ svenska _ engelska
Teater
De flesta städer i Finland har minst en teater.
En del teatrar är professionella, andra är amatörteatrar.
På webbplatsen för Informationscentralen för teater i Finland kan du söka teatrar på olika orter på finska.
Centralen har också ett arkiv där du kan låna översättningar av finska pjäser på olika språk.
Du kan söka information om teatrarnas repertoar och tillgängligheten av biljetter och biljettpriserna till exempel på biljettjänstens eller teatrarnas webbplatser.
I Finland ordnas också många teaterfestivaler.
Information om dessa hittar du på webbplatserna för Informationscentralen för teater i Finland på finska, svenska och på engelska.
linkkiInformationscentralen för teater i Finland:
Kontaktuppgifter till teatrarfinska
linkkiTeaterinfo Finland:
Teaterfestivalerfinska _ svenska _ engelska
Film
I de flesta städer finns en biograf.
Enklast hittar du information om biograferna i ditt område, bioprogrammet och biljettpriserna på internet.
Veckans bioprogram publiceras ofta också i lokaltidningen.
Finnkino är den största biografkedjan i Finland.
På Finnkinos webbplats kan du söka biografer enligt stad på engelska och finska och se vilka filmer som visas.
Om bioprogrammet på andra biografer kan du fråga direkt på biografen eller söka information på internet och i tidningar.
Biobiljetternas priser varierar något i Finland.
Som billigast kostar biljetten ungefär fem euro, som dyrast över tio euro.
Du kan ta reda på biljettpriset på förhand på biografens webbplats.
I Finland visas filmerna oftast på originalspråket.
Dessutom är de textade till finska och svenska.
Barnfilmerna är ett undantag. De kan vara dubbade till finska även om filmens originalspråk är något annat.
Biografer
Nationella audiovisuella arkivet visar nya och gamla filmer från hela världen.
Information om visningarna finns på finska på arkivets webbplats.
Visningar ordnas på flera orter.
Filmer på främmande språk har vanligen finsk- och svenskspråkig textning.
Filmfestivaler
I Finland ordnas årligen högklassiga filmfestivaler, varav de bäst kända är Kärlek och anarki-festivalen, som ordnas varje höst i Helsingfors, och Sodankylä filmfestival som ordnas på sommaren.
linkkiFinnkino:
Filmerfinska _ engelska
linkkiKärlek och anarki:
Filmfestivalfinska _ svenska _ engelska
Filmfestivalfinska _ engelska
Information om filmer och filmvisningarfinska _ svenska _ engelska
Teater
De flesta städer i Finland har minst en teater.
En del teatrar är professionella, andra är amatörteatrar.
På webbplatsen för Informationscentralen för teater i Finland kan du söka teatrar på olika orter på finska.
Centralen har också ett arkiv där du kan låna översättningar av finska pjäser på olika språk.
Du kan söka information om teatrarnas repertoar och tillgängligheten av biljetter och biljettpriserna till exempel på biljettjänstens eller teatrarnas webbplatser.
I Finland ordnas också många teaterfestivaler.
Information om dessa hittar du på webbplatserna för Informationscentralen för teater i Finland på finska, svenska och på engelska.
linkkiInformationscentralen för teater i Finland:
Kontaktuppgifter till teatrarfinska
linkkiTeaterinfo Finland:
Teaterfestivalerfinska _ svenska _ engelska
Film
I de flesta städer finns en biograf.
Enklast hittar du information om biograferna i ditt område, bioprogrammet och biljettpriserna på internet.
Veckans bioprogram publiceras ofta också i lokaltidningen.
Finnkino är den största biografkedjan i Finland.
På Finnkinos webbplats kan du söka biografer enligt stad på engelska och finska och se vilka filmer som visas.
Om bioprogrammet på andra biografer kan du fråga direkt på biografen eller söka information på internet och i tidningar.
Biobiljetternas priser varierar något i Finland.
Som billigast kostar biljetten ungefär fem euro, som dyrast över tio euro.
Du kan ta reda på biljettpriset på förhand på biografens webbplats.
I Finland visas filmerna oftast på originalspråket.
Dessutom är de textade till finska och svenska.
Barnfilmerna är ett undantag. De kan vara dubbade till finska även om filmens originalspråk är något annat.
Biografer
Nationella audiovisuella arkivet visar nya och gamla filmer från hela världen.
Information om visningarna finns på finska på arkivets webbplats.
Visningar ordnas på flera orter.
Filmer på främmande språk har vanligen finsk- och svenskspråkig textning.
Filmfestivaler
I Finland ordnas årligen högklassiga filmfestivaler, varav de bäst kända är Kärlek och anarki-festivalen, som ordnas varje höst i Helsingfors, och Sodankylä filmfestival som ordnas på sommaren.
linkkiFinnkino:
Filmerfinska _ engelska
linkkiKärlek och anarki:
Filmfestivalfinska _ svenska _ engelska
Filmfestivalfinska _ engelska
Information om filmer och filmvisningarfinska _ svenska _ engelska
Teater
De flesta städer i Finland har minst en teater.
En del teatrar är professionella, andra är amatörteatrar.
På webbplatsen för Informationscentralen för teater i Finland kan du söka teatrar på olika orter på finska.
Centralen har också ett arkiv där du kan låna översättningar av finska pjäser på olika språk.
Du kan söka information om teatrarnas repertoar och tillgängligheten av biljetter och biljettpriserna till exempel på biljettjänstens eller teatrarnas webbplatser.
I Finland ordnas också många teaterfestivaler.
Information om dessa hittar du på webbplatserna för Informationscentralen för teater i Finland på finska, svenska och på engelska.
linkkiInformationscentralen för teater i Finland:
Kontaktuppgifter till teatrarfinska
linkkiTeaterinfo Finland:
Teaterfestivalerfinska _ svenska _ engelska
Film
I de flesta städer finns en biograf.
Enklast hittar du information om biograferna i ditt område, bioprogrammet och biljettpriserna på internet.
Veckans bioprogram publiceras ofta också i lokaltidningen.
Finnkino är den största biografkedjan i Finland.
På Finnkinos webbplats kan du söka biografer enligt stad på engelska och finska och se vilka filmer som visas.
Om bioprogrammet på andra biografer kan du fråga direkt på biografen eller söka information på internet och i tidningar.
Biobiljetternas priser varierar något i Finland.
Som billigast kostar biljetten ungefär fem euro, som dyrast över tio euro.
Du kan ta reda på biljettpriset på förhand på biografens webbplats.
I Finland visas filmerna oftast på originalspråket.
Dessutom är de textade till finska och svenska.
Barnfilmerna är ett undantag. De kan vara dubbade till finska även om filmens originalspråk är något annat.
Biografer
Nationella audiovisuella arkivet visar nya och gamla filmer från hela världen.
Information om visningarna finns på finska på arkivets webbplats.
Visningar ordnas på flera orter.
Filmer på främmande språk har vanligen finsk- och svenskspråkig textning.
Filmfestivaler
I Finland ordnas årligen högklassiga filmfestivaler, varav de bäst kända är Kärlek och anarki-festivalen, som ordnas varje höst i Helsingfors, och Sodankylä filmfestival som ordnas på sommaren.
linkkiFinnkino:
Filmerfinska _ engelska
linkkiKärlek och anarki:
Filmfestivalfinska _ svenska _ engelska
Filmfestivalfinska _ engelska
Information om filmer och filmvisningarfinska _ svenska _ engelska
På den här sidan finns information om tjänsterna i Rovaniemi.
Sjukanfall och olyckor
Familjerådgivning
Rovaniemi stads familjerådgivning
Familjerådgivningscentralen vid Rovaniemi församling
Kriscentret vid Lapplands mödra- och skyddshem
Ekonomi- och skuldrådgivning
Missbrukararbete
Missbruksproblem hos ungdomar
Våld i familjen
Brottsofferjouren
Rättshjälpsbyrån i Rovaniemi
Sjukanfall och olyckor
Vid akuta och livshotande sjukfall kan du tillkalla ambulans genom att ringa numret 112.
På samma nummer kan du även tillkalla brandkår eller polis.
Familjerådgivning
Om du har problem i familjen eller i parförhållandet och vill diskutera situationen med en utomstående person, kan du ta kontakt med följande instanser::
Rovaniemi stads familjerådgivning
Familjerådgivningen i Rovaniemi betjänar barnfamiljer med under 16-åriga barn.
Du kan kontakta rådgivningen om ditt barn har problem eller om ni har problem i familjen och du vill ha hjälp.
Kontaktuppgifter
tfn 016 322 2538
Öppet
mån–tors kl. 8–16
fre kl. 8–15.30
Familjerådgivningscentralen vid Rovaniemi församling
På familjerådgivningscentralen får du hjälp om ni har problem i familjen eller i parförhållandet.
Kontaktuppgifter
tfn 016 335 5250
Tidsbeställning mån–fre 9–11
Läs mer linkkiFörsamlingen:
Familjerådgivningscentralenfinska
Kriscentret vid Lapplands mödra- och skyddshem
Du kan kontakta kriscentret i alla slags situationer där du eller din familj behöver stöd eller hjälp; till exempel vid skilsmässa, svårigheter hos barn och unga, våld med mera.
Kontaktuppgifter:
tfn 020 741 4732
Jourtelefon med dygnet runt-bemanning (24 h), tfn 040 553 7508
Läs mer på webbplatsen för linkkiFörbundet för mödra- och skyddshem:
Kriscentret vid Lapplands mödra- och skyddshemfinska _ svenska _ engelska
Ekonomi- och skuldrådgivning
Om du har svårt att sköta din ekonomi, betalningssvårigheter eller skulder kan du få råd av en ekonomi- och skuldrådgivare.
Rådgivningen är avgiftsfri.
Läs mer på linkkiRovaniemi stad:
Ekonomi- och skuldrådgivningfinska.
Missbrukararbete
Om du har problem med alkohol eller andra droger eller spelproblem kan du ta kontakt med A-klinikkaan.
Också familjemedlemmar kan ringa eller besöka A-kliniken.
A-klinikens tjänster är avsedda för personer som har fyllt 25 år.
Kontaktuppgifter:
Öppet
mån–ons kl. 8–16
tors–fre kl. 8–15
Du kan besöka sjukskötarmottagningen utan tidsbeställning mån–fre kl. 8.30–11.
Du kan ringa A-klinikens medarbetare mån–fre kl. 8.30–10, tfn 040 195 3981
Missbruksproblem hos ungdomar
Romppu är settlementföreningen Rovalan Setlementti ry:s drog- och rusmedelsmottagning för ungdomar i Lappland.
Ungdomar som oroar sig för sitt eget eller sina föräldrars alkohol- eller drogbruk eller spelande kan kontakta Romppu.
Också föräldrar kan kontakta Romppu.
Du kan besöka kliniken utan tidsbeställning torsdagar kl. 14–15.30 eller boka en tid.
Tidsbeställning per telefon mån–ons kl. 9–10.
Kontaktuppgifter:
tfn 040 487 3030
Öppet
mån–tors kl. 8–16
fre kl. 8–14
Läs mer:
Romppu
Våld i familjen
Du kan komma till *Lapplands mödra- och skyddshem om någon i din familj är våldsam eller om du på grund av hot om våld inte vågar stanna hemma.
Du kan ta med dig barnen till skyddshemmet.
Du kan komma till skyddshemmet dygnet runt.
Kontaktuppgifter:
Jourtelefon med dygnet runt-bemanning (24 h), tfn 040 553 7508
Brottsofferjouren
Om du råkar ut för ett brott kan du be om hjälp vid *Brottsofferjouren.
Du kan få en stödperson som hjälper dig och stöder dig i skötseln av praktiska ärenden..
Kontaktuppgifter:
Lapplands regionkontor/ Rovaniemi serviceställe
tfn 0400 979 175
Hjälptelefon: 020 316 116
mån–tis kl. 13–21
ons–fre kl. 17–21
Juristens rådgivning per telefon 020 316 117
mån–tors kl. 17–19
Rättshjälpsbyrån i Rovaniemi
Om du behöver rättshjälpsbyråns tjänster ska du boka tid för ett besök.
Kontaktuppgifter:
tfn 010 366 1560
Läs mer: linkkiJustitieministeriet:
Rättshjälpfinska
På den här sidan finns information om tjänsterna i Rovaniemi.
Sjukanfall och olyckor
Familjerådgivning
Rovaniemi stads familjerådgivning
Familjerådgivningscentralen vid Rovaniemi församling
Kriscentret vid Lapplands mödra- och skyddshem
Ekonomi- och skuldrådgivning
Missbrukararbete
Missbruksproblem hos ungdomar
Våld i familjen
Brottsofferjouren
Rättshjälpsbyrån i Rovaniemi
Sjukanfall och olyckor
Vid akuta och livshotande sjukfall kan du tillkalla ambulans genom att ringa numret 112.
På samma nummer kan du även tillkalla brandkår eller polis.
Familjerådgivning
Om du har problem i familjen eller i parförhållandet och vill diskutera situationen med en utomstående person, kan du ta kontakt med följande instanser::
Rovaniemi stads familjerådgivning
Familjerådgivningen i Rovaniemi betjänar barnfamiljer med under 16-åriga barn.
Du kan kontakta rådgivningen om ditt barn har problem eller om ni har problem i familjen och du vill ha hjälp.
Kontaktuppgifter
tfn 016 322 2538
Öppet
mån–tors kl. 8–16
fre kl. 8–15.30
Familjerådgivningscentralen vid Rovaniemi församling
På familjerådgivningscentralen får du hjälp om ni har problem i familjen eller i parförhållandet.
Kontaktuppgifter
tfn 016 335 5250
Tidsbeställning mån–fre 9–11
Läs mer linkkiFörsamlingen:
Familjerådgivningscentralenfinska
Kriscentret vid Lapplands mödra- och skyddshem
Du kan kontakta kriscentret i alla slags situationer där du eller din familj behöver stöd eller hjälp; till exempel vid skilsmässa, svårigheter hos barn och unga, våld med mera.
Kontaktuppgifter:
tfn 020 741 4732
Jourtelefon med dygnet runt-bemanning (24 h), tfn 040 553 7508
Läs mer på webbplatsen för linkkiFörbundet för mödra- och skyddshem:
Kriscentret vid Lapplands mödra- och skyddshemfinska _ svenska _ engelska
Ekonomi- och skuldrådgivning
Om du har svårt att sköta din ekonomi, betalningssvårigheter eller skulder kan du få råd av en ekonomi- och skuldrådgivare.
Rådgivningen är avgiftsfri.
Läs mer på linkkiRovaniemi stad:
Ekonomi- och skuldrådgivningfinska.
Missbrukararbete
Om du har problem med alkohol eller andra droger eller spelproblem kan du ta kontakt med A-klinikkaan.
Också familjemedlemmar kan ringa eller besöka A-kliniken.
A-klinikens tjänster är avsedda för personer som har fyllt 25 år.
Kontaktuppgifter:
Öppet
mån–ons kl. 8–16
tors–fre kl. 8–15
Du kan besöka sjukskötarmottagningen utan tidsbeställning mån–fre kl. 8.30–11.
Du kan ringa A-klinikens medarbetare mån–fre kl. 8.30–10, tfn 040 195 3981
Missbruksproblem hos ungdomar
Romppu är settlementföreningen Rovalan Setlementti ry:s drog- och rusmedelsmottagning för ungdomar i Lappland.
Ungdomar som oroar sig för sitt eget eller sina föräldrars alkohol- eller drogbruk eller spelande kan kontakta Romppu.
Också föräldrar kan kontakta Romppu.
Du kan besöka kliniken utan tidsbeställning torsdagar kl. 14–15.30 eller boka en tid.
Tidsbeställning per telefon mån–ons kl. 9–10.
Kontaktuppgifter:
tfn 040 487 3030
Öppet
mån–tors kl. 8–16
fre kl. 8–14
Läs mer:
Romppu
Våld i familjen
Du kan komma till *Lapplands mödra- och skyddshem om någon i din familj är våldsam eller om du på grund av hot om våld inte vågar stanna hemma.
Du kan ta med dig barnen till skyddshemmet.
Du kan komma till skyddshemmet dygnet runt.
Kontaktuppgifter:
Jourtelefon med dygnet runt-bemanning (24 h), tfn 040 553 7508
Brottsofferjouren
Om du råkar ut för ett brott kan du be om hjälp vid *Brottsofferjouren.
Du kan få en stödperson som hjälper dig och stöder dig i skötseln av praktiska ärenden..
Kontaktuppgifter:
Lapplands regionkontor/ Rovaniemi serviceställe
tfn 0400 979 175
Hjälptelefon: 020 316 116
mån–tis kl. 13–21
ons–fre kl. 17–21
Juristens rådgivning per telefon 020 316 117
mån–tors kl. 17–19
Rättshjälpsbyrån i Rovaniemi
Om du behöver rättshjälpsbyråns tjänster ska du boka tid för ett besök.
Kontaktuppgifter:
tfn 010 366 1560
Läs mer: linkkiJustitieministeriet:
Rättshjälpfinska
På den här sidan finns information om tjänsterna i Rovaniemi.
Sjukanfall och olyckor
Familjerådgivning
Rovaniemi stads familjerådgivning
Familjerådgivningscentralen vid Rovaniemi församling
Kriscentret vid Lapplands mödra- och skyddshem
Ekonomi- och skuldrådgivning
Missbrukararbete
Missbruksproblem hos ungdomar
Våld i familjen
Brottsofferjouren
Rättshjälpsbyrån i Rovaniemi
Sjukanfall och olyckor
Vid akuta och livshotande sjukfall kan du tillkalla ambulans genom att ringa numret 112.
På samma nummer kan du även tillkalla brandkår eller polis.
Familjerådgivning
Om du har problem i familjen eller i parförhållandet och vill diskutera situationen med en utomstående person, kan du ta kontakt med följande instanser::
Rovaniemi stads familjerådgivning
Familjerådgivningen i Rovaniemi betjänar barnfamiljer med under 16-åriga barn.
Du kan kontakta rådgivningen om ditt barn har problem eller om ni har problem i familjen och du vill ha hjälp.
Kontaktuppgifter
tfn 016 322 2538
Öppet
mån–tors kl. 8–16
fre kl. 8–15.30
Familjerådgivningscentralen vid Rovaniemi församling
På familjerådgivningscentralen får du hjälp om ni har problem i familjen eller i parförhållandet.
Kontaktuppgifter
tfn 016 335 5250
Tidsbeställning mån–fre 9–11
Läs mer linkkiFörsamlingen:
Familjerådgivningscentralenfinska
Kriscentret vid Lapplands mödra- och skyddshem
Du kan kontakta kriscentret i alla slags situationer där du eller din familj behöver stöd eller hjälp; till exempel vid skilsmässa, svårigheter hos barn och unga, våld med mera.
Kontaktuppgifter:
tfn 020 741 4732
Jourtelefon med dygnet runt-bemanning (24 h), tfn 040 553 7508
Läs mer på webbplatsen för linkkiFörbundet för mödra- och skyddshem:
Kriscentret vid Lapplands mödra- och skyddshemfinska _ svenska _ engelska
Ekonomi- och skuldrådgivning
Om du har svårt att sköta din ekonomi, betalningssvårigheter eller skulder kan du få råd av en ekonomi- och skuldrådgivare.
Rådgivningen är avgiftsfri.
Läs mer på linkkiRovaniemi stad:
Ekonomi- och skuldrådgivningfinska.
Missbrukararbete
Om du har problem med alkohol eller andra droger eller spelproblem kan du ta kontakt med A-klinikkaan.
Också familjemedlemmar kan ringa eller besöka A-kliniken.
A-klinikens tjänster är avsedda för personer som har fyllt 25 år.
Kontaktuppgifter:
Öppet
mån–ons kl. 8–16
tors–fre kl. 8–15
Du kan besöka sjukskötarmottagningen utan tidsbeställning mån–fre kl. 8.30–11.
Du kan ringa A-klinikens medarbetare mån–fre kl. 8.30–10, tfn 040 195 3981
Missbruksproblem hos ungdomar
Romppu är settlementföreningen Rovalan Setlementti ry:s drog- och rusmedelsmottagning för ungdomar i Lappland.
Ungdomar som oroar sig för sitt eget eller sina föräldrars alkohol- eller drogbruk eller spelande kan kontakta Romppu.
Också föräldrar kan kontakta Romppu.
Du kan besöka kliniken utan tidsbeställning torsdagar kl. 14–15.30 eller boka en tid.
Tidsbeställning per telefon mån–ons kl. 9–10.
Kontaktuppgifter:
tfn 040 487 3030
Öppet
mån–tors kl. 8–16
fre kl. 8–14
Läs mer:
Romppu
Våld i familjen
Du kan komma till *Lapplands mödra- och skyddshem om någon i din familj är våldsam eller om du på grund av hot om våld inte vågar stanna hemma.
Du kan ta med dig barnen till skyddshemmet.
Du kan komma till skyddshemmet dygnet runt.
Kontaktuppgifter:
Jourtelefon med dygnet runt-bemanning (24 h), tfn 040 553 7508
Brottsofferjouren
Om du råkar ut för ett brott kan du be om hjälp vid *Brottsofferjouren.
Du kan få en stödperson som hjälper dig och stöder dig i skötseln av praktiska ärenden..
Kontaktuppgifter:
Lapplands regionkontor/ Rovaniemi serviceställe
tfn 0400 979 175
Hjälptelefon: 020 316 116
mån–tis kl. 13–21
ons–fre kl. 17–21
Juristens rådgivning per telefon 020 316 117
mån–tors kl. 17–19
Rättshjälpsbyrån i Rovaniemi
Om du behöver rättshjälpsbyråns tjänster ska du boka tid för ett besök.
Kontaktuppgifter:
tfn 010 366 1560
Läs mer: linkkiJustitieministeriet:
Rättshjälpfinska
Naturen i Finland är mångsidig.
Det är roligt och tryggt att röra sig i naturen när du väljer rutter som passar dig med hänsyn till din kondition och dina kunskaper och följer anvisningar.
I Finland har vi fyra mycket olika årstider.
Beroende på årstiden och området finns det olika aktivitetsmöjligheter.
Läs mer om årstiderna i Finland på InfoFinlands sida Klimatet i Finland.
Friluftsliv och vandring
Vandring och friluftsliv är hobbyer som kan idkas alla årstider.
Om du inte har tidigare erfarenhet av friluftsliv eller vandring är det bra att börja med korta och enkla rutter som ligger nära bosättningen.
Korta turer kan du göra utan speciell utrustning.
Det är dock bra att ta med sig något att dricka, telefonen och en karta.
Det är bäst att börja med en rutt som märkts ut.
Ruttkartor säljs i bokhandlar och på internet.
Längre utflykter och vandringar kräver mer planering och förberedelser.
Norrsken
Finland är en av de bästa länderna i världen om man vill se norrsken (aurora borealis).
Oftast kan de ses på himlen i norra Lappland från september till mars.
Ibland kan norrsken ses också i södra Finland.
För att norrsken ska synas bra ska natten vara klar och mörk och man ska befinna sig långt från belysta tätorter.
Det lönar sig att klä sig varmt eftersom klara nätter vanligtvis också är kalla.
På sommaren är nätterna för ljusa för att man ska kunna se norrsken.
Norrskenfinska _ engelska
Skidåkning
Att åka skidor är en av de populäraste vintersporterna i Finland.
Den är en hälsosam och nästan gratis motionsform.
Information om kurser i skidåkning, om att hyra skidor och om skidspår finns till exempel på Suomen Latu ry:s webbplats på finska.
Information om skidåkningfinska
Att röra sig till sjöss
Finländarna rör sig mycket till sjöss.
Finländarna är också aktiva paddlare och seglare.
Säkerheten är viktig till sjöss.
Följ väderleksrapporterna och använd alltid en flytväst i rätt storlek.
Att färdas på isen
På vintern fryser de flesta vattendrag till i Finland.
På isen kan du till exempel promenera, åka skridskor eller skidor eller pimpla.
När isen är mycket tjock kan man också köra med motorkälke eller bil på den.
Man är alltid utsatt för risker när man färdas på isen och det är viktigt att iaktta säkerheten.
Checklista för den som ska färdas på isen:
Då isen fryser håller den inte genast för att gå på.
Isens tjocklek kan variera även på korta sträckor.
På våren är det mycket svårt att bedöma isens bärkraft och då är det bäst att undvika att färdas på isen.
Det viktigaste redskapet för den som färdas på isen är isdubbar.
Utan dem är det mycket svårt att ta sig upp ur en vak.
Om du inte är säker på att isen håller, gå inte ut på isen.
Fiske
Mete (med metspö) och pimpelfiske omfattas, med vissa undantag, av allemansrätten och du behöver inte skaffa dig ett fisketillstånd för dessa.
För allt annat fiske och kräftfiske ska du betala:
Den länsbaserade handredskapsavgiften är personlig och ska betalas innan fisket påbörjas.
Du kan betala avgiften antingen för ett kalenderår eller för sju dygn.
Information om fisketillståndfinska _ svenska _ engelska
Allemansrätten
Allemansrätten (jokamiehen oikeudet) är en väsentlig del av den finländska kulturen och lagstiftningen.
Allemansrätten i ett nötskal
Du får:
röra dig till fots, cykla och åka skidor överallt i naturen utom på gårdsplaner eller över åkrar, ängar eller planteringar som kan ta skada
tillfälligt vistas på marker där det är tillåtet att röra sig enligt ovan. Du kan till exempel tälta relativt fritt bara du håller ett tillräckligt avstånd till andras bostäder.
plocka vilda bär och blommor samt svamp
meta och pimpelfiska
ägna dig åt båtliv, simma och tvätta dig i sjöar och vattendrag samt färdas på isen.
Du får inte:
störa andra eller orsaka olägenhet för andra
störa eller skada fågelbon eller fågelungar
störa renar eller vilt
fälla eller skada växande träd
ta torra eller kullfallna träd, ris, mossa eller liknande på annans mark utan tillstånd
utan tvingande skäl göra upp öppen eld på annans mark
störa hemfriden till exempel genom att slå läger alltför nära en bostad eller genom att föra oväsen
skräpa ner i naturen
köra ett motorfordon i terrängen utan tillstånd av markägaren
fiska eller jaga utan de tillstånd som krävs.
linkkiMiljöministeriet:
Broschyren Allemansrättenfinska _ svenska _ engelska _ ryska
Friluftsliv och vandringfinska _ svenska _ engelska
Friluftskartor på Internetfinska _ svenska _ engelska
Tillståndfinska _ svenska
Nationalparker och naturskyddsområden
I Finland finns 40 nationalparker.
Med nationalpark avses ett över 1 000 hektar stort naturskyddsområde.
Det främsta syftet med nationalparker är att trygga naturens mångfald men samtidigt är de sevärdheter som är öppna för alla.
Nationalparkernas vackra landskap är ett bra resemål.
I de större parkerna kan man övernatta och göra längre utflykter.
I många nationalparker finns forststyrelsens naturcenter där man får aktuell information om områdets natur och om hur man ska röra sig i området.
Det är ett bra ställe att börja besöket på.
Nationalparkerna är populära utflyktsmål.
Friluftskartor på Internetfinska _ svenska _ engelska
Nationalparkerfinska _ svenska _ engelska _ ryska _ kinesiska
Fritidsobjekt på kartanfinska _ svenska _ engelska _ ryska _ estniska _ franska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ tyska _ vietnamesiska _ portugisiska _ polska _ holländska _ japanska _ italienska
_ isländska
Naturen i Finland är mångsidig.
Det är roligt och tryggt att röra sig i naturen när du väljer rutter som passar dig med hänsyn till din kondition och dina kunskaper och följer anvisningar.
I Finland har vi fyra mycket olika årstider.
Beroende på årstiden och området finns det olika aktivitetsmöjligheter.
Läs mer om årstiderna i Finland på InfoFinlands sida Klimatet i Finland.
Friluftsliv och vandring
Vandring och friluftsliv är hobbyer som kan idkas alla årstider.
Om du inte har tidigare erfarenhet av friluftsliv eller vandring är det bra att börja med korta och enkla rutter som ligger nära bosättningen.
Korta turer kan du göra utan speciell utrustning.
Det är dock bra att ta med sig något att dricka, telefonen och en karta.
Det är bäst att börja med en rutt som märkts ut.
Ruttkartor säljs i bokhandlar och på internet.
Längre utflykter och vandringar kräver mer planering och förberedelser.
Norrsken
Finland är en av de bästa länderna i världen om man vill se norrsken (aurora borealis).
Oftast kan de ses på himlen i norra Lappland från september till mars.
Ibland kan norrsken ses också i södra Finland.
För att norrsken ska synas bra ska natten vara klar och mörk och man ska befinna sig långt från belysta tätorter.
Det lönar sig att klä sig varmt eftersom klara nätter vanligtvis också är kalla.
På sommaren är nätterna för ljusa för att man ska kunna se norrsken.
Norrskenfinska _ engelska
Skidåkning
Att åka skidor är en av de populäraste vintersporterna i Finland.
Den är en hälsosam och nästan gratis motionsform.
Information om kurser i skidåkning, om att hyra skidor och om skidspår finns till exempel på Suomen Latu ry:s webbplats på finska.
Information om skidåkningfinska
Att röra sig till sjöss
Finländarna rör sig mycket till sjöss.
Finländarna är också aktiva paddlare och seglare.
Säkerheten är viktig till sjöss.
Följ väderleksrapporterna och använd alltid en flytväst i rätt storlek.
Att färdas på isen
På vintern fryser de flesta vattendrag till i Finland.
På isen kan du till exempel promenera, åka skridskor eller skidor eller pimpla.
När isen är mycket tjock kan man också köra med motorkälke eller bil på den.
Man är alltid utsatt för risker när man färdas på isen och det är viktigt att iaktta säkerheten.
Checklista för den som ska färdas på isen:
Då isen fryser håller den inte genast för att gå på.
Isens tjocklek kan variera även på korta sträckor.
På våren är det mycket svårt att bedöma isens bärkraft och då är det bäst att undvika att färdas på isen.
Det viktigaste redskapet för den som färdas på isen är isdubbar.
Utan dem är det mycket svårt att ta sig upp ur en vak.
Om du inte är säker på att isen håller, gå inte ut på isen.
Fiske
Mete (med metspö) och pimpelfiske omfattas, med vissa undantag, av allemansrätten och du behöver inte skaffa dig ett fisketillstånd för dessa.
För allt annat fiske och kräftfiske ska du betala:
Den länsbaserade handredskapsavgiften är personlig och ska betalas innan fisket påbörjas.
Du kan betala avgiften antingen för ett kalenderår eller för sju dygn.
Information om fisketillståndfinska _ svenska _ engelska
Allemansrätten
Allemansrätten (jokamiehen oikeudet) är en väsentlig del av den finländska kulturen och lagstiftningen.
Allemansrätten i ett nötskal
Du får:
röra dig till fots, cykla och åka skidor överallt i naturen utom på gårdsplaner eller över åkrar, ängar eller planteringar som kan ta skada
tillfälligt vistas på marker där det är tillåtet att röra sig enligt ovan. Du kan till exempel tälta relativt fritt bara du håller ett tillräckligt avstånd till andras bostäder.
plocka vilda bär och blommor samt svamp
meta och pimpelfiska
ägna dig åt båtliv, simma och tvätta dig i sjöar och vattendrag samt färdas på isen.
Du får inte:
störa andra eller orsaka olägenhet för andra
störa eller skada fågelbon eller fågelungar
störa renar eller vilt
fälla eller skada växande träd
ta torra eller kullfallna träd, ris, mossa eller liknande på annans mark utan tillstånd
utan tvingande skäl göra upp öppen eld på annans mark
störa hemfriden till exempel genom att slå läger alltför nära en bostad eller genom att föra oväsen
skräpa ner i naturen
köra ett motorfordon i terrängen utan tillstånd av markägaren
fiska eller jaga utan de tillstånd som krävs.
linkkiMiljöministeriet:
Broschyren Allemansrättenfinska _ svenska _ engelska _ ryska
Friluftsliv och vandringfinska _ svenska _ engelska
Friluftskartor på Internetfinska _ svenska _ engelska
Tillståndfinska _ svenska
Nationalparker och naturskyddsområden
I Finland finns 40 nationalparker.
Med nationalpark avses ett över 1 000 hektar stort naturskyddsområde.
Det främsta syftet med nationalparker är att trygga naturens mångfald men samtidigt är de sevärdheter som är öppna för alla.
Nationalparkernas vackra landskap är ett bra resemål.
I de större parkerna kan man övernatta och göra längre utflykter.
I många nationalparker finns forststyrelsens naturcenter där man får aktuell information om områdets natur och om hur man ska röra sig i området.
Det är ett bra ställe att börja besöket på.
Nationalparkerna är populära utflyktsmål.
Friluftskartor på Internetfinska _ svenska _ engelska
Nationalparkerfinska _ svenska _ engelska _ ryska _ kinesiska
Fritidsobjekt på kartanfinska _ svenska _ engelska _ ryska _ estniska _ franska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ tyska _ vietnamesiska _ portugisiska _ polska _ holländska _ japanska _ italienska
_ isländska
Naturen i Finland är mångsidig.
Det är roligt och tryggt att röra sig i naturen när du väljer rutter som passar dig med hänsyn till din kondition och dina kunskaper och följer anvisningar.
I Finland har vi fyra mycket olika årstider.
Beroende på årstiden och området finns det olika aktivitetsmöjligheter.
Läs mer om årstiderna i Finland på InfoFinlands sida Klimatet i Finland.
Friluftsliv och vandring
Vandring och friluftsliv är hobbyer som kan idkas alla årstider.
Om du inte har tidigare erfarenhet av friluftsliv eller vandring är det bra att börja med korta och enkla rutter som ligger nära bosättningen.
Korta turer kan du göra utan speciell utrustning.
Det är dock bra att ta med sig något att dricka, telefonen och en karta.
Det är bäst att börja med en rutt som märkts ut.
Ruttkartor säljs i bokhandlar och på internet.
Längre utflykter och vandringar kräver mer planering och förberedelser.
Norrsken
Finland är en av de bästa länderna i världen om man vill se norrsken (aurora borealis).
Oftast kan de ses på himlen i norra Lappland från september till mars.
Ibland kan norrsken ses också i södra Finland.
För att norrsken ska synas bra ska natten vara klar och mörk och man ska befinna sig långt från belysta tätorter.
Det lönar sig att klä sig varmt eftersom klara nätter vanligtvis också är kalla.
På sommaren är nätterna för ljusa för att man ska kunna se norrsken.
Norrskenfinska _ engelska
Skidåkning
Att åka skidor är en av de populäraste vintersporterna i Finland.
Den är en hälsosam och nästan gratis motionsform.
Information om kurser i skidåkning, om att hyra skidor och om skidspår finns till exempel på Suomen Latu ry:s webbplats på finska.
Information om skidåkningfinska
Att röra sig till sjöss
Finländarna rör sig mycket till sjöss.
Finländarna är också aktiva paddlare och seglare.
Säkerheten är viktig till sjöss.
Följ väderleksrapporterna och använd alltid en flytväst i rätt storlek.
Att färdas på isen
På vintern fryser de flesta vattendrag till i Finland.
På isen kan du till exempel promenera, åka skridskor eller skidor eller pimpla.
När isen är mycket tjock kan man också köra med motorkälke eller bil på den.
Man är alltid utsatt för risker när man färdas på isen och det är viktigt att iaktta säkerheten.
Checklista för den som ska färdas på isen:
Då isen fryser håller den inte genast för att gå på.
Isens tjocklek kan variera även på korta sträckor.
På våren är det mycket svårt att bedöma isens bärkraft och då är det bäst att undvika att färdas på isen.
Det viktigaste redskapet för den som färdas på isen är isdubbar.
Utan dem är det mycket svårt att ta sig upp ur en vak.
Om du inte är säker på att isen håller, gå inte ut på isen.
Fiske
Mete (med metspö) och pimpelfiske omfattas, med vissa undantag, av allemansrätten och du behöver inte skaffa dig ett fisketillstånd för dessa.
För allt annat fiske och kräftfiske ska du betala:
Den länsbaserade handredskapsavgiften är personlig och ska betalas innan fisket påbörjas.
Du kan betala avgiften antingen för ett kalenderår eller för sju dygn.
Information om fisketillståndfinska _ svenska _ engelska
Allemansrätten
Allemansrätten (jokamiehen oikeudet) är en väsentlig del av den finländska kulturen och lagstiftningen.
Allemansrätten i ett nötskal
Du får:
röra dig till fots, cykla och åka skidor överallt i naturen utom på gårdsplaner eller över åkrar, ängar eller planteringar som kan ta skada
tillfälligt vistas på marker där det är tillåtet att röra sig enligt ovan. Du kan till exempel tälta relativt fritt bara du håller ett tillräckligt avstånd till andras bostäder.
plocka vilda bär och blommor samt svamp
meta och pimpelfiska
ägna dig åt båtliv, simma och tvätta dig i sjöar och vattendrag samt färdas på isen.
Du får inte:
störa andra eller orsaka olägenhet för andra
störa eller skada fågelbon eller fågelungar
störa renar eller vilt
fälla eller skada växande träd
ta torra eller kullfallna träd, ris, mossa eller liknande på annans mark utan tillstånd
utan tvingande skäl göra upp öppen eld på annans mark
störa hemfriden till exempel genom att slå läger alltför nära en bostad eller genom att föra oväsen
skräpa ner i naturen
köra ett motorfordon i terrängen utan tillstånd av markägaren
fiska eller jaga utan de tillstånd som krävs.
linkkiMiljöministeriet:
Broschyren Allemansrättenfinska _ svenska _ engelska _ ryska
Friluftsliv och vandringfinska _ svenska _ engelska
Friluftskartor på Internetfinska _ svenska _ engelska
Tillståndfinska _ svenska
Nationalparker och naturskyddsområden
I Finland finns 40 nationalparker.
Med nationalpark avses ett över 1 000 hektar stort naturskyddsområde.
Det främsta syftet med nationalparker är att trygga naturens mångfald men samtidigt är de sevärdheter som är öppna för alla.
Nationalparkernas vackra landskap är ett bra resemål.
I de större parkerna kan man övernatta och göra längre utflykter.
I många nationalparker finns forststyrelsens naturcenter där man får aktuell information om områdets natur och om hur man ska röra sig i området.
Det är ett bra ställe att börja besöket på.
Nationalparkerna är populära utflyktsmål.
Friluftskartor på Internetfinska _ svenska _ engelska
Nationalparkerfinska _ svenska _ engelska _ ryska _ kinesiska
Fritidsobjekt på kartanfinska _ svenska _ engelska _ ryska _ estniska _ franska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ tyska _ vietnamesiska _ portugisiska _ polska _ holländska _ japanska _ italienska
_ isländska
Folk i Finland är aktiva motionärer och olika motionshobbyer kan hjälpa dig att bli bekant med människor och få nya vänner.
Ledd motion ordnas till exempel av olika idrottssällskap som ofta drivs med frivilligarbete.
Lätt motion kan även vara till exempel trädgårdsskötsel, städning eller snöskottande, d.v.s. så kallad vardagsmotion (hyötyliikunta).
Att ta sig till arbetet eller butiken till fots eller med cykeln är ett lätt sätt att få den dagliga motionsdosen.
Också äldre människor har nytta av att röra på sig, eftersom motion upprätthåller den fysiska konditionen och funktionsförmågan.
Motion är även viktigt för barn.
Läs mer på Infobankens sida Barn och ungas hobbyer.
Ledd motion
Ledd motion ordnas till exempel av kommuner och idrottsklubbar.
På några orter finns det dessutom ledd motion som är avsedd endast för invandrare, exempelvis egna grupper för kvinnor eller för personer som vill bekanta sig med nya idrottsgrenar.
Ledd motion är tillgänglig för alla.
Alla kan delta i idrottsklubbarnas verksamhet.
Ledd motion kan vara till exempel jympa eller promenader, löpning eller skidåkning i grupp.
Val av gren och grupp
När du väljer en motionshobby är det klokt att beakta den egna konditionen.
Hobbygrupper finns både för nybörjare och mer avancerade.
Simning och skidåkning är mycket populära grenar i Finland och i dem ordnas nybörjarkurser även för vuxna.
Du kan idka båda grenarna på egen hand när du väl lärt dig grunderna.
Idrottsanläggningar
I Finland ägs cirka 70 procent av idrottsanläggningarna av kommunerna.
Sådana är till exempel många idrotts- och simhallar och andra idrottsanläggningar, såsom fotbollsplaner och skridskobanor.
Kommunernas idrottsplatser får användas av alla invånare.
Bästa stället att fråga mer om kommunernas idrottsplatser är vid idrottsväsendet i den egna kommunen.
Kontaktuppgifterna hittar på din kommuns hemsida.
I stora städer finns också privata idrottsanläggningar.
Fråga mer om utbudet och priserna direkt på idrottscentret.
För studerande och förvärvsarbetande lönar det sig att ta reda på om läroanstalten eller arbetsplatsen erbjuder motionsmöjligheter.
linkkiFinlands Simundervisnings- och Livräddningsförbund rf:
Kom till simhallen!(pdf, 2 MB)finska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ arabiska _ kurdiska _ thai
Motionsföreningfinska _ engelska
Motionsrekommendationerfinska _ engelska
Folk i Finland är aktiva motionärer och olika motionshobbyer kan hjälpa dig att bli bekant med människor och få nya vänner.
Ledd motion ordnas till exempel av olika idrottssällskap som ofta drivs med frivilligarbete.
Lätt motion kan även vara till exempel trädgårdsskötsel, städning eller snöskottande, d.v.s. så kallad vardagsmotion (hyötyliikunta).
Att ta sig till arbetet eller butiken till fots eller med cykeln är ett lätt sätt att få den dagliga motionsdosen.
Också äldre människor har nytta av att röra på sig, eftersom motion upprätthåller den fysiska konditionen och funktionsförmågan.
Motion är även viktigt för barn.
Läs mer på Infobankens sida Barn och ungas hobbyer.
Ledd motion
Ledd motion ordnas till exempel av kommuner och idrottsklubbar.
På några orter finns det dessutom ledd motion som är avsedd endast för invandrare, exempelvis egna grupper för kvinnor eller för personer som vill bekanta sig med nya idrottsgrenar.
Ledd motion är tillgänglig för alla.
Alla kan delta i idrottsklubbarnas verksamhet.
Ledd motion kan vara till exempel jympa eller promenader, löpning eller skidåkning i grupp.
Val av gren och grupp
När du väljer en motionshobby är det klokt att beakta den egna konditionen.
Hobbygrupper finns både för nybörjare och mer avancerade.
Simning och skidåkning är mycket populära grenar i Finland och i dem ordnas nybörjarkurser även för vuxna.
Du kan idka båda grenarna på egen hand när du väl lärt dig grunderna.
Idrottsanläggningar
I Finland ägs cirka 70 procent av idrottsanläggningarna av kommunerna.
Sådana är till exempel många idrotts- och simhallar och andra idrottsanläggningar, såsom fotbollsplaner och skridskobanor.
Kommunernas idrottsplatser får användas av alla invånare.
Bästa stället att fråga mer om kommunernas idrottsplatser är vid idrottsväsendet i den egna kommunen.
Kontaktuppgifterna hittar på din kommuns hemsida.
I stora städer finns också privata idrottsanläggningar.
Fråga mer om utbudet och priserna direkt på idrottscentret.
För studerande och förvärvsarbetande lönar det sig att ta reda på om läroanstalten eller arbetsplatsen erbjuder motionsmöjligheter.
linkkiFinlands Simundervisnings- och Livräddningsförbund rf:
Kom till simhallen!(pdf, 2 MB)finska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ arabiska _ kurdiska _ thai
Motionsföreningfinska _ engelska
Motionsrekommendationerfinska _ engelska
Folk i Finland är aktiva motionärer och olika motionshobbyer kan hjälpa dig att bli bekant med människor och få nya vänner.
Ledd motion ordnas till exempel av olika idrottssällskap som ofta drivs med frivilligarbete.
Lätt motion kan även vara till exempel trädgårdsskötsel, städning eller snöskottande, d.v.s. så kallad vardagsmotion (hyötyliikunta).
Att ta sig till arbetet eller butiken till fots eller med cykeln är ett lätt sätt att få den dagliga motionsdosen.
Också äldre människor har nytta av att röra på sig, eftersom motion upprätthåller den fysiska konditionen och funktionsförmågan.
Motion är även viktigt för barn.
Läs mer på Infobankens sida Barn och ungas hobbyer.
Ledd motion
Ledd motion ordnas till exempel av kommuner och idrottsklubbar.
På några orter finns det dessutom ledd motion som är avsedd endast för invandrare, exempelvis egna grupper för kvinnor eller för personer som vill bekanta sig med nya idrottsgrenar.
Ledd motion är tillgänglig för alla.
Alla kan delta i idrottsklubbarnas verksamhet.
Ledd motion kan vara till exempel jympa eller promenader, löpning eller skidåkning i grupp.
Val av gren och grupp
När du väljer en motionshobby är det klokt att beakta den egna konditionen.
Hobbygrupper finns både för nybörjare och mer avancerade.
Simning och skidåkning är mycket populära grenar i Finland och i dem ordnas nybörjarkurser även för vuxna.
Du kan idka båda grenarna på egen hand när du väl lärt dig grunderna.
Idrottsanläggningar
I Finland ägs cirka 70 procent av idrottsanläggningarna av kommunerna.
Sådana är till exempel många idrotts- och simhallar och andra idrottsanläggningar, såsom fotbollsplaner och skridskobanor.
Kommunernas idrottsplatser får användas av alla invånare.
Bästa stället att fråga mer om kommunernas idrottsplatser är vid idrottsväsendet i den egna kommunen.
Kontaktuppgifterna hittar på din kommuns hemsida.
I stora städer finns också privata idrottsanläggningar.
Fråga mer om utbudet och priserna direkt på idrottscentret.
För studerande och förvärvsarbetande lönar det sig att ta reda på om läroanstalten eller arbetsplatsen erbjuder motionsmöjligheter.
linkkiFinlands Simundervisnings- och Livräddningsförbund rf:
Kom till simhallen!(pdf, 2 MB)finska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ arabiska _ kurdiska _ thai
Motionsföreningfinska
Motionsrekommendationerfinska _ engelska
I Finland finns ett kommunalt bibliotek eller stadsbibliotek på alla orter.
Biblioteket är en plats där du kan låna böcker, läsa tidningar, använda datorn, studera eller delta i olika evenemang.
På biblioteket kan det även finnas sagotimmar och spel för barn.
I de flesta biblioteken finns en läsesal.
Läsesalen är ett tyst rum som passar för läsning eller till exempel tyst läxläsning.
Du kan också få handledning i datoranvändningen och på vissa bibliotek ordnas finska språkcaféer.
Du hittar bibliotekens kontaktuppgifter i webbtjänsten kirjastot.fi.
linkkiBiblioteken.fi:
Bibliotekets webbtjänstfinska _ svenska _ engelska
I Finland finns även vetenskapsbibliotek och läroanstalternas bibliotek samt olika slags specialbibliotek.
Användningen av dem kan vara begränsad, men oftast är de öppna för alla.
Bibliotekskort
För att låna material behöver du ett bibliotekskort.
Ett sådant får du på biblioteket.
Om du inte har en finländsk personbeteckning, kan du få ett bibliotekskort som är giltigt en bestämd tid.
Bibliotekskortet är avgiftsfritt.
Om du tappar bort kortet, måste du betala för ett nytt kort.
När du flyttar ska du meddela din nya adress till biblioteket.
Om du flyttar till en kommun där ditt bibliotekskort inte gäller, måste du skaffa dig ett nytt bibliotekskort vid biblioteket på din nya hemort.
Att låna material
Alla bibliotek har en webbplats där du kan söka information om bibliotekets samlingar och förnya dina lån samt reservera material.
Om du letar efter en viss bok, kan du också be om hjälp av personalen på biblioteket.
Du kan även låna böcker på bokbussarna.
Lånetiden för böckerna är vanligtvis en månad.
Kom ihåg att returnera eller förnya dina lån i tid.
För försenade lån måste du betala en förseningsavgift.
Avgiftens storlek beror på hur många böcker som är försenade och hur många dagar de är försenade.
På biblioteket kan du låna böcker på klarspråk som är skrivna på lättläst finska.
De är även lämpliga för studier i det finska språket.
På biblioteket kan du även låna tidskrifter, e-böcker samt CD- och DVD-skivor.
Flerspråkiga biblioteket
Flerspråkiga biblioteket har material på över 60 språk.
Biblioteket ligger i Böle i Helsingfors.
Material från Flerspråkiga bibliotekets samlingar kan lånas från hela Finland.
Du kan be bibliotekarien på ditt eget bibliotek att beställa det material du vill ha åt dig.
Mer information om Flerspråkiga biblioteket får du på Helmet.fi som är en gemensam webbplats för biblioteken i huvudstadsregionen.
linkkiHelsingfors stadsbibliotek:
Flerspråkiga biblioteketfinska _ svenska _ engelska
Webbaserat material
eBiblioteket (eKirjasto) tillhandahåller elektroniska material, såsom böcker, tidskrifter och filmer.
En del av eBibliotekets material kan användas fritt på internet och för en del av materialen behöver du ett bibliotekskort och en PIN-kod för kortet.
eBiblioteketfinska _ svenska _ engelska
Fråga bibliotekarien-tjänsten
Fråga bibliotekarien-tjänsten svarar på alla slags frågor.
Du kan skicka in din fråga via webblanketten på finska, svenska eller engelska.
Svaret skickas till din e-post och publiceras på tjänstens webbplats.
Fråga bibliotekarienfinska _ svenska _ engelska
I Finland finns ett kommunalt bibliotek eller stadsbibliotek på alla orter.
Biblioteket är en plats där du kan låna böcker, läsa tidningar, använda datorn, studera eller delta i olika evenemang.
På biblioteket kan det även finnas sagotimmar och spel för barn.
I de flesta biblioteken finns en läsesal.
Läsesalen är ett tyst rum som passar för läsning eller till exempel tyst läxläsning.
Du kan också få handledning i datoranvändningen och på vissa bibliotek ordnas finska språkcaféer.
Du hittar bibliotekens kontaktuppgifter i webbtjänsten kirjastot.fi.
linkkiBiblioteken.fi:
Bibliotekets webbtjänstfinska _ svenska _ engelska
I Finland finns även vetenskapsbibliotek och läroanstalternas bibliotek samt olika slags specialbibliotek.
Användningen av dem kan vara begränsad, men oftast är de öppna för alla.
Bibliotekskort
För att låna material behöver du ett bibliotekskort.
Ett sådant får du på biblioteket.
Om du inte har en finländsk personbeteckning, kan du få ett bibliotekskort som är giltigt en bestämd tid.
Bibliotekskortet är avgiftsfritt.
Om du tappar bort kortet, måste du betala för ett nytt kort.
När du flyttar ska du meddela din nya adress till biblioteket.
Om du flyttar till en kommun där ditt bibliotekskort inte gäller, måste du skaffa dig ett nytt bibliotekskort vid biblioteket på din nya hemort.
Att låna material
Alla bibliotek har en webbplats där du kan söka information om bibliotekets samlingar och förnya dina lån samt reservera material.
Om du letar efter en viss bok, kan du också be om hjälp av personalen på biblioteket.
Du kan även låna böcker på bokbussarna.
Lånetiden för böckerna är vanligtvis en månad.
Kom ihåg att returnera eller förnya dina lån i tid.
För försenade lån måste du betala en förseningsavgift.
Avgiftens storlek beror på hur många böcker som är försenade och hur många dagar de är försenade.
På biblioteket kan du låna böcker på klarspråk som är skrivna på lättläst finska.
De är även lämpliga för studier i det finska språket.
På biblioteket kan du även låna tidskrifter, e-böcker samt CD- och DVD-skivor.
Flerspråkiga biblioteket
Flerspråkiga biblioteket har material på över 60 språk.
Biblioteket ligger i Böle i Helsingfors.
Material från Flerspråkiga bibliotekets samlingar kan lånas från hela Finland.
Du kan be bibliotekarien på ditt eget bibliotek att beställa det material du vill ha åt dig.
Mer information om Flerspråkiga biblioteket får du på Helmet.fi som är en gemensam webbplats för biblioteken i huvudstadsregionen.
linkkiHelsingfors stadsbibliotek:
Flerspråkiga biblioteketfinska _ svenska _ engelska
Webbaserat material
eBiblioteket (eKirjasto) tillhandahåller elektroniska material, såsom böcker, tidskrifter och filmer.
En del av eBibliotekets material kan användas fritt på internet och för en del av materialen behöver du ett bibliotekskort och en PIN-kod för kortet.
eBiblioteketfinska _ svenska _ engelska
Fråga bibliotekarien-tjänsten
Fråga bibliotekarien-tjänsten svarar på alla slags frågor.
Du kan skicka in din fråga via webblanketten på finska, svenska eller engelska.
Svaret skickas till din e-post och publiceras på tjänstens webbplats.
Fråga bibliotekarienfinska _ svenska _ engelska
I Finland finns ett kommunalt bibliotek eller stadsbibliotek på alla orter.
Biblioteket är en plats där du kan låna böcker, läsa tidningar, använda datorn, studera eller delta i olika evenemang.
På biblioteket kan det även finnas sagotimmar och spel för barn.
I de flesta biblioteken finns en läsesal.
Läsesalen är ett tyst rum som passar för läsning eller till exempel tyst läxläsning.
Du kan också få handledning i datoranvändningen och på vissa bibliotek ordnas finska språkcaféer.
Du hittar bibliotekens kontaktuppgifter i webbtjänsten kirjastot.fi.
linkkiBiblioteken.fi:
Bibliotekets webbtjänstfinska _ svenska _ engelska
I Finland finns även vetenskapsbibliotek och läroanstalternas bibliotek samt olika slags specialbibliotek.
Användningen av dem kan vara begränsad, men oftast är de öppna för alla.
Bibliotekskort
För att låna material behöver du ett bibliotekskort.
Ett sådant får du på biblioteket.
Om du inte har en finländsk personbeteckning, kan du få ett bibliotekskort som är giltigt en bestämd tid.
Bibliotekskortet är avgiftsfritt.
Om du tappar bort kortet, måste du betala för ett nytt kort.
När du flyttar ska du meddela din nya adress till biblioteket.
Om du flyttar till en kommun där ditt bibliotekskort inte gäller, måste du skaffa dig ett nytt bibliotekskort vid biblioteket på din nya hemort.
Att låna material
Alla bibliotek har en webbplats där du kan söka information om bibliotekets samlingar och förnya dina lån samt reservera material.
Om du letar efter en viss bok, kan du också be om hjälp av personalen på biblioteket.
Du kan även låna böcker på bokbussarna.
Lånetiden för böckerna är vanligtvis en månad.
Kom ihåg att returnera eller förnya dina lån i tid.
För försenade lån måste du betala en förseningsavgift.
Avgiftens storlek beror på hur många böcker som är försenade och hur många dagar de är försenade.
På biblioteket kan du låna böcker på klarspråk som är skrivna på lättläst finska.
De är även lämpliga för studier i det finska språket.
På biblioteket kan du även låna tidskrifter, e-böcker samt CD- och DVD-skivor.
Flerspråkiga biblioteket
Flerspråkiga biblioteket har material på över 60 språk.
Biblioteket ligger i Böle i Helsingfors.
Material från Flerspråkiga bibliotekets samlingar kan lånas från hela Finland.
Du kan be bibliotekarien på ditt eget bibliotek att beställa det material du vill ha åt dig.
Mer information om Flerspråkiga biblioteket får du på Helmet.fi som är en gemensam webbplats för biblioteken i huvudstadsregionen.
linkkiHelsingfors stadsbibliotek:
Flerspråkiga biblioteketfinska _ svenska _ engelska
Webbaserat material
eBiblioteket (eKirjasto) tillhandahåller elektroniska material, såsom böcker, tidskrifter och filmer.
En del av eBibliotekets material kan användas fritt på internet och för en del av materialen behöver du ett bibliotekskort och en PIN-kod för kortet.
eBiblioteketfinska _ svenska _ engelska
Fråga bibliotekarien-tjänsten
Fråga bibliotekarien-tjänsten svarar på alla slags frågor.
Du kan skicka in din fråga via webblanketten på finska, svenska eller engelska.
Svaret skickas till din e-post och publiceras på tjänstens webbplats.
Fråga bibliotekarienfinska _ svenska _ engelska
Om en person dör utanför sjukhuset ska du genast anmäla ärendet till polisen eller en läkare.
Polisen ser till att dödsorsaken fastställs och anmäler dödsfallet till Befolkningsregistercentralen (Väestörekisterikeskus).
När en person dör på sjukhuset anmäls dödsfallet automatiskt till Befolkningsregistercentralen, Fpa (Kela) och pensionsanstalter.
När en närstående person avlider kan du få stöd och hjälp med din sorg vid hälsostationerna (terveysasema), på familjerådgivningen (perheneuvola), SOS-kriscentret för utlänningar inom Föreningen för mental hälsa i Finland (Suomen mielenterveysseuran ulkomaalaisten kriisipalvelu) samt hos församlingarna.
Du får hjälp på finska och svenska, och på de flesta ställena även på engelska.
Om det behövs kan du också anlita en tolk.
När en närstående har avliditfinska _ svenska _ engelska
Information om krissituationer och sorgfinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
linkkiFöreningen för mental hälsa i Finland:
Krishjälpfinska _ svenska _ engelska
Begravningstillstånd
För att den avlidne ska kunna begravas, behövs en dödsattest (kuolintodistus) som alltid skrivs av en läkare.
Dödsattesten kan fås när dödsorsaken har fastställts.
Om det är fråga om ett akut, oklart dödsfall, en olycka eller ett brott, utförs en obduktion för att utreda dödsorsaken.
Också polisen kan undersöka orsaken till dödsfallet.
Ibland kan begravningen fördröjas på grund av att utredningen av dödsorsaken räcker länge.
Begravning
Religiösa samfund kan hjälpa dig med att ordna begravningen.
Fråga mer hos din egen samfällighet.
På webbplatsen för evangelisk-lutherska kyrkan i Finland hittar du information om kyrkans tjänster.
Man kan också ordna en civil begravning utan religiösa inslag.Om civil begravning får du information hos servicecentret Pro-Ceremonier (Pro-Seremoniat).
Begravningsbyråernas tjänster är avgiftsbelagda.
De sköter begravningsarrangemangen, som till exempel transporten av den avlidne.
Begravningsbyråerna säljer också kistor och sköter enligt avtal och de anhörigas önskemål även allt annat som rör begravningen.
Om begravningsbyråer får du information till exempel från Finlands Begravningsbyråers Förbund (Suomen Hautaustoimistojen Liitto).
Många begravningsbyråer betjänar även på engelska.
Civil begravningfinska _ svenska _ engelska
linkkiEvangelisk-lutherska kyrkan i Finland:
Information om kyrklig begravningfinska _ svenska _ engelska
Gravplats
Nästan alla begravningsplatser i Finland ägs av evangelisk-lutherska församlingar men man kan få en gravplats även om man inte är medlem i den evangelisk-lutherska kyrkan.
Gravplatserna är avgiftsbelagda och förfrågningar om dessa kan ställas till församlingarna.
Om en person inte var medlem i kyrkan och inte ville ha en religiös begravning, förrättas en sådan inte.
Den avlidne kan begravas i kista eller kremeras.
På många orter finns också andra religionssamfunds begravningsplatser.
I de största städerna finns till exempel ortodoxa, islamska och judiska begravningsplatser.
På många orter finns även gravområden för avlidna personer som inte har varit medlemmar i något religionssamfund.
Den avlidnes aska kan också strös ut i naturen eller i ett vattendrag om markägaren ger tillstånd till detta.
Begravningsbidrag
Den avlidne kan ibland ha rätt till begravningsbidrag (hautausavustus) genom sitt senaste anställningsförhållande eller medlemskap i ett fackförbund.
Fråga den senaste arbetsgivaren eller fackförbundet om detta.
För begravningskostnaderna för en medellös avliden kan du ansöka om utkomststöd från hemortens socialbyrå (sosiaalitoimisto).
Efter att en person dött kan dennes änka eller änkling och barn få familjepension (perhe-eläke).
Syftet med familjepensionen är att trygga de efterlevandes utkomst.
I Finland finns två olika familjepensioner, Fpa:s familjepension och arbetspensionssystemets familjepension.
Om den avlidne har arbetat eller varit företagare i Finland kan dennes efterlevande få familjepension från arbetspensionssystemet.
Båda pensionerna kan sökas hos Fpa.
Om den avlidne har bott eller arbetat utomlands en lång tid innan flytten till Finland, kan de efterlevande även ha rätt till familjepension från det landet.
Information om familjepensionfinska _ svenska _ engelska
Testamente
Vem som ärver egendomen efter en avliden person stadgas i lagen.
Du kan också själv påverka vem din förmögenhet delas till.
Du kan skriva ett testamente (testamentti), d.v.s. en skriftlig utredning över vem som ska ärva din egendom efter din bortgång.
Det är bra att ta hjälp av en jurist när du skriver ditt testamente för att det ska vara lagligt.
Bouppteckning
Bouppteckningen (perunkirjoitus) är ett möte där man upprättar en skriftlig utredning över den avlidnes förmögenhet och skulder.Bouppteckningen måste göras inom tre månader från dödsfallet.
För bouppteckningen behövs en släktutredning över den avlidne.
Det krävs även ämbetsbevis (virkatodistus), som du får från magistraten eller kyrkoherdeämbetet.
Därtill behövs uppgifter om dödsbodelägarna, det vill säga om dem som ärver den avlidnes egendom.
Bouppteckningshandlingen (perukirja) ska lämnas till skattebyrån senast en månad efter bouppteckningen.
Mer information om bouppteckningen får du från rättsväsendet och skatteförvaltningen.
Bouppteckningen ordnas av den person som bäst känner till den avlidnes egendom och skulder.
Bouppteckningshandlingen undertecknas av två personer som bedömer den avlidnes egendom.
Det är bra att anlita en jurist för upprättandet av bouppteckningen.
Att inte göra bouppteckningen inom utsatt tid kan ha ofördelaktiga följder, till exempel större arvsskatt.
Arvsskatt
Om du ärver egendom av en avliden person måste du betala arvsskatt (perintövero) för egendomen.
Skattebeloppet beror på hur stor förmögenhet du har ärvt och hur nära släkt du är till den avlidne.
Arv vilkas värde understiger 20 000 euro är skattefria.
linkkiSkatteförvaltningen:
Information om bouppteckningfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Information om arvsskattfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Information till en avlidnes anhörigfinska _ svenska
Om en person dör utanför sjukhuset ska du genast anmäla ärendet till polisen eller en läkare.
Polisen ser till att dödsorsaken fastställs och anmäler dödsfallet till Befolkningsregistercentralen (Väestörekisterikeskus).
När en person dör på sjukhuset anmäls dödsfallet automatiskt till Befolkningsregistercentralen, Fpa (Kela) och pensionsanstalter.
När en närstående person avlider kan du få stöd och hjälp med din sorg vid hälsostationerna (terveysasema), på familjerådgivningen (perheneuvola), SOS-kriscentret för utlänningar inom Föreningen för mental hälsa i Finland (Suomen mielenterveysseuran ulkomaalaisten kriisipalvelu) samt hos församlingarna.
Du får hjälp på finska och svenska, och på de flesta ställena även på engelska.
Om det behövs kan du också anlita en tolk.
När en närstående har avliditfinska _ svenska _ engelska
Information om krissituationer och sorgfinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
linkkiFöreningen för mental hälsa i Finland:
Krishjälpfinska _ svenska _ engelska
Begravningstillstånd
För att den avlidne ska kunna begravas, behövs en dödsattest (kuolintodistus) som alltid skrivs av en läkare.
Dödsattesten kan fås när dödsorsaken har fastställts.
Om det är fråga om ett akut, oklart dödsfall, en olycka eller ett brott, utförs en obduktion för att utreda dödsorsaken.
Också polisen kan undersöka orsaken till dödsfallet.
Ibland kan begravningen fördröjas på grund av att utredningen av dödsorsaken räcker länge.
Begravning
Religiösa samfund kan hjälpa dig med att ordna begravningen.
Fråga mer hos din egen samfällighet.
På webbplatsen för evangelisk-lutherska kyrkan i Finland hittar du information om kyrkans tjänster.
Man kan också ordna en civil begravning utan religiösa inslag.Om civil begravning får du information hos servicecentret Pro-Ceremonier (Pro-Seremoniat).
Begravningsbyråernas tjänster är avgiftsbelagda.
De sköter begravningsarrangemangen, som till exempel transporten av den avlidne.
Begravningsbyråerna säljer också kistor och sköter enligt avtal och de anhörigas önskemål även allt annat som rör begravningen.
Om begravningsbyråer får du information till exempel från Finlands Begravningsbyråers Förbund (Suomen Hautaustoimistojen Liitto).
Många begravningsbyråer betjänar även på engelska.
Civil begravningfinska _ svenska _ engelska
linkkiEvangelisk-lutherska kyrkan i Finland:
Information om kyrklig begravningfinska _ svenska _ engelska
Gravplats
Nästan alla begravningsplatser i Finland ägs av evangelisk-lutherska församlingar men man kan få en gravplats även om man inte är medlem i den evangelisk-lutherska kyrkan.
Gravplatserna är avgiftsbelagda och förfrågningar om dessa kan ställas till församlingarna.
Om en person inte var medlem i kyrkan och inte ville ha en religiös begravning, förrättas en sådan inte.
Den avlidne kan begravas i kista eller kremeras.
På många orter finns också andra religionssamfunds begravningsplatser.
I de största städerna finns till exempel ortodoxa, islamska och judiska begravningsplatser.
På många orter finns även gravområden för avlidna personer som inte har varit medlemmar i något religionssamfund.
Den avlidnes aska kan också strös ut i naturen eller i ett vattendrag om markägaren ger tillstånd till detta.
Begravningsbidrag
Den avlidne kan ibland ha rätt till begravningsbidrag (hautausavustus) genom sitt senaste anställningsförhållande eller medlemskap i ett fackförbund.
Fråga den senaste arbetsgivaren eller fackförbundet om detta.
För begravningskostnaderna för en medellös avliden kan du ansöka om utkomststöd från hemortens socialbyrå (sosiaalitoimisto).
Efter att en person dött kan dennes änka eller änkling och barn få familjepension (perhe-eläke).
Syftet med familjepensionen är att trygga de efterlevandes utkomst.
I Finland finns två olika familjepensioner, Fpa:s familjepension och arbetspensionssystemets familjepension.
Om den avlidne har arbetat eller varit företagare i Finland kan dennes efterlevande få familjepension från arbetspensionssystemet.
Båda pensionerna kan sökas hos Fpa.
Om den avlidne har bott eller arbetat utomlands en lång tid innan flytten till Finland, kan de efterlevande även ha rätt till familjepension från det landet.
Information om familjepensionfinska _ svenska _ engelska
Testamente
Vem som ärver egendomen efter en avliden person stadgas i lagen.
Du kan också själv påverka vem din förmögenhet delas till.
Du kan skriva ett testamente (testamentti), d.v.s. en skriftlig utredning över vem som ska ärva din egendom efter din bortgång.
Det är bra att ta hjälp av en jurist när du skriver ditt testamente för att det ska vara lagligt.
Bouppteckning
Bouppteckningen (perunkirjoitus) är ett möte där man upprättar en skriftlig utredning över den avlidnes förmögenhet och skulder.Bouppteckningen måste göras inom tre månader från dödsfallet.
För bouppteckningen behövs en släktutredning över den avlidne.
Det krävs även ämbetsbevis (virkatodistus), som du får från magistraten eller kyrkoherdeämbetet.
Därtill behövs uppgifter om dödsbodelägarna, det vill säga om dem som ärver den avlidnes egendom.
Bouppteckningshandlingen (perukirja) ska lämnas till skattebyrån senast en månad efter bouppteckningen.
Mer information om bouppteckningen får du från rättsväsendet och skatteförvaltningen.
Bouppteckningen ordnas av den person som bäst känner till den avlidnes egendom och skulder.
Bouppteckningshandlingen undertecknas av två personer som bedömer den avlidnes egendom.
Det är bra att anlita en jurist för upprättandet av bouppteckningen.
Att inte göra bouppteckningen inom utsatt tid kan ha ofördelaktiga följder, till exempel större arvsskatt.
Arvsskatt
Om du ärver egendom av en avliden person måste du betala arvsskatt (perintövero) för egendomen.
Skattebeloppet beror på hur stor förmögenhet du har ärvt och hur nära släkt du är till den avlidne.
Arv vilkas värde understiger 20 000 euro är skattefria.
linkkiSkatteförvaltningen:
Information om bouppteckningfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Information om arvsskattfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Information till en avlidnes anhörigfinska _ svenska
Om en person dör utanför sjukhuset ska du genast anmäla ärendet till polisen eller en läkare.
Polisen ser till att dödsorsaken fastställs och anmäler dödsfallet till Befolkningsregistercentralen (Väestörekisterikeskus).
När en person dör på sjukhuset anmäls dödsfallet automatiskt till Befolkningsregistercentralen, Fpa (Kela) och pensionsanstalter.
När en närstående person avlider kan du få stöd och hjälp med din sorg vid hälsostationerna (terveysasema), på familjerådgivningen (perheneuvola), SOS-kriscentret för utlänningar inom Föreningen för mental hälsa i Finland (Suomen mielenterveysseuran ulkomaalaisten kriisipalvelu) samt hos församlingarna.
Du får hjälp på finska och svenska, och på de flesta ställena även på engelska.
Om det behövs kan du också anlita en tolk.
När en närstående har avliditfinska _ svenska _ engelska
Information om krissituationer och sorgfinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
linkkiFöreningen för mental hälsa i Finland:
Krishjälpfinska _ svenska _ engelska
Begravningstillstånd
För att den avlidne ska kunna begravas, behövs en dödsattest (kuolintodistus) som alltid skrivs av en läkare.
Dödsattesten kan fås när dödsorsaken har fastställts.
Om det är fråga om ett akut, oklart dödsfall, en olycka eller ett brott, utförs en obduktion för att utreda dödsorsaken.
Också polisen kan undersöka orsaken till dödsfallet.
Ibland kan begravningen fördröjas på grund av att utredningen av dödsorsaken räcker länge.
Begravning
Religiösa samfund kan hjälpa dig med att ordna begravningen.
Fråga mer hos din egen samfällighet.
På webbplatsen för evangelisk-lutherska kyrkan i Finland hittar du information om kyrkans tjänster.
Man kan också ordna en civil begravning utan religiösa inslag.Om civil begravning får du information hos servicecentret Pro-Ceremonier (Pro-Seremoniat).
Begravningsbyråernas tjänster är avgiftsbelagda.
De sköter begravningsarrangemangen, som till exempel transporten av den avlidne.
Begravningsbyråerna säljer också kistor och sköter enligt avtal och de anhörigas önskemål även allt annat som rör begravningen.
Om begravningsbyråer får du information till exempel från Finlands Begravningsbyråers Förbund (Suomen Hautaustoimistojen Liitto).
Många begravningsbyråer betjänar även på engelska.
Civil begravningfinska _ svenska _ engelska
linkkiEvangelisk-lutherska kyrkan i Finland:
Information om kyrklig begravningfinska _ svenska _ engelska
Gravplats
Nästan alla begravningsplatser i Finland ägs av evangelisk-lutherska församlingar men man kan få en gravplats även om man inte är medlem i den evangelisk-lutherska kyrkan.
Gravplatserna är avgiftsbelagda och förfrågningar om dessa kan ställas till församlingarna.
Om en person inte var medlem i kyrkan och inte ville ha en religiös begravning, förrättas en sådan inte.
Den avlidne kan begravas i kista eller kremeras.
På många orter finns också andra religionssamfunds begravningsplatser.
I de största städerna finns till exempel ortodoxa, islamska och judiska begravningsplatser.
På många orter finns även gravområden för avlidna personer som inte har varit medlemmar i något religionssamfund.
Den avlidnes aska kan också strös ut i naturen eller i ett vattendrag om markägaren ger tillstånd till detta.
Begravningsbidrag
Den avlidne kan ibland ha rätt till begravningsbidrag (hautausavustus) genom sitt senaste anställningsförhållande eller medlemskap i ett fackförbund.
Fråga den senaste arbetsgivaren eller fackförbundet om detta.
För begravningskostnaderna för en medellös avliden kan du ansöka om utkomststöd från hemortens socialbyrå (sosiaalitoimisto).
Efter att en person dött kan dennes änka eller änkling och barn få familjepension (perhe-eläke).
Syftet med familjepensionen är att trygga de efterlevandes utkomst.
I Finland finns två olika familjepensioner, Fpa:s familjepension och arbetspensionssystemets familjepension.
Om den avlidne har arbetat eller varit företagare i Finland kan dennes efterlevande få familjepension från arbetspensionssystemet.
Båda pensionerna kan sökas hos Fpa.
Om den avlidne har bott eller arbetat utomlands en lång tid innan flytten till Finland, kan de efterlevande även ha rätt till familjepension från det landet.
Information om familjepensionfinska _ svenska _ engelska
Testamente
Vem som ärver egendomen efter en avliden person stadgas i lagen.
Du kan också själv påverka vem din förmögenhet delas till.
Du kan skriva ett testamente (testamentti), d.v.s. en skriftlig utredning över vem som ska ärva din egendom efter din bortgång.
Det är bra att ta hjälp av en jurist när du skriver ditt testamente för att det ska vara lagligt.
Bouppteckning
Bouppteckningen (perunkirjoitus) är ett möte där man upprättar en skriftlig utredning över den avlidnes förmögenhet och skulder.Bouppteckningen måste göras inom tre månader från dödsfallet.
För bouppteckningen behövs en släktutredning över den avlidne.
Det krävs även ämbetsbevis (virkatodistus), som du får från magistraten eller kyrkoherdeämbetet.
Därtill behövs uppgifter om dödsbodelägarna, det vill säga om dem som ärver den avlidnes egendom.
Bouppteckningshandlingen (perukirja) ska lämnas till skattebyrån senast en månad efter bouppteckningen.
Mer information om bouppteckningen får du från rättsväsendet och skatteförvaltningen.
Bouppteckningen ordnas av den person som bäst känner till den avlidnes egendom och skulder.
Bouppteckningshandlingen undertecknas av två personer som bedömer den avlidnes egendom.
Det är bra att anlita en jurist för upprättandet av bouppteckningen.
Att inte göra bouppteckningen inom utsatt tid kan ha ofördelaktiga följder, till exempel större arvsskatt.
Arvsskatt
Om du ärver egendom av en avliden person måste du betala arvsskatt (perintövero) för egendomen.
Skattebeloppet beror på hur stor förmögenhet du har ärvt och hur nära släkt du är till den avlidne.
Arv vilkas värde understiger 20 000 euro är skattefria.
linkkiSkatteförvaltningen:
Information om bouppteckningfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Information om arvsskattfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Information till en avlidnes anhörigfinska _ svenska
Du kan söka hjälp vid alkohol- och drogproblem på följande ställen:
Hälsovårdscentralen
Du kan kontakta den närmaste hälsovårdscentralen (terveysasema), om du har problem med alkohol eller droger.
A-klinikerna (A-klinikka) är vårdenheter där personer med missbruks- och beroendeproblem och deras närstående får stöd och hjälp. På A-klinikstiftelsens webbplats hittar du kontaktuppgifterna till A-kliniker runtom i Finland.
Du behöver ingen remiss till A-kliniken, utan kan själv boka en tid.
Många kliniker har även en jourtid, då man kan komma för vård utan en tidsbokning.
Tjänsterna vid A-kliniken i den egna kommunen är kostnadsfria för klienter som bor stadigvarande i Finland.
Behandlingen på A-kliniken är konfidentiell.
linkkiA-klinikstiftelsen:
Hjälp med rusmedelsberoendefinska _ engelska
Webbtjänsten Päihdelinkki
I A-klinikstiftelsens webbtjänst Päihdelinkki får du information om missbruk och beroende.
En del av tjänsterna i Päihdelinkki finns även på svenska, engelska och ryska.
linkkiDroglänken:
Information och hjälp för rusmedelsberoendefinska _ svenska _ engelska _ ryska
Anonyma Alkoholister
Anonyma Alkoholister (Anonyymit Alkoholistit) AA on är en kamratförening för män och kvinnor, där de delar med sig av sina erfarenheter av alkoholism och försöker hjälpa varandra att bli friska.
AA-grupper finns på många orter och i de större städerna finns även grupper på engelska.
Al-Anon erbjuder stöd till närstående personer till en alkoholist.
I Helsingfors finns en engelskspråkig Al-Anon-grupp.
linkkiAnonyma alkoholister, AA:
Stöd för alkoholisterfinska _ svenska _ engelska
Stöd för närstående till rusmedelsberoende personerfinska _ svenska
Anonyma narkomaner
Anonyma narkomaner (Nimettömät narkomaanit NA) erbjuder stöd och information samt gruppmöten.
Den som vill sluta använda droger kan bli medlem.
Du kan söka information om möten på webbplatsen på finska, engelska och svenska.
linkkiAnonyma Narkomaner:
Hjälp vid drogproblemfinska _ svenska _ engelska
linkkiSäg nej till droger -projektet:
Information om droger och faror som anknyter till dem särskilt för ungafinska _ somaliska _ arabiska _ kurdiska _ albanska
Du kan söka hjälp vid alkohol- och drogproblem på följande ställen:
Hälsovårdscentralen
Du kan kontakta den närmaste hälsovårdscentralen (terveysasema), om du har problem med alkohol eller droger.
A-klinikerna (A-klinikka) är vårdenheter där personer med missbruks- och beroendeproblem och deras närstående får stöd och hjälp. På A-klinikstiftelsens webbplats hittar du kontaktuppgifterna till A-kliniker runtom i Finland.
Du behöver ingen remiss till A-kliniken, utan kan själv boka en tid.
Många kliniker har även en jourtid, då man kan komma för vård utan en tidsbokning.
Tjänsterna vid A-kliniken i den egna kommunen är kostnadsfria för klienter som bor stadigvarande i Finland.
Behandlingen på A-kliniken är konfidentiell.
linkkiA-klinikstiftelsen:
Hjälp med rusmedelsberoendefinska _ engelska
Webbtjänsten Päihdelinkki
I A-klinikstiftelsens webbtjänst Päihdelinkki får du information om missbruk och beroende.
En del av tjänsterna i Päihdelinkki finns även på svenska, engelska och ryska.
linkkiDroglänken:
Information och hjälp för rusmedelsberoendefinska _ svenska _ engelska _ ryska
Anonyma Alkoholister
Anonyma Alkoholister (Anonyymit Alkoholistit) AA on är en kamratförening för män och kvinnor, där de delar med sig av sina erfarenheter av alkoholism och försöker hjälpa varandra att bli friska.
AA-grupper finns på många orter och i de större städerna finns även grupper på engelska.
Al-Anon erbjuder stöd till närstående personer till en alkoholist.
I Helsingfors finns en engelskspråkig Al-Anon-grupp.
linkkiAnonyma alkoholister, AA:
Stöd för alkoholisterfinska _ svenska _ engelska
Stöd för närstående till rusmedelsberoende personerfinska _ svenska
Anonyma narkomaner
Anonyma narkomaner (Nimettömät narkomaanit NA) erbjuder stöd och information samt gruppmöten.
Den som vill sluta använda droger kan bli medlem.
Du kan söka information om möten på webbplatsen på finska, engelska och svenska.
linkkiAnonyma Narkomaner:
Hjälp vid drogproblemfinska _ svenska _ engelska
linkkiSäg nej till droger -projektet:
Information om droger och faror som anknyter till dem särskilt för ungafinska _ somaliska _ arabiska _ kurdiska _ albanska
Du kan söka hjälp vid alkohol- och drogproblem på följande ställen:
Hälsovårdscentralen
Du kan kontakta den närmaste hälsovårdscentralen (terveysasema), om du har problem med alkohol eller droger.
A-klinikerna (A-klinikka) är vårdenheter där personer med missbruks- och beroendeproblem och deras närstående får stöd och hjälp. På A-klinikstiftelsens webbplats hittar du kontaktuppgifterna till A-kliniker runtom i Finland.
Du behöver ingen remiss till A-kliniken, utan kan själv boka en tid.
Många kliniker har även en jourtid, då man kan komma för vård utan en tidsbokning.
Tjänsterna vid A-kliniken i den egna kommunen är kostnadsfria för klienter som bor stadigvarande i Finland.
Behandlingen på A-kliniken är konfidentiell.
linkkiA-klinikstiftelsen:
Hjälp med rusmedelsberoendefinska _ engelska
Webbtjänsten Päihdelinkki
I A-klinikstiftelsens webbtjänst Päihdelinkki får du information om missbruk och beroende.
En del av tjänsterna i Päihdelinkki finns även på svenska, engelska och ryska.
linkkiDroglänken:
Information och hjälp för rusmedelsberoendefinska _ svenska _ engelska _ ryska
Anonyma Alkoholister
Anonyma Alkoholister (Anonyymit Alkoholistit) AA on är en kamratförening för män och kvinnor, där de delar med sig av sina erfarenheter av alkoholism och försöker hjälpa varandra att bli friska.
AA-grupper finns på många orter och i de större städerna finns även grupper på engelska.
Al-Anon erbjuder stöd till närstående personer till en alkoholist.
I Helsingfors finns en engelskspråkig Al-Anon-grupp.
linkkiAnonyma alkoholister, AA:
Stöd för alkoholisterfinska _ svenska _ engelska
Stöd för närstående till rusmedelsberoende personerfinska _ svenska
Anonyma narkomaner
Anonyma narkomaner (Nimettömät narkomaanit NA) erbjuder stöd och information samt gruppmöten.
Den som vill sluta använda droger kan bli medlem.
Du kan söka information om möten på webbplatsen på finska, engelska och svenska.
linkkiAnonyma Narkomaner:
Hjälp vid drogproblemfinska _ svenska _ engelska
linkkiSäg nej till droger -projektet:
Information om droger och faror som anknyter till dem särskilt för ungafinska _ somaliska _ arabiska _ kurdiska _ albanska
Människohandel är ett brott i Finland.
Människohandel är till exempel:
att tvinga någon till arbete, för vilket man betalar för lite eller ingen lön alls
att tvinga någon att sälja sex
att tvinga någon att tigga eller begå brott
att tvinga någon till äktenskap.
Den vanligaste formen av människohandel är att tvinga någon till arbete utan lön eller under annars dåliga förhållanden.
På InfoFinlands sidor Arbetstagarens rättigheter och skyldigheter samt Problem i arbetslivet hittar du information om arbetstagarens rättigheter i Finland.
Är jag offer för människohandel?
Du kan vara offer för människohandel, om
någon tvingar dig att göra saker som du inte vill göra
någon hotar dig eller din familj med våld
någon hotar med att ange dig till myndigheter om du inte gör som hen säger
någon hindrar eller övervakar dina rörelser
du inte kan fritt prata om din situation för andra.
Såväl män som kvinnor och barn kan vara offer till människohandel.
Förövarna kan vara yrkesbrottslingar men även offrets bekanta, vänner eller släktingar.
Hjälp till människohandelns offer
Människohandelns offer kan få hjälp.
Om du misstänker att du är offer för människohandel, kontakta systemet för hjälp till människohandelns offer (Ihmiskaupan uhrien auttamisjärjestelmä).
Du hittar kontaktuppgifterna på webbplatsen ihmiskauppa.fi.
Om du har tvingats att sälja sex, kan du även få hjälp vid Pro-tukipiste.
Pro-tukipiste har verksamhetsställen i Helsingfors, Tammerfors och Åbo.
Du hittar kontaktuppgifterna på Pro-tukipistes webbplats.
Hjälp till offer för människohandelfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska _ polska _ rumänska _ bulgariska
Rådgivning för personer som säljer sexuella tjänsterfinska _ engelska
Människohandel är ett brott i Finland.
Människohandel är till exempel:
att tvinga någon till arbete, för vilket man betalar för lite eller ingen lön alls
att tvinga någon att sälja sex
att tvinga någon att tigga eller begå brott
att tvinga någon till äktenskap.
Den vanligaste formen av människohandel är att tvinga någon till arbete utan lön eller under annars dåliga förhållanden.
På InfoFinlands sidor Arbetstagarens rättigheter och skyldigheter samt Problem i arbetslivet hittar du information om arbetstagarens rättigheter i Finland.
Är jag offer för människohandel?
Du kan vara offer för människohandel, om
någon tvingar dig att göra saker som du inte vill göra
någon hotar dig eller din familj med våld
någon hotar med att ange dig till myndigheter om du inte gör som hen säger
någon hindrar eller övervakar dina rörelser
du inte kan fritt prata om din situation för andra.
Såväl män som kvinnor och barn kan vara offer till människohandel.
Förövarna kan vara yrkesbrottslingar men även offrets bekanta, vänner eller släktingar.
Hjälp till människohandelns offer
Människohandelns offer kan få hjälp.
Om du misstänker att du är offer för människohandel, kontakta systemet för hjälp till människohandelns offer (Ihmiskaupan uhrien auttamisjärjestelmä).
Du hittar kontaktuppgifterna på webbplatsen ihmiskauppa.fi.
Om du har tvingats att sälja sex, kan du även få hjälp vid Pro-tukipiste.
Pro-tukipiste har verksamhetsställen i Helsingfors, Tammerfors och Åbo.
Du hittar kontaktuppgifterna på Pro-tukipistes webbplats.
Hjälp till offer för människohandelfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska _ polska _ rumänska _ bulgariska
Rådgivning för personer som säljer sexuella tjänsterfinska _ engelska
Människohandel är ett brott i Finland.
Människohandel är till exempel:
att tvinga någon till arbete, för vilket man betalar för lite eller ingen lön alls
att tvinga någon att sälja sex
att tvinga någon att tigga eller begå brott
att tvinga någon till äktenskap.
Den vanligaste formen av människohandel är att tvinga någon till arbete utan lön eller under annars dåliga förhållanden.
På InfoFinlands sidor Arbetstagarens rättigheter och skyldigheter samt Problem i arbetslivet hittar du information om arbetstagarens rättigheter i Finland.
Är jag offer för människohandel?
Du kan vara offer för människohandel, om
någon tvingar dig att göra saker som du inte vill göra
någon hotar dig eller din familj med våld
någon hotar med att ange dig till myndigheter om du inte gör som hen säger
någon hindrar eller övervakar dina rörelser
du inte kan fritt prata om din situation för andra.
Såväl män som kvinnor och barn kan vara offer till människohandel.
Förövarna kan vara yrkesbrottslingar men även offrets bekanta, vänner eller släktingar.
Hjälp till människohandelns offer
Människohandelns offer kan få hjälp.
Om du misstänker att du är offer för människohandel, kontakta systemet för hjälp till människohandelns offer (Ihmiskaupan uhrien auttamisjärjestelmä).
Du hittar kontaktuppgifterna på webbplatsen ihmiskauppa.fi.
Om du har tvingats att sälja sex, kan du även få hjälp vid Pro-tukipiste.
Pro-tukipiste har verksamhetsställen i Helsingfors, Tammerfors och Åbo.
Du hittar kontaktuppgifterna på Pro-tukipistes webbplats.
Hjälp till offer för människohandelfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska _ polska _ rumänska _ bulgariska
Rådgivning för personer som säljer sexuella tjänsterfinska _ engelska
Problem i skolan eller med studierna
Om ett barn eller en ung har problem i skolan eller med studierna är det bra att diskutera dessa med skolans eller läroanstaltens studievägledare.
I skolan arbetar även en psykolog eller en kurator.
Hen hjälper elever som har det svårt i skolan.
Om ett barn eller en ung blir mobbad i skolan är det skolans skyldighet att ingripa i detta.
Berätta om mobbning för läraren eller rektorn.
Ibland kan mobbning även vara ett brott enligt lagen, som kan anmälas till polisen.
Till exempel fysiskt våld eller stjälande är brott.
Råd vid mobbningfinska _ svenska _ engelska
Rusmedelsbruk
Om en ung har problem med alkohol, droger eller spelande, kan hen få hjälp vid ungdomsstationen.
Ungdomsstationer finns i många städer.
Den unga kan komma till ungdomsstationen ensam eller med sina föräldrar.
Kulturkonflikter hemma
Ibland kan konflikterna mellan olika kulturer skapa problem mellan barnen och föräldrarna.
Problemen kan gälla till exempel flick- och pojkvänner eller klädstilen.
Föräldrarna kan förvänta att flickor beter sig på ett annat sätt än pojkar.
Det är viktigt att kunna diskutera konflikterna inom familjen.
Den unga har rätt att veta varför föräldrarna vill att hen ska bete sig på ett visst sätt.
Ingen kultur eller religion får begränsa barns och ungas grundläggande rättigheter.
Läs mer om de grundläggande rättigheterna på InfoFinlands sida Barns och ungdomars rättigheter och skyldigheter.
Man kan be om hjälp med sina problem.
Unga flickor kan söka hjälp vid Flickornas hus som finns på många orter.
I Helsingfors finns Sopu-arbetet och i Tammerfors Didar.
De hjälper både ungdomarna och föräldrarna i hedersrelaterade konflikter.
linkkiSopu-arbetet:
Hedersrelaterade konflikterfinska _ engelska _ somaliska _ turkiska _ persiska
linkkiDidar:
Hedersrelaterade konflikterfinska _ engelska _ ryska _ somaliska _ turkiska _ persiska _ arabiska _ thai
linkkiSettlementförbundet i Finland:
Flickornas husfinska
Våld i familjen
Kroppslig bestraffning av barn är ett brott i Finland.
Detta betyder att man inte till exempel får slå eller lugga barn när de är olydiga.
Om föräldrarna utövar våld mot ett barn eller en ung, kan denne söka hjälp till exempel hos skolans hälsovårdare, vid familjerådgivningen eller FRK:s De ungas skyddshus.
På InfoFinlands sida Fostran av barn i Finland finns information om hur barn fostras i Finland.
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Brott
Ungdomar under 15 år bestraffas inte för brott.
Att begå ett brott har dock påföljder även för personer under 15 år.
Personen är skyldig att ersätta de skador som hen orsakat.
Polisen anmäler brott som begåtts av barn under 18 år till barnskyddsmyndigheten.
Mer information om barnskyddet finns på InfoFinlands sida Barnskydd.
Hjälp med fostran av barn
Familjerådgivningen
Hos familjerådgivningen får barn, unga och familjer hjälp med problem som rör fostran av barn och barns utveckling.
Du kan själv kontakta familjerådgivningen och komma överens om ett möte.
Familjerådgivningar finns på många orter.
Familjerådgivningen är en kommunal tjänst.
Du hittar kontaktuppgifterna via din hemkommuns webbplats.
Vid Väestöliitto får du information om föräldraskap.
Du kan kontakta Väestöliitto när du har funderingar kring problem i parförhållandet, fostran av barn eller skilsmässa.
Väestöliittos mångkulturella kunskapscenter stödjer invandrafamiljer.
Från kunskapscentret får du även rådgivning på telefon eller via e-post när du behöver råd om fostran av barn eller relationerna i familjen.
Du kan skriva till Väestöliittos mångkulturella kunskapscenter på dari, kurdiska (sorani), persiska, finska, ryska, engelska eller svenska.
Du hittar kontaktuppgifterna på Väestöliittos webbplats.
Stöd för mångkulturella familjerfinska _ svenska _ engelska
linkkiMannerheims barnskyddsförbund:
Stöd för barnfamiljerfinska _ svenska _ engelska
linkkiBarnombudsmannen:
Broschyren Barnets rättigheterfinska _ svenska _ engelska _ ryska
Information om barnskyddfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
Problem i skolan eller med studierna
Om ett barn eller en ung har problem i skolan eller med studierna är det bra att diskutera dessa med skolans eller läroanstaltens studievägledare.
I skolan arbetar även en psykolog eller en kurator.
Hen hjälper elever som har det svårt i skolan.
Om ett barn eller en ung blir mobbad i skolan är det skolans skyldighet att ingripa i detta.
Berätta om mobbning för läraren eller rektorn.
Ibland kan mobbning även vara ett brott enligt lagen, som kan anmälas till polisen.
Till exempel fysiskt våld eller stjälande är brott.
Råd vid mobbningfinska _ svenska _ engelska
Rusmedelsbruk
Om en ung har problem med alkohol, droger eller spelande, kan hen få hjälp vid ungdomsstationen.
Ungdomsstationer finns i många städer.
Den unga kan komma till ungdomsstationen ensam eller med sina föräldrar.
Kulturkonflikter hemma
Ibland kan konflikterna mellan olika kulturer skapa problem mellan barnen och föräldrarna.
Problemen kan gälla till exempel flick- och pojkvänner eller klädstilen.
Det kan hända att föräldrarna förväntar sig att flickor beter sig på ett annat sätt än pojkar.
Det är viktigt att kunna diskutera konflikterna inom familjen.
Den unga har rätt att veta varför föräldrarna vill att hen ska bete sig på ett visst sätt.
Ingen kultur eller religion får begränsa barns och ungas grundläggande rättigheter.
Läs mer om de grundläggande rättigheterna på InfoFinlands sida Barns och ungdomars rättigheter och skyldigheter.
Man kan be om hjälp med sina problem.
Unga flickor kan söka hjälp vid Flickornas hus som finns på många orter.
I Helsingfors och Uleåborg finns för ungdomar även Pojkarnas hus där pojkar kan söka hjälp.
I Helsingfors finns Sopu-arbetet och i Tammerfors Didar.
De hjälper både ungdomarna och föräldrarna i hedersrelaterade konflikter.
linkkiSopu-arbetet:
Hedersrelaterade konflikterfinska _ engelska _ somaliska _ turkiska _ persiska
linkkiDidar:
Hedersrelaterade konflikterfinska _ engelska _ ryska _ somaliska _ turkiska _ persiska _ arabiska _ thai
Våld i familjen
Kroppslig bestraffning av barn är ett brott i Finland.
Detta betyder att man inte till exempel får slå eller lugga barn när de är olydiga.
Om föräldrarna utövar våld mot ett barn eller en ung, kan denne söka hjälp till exempel hos skolans hälsovårdare, vid familjerådgivningen eller FRK:s De ungas skyddshus.
På InfoFinlands sida Fostran av barn i Finland finns information om hur barn fostras i Finland.
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Brott
Ungdomar under 15 år bestraffas inte för brott.
Att begå ett brott har dock påföljder även för personer under 15 år.
Personen är skyldig att ersätta de skador som hen orsakat.
Polisen anmäler brott som begåtts av barn under 18 år till föräldrarna och barnskyddsmyndigheten.
Mer information om barnskyddet finns på InfoFinlands sida Barnskydd.
Hjälp med fostran av barn
Familjerådgivningen/familjecentret
Hos familjerådgivningen eller vid familjecentret får barn, unga och familjer hjälp med problem som rör fostran av barn och barns utveckling.
Du kan själv kontakta familjerådgivningen och komma överens om ett möte.
Familjerådgivningar och familjecenter finns på många orter.
Familjerådgivningen är en kommunal tjänst.
Du hittar kontaktuppgifterna via din hemkommuns webbplats.
Mannerheims barnskyddsförbund MLL
Mannerheims barnskyddsförbund ordnar familjekaféer och barnklubbar för barnfamiljer på många orter i Finland.
Förbundet erbjuder även fostringsråd för föräldrar.
Vid Väestöliitto får du information om föräldraskap.
Du kan kontakta Väestöliitto när du har funderingar kring problem i parförhållandet, fostran av barn eller skilsmässa.
Väestöliittos mångkulturella arbete stödjer invandrafamiljer.
Vid Väestöliitto får du även rådgivning på telefon eller via e-post när du behöver råd om fostran av barn eller relationerna i familjen.
Du kan skriva till Väestöliitto på dari, kurdiska (sorani), persiska, finska, ryska, engelska eller svenska.
Du hittar kontaktuppgifterna på Väestöliittos webbplats.
Stöd för mångkulturella familjerfinska _ svenska _ engelska
linkkiMannerheims barnskyddsförbund:
Stöd för barnfamiljerfinska _ svenska _ engelska
linkkiBarnombudsmannen:
Broschyren Barnets rättigheterfinska _ svenska _ engelska _ ryska
Information om barnskyddfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
Problem i skolan eller med studierna
Om ett barn eller en ung har problem i skolan eller med studierna är det bra att diskutera dessa med skolans eller läroanstaltens studievägledare.
I skolan arbetar även en psykolog eller en kurator.
Hen hjälper elever som har det svårt i skolan.
Om ett barn eller en ung blir mobbad i skolan är det skolans skyldighet att ingripa i detta.
Berätta om mobbning för läraren eller rektorn.
Ibland kan mobbning även vara ett brott enligt lagen, som kan anmälas till polisen.
Till exempel fysiskt våld eller stjälande är brott.
Råd vid mobbningfinska _ svenska _ engelska
Rusmedelsbruk
Om en ung har problem med alkohol, droger eller spelande, kan hen få hjälp vid ungdomsstationen.
Ungdomsstationer finns i många städer.
Den unga kan komma till ungdomsstationen ensam eller med sina föräldrar.
Kulturkonflikter hemma
Ibland kan konflikterna mellan olika kulturer skapa problem mellan barnen och föräldrarna.
Problemen kan gälla till exempel flick- och pojkvänner eller klädstilen.
Det kan hända att föräldrarna förväntar sig att flickor beter sig på ett annat sätt än pojkar.
Det är viktigt att kunna diskutera konflikterna inom familjen.
Den unga har rätt att veta varför föräldrarna vill att hen ska bete sig på ett visst sätt.
Ingen kultur eller religion får begränsa barns och ungas grundläggande rättigheter.
Läs mer om de grundläggande rättigheterna på InfoFinlands sida Barns och ungdomars rättigheter och skyldigheter.
Man kan be om hjälp med sina problem.
Unga flickor kan söka hjälp vid Flickornas hus som finns på många orter.
I Helsingfors och Uleåborg finns för ungdomar även Pojkarnas hus där pojkar kan söka hjälp.
I Helsingfors finns Sopu-arbetet och i Tammerfors Didar.
De hjälper både ungdomarna och föräldrarna i hedersrelaterade konflikter.
linkkiSopu-arbetet:
Hedersrelaterade konflikterfinska _ engelska _ somaliska _ turkiska _ persiska
linkkiDidar:
Hedersrelaterade konflikterfinska _ engelska _ ryska _ somaliska _ turkiska _ persiska _ arabiska _ thai
Våld i familjen
Kroppslig bestraffning av barn är ett brott i Finland.
Detta betyder att man inte till exempel får slå eller lugga barn när de är olydiga.
Om föräldrarna utövar våld mot ett barn eller en ung, kan denne söka hjälp till exempel hos skolans hälsovårdare, vid familjerådgivningen eller FRK:s De ungas skyddshus.
På InfoFinlands sida Fostran av barn i Finland finns information om hur barn fostras i Finland.
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Brott
Ungdomar under 15 år bestraffas inte för brott.
Att begå ett brott har dock påföljder även för personer under 15 år.
Personen är skyldig att ersätta de skador som hen orsakat.
Polisen anmäler brott som begåtts av barn under 18 år till föräldrarna och barnskyddsmyndigheten.
Mer information om barnskyddet finns på InfoFinlands sida Barnskydd.
Hjälp med fostran av barn
Familjerådgivningen/familjecentret
Hos familjerådgivningen eller vid familjecentret får barn, unga och familjer hjälp med problem som rör fostran av barn och barns utveckling.
Du kan själv kontakta familjerådgivningen och komma överens om ett möte.
Familjerådgivningar och familjecenter finns på många orter.
Familjerådgivningen är en kommunal tjänst.
Du hittar kontaktuppgifterna via din hemkommuns webbplats.
Mannerheims barnskyddsförbund MLL
Mannerheims barnskyddsförbund ordnar familjekaféer och barnklubbar för barnfamiljer på många orter i Finland.
Förbundet erbjuder även fostringsråd för föräldrar.
Vid Väestöliitto får du information om föräldraskap.
Du kan kontakta Väestöliitto när du har funderingar kring problem i parförhållandet, fostran av barn eller skilsmässa.
Väestöliittos mångkulturella arbete stödjer invandrafamiljer.
Vid Väestöliitto får du även rådgivning på telefon eller via e-post när du behöver råd om fostran av barn eller relationerna i familjen.
Du kan skriva till Väestöliitto på dari, kurdiska (sorani), persiska, finska, ryska, engelska eller svenska.
Du hittar kontaktuppgifterna på Väestöliittos webbplats.
Stöd för mångkulturella familjerfinska _ svenska _ engelska
linkkiMannerheims barnskyddsförbund:
Stöd för barnfamiljerfinska _ svenska _ engelska
linkkiBarnombudsmannen:
Broschyren Barnets rättigheterfinska _ svenska _ engelska _ ryska
Information om barnskyddfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
Problem i parförhållandet
Problem i parförhållandet kan behandlas i par- och familjeterapi.
Problemen kan vara till exempel kommunikationssvårigheter, otrogenhet, eller svartsjuka, d.v.s. rädsla för att förlora den andra.
Par- och familjeterapi ges på familjerådgivningen (perheneuvola), av medlare i familjefrågor (perheasiain sovittelija), på psykiatriska polikliniker, vid Kyrkans familjerådgivningscentral (Kirkon perheasiain neuvottelukeskus) och Föreningen för mental hälsa i Finland (Suomen mielenterveysseura).
Du kan få kostnadsfri hjälp vid Kyrkans familjerådgivningscentral även på engelska och svenska, även om du inte är medlem i kyrkan.
Information om våld i familjen eller parförhållandet hittar du på InfoFinlands sida Våld.
linkkiEvangelisk-lutherska kyrkan i Finland:
Information om kyrkans familjerådgivningfinska _ svenska
Hjälp med problem i parförhållandetfinska
Information om förmedling i familjefrågorfinska _ svenska _ engelska
Skilsmässa och vårdnad om barn
Du kan lämna in ansökan om skilsmässa till tingsrätten i din egen eller din makas/makes hemkommun.
Du kan söka skilsmässa ensam eller tillsammans med din maka/make.
Ansökan om skilsmässa görs i två skeden.
När du har lämnat in din ansökan om skilsmässa till tingsrätten (käräjäoikeus) börjar en betänketid på ett halvt år.
Efter att betänketiden gått ut ska du eller ni ansöka om slutlig äktenskapsskillnad inom ett halvt år.
Skilsmässan är officiell först när den andra ansökan har godkänts.
Om du och din maka/make har minderåriga barn, kan barnens situation avgöras samtidigt som ni ansöker om skilsmässa.
Ni kan komma överens om vem som blir barnens vårdnadshavare, var barnen bor och när vardera föräldern får träffa barnen.
Samtidigt kan ni också komma överens om underhållsbidraget, d.v.s. det ekonomiska stöd som den ena föräldern betalar för barnet.
Ni kan komma överens om allt detta på egen hand eller vända er till kommunens socialbyrå (sosiaalitoimisto).
Om ditt äktenskap upphör kan du eventuellt ha behov av både psykisk och juridisk hjälp.
Juridisk hjälp kan du be om vid rättshjälpsbyrån (oikeusaputoimisto).
Psykisk hjälp vid skilsmässa kan du få till exempel i olika stödgrupper avsedda för dem som genomgått skilsmässa.
Sådan verksamhet ordnas till exempel av församlingar och organisationer.
Läs mer om vårdnaden om barn på InfoFinlands sidor Skilsmässa, Familjer med en förälder och Vad är en familj?.
linkkiRättsväsendet:
Att ansöka om skilsmässafinska _ svenska _ engelska
linkkiRättsväsendet:
Rättshjälpsbyråerfinska _ svenska _ engelska
linkkiFinlands Advokatförbund:
Advokaterfinska _ svenska _ engelska
Problem i parförhållandet
Problem i parförhållandet kan behandlas i par- och familjeterapi.
Problemen kan vara till exempel kommunikationssvårigheter, otrogenhet, eller svartsjuka, d.v.s. rädsla för att förlora den andra.
Par- och familjeterapi ges på familjerådgivningen (perheneuvola), av medlare i familjefrågor (perheasiain sovittelija), på psykiatriska polikliniker, vid Kyrkans familjerådgivningscentral (Kirkon perheasiain neuvottelukeskus) och Föreningen för mental hälsa i Finland (Suomen mielenterveysseura).
Du kan få kostnadsfri hjälp vid Kyrkans familjerådgivningscentral även på engelska och svenska, även om du inte är medlem i kyrkan.
Information om våld i familjen eller parförhållandet hittar du på InfoFinlands sida Våld.
linkkiEvangelisk-lutherska kyrkan i Finland:
Information om kyrkans familjerådgivningfinska _ svenska
Hjälp med problem i parförhållandetfinska
Information om förmedling i familjefrågorfinska _ svenska _ engelska
Skilsmässa och vårdnad om barn
Du kan lämna in ansökan om skilsmässa till tingsrätten i din egen eller din makas/makes hemkommun.
Du kan söka skilsmässa ensam eller tillsammans med din maka/make.
Ansökan om skilsmässa görs i två skeden.
När du har lämnat in din ansökan om skilsmässa till tingsrätten (käräjäoikeus) börjar en betänketid på ett halvt år.
Efter att betänketiden gått ut ska du eller ni ansöka om slutlig äktenskapsskillnad inom ett halvt år.
Skilsmässan är officiell först när den andra ansökan har godkänts.
Om du och din maka/make har minderåriga barn, kan barnens situation avgöras samtidigt som ni ansöker om skilsmässa.
Ni kan komma överens om vem som blir barnens vårdnadshavare, var barnen bor och när vardera föräldern får träffa barnen.
Samtidigt kan ni också komma överens om underhållsbidraget, d.v.s. det ekonomiska stöd som den ena föräldern betalar för barnet.
Ni kan komma överens om allt detta på egen hand eller vända er till kommunens socialbyrå (sosiaalitoimisto).
Om ditt äktenskap upphör kan du eventuellt ha behov av både psykisk och juridisk hjälp.
Juridisk hjälp kan du be om vid rättshjälpsbyrån (oikeusaputoimisto).
Psykisk hjälp vid skilsmässa kan du få till exempel i olika stödgrupper avsedda för dem som genomgått skilsmässa.
Sådan verksamhet ordnas till exempel av församlingar och organisationer.
Läs mer om vårdnaden om barn på InfoFinlands sidor Skilsmässa, Familjer med en förälder och Vad är en familj?.
linkkiRättsväsendet:
Att ansöka om skilsmässafinska _ svenska _ engelska
linkkiRättsväsendet:
Rättshjälpsbyråerfinska _ svenska _ engelska
linkkiFinlands Advokatförbund:
Advokaterfinska _ svenska _ engelska
Problem i parförhållandet
Problem i parförhållandet kan behandlas i par- och familjeterapi.
Problemen kan vara till exempel kommunikationssvårigheter, otrogenhet, eller svartsjuka, d.v.s. rädsla för att förlora den andra.
Par- och familjeterapi ges på familjerådgivningen (perheneuvola), av medlare i familjefrågor (perheasiain sovittelija), på psykiatriska polikliniker, vid Kyrkans familjerådgivningscentral (Kirkon perheasiain neuvottelukeskus) och Föreningen för mental hälsa i Finland (Suomen mielenterveysseura).
Du kan få kostnadsfri hjälp vid Kyrkans familjerådgivningscentral även på engelska och svenska, även om du inte är medlem i kyrkan.
Information om våld i familjen eller parförhållandet hittar du på InfoFinlands sida Våld.
linkkiEvangelisk-lutherska kyrkan i Finland:
Information om kyrkans familjerådgivningfinska _ svenska
Hjälp med problem i parförhållandetfinska
Information om förmedling i familjefrågorfinska _ svenska _ engelska
Skilsmässa och vårdnad om barn
Du kan lämna in ansökan om skilsmässa till tingsrätten i din egen eller din makas/makes hemkommun.
Du kan söka skilsmässa ensam eller tillsammans med din maka/make.
Ansökan om skilsmässa görs i två skeden.
När du har lämnat in din ansökan om skilsmässa till tingsrätten (käräjäoikeus) börjar en betänketid på ett halvt år.
Efter att betänketiden gått ut ska du eller ni ansöka om slutlig äktenskapsskillnad inom ett halvt år.
Skilsmässan är officiell först när den andra ansökan har godkänts.
Om du och din maka/make har minderåriga barn, kan barnens situation avgöras samtidigt som ni ansöker om skilsmässa.
Ni kan komma överens om vem som blir barnens vårdnadshavare, var barnen bor och när vardera föräldern får träffa barnen.
Samtidigt kan ni också komma överens om underhållsbidraget, d.v.s. det ekonomiska stöd som den ena föräldern betalar för barnet.
Ni kan komma överens om allt detta på egen hand eller vända er till kommunens socialbyrå (sosiaalitoimisto).
Om ditt äktenskap upphör kan du eventuellt ha behov av både psykisk och juridisk hjälp.
Juridisk hjälp kan du be om vid rättshjälpsbyrån (oikeusaputoimisto).
Psykisk hjälp vid skilsmässa kan du få till exempel i olika stödgrupper avsedda för dem som genomgått skilsmässa.
Sådan verksamhet ordnas till exempel av församlingar och organisationer.
Läs mer om vårdnaden om barn på InfoFinlands sidor Skilsmässa, Familjer med en förälder och Vad är en familj?.
linkkiRättsväsendet:
Att ansöka om skilsmässafinska _ svenska _ engelska
linkkiRättsväsendet:
Rättshjälpsbyråerfinska _ svenska _ engelska
linkkiFinlands Advokatförbund:
Advokaterfinska _ svenska _ engelska
Vad är våld?
Våld kan vara till exempel
att skrämma, följa eller observera någon
att undertrycka och tvinga
att slå, sparka och knuffa
sexuellt våld.
I Finland är våld brottsligt.
Även våld mot familjemedlemmarna är ett brott.
Barnaga, till exempel att slå barnen, är likaså ett brott.
Både offret och förövaren kan få hjälp.
Sexuellt våld
Sexuellt våld är
våldtäkt
att tvinga till sexuella handlingar
sexuellt utnyttjande
att köpa sex av barn under 18 år eller ett offer till människohandel
koppleri.
Sexuellt våld kan även förekomma i parförhållanden och äktenskap.
Sexuellt våld är alltid ett brott, även i äktenskap.
Hedersrelaterat våld
Hedersrelaterat våld är våld som syftar till att försvara familjens eller släktens heder när man misstänker att en familjemedlem kränkt familjens eller släktens heder.
I Finland är försvarandet av familjens eller släktens heder inte en godtagbar anledning till hot, påtryckningar eller våld.
Våld och hot är brott oavsett offrets och förövarens kultur.
Hedersrelaterat våld kan vara till exempel
påtryckningar
inskränkningar, till exempel ingripande i klädstil, sällskapande eller hobbyer
hot, till exempel att hota med att skicka till hemlandet
att tvinga till äktenskap eller förhindra skilsmässa.
Hjälp vid våld
När du behöver hjälp av polisen i en nödsituation, ring det allmänna nödnumret 112.
Ring inte nödnumret om det inte är en brådskande nödsituation.
Mer information om nödsituationer finns på sidan Nödsituationer.
Hjälptelefoner
Nollalinja
Tfn 080 005 005
Öppet: varje dag
Nollalinja är en hjälptelefon som du kan ringa om du har blivit utsatt för våld i familjen, sexuellt våld eller hot om våld.
Du kan ringa när som helst.
Medarbetarna pratar finska, svenska och engelska.
Samtal till Nollalinja är kostnadsfria och de syns inte i telefonräkningen.
Du behöver inte uppge ditt namn när du ringer.
Nollalinja är avsedd för både kvinnor och män.
Tfn 0800 05058
Öppet: vardagar
Kriscentret Monikas hjälptelefon är avsedd för invandrarkvinnor.
Hjälptelefonen betjänar på många olika språk.
Du kan ringa om du har blivit utsatt för våld i familjen, sexuellt våld eller hot om våld.
Samtalet är kostnadsfritt.
Du kan även kontakta Kriscentret Monika via chatten.
Chatten betjänar på finska, engelska, ryska och arabiska.
Hjälptelefonfinska _ svenska _ engelska
Hjälptelefonfinska _ engelska _ ryska _ arabiska
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Skyddshem
Om dina make eller maka eller någon annan familjemedlem utövar våld mot dig kan du ta dig till ett skyddshem (turvakoti).
I skyddshemmet är du i säkerhet och där finns personal på plats hela tiden.
Du får hjälp med att göra ett slut på våldet och råd som hjälper dig att hantera situationen.
Vistelse i skyddshemmet är kostnadsfritt.
Du kan kontakta skyddshemmet även när en familjemedlem har hotat dig med våld.
Skyddshemmet Mona är endast avsett för invandrarkvinnor och deras barn.
Ring journumret 045 639 6274 om du behöver en plats på skyddshemmet.
linkkiInstitutet för hälsa och välfärd:
Kontaktuppgifter till skyddshemfinska _ svenska
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Hjälp vid sexuellt våld
Tukinainen
Tfn 0800 97899
Tukinainen är ett kriscenter för våldtäktsoffer där du får stöd och hjälp om du har blivit utsatt för sexuellt våld.
Du får hjälp på finska och engelska.
SERI-stödcentret
Tfn 040 701 8446
I Helsingfors finns SERI-stödcentret som är avsett för offer för sexuellt våld.
SERI-stödcentret hjälper och ger råd till offer för sexuellt våld.
Centret erbjuder bland annat medicinsk undersökning och psykologhjälp.
Stödcentret betjänar alla, oavsett kön.
Du kan komma direkt till SERI-stödcentret på egen hand, men det rekommenderas att man ringer i förväg.
Du kan även alltid söka hjälp vid hälsovårdscentralen i din hemkommun.
linkkiVåldtäktskriscentralen Tukinainen:
Stöd till offer för sexuellt våldfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
SERI-stödcentretfinska _ svenska _ engelska
Hjälp vid hedersrelaterade konflikter
Om du har upplevt hedersrelaterat våld eller hot om det i din familj, kan du kontakta Sopu-arbetet.
Du hittar kontaktuppgifterna på Sopu-arbetets webbplats.
linkkiSopu-arbetet:
Hedersrelaterade konflikterfinska _ engelska _ somaliska _ turkiska _ persiska
Hjälp med att få slut på våld
Tfn 09 276 62 899
Miehen Linja är en tjänst för invandrarmän som har utövat våld eller fruktar att de kommer att utöva våld mot sin maka eller någon annan familjemedlem.
Miehen Linja betjänar på finska, engelska, svenska, franska och grekiska.
Betjäning kan även fås via tolk på det egna modersmålet.
Maria Akatemia
Tfn 09 7562 2260
Maria Akatemia hjälper kvinnor som har utövat våld eller fruktar att de kommer att utöva våld mot en familjemedlem.
Hjälp för invandrarmänfinska _ engelska
linkkiMaria Akademi:
Hjälp för kvinnor för att sluta med våldsamt beteendefinska _ svenska _ engelska
Besöksförbud
Om någon upprepade gånger hotar eller trakasserar dig och du vill ha skydd, kan du ansöka om besöksförbud (lähestymiskielto) för denna person.
Besöksförbudet innebär att personen inte får ta kontakt med dig.
Du kan ansöka om besöksförbud hos polisen eller i tingsrätten (käräjäoikeus).
Du kan fråga om råd vid socialbyrån (sosiaalitoimisto) eller rättshjälpsbyrån (oikeusaputoimisto) i din hemkommun.
Om du har bevis på hot och trakasserier är det bra att spara dem.
Information om besöksförbudfinska _ svenska _ engelska
linkkiAndra ämbetsverk:
Broschyr om besöksförbud(pdf, 418,92 kt)finska _ svenska _ engelska
Vad är våld?
Våld kan vara till exempel
att skrämma, följa eller observera någon
att undertrycka och tvinga
att slå, sparka och knuffa
sexuellt våld.
I Finland är våld brottsligt.
Även våld mot familjemedlemmarna är ett brott.
Barnaga, till exempel att slå barnen, är likaså ett brott.
Både offret och förövaren kan få hjälp.
Sexuellt våld
Sexuellt våld är
våldtäkt
att tvinga till sexuella handlingar
sexuellt utnyttjande
att köpa sex av barn under 18 år eller ett offer till människohandel
koppleri.
Sexuellt våld kan även förekomma i parförhållanden och äktenskap.
Sexuellt våld är alltid ett brott, även i äktenskap.
Hedersrelaterat våld
Hedersrelaterat våld är våld som syftar till att försvara familjens eller släktens heder när man misstänker att en familjemedlem kränkt familjens eller släktens heder.
I Finland är försvarandet av familjens eller släktens heder inte en godtagbar anledning till hot, påtryckningar eller våld.
Våld och hot är brott oavsett offrets och förövarens kultur.
Hedersrelaterat våld kan vara till exempel
påtryckningar
inskränkningar, till exempel ingripande i klädstil, sällskapande eller hobbyer
hot, till exempel att hota med att skicka till hemlandet
att tvinga till äktenskap eller förhindra skilsmässa.
Hjälp vid våld
När du behöver hjälp av polisen i en nödsituation, ring det allmänna nödnumret 112.
Ring inte nödnumret om det inte är en brådskande nödsituation.
Mer information om nödsituationer finns på sidan Nödsituationer.
Hjälptelefoner
Nollalinja
Tfn 080 005 005
Öppet: varje dag
Nollalinja är en hjälptelefon som du kan ringa om du har blivit utsatt för våld i familjen, sexuellt våld eller hot om våld.
Du kan ringa när som helst.
Medarbetarna pratar finska, svenska och engelska.
Samtal till Nollalinja är kostnadsfria och de syns inte i telefonräkningen.
Du behöver inte uppge ditt namn när du ringer.
Nollalinja är avsedd för både kvinnor och män.
Tfn 0800 05058
Öppet: vardagar
Kriscentret Monikas hjälptelefon är avsedd för invandrarkvinnor.
Hjälptelefonen betjänar på många olika språk.
Du kan ringa om du har blivit utsatt för våld i familjen, sexuellt våld eller hot om våld.
Samtalet är kostnadsfritt.
Du kan även kontakta Kriscentret Monika via chatten.
Chatten betjänar på finska, engelska, ryska och arabiska.
Hjälptelefonfinska _ svenska _ engelska
Hjälptelefonfinska _ engelska _ ryska _ arabiska
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Skyddshem
Om dina make eller maka eller någon annan familjemedlem utövar våld mot dig kan du ta dig till ett skyddshem (turvakoti).
I skyddshemmet är du i säkerhet och där finns personal på plats hela tiden.
Du får hjälp med att göra ett slut på våldet och råd som hjälper dig att hantera situationen.
Vistelse i skyddshemmet är kostnadsfritt.
Du kan kontakta skyddshemmet även när en familjemedlem har hotat dig med våld.
Skyddshemmet Mona är endast avsett för invandrarkvinnor och deras barn.
Ring journumret 045 639 6274 om du behöver en plats på skyddshemmet.
linkkiInstitutet för hälsa och välfärd:
Kontaktuppgifter till skyddshemfinska _ svenska
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Hjälp vid sexuellt våld
Tukinainen
Tfn 0800 97899
Tukinainen är ett kriscenter för våldtäktsoffer där du får stöd och hjälp om du har blivit utsatt för sexuellt våld.
Du får hjälp på finska och engelska.
SERI-stödcentret
Tfn 040 701 8446
I Helsingfors finns SERI-stödcentret som är avsett för offer för sexuellt våld.
SERI-stödcentret hjälper och ger råd till offer för sexuellt våld.
Centret erbjuder bland annat medicinsk undersökning och psykologhjälp.
Stödcentret betjänar alla, oavsett kön.
Du kan komma direkt till SERI-stödcentret på egen hand, men det rekommenderas att man ringer i förväg.
Du kan även alltid söka hjälp vid hälsovårdscentralen i din hemkommun.
linkkiVåldtäktskriscentralen Tukinainen:
Stöd till offer för sexuellt våldfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
SERI-stödcentretfinska _ svenska _ engelska
Hjälp vid hedersrelaterade konflikter
Om du har upplevt hedersrelaterat våld eller hot om det i din familj, kan du kontakta Sopu-arbetet.
Du hittar kontaktuppgifterna på Sopu-arbetets webbplats.
linkkiSopu-arbetet:
Hedersrelaterade konflikterfinska _ engelska _ somaliska _ turkiska _ persiska
Hjälp med att få slut på våld
Tfn 09 276 62 899
Miehen Linja är en tjänst för invandrarmän som har utövat våld eller fruktar att de kommer att utöva våld mot sin maka eller någon annan familjemedlem.
Miehen Linja betjänar på finska, engelska, svenska, franska och grekiska.
Betjäning kan även fås via tolk på det egna modersmålet.
Maria Akatemia
Tfn 09 7562 2260
Maria Akatemia hjälper kvinnor som har utövat våld eller fruktar att de kommer att utöva våld mot en familjemedlem.
Hjälp för invandrarmänfinska _ engelska
linkkiMaria Akademi:
Hjälp för kvinnor för att sluta med våldsamt beteendefinska _ svenska _ engelska
Besöksförbud
Om någon upprepade gånger hotar eller trakasserar dig och du vill ha skydd, kan du ansöka om besöksförbud (lähestymiskielto) för denna person.
Besöksförbudet innebär att personen inte får ta kontakt med dig.
Du kan ansöka om besöksförbud hos polisen eller i tingsrätten (käräjäoikeus).
Du kan fråga om råd vid socialbyrån (sosiaalitoimisto) eller rättshjälpsbyrån (oikeusaputoimisto) i din hemkommun.
Om du har bevis på hot och trakasserier är det bra att spara dem.
Information om besöksförbudfinska _ svenska _ engelska
linkkiAndra ämbetsverk:
Broschyr om besöksförbud(pdf, 418,92 kt)finska _ svenska _ engelska
Vad är våld?
Våld kan vara till exempel
att skrämma, följa eller observera någon
att undertrycka och tvinga
att slå, sparka och knuffa
sexuellt våld.
I Finland är våld brottsligt.
Även våld mot familjemedlemmarna är ett brott.
Barnaga, till exempel att slå barnen, är likaså ett brott.
Både offret och förövaren kan få hjälp.
Sexuellt våld
Sexuellt våld är
våldtäkt
att tvinga till sexuella handlingar
sexuellt utnyttjande
att köpa sex av barn under 18 år eller ett offer till människohandel
koppleri.
Sexuellt våld kan även förekomma i parförhållanden och äktenskap.
Sexuellt våld är alltid ett brott, även i äktenskap.
Hedersrelaterat våld
Hedersrelaterat våld är våld som syftar till att försvara familjens eller släktens heder när man misstänker att en familjemedlem kränkt familjens eller släktens heder.
I Finland är försvarandet av familjens eller släktens heder inte en godtagbar anledning till hot, påtryckningar eller våld.
Våld och hot är brott oavsett offrets och förövarens kultur.
Hedersrelaterat våld kan vara till exempel
påtryckningar
inskränkningar, till exempel ingripande i klädstil, sällskapande eller hobbyer
hot, till exempel att hota med att skicka till hemlandet
att tvinga till äktenskap eller förhindra skilsmässa.
Hjälp vid våld
När du behöver hjälp av polisen i en nödsituation, ring det allmänna nödnumret 112.
Ring inte nödnumret om det inte är en brådskande nödsituation.
Mer information om nödsituationer finns på sidan Nödsituationer.
Hjälptelefoner
Nollalinja
Tfn 080 005 005
Öppet: varje dag
Nollalinja är en hjälptelefon som du kan ringa om du har blivit utsatt för våld i familjen, sexuellt våld eller hot om våld.
Du kan ringa när som helst.
Medarbetarna pratar finska, svenska och engelska.
Samtal till Nollalinja är kostnadsfria och de syns inte i telefonräkningen.
Du behöver inte uppge ditt namn när du ringer.
Nollalinja är avsedd för både kvinnor och män.
Tfn 0800 05058
Öppet: vardagar
Kriscentret Monikas hjälptelefon är avsedd för invandrarkvinnor.
Hjälptelefonen betjänar på många olika språk.
Du kan ringa om du har blivit utsatt för våld i familjen, sexuellt våld eller hot om våld.
Samtalet är kostnadsfritt.
Du kan även kontakta Kriscentret Monika via chatten.
Chatten betjänar på finska, engelska, ryska och arabiska.
Hjälptelefonfinska _ svenska _ engelska
Hjälptelefonfinska _ engelska _ ryska _ arabiska
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Skyddshem
Om dina make eller maka eller någon annan familjemedlem utövar våld mot dig kan du ta dig till ett skyddshem (turvakoti).
I skyddshemmet är du i säkerhet och där finns personal på plats hela tiden.
Du får hjälp med att göra ett slut på våldet och råd som hjälper dig att hantera situationen.
Vistelse i skyddshemmet är kostnadsfritt.
Du kan kontakta skyddshemmet även när en familjemedlem har hotat dig med våld.
Skyddshemmet Mona är endast avsett för invandrarkvinnor och deras barn.
Ring journumret 045 639 6274 om du behöver en plats på skyddshemmet.
linkkiInstitutet för hälsa och välfärd:
Kontaktuppgifter till skyddshemfinska _ svenska
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Hjälp vid sexuellt våld
Tukinainen
Tfn 0800 97899
Tukinainen är ett kriscenter för våldtäktsoffer där du får stöd och hjälp om du har blivit utsatt för sexuellt våld.
Du får hjälp på finska och engelska.
SERI-stödcentret
Tfn 040 701 8446
I Helsingfors finns SERI-stödcentret som är avsett för offer för sexuellt våld.
SERI-stödcentret hjälper och ger råd till offer för sexuellt våld.
Centret erbjuder bland annat medicinsk undersökning och psykologhjälp.
Stödcentret betjänar alla, oavsett kön.
Du kan komma direkt till SERI-stödcentret på egen hand, men det rekommenderas att man ringer i förväg.
Du kan även alltid söka hjälp vid hälsovårdscentralen i din hemkommun.
linkkiVåldtäktskriscentralen Tukinainen:
Stöd till offer för sexuellt våldfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
SERI-stödcentretfinska _ svenska _ engelska
Hjälp vid hedersrelaterade konflikter
Om du har upplevt hedersrelaterat våld eller hot om det i din familj, kan du kontakta Sopu-arbetet.
Du hittar kontaktuppgifterna på Sopu-arbetets webbplats.
linkkiSopu-arbetet:
Hedersrelaterade konflikterfinska _ engelska _ somaliska _ turkiska _ persiska
Hjälp med att få slut på våld
Tfn 09 276 62 899
Miehen Linja är en tjänst för invandrarmän som har utövat våld eller fruktar att de kommer att utöva våld mot sin maka eller någon annan familjemedlem.
Miehen Linja betjänar på finska, engelska, svenska, franska och grekiska.
Betjäning kan även fås via tolk på det egna modersmålet.
Maria Akatemia
Tfn 09 7562 2260
Maria Akatemia hjälper kvinnor som har utövat våld eller fruktar att de kommer att utöva våld mot en familjemedlem.
Hjälp för invandrarmänfinska _ engelska
linkkiMaria Akademi:
Hjälp för kvinnor för att sluta med våldsamt beteendefinska _ svenska _ engelska
Besöksförbud
Om någon upprepade gånger hotar eller trakasserar dig och du vill ha skydd, kan du ansöka om besöksförbud (lähestymiskielto) för denna person.
Besöksförbudet innebär att personen inte får ta kontakt med dig.
Du kan ansöka om besöksförbud hos polisen eller i tingsrätten (käräjäoikeus).
Du kan fråga om råd vid socialbyrån (sosiaalitoimisto) eller rättshjälpsbyrån (oikeusaputoimisto) i din hemkommun.
Om du har bevis på hot och trakasserier är det bra att spara dem.
Information om besöksförbudfinska _ svenska _ engelska
linkkiAndra ämbetsverk:
Broschyr om besöksförbud(pdf, 418,92 kt)finska _ svenska _ engelska
I juridiska ärenden får du hjälp av en jurist.
Hen ger dig råd och ser till att dina rättigheter förverkligas.
När du söker hjälp hos en jurist, är det bra att säkerställa att juristen har sakkunskap i det område där du behöver hjälp.
Inte alla företag eller personer som erbjuder hjälp med juridiska ärenden är nödvändigtvis sakkunniga.
Offentlig rättshjälp
Juristtjänsterna är avgiftsbelagda men om du har låg eller medelhög inkomst, kan du få gratis eller delvis ersättningsgill juridisk hjälp vid statens rättshjälpsbyrå (oikeusaputoimisto).
Den offentliga rättshjälpen finns även tillgänglig på engelska och vid behov kan man använda tolktjänster.
Offentlig rättshjälp söks vid statens rättshjälpsbyråer.
Om du har en rättsskyddsförsäkring (oikeusturvavakuutus), som ersätter dina utgifter, kan du inte få offentlig rättshjälp.
Ofta ingår rättsskyddsförsäkringen i hemförsäkringen.
Rättshjälpfinska _ svenska _ engelska _ ryska _ arabiska
linkkiStatens rättshjälpsbyrå:
Information om rättshjälpfinska _ svenska _ engelska
linkkiRättsväsendet:
Rättshjälpsbyråerfinska _ svenska _ engelska
Privata jurister och advokater
Du kan söka en jurist till exempel på Finlands advokatförbunds webbplats, via tjänsten Etsi asianajaja.
Om du behöver juristens hjälp med något som har med uppehållstillstånd eller ansökan om finskt medborgarskap att göra kan du kontakta Flyktingrådgivningen som har jurister specialiserade på tillståndsärenden.
linkkiFinlands Advokatförbund:
Advokaterfinska _ svenska _ engelska
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Juridisk rådgivning
Flyktingrådgivningen
Flyktingrådgivningen (Pakolaisneuvonta) ger kostnadsfri juridisk rådgivning till asylsökande, flyktingar och andra utlänningar.
Du får rådgivning på finska och engelska.
Du kan även skicka e-post.
09 2313 9325 (mån.–fre. kl. 10–12)
Rådgivning för papperslösa utlänningar: 045 2377 104 (måndagar kl. 14–16).
Brottsofferjouren
På InfoFinlands sida Brott hittar du information om vad du kan göra om du blir utsatt för ett brott.
Broschyren Om du faller offer för ett brottfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ arabiska
linkkiBrottsofferjouren:
Juridisk rådgivning till brottsofferfinska _ svenska _ engelska
Övriga rådgivningstjänster
På InfoFinlands sida Ring och fråga om råd hittar du mer rådgivningstjänster.
I juridiska ärenden får du hjälp av en jurist.
Hen ger dig råd och ser till att dina rättigheter förverkligas.
När du söker hjälp hos en jurist, är det bra att säkerställa att juristen har sakkunskap i det område där du behöver hjälp.
Inte alla företag eller personer som erbjuder hjälp med juridiska ärenden är nödvändigtvis sakkunniga.
Offentlig rättshjälp
Juristtjänsterna är avgiftsbelagda men om du har låg eller medelhög inkomst, kan du få gratis eller delvis ersättningsgill juridisk hjälp vid statens rättshjälpsbyrå (oikeusaputoimisto).
Den offentliga rättshjälpen finns även tillgänglig på engelska och vid behov kan man använda tolktjänster.
Offentlig rättshjälp söks vid statens rättshjälpsbyråer.
Om du har en rättsskyddsförsäkring (oikeusturvavakuutus), som ersätter dina utgifter, kan du inte få offentlig rättshjälp.
Ofta ingår rättsskyddsförsäkringen i hemförsäkringen.
Rättshjälpfinska _ svenska _ engelska _ ryska _ arabiska
linkkiStatens rättshjälpsbyrå:
Information om rättshjälpfinska _ svenska _ engelska
linkkiRättsväsendet:
Rättshjälpsbyråerfinska _ svenska _ engelska
Privata jurister och advokater
Du kan söka en jurist till exempel på Finlands advokatförbunds webbplats, via tjänsten Etsi asianajaja.
Om du behöver juristens hjälp med något som har med uppehållstillstånd eller ansökan om finskt medborgarskap att göra kan du kontakta Flyktingrådgivningen som har jurister specialiserade på tillståndsärenden.
linkkiFinlands Advokatförbund:
Advokaterfinska _ svenska _ engelska
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Juridisk rådgivning
Flyktingrådgivningen
Flyktingrådgivningen (Pakolaisneuvonta) ger kostnadsfri juridisk rådgivning till asylsökande, flyktingar och andra utlänningar.
Du får rådgivning på finska och engelska.
Du kan även skicka e-post.
09 2313 9325 (mån.–fre. kl. 10–12)
Rådgivning för papperslösa utlänningar: 045 2377 104 (måndagar kl. 14–16).
Brottsofferjouren
På InfoFinlands sida Brott hittar du information om vad du kan göra om du blir utsatt för ett brott.
Broschyren Om du faller offer för ett brottfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ arabiska
linkkiBrottsofferjouren:
Juridisk rådgivning till brottsofferfinska _ svenska _ engelska
Övriga rådgivningstjänster
På InfoFinlands sida Ring och fråga om råd hittar du mer rådgivningstjänster.
I juridiska ärenden får du hjälp av en jurist.
Hen ger dig råd och ser till att dina rättigheter förverkligas.
När du söker hjälp hos en jurist, är det bra att säkerställa att juristen har sakkunskap i det område där du behöver hjälp.
Inte alla företag eller personer som erbjuder hjälp med juridiska ärenden är nödvändigtvis sakkunniga.
Offentlig rättshjälp
Juristtjänsterna är avgiftsbelagda men om du har låg eller medelhög inkomst, kan du få gratis eller delvis ersättningsgill juridisk hjälp vid statens rättshjälpsbyrå (oikeusaputoimisto).
Den offentliga rättshjälpen finns även tillgänglig på engelska och vid behov kan man använda tolktjänster.
Offentlig rättshjälp söks vid statens rättshjälpsbyråer.
Om du har en rättsskyddsförsäkring (oikeusturvavakuutus), som ersätter dina utgifter, kan du inte få offentlig rättshjälp.
Ofta ingår rättsskyddsförsäkringen i hemförsäkringen.
Rättshjälpfinska _ svenska _ engelska _ ryska _ arabiska
linkkiStatens rättshjälpsbyrå:
Information om rättshjälpfinska _ svenska _ engelska
linkkiRättsväsendet:
Rättshjälpsbyråerfinska _ svenska _ engelska
Privata jurister och advokater
Du kan söka en jurist till exempel på Finlands advokatförbunds webbplats, via tjänsten Etsi asianajaja.
Om du behöver juristens hjälp med något som har med uppehållstillstånd eller ansökan om finskt medborgarskap att göra kan du kontakta Flyktingrådgivningen som har jurister specialiserade på tillståndsärenden.
linkkiFinlands Advokatförbund:
Advokaterfinska _ svenska _ engelska
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Juridisk rådgivning
Flyktingrådgivningen
Flyktingrådgivningen (Pakolaisneuvonta) ger kostnadsfri juridisk rådgivning till asylsökande, flyktingar och andra utlänningar.
Du får rådgivning på finska och engelska.
Du kan även skicka e-post.
09 2313 9325 (mån.–fre. kl. 10–12)
Rådgivning för papperslösa utlänningar: 045 2377 104 (måndagar kl. 14–16).
Brottsofferjouren
På InfoFinlands sida Brott hittar du information om vad du kan göra om du blir utsatt för ett brott.
Broschyren Om du faller offer för ett brottfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ arabiska
linkkiBrottsofferjouren:
Juridisk rådgivning till brottsofferfinska _ svenska _ engelska
Övriga rådgivningstjänster
På InfoFinlands sida Ring och fråga om råd hittar du mer rådgivningstjänster.
Äktenskap
Registrerat parförhållande
Skilsmässa
Familjeplanering
När du är gravid
Barndagvård
Äktenskap
Före äktenskap måste man skriftligt begära prövning av äktenskapshinder.
Hindersprövningen görs på magistraten.
Begäran om prövning kan ställas på vilken magistrat som helst.
Mer information finns på magistratens webbplats.
Också borgerliga vigslar förrättas på magistraten.
Läs mer:
Samboförhållande, äktenskap och separation
Registrerat parförhållande
Parförhållandet registreras på magistraten.
Före registrering av parförhållandet måste man skriftligt begära prövning av hinder för registreringen.
Hindersprövningen görs på magistraten.
Begäran om prövning kan ställas på vilken magistrat som helst.
Mer information finns på magistratens webbplats.
Läs mer:
Registrerat parförhållande
Skilsmässa
Kvinnan eller mannen kan lämna in skilsmässoansökan på Lapplands tingsrätts kansli i Rovaniemi.
Man kan också söka skilsmässa ensam.
Ansökan kan även skickas till tingsrättens kansli per post eller via e-post.
Ett registrerat parförhållande upplöses på samma sätt som ett äktenskap.
Läs mer:
Barn vid skilsmässa
Barnatillsyningsmannens tjänster hjälper föräldrarna att vid skilsmässa komma överens om avtal som är i barnets intresse.
I tjänsten ingår hjälp under avtalsförhandlingar i fråga om vårdnaden om barnet samt dess boende, umgänge och underhåll och med att bestyrka avtalen.
Det finns även stödtjänster i grupp och en möjlighet till umgänge med stöd eller under tillsyn av barnatillsyningsmannen och till sömnskola.
Familjeplanering
Familjeplanering är helhetsbetonat främjande och upprätthållande av kvinnans och mannens sexuella hälsa.
Rådgivningsbyrån för familjeplanering ger stöd i frågor om familjeplanering och graviditetsprevention.
Tjänsten är avsedd för personer under 35 år.
De som har fyllt 35 år kan söka sig till hälsocentralläkarens mottagning i sitt eget område.
För att träffa en hälsovårdare på rådgivningsbyrån för familjeplanering krävs tidsbokning.
Läs mer:
När du är gravid
Mödrarådgivningen
Kontakta mödrarådgivningen direkt i början av graviditeten.
Målet med mödravården är att trygga bästa möjliga hälsa för den gravida modern, fostret, den nyfödda och familjen, förebygga problem under graviditeten och upptäcka dem i ett tidigt skede och vid behov anvisa till fortsatt vård.
Målet är att främja hälsan och välbefinnandet för de blivande föräldrarna och hela familjen och att stöda familjen inför deras nya uppgift som föräldrar och i växelverkan.
Läs mer:
Kontaktuppgifter till rådgivningsbyråerna
Stöd under graviditeten
Om du har rätt till moderskapsunderstöd, moderskapspenning eller andra understöd, ska du ansöka om dem vid FPA.
Du kan fylla i ansökan på Internet, skicka den till FPA per post eller besöka FPA:s kontor.
Läs mer:
InfoFinland
Stöd för den blivande modern
Barnrådgivningen
Barnrådgivningens arbete omfattar hälsofrämjande arbete, förebyggande av sjukdomar och upptäckande av dem i ett tidigt skede samt uppföljning av och stöd för barnets helhetsbetonade psykiska, fysiska och sociala utveckling.
I hälsorådgivningen beaktas hela familjen och ges särskilt stöd till den tidiga växelverkan.
Barnrådgivningens arbete omfattar barn under skolåldern och deras familjer.
På barnrådgivningsbyrån följer man barnets uppväxt och utveckling på ett helhetsbetonat sätt med regelbundna hälsokontroller.
Vaccinationer är en central del av förebyggandet av smittsamma sjukdomar hos barn. Barnrådgivningen ger barnet de vanliga vaccinationerna.
Läs mer:
Barnrådgivningen
Barndagvård
Rovaniemi stads barndagvård erbjuder dagvårdstjänster för barnfamiljer. Verksamhetsformerna och -tiderna är i linje med barnens och familjernas behov och i enlighet med lagen om barndagvård.
I Rovaniemi finns kommunala daghem och privata daghem.
I staden finns även möjlighet till mångkulturell dagvård, familjedagvård och specialdagvård.
Man kan ansöka om en plats inom den kommunala dagvården året runt.
Ansökan ska ställas fyra månader innan dagvårdsbehovet börjar.
Till dagvårdsplatser för verksamhetsåret som börjar i augusti ansöker man senast i slutet av mars.
Målet är att familjen meddelas om dagvårdsplatsen senast två veckor innan dagvården inleds.
Läs mer:
Dagvård och förskoleundervisning
Daghem
Familjedagvård
Privat dagvård och hemvårdsstöd
Om du har rätt till hemvårdsstöd kan du ansöka om det vid FPA.
Du kan fylla i ansökan på Internet eller posta den till FPA.
Du kan även besöka FPA:s kontor.
Läs mer:
Äktenskap
Registrerat parförhållande
Skilsmässa
Familjeplanering
När du är gravid
Barndagvård
Äktenskap
Före äktenskap måste man skriftligt begära prövning av äktenskapshinder.
Hindersprövningen görs på magistraten.
Begäran om prövning kan ställas på vilken magistrat som helst.
Mer information finns på magistratens webbplats.
Också borgerliga vigslar förrättas på magistraten.
Läs mer:
Samboförhållande, äktenskap och separation
Registrerat parförhållande
Parförhållandet registreras på magistraten.
Före registrering av parförhållandet måste man skriftligt begära prövning av hinder för registreringen.
Hindersprövningen görs på magistraten.
Begäran om prövning kan ställas på vilken magistrat som helst.
Mer information finns på magistratens webbplats.
Läs mer:
Registrerat parförhållande
Skilsmässa
Kvinnan eller mannen kan lämna in skilsmässoansökan på Lapplands tingsrätts kansli i Rovaniemi.
Man kan också söka skilsmässa ensam.
Ansökan kan även skickas till tingsrättens kansli per post eller via e-post.
Ett registrerat parförhållande upplöses på samma sätt som ett äktenskap.
Läs mer:
Barn vid skilsmässa
Barnatillsyningsmannens tjänster hjälper föräldrarna att vid skilsmässa komma överens om avtal som är i barnets intresse.
I tjänsten ingår hjälp under avtalsförhandlingar i fråga om vårdnaden om barnet samt dess boende, umgänge och underhåll och med att bestyrka avtalen.
Det finns även stödtjänster i grupp och en möjlighet till umgänge med stöd eller under tillsyn av barnatillsyningsmannen och till sömnskola.
Familjeplanering
Familjeplanering är helhetsbetonat främjande och upprätthållande av kvinnans och mannens sexuella hälsa.
Rådgivningsbyrån för familjeplanering ger stöd i frågor om familjeplanering och graviditetsprevention.
Tjänsten är avsedd för personer under 35 år.
De som har fyllt 35 år kan söka sig till hälsocentralläkarens mottagning i sitt eget område.
För att träffa en hälsovårdare på rådgivningsbyrån för familjeplanering krävs tidsbokning.
Läs mer:
När du är gravid
Mödrarådgivningen
Kontakta mödrarådgivningen direkt i början av graviditeten.
Målet med mödravården är att trygga bästa möjliga hälsa för den gravida modern, fostret, den nyfödda och familjen, förebygga problem under graviditeten och upptäcka dem i ett tidigt skede och vid behov anvisa till fortsatt vård.
Målet är att främja hälsan och välbefinnandet för de blivande föräldrarna och hela familjen och att stöda familjen inför deras nya uppgift som föräldrar och i växelverkan.
Läs mer:
Kontaktuppgifter till rådgivningsbyråerna
Stöd under graviditeten
Om du har rätt till moderskapsunderstöd, moderskapspenning eller andra understöd, ska du ansöka om dem vid FPA.
Du kan fylla i ansökan på Internet, skicka den till FPA per post eller besöka FPA:s kontor.
Läs mer:
InfoFinland
Stöd för den blivande modern
Barnrådgivningen
Barnrådgivningens arbete omfattar hälsofrämjande arbete, förebyggande av sjukdomar och upptäckande av dem i ett tidigt skede samt uppföljning av och stöd för barnets helhetsbetonade psykiska, fysiska och sociala utveckling.
I hälsorådgivningen beaktas hela familjen och ges särskilt stöd till den tidiga växelverkan.
Barnrådgivningens arbete omfattar barn under skolåldern och deras familjer.
På barnrådgivningsbyrån följer man barnets uppväxt och utveckling på ett helhetsbetonat sätt med regelbundna hälsokontroller.
Vaccinationer är en central del av förebyggandet av smittsamma sjukdomar hos barn. Barnrådgivningen ger barnet de vanliga vaccinationerna.
Läs mer:
Barnrådgivningen
Barndagvård
Rovaniemi stads barndagvård erbjuder dagvårdstjänster för barnfamiljer. Verksamhetsformerna och -tiderna är i linje med barnens och familjernas behov och i enlighet med lagen om barndagvård.
I Rovaniemi finns kommunala daghem och privata daghem.
I staden finns även möjlighet till mångkulturell dagvård, familjedagvård och specialdagvård.
Man kan ansöka om en plats inom den kommunala dagvården året runt.
Ansökan ska ställas fyra månader innan dagvårdsbehovet börjar.
Till dagvårdsplatser för verksamhetsåret som börjar i augusti ansöker man senast i slutet av mars.
Målet är att familjen meddelas om dagvårdsplatsen senast två veckor innan dagvården inleds.
Läs mer:
Dagvård och förskoleundervisning
Daghem
Familjedagvård
Privat dagvård och hemvårdsstöd
Om du har rätt till hemvårdsstöd kan du ansöka om det vid FPA.
Du kan fylla i ansökan på Internet eller posta den till FPA.
Du kan även besöka FPA:s kontor.
Läs mer:
Äktenskap
Registrerat parförhållande
Skilsmässa
Familjeplanering
När du är gravid
Barndagvård
Äktenskap
Före äktenskap måste man skriftligt begära prövning av äktenskapshinder.
Hindersprövningen görs på magistraten.
Begäran om prövning kan ställas på vilken magistrat som helst.
Mer information finns på magistratens webbplats.
Också borgerliga vigslar förrättas på magistraten.
Läs mer:
Samboförhållande, äktenskap och separation
Registrerat parförhållande
Parförhållandet registreras på magistraten.
Före registrering av parförhållandet måste man skriftligt begära prövning av hinder för registreringen.
Hindersprövningen görs på magistraten.
Begäran om prövning kan ställas på vilken magistrat som helst.
Mer information finns på magistratens webbplats.
Läs mer:
Registrerat parförhållande
Skilsmässa
Kvinnan eller mannen kan lämna in skilsmässoansökan på Lapplands tingsrätts kansli i Rovaniemi.
Man kan också söka skilsmässa ensam.
Ansökan kan även skickas till tingsrättens kansli per post eller via e-post.
Ett registrerat parförhållande upplöses på samma sätt som ett äktenskap.
Läs mer:
Barn vid skilsmässa
Barnatillsyningsmannens tjänster hjälper föräldrarna att vid skilsmässa komma överens om avtal som är i barnets intresse.
I tjänsten ingår hjälp under avtalsförhandlingar i fråga om vårdnaden om barnet samt dess boende, umgänge och underhåll och med att bestyrka avtalen.
Det finns även stödtjänster i grupp och en möjlighet till umgänge med stöd eller under tillsyn av barnatillsyningsmannen och till sömnskola.
Familjeplanering
Familjeplanering är helhetsbetonat främjande och upprätthållande av kvinnans och mannens sexuella hälsa.
Rådgivningsbyrån för familjeplanering ger stöd i frågor om familjeplanering och graviditetsprevention.
Tjänsten är avsedd för personer under 35 år.
De som har fyllt 35 år kan söka sig till hälsocentralläkarens mottagning i sitt eget område.
För att träffa en hälsovårdare på rådgivningsbyrån för familjeplanering krävs tidsbokning.
Läs mer:
När du är gravid
Mödrarådgivningen
Kontakta mödrarådgivningen direkt i början av graviditeten.
Målet med mödravården är att trygga bästa möjliga hälsa för den gravida modern, fostret, den nyfödda och familjen, förebygga problem under graviditeten och upptäcka dem i ett tidigt skede och vid behov anvisa till fortsatt vård.
Målet är att främja hälsan och välbefinnandet för de blivande föräldrarna och hela familjen och att stöda familjen inför deras nya uppgift som föräldrar och i växelverkan.
Läs mer:
Kontaktuppgifter till rådgivningsbyråerna
Stöd under graviditeten
Om du har rätt till moderskapsunderstöd, moderskapspenning eller andra understöd, ska du ansöka om dem vid FPA.
Du kan fylla i ansökan på Internet, skicka den till FPA per post eller besöka FPA:s kontor.
Läs mer:
InfoFinland
Stöd för den blivande modern
Barnrådgivningen
Barnrådgivningens arbete omfattar hälsofrämjande arbete, förebyggande av sjukdomar och upptäckande av dem i ett tidigt skede samt uppföljning av och stöd för barnets helhetsbetonade psykiska, fysiska och sociala utveckling.
I hälsorådgivningen beaktas hela familjen och ges särskilt stöd till den tidiga växelverkan.
Barnrådgivningens arbete omfattar barn under skolåldern och deras familjer.
På barnrådgivningsbyrån följer man barnets uppväxt och utveckling på ett helhetsbetonat sätt med regelbundna hälsokontroller.
Vaccinationer är en central del av förebyggandet av smittsamma sjukdomar hos barn. Barnrådgivningen ger barnet de vanliga vaccinationerna.
Läs mer:
Barnrådgivningen
Barndagvård
Rovaniemi stads barndagvård erbjuder dagvårdstjänster för barnfamiljer. Verksamhetsformerna och -tiderna är i linje med barnens och familjernas behov och i enlighet med lagen om barndagvård.
I Rovaniemi finns kommunala daghem och privata daghem.
I staden finns även möjlighet till mångkulturell dagvård, familjedagvård och specialdagvård.
Man kan ansöka om en plats inom den kommunala dagvården året runt.
Ansökan ska ställas fyra månader innan dagvårdsbehovet börjar.
Till dagvårdsplatser för verksamhetsåret som börjar i augusti ansöker man senast i slutet av mars.
Målet är att familjen meddelas om dagvårdsplatsen senast två veckor innan dagvården inleds.
Läs mer:
Dagvård och förskoleundervisning
Daghem
Familjedagvård
Privat dagvård och hemvårdsstöd
Om du har rätt till hemvårdsstöd kan du ansöka om det vid FPA.
Du kan fylla i ansökan på Internet eller posta den till FPA.
Du kan även besöka FPA:s kontor.
Läs mer:
Om du blir utsatt för ett brott
Om du behöver brådskande hjälp av polisen, ring nödnumret 112.
Du ska ringa nödnumret endast i brådskande fall där livet, hälsan, egendomen eller miljön är i fara.
Läs mer på InfoFinlands sida Nödsituationer.
Brottsanmälan
Var och en har rätt att anmäla till polisen ett brott som ägt rum, alltså göra en brottsanmälan.
Brottsanmälan kan göras per telefon, personligen på polisstationen eller via polisens webbplats.
Gör brottsanmälan så snabbt som möjligt.
Elektronisk polisanmälanfinska _ svenska _ engelska
Anvisning om brottsanmälanfinska _ svenska _ engelska
Broschyren Om du faller offer för ett brottfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ arabiska
Brottsofferjouren
Om du har blivit utsatt för ett brott, kan du få hjälp och råd vid Brottsofferjouren.
Du kan kontakta Brottsofferjouren per telefon eller via chatten eller besöka servicepunkten.
Brottsofferjouren erbjuder även kostnadsfri rådgivning av en jurist.
Brottsofferjouren ger även rådgivning för att motarbeta diskriminering.
Du kan kontakta rådgivningen om du tror att du har blivit utsatt för diskriminering.
Du hittar kontaktuppgifterna till Brottsofferjouren på webbplatsen.
linkkiBrottsofferjouren:
Hjälp för brottsofferfinska _ svenska _ engelska
Hjälp till brottsofferfinska _ svenska _ engelska
linkkiBrottsofferjouren:
Juridisk rådgivning till brottsofferfinska _ svenska _ engelska
Rättshjälp till brottsoffer
Rättshjälp betyder att du kan få en advokat helt eller delvis för statliga medel.
Du hittar mer information om juridisk hjälp på InfoFinlands sida Behöver du en jurist?
linkkiStatens rättshjälpsbyrå:
Information om rättshjälpfinska _ svenska _ engelska
Om du misstänks för ett brott
Om polisen misstänker att du är skyldig till ett brott, kallar den dig för förhör till polisstationen.
Om det är fråga om ett allvarligt brott, kan polisen gripa eller anhålla den brottsmisstänkta.
Även en brottsmisstänkt har rätt till juridisk hjälp.
Du hittar mer information om juridisk hjälp på InfoFinlands sida Behöver du en jurist?
Behandling av brottmål i Finland
Om polisen misstänker ett brott, inleder den en förundersökning.
När polisen är klar med förundersökningen, övergår brottmålet till åklagaren.
Åklagaren överväger om hen väcker åtal.
Om åklagaren beslutar att väcka åtal, övergår brottmålet till domstolen för behandling.
Åklagaren kan även besluta att inte väcka åtal.
När brottmålet övergår till domstolen, hålls en rättegång i tingsrätten.
Dit kallas brottsoffret, den brottsmisstänkta och vittnen.
Man måste delta i rättegången.
Vissa brottmål kan behandlas skriftligt i domstolen, och då behöver man inte delta i rättegången.
I slutet av rättegången fäller domstolen sin dom.
Inte alla brottmål behandlas i domstolen.
Ett brottmål kan även medlas, om offret och den brottsmisstänkta samtycker till detta.
Syftet med medlingen är att komma överens om hur skadan som uppstått ska ersättas.
Handläggning av brottsmål i tingsrättenfinska _ svenska _ ryska _ arabiska
Om du blir utsatt för ett brott
Om du behöver brådskande hjälp av polisen, ring nödnumret 112.
Du ska ringa nödnumret endast i brådskande fall där livet, hälsan, egendomen eller miljön är i fara.
Läs mer på InfoFinlands sida Nödsituationer.
Brottsanmälan
Var och en har rätt att anmäla till polisen ett brott som ägt rum, alltså göra en brottsanmälan.
Brottsanmälan kan göras per telefon, personligen på polisstationen eller via polisens webbplats.
Gör brottsanmälan så snabbt som möjligt.
Elektronisk polisanmälanfinska _ svenska _ engelska
Anvisning om brottsanmälanfinska _ svenska _ engelska
Broschyren Om du faller offer för ett brottfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ arabiska
Brottsofferjouren
Om du har blivit utsatt för ett brott, kan du få hjälp och råd vid Brottsofferjouren.
Du kan kontakta Brottsofferjouren per telefon eller via chatten eller besöka servicepunkten.
Brottsofferjouren erbjuder även kostnadsfri rådgivning av en jurist.
Brottsofferjouren ger även rådgivning för att motarbeta diskriminering.
Du kan kontakta rådgivningen om du tror att du har blivit utsatt för diskriminering.
Du hittar kontaktuppgifterna till Brottsofferjouren på webbplatsen.
linkkiBrottsofferjouren:
Hjälp för brottsofferfinska _ svenska _ engelska
Hjälp till brottsofferfinska _ svenska _ engelska
linkkiBrottsofferjouren:
Juridisk rådgivning till brottsofferfinska _ svenska _ engelska
Rättshjälp till brottsoffer
Rättshjälp betyder att du kan få en advokat helt eller delvis för statliga medel.
Du hittar mer information om juridisk hjälp på InfoFinlands sida Behöver du en jurist?
linkkiStatens rättshjälpsbyrå:
Information om rättshjälpfinska _ svenska _ engelska
Om du misstänks för ett brott
Om polisen misstänker att du är skyldig till ett brott, kallar den dig för förhör till polisstationen.
Om det är fråga om ett allvarligt brott, kan polisen gripa eller anhålla den brottsmisstänkta.
Även en brottsmisstänkt har rätt till juridisk hjälp.
Du hittar mer information om juridisk hjälp på InfoFinlands sida Behöver du en jurist?
Behandling av brottmål i Finland
Om polisen misstänker ett brott, inleder den en förundersökning.
När polisen är klar med förundersökningen, övergår brottmålet till åklagaren.
Åklagaren överväger om hen väcker åtal.
Om åklagaren beslutar att väcka åtal, övergår brottmålet till domstolen för behandling.
Åklagaren kan även besluta att inte väcka åtal.
När brottmålet övergår till domstolen, hålls en rättegång i tingsrätten.
Dit kallas brottsoffret, den brottsmisstänkta och vittnen.
Man måste delta i rättegången.
Vissa brottmål kan behandlas skriftligt i domstolen, och då behöver man inte delta i rättegången.
I slutet av rättegången fäller domstolen sin dom.
Inte alla brottmål behandlas i domstolen.
Ett brottmål kan även medlas, om offret och den brottsmisstänkta samtycker till detta.
Syftet med medlingen är att komma överens om hur skadan som uppstått ska ersättas.
Handläggning av brottsmål i tingsrättenfinska _ svenska _ ryska _ arabiska
Om du blir utsatt för ett brott
Om du behöver brådskande hjälp av polisen, ring nödnumret 112.
Du ska ringa nödnumret endast i brådskande fall där livet, hälsan, egendomen eller miljön är i fara.
Läs mer på InfoFinlands sida Nödsituationer.
Brottsanmälan
Var och en har rätt att anmäla till polisen ett brott som ägt rum, alltså göra en brottsanmälan.
Brottsanmälan kan göras per telefon, personligen på polisstationen eller via polisens webbplats.
Gör brottsanmälan så snabbt som möjligt.
Elektronisk polisanmälanfinska _ svenska _ engelska
Anvisning om brottsanmälanfinska _ svenska _ engelska
Broschyren Om du faller offer för ett brottfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ arabiska
Brottsofferjouren
Om du har blivit utsatt för ett brott, kan du få hjälp och råd vid Brottsofferjouren.
Du kan kontakta Brottsofferjouren per telefon eller via chatten eller besöka servicepunkten.
Brottsofferjouren erbjuder även kostnadsfri rådgivning av en jurist.
Brottsofferjouren ger även rådgivning för att motarbeta diskriminering.
Du kan kontakta rådgivningen om du tror att du har blivit utsatt för diskriminering.
Du hittar kontaktuppgifterna till Brottsofferjouren på webbplatsen.
linkkiBrottsofferjouren:
Hjälp för brottsofferfinska _ svenska _ engelska
Hjälp till brottsofferfinska _ svenska _ engelska
linkkiBrottsofferjouren:
Juridisk rådgivning till brottsofferfinska _ svenska _ engelska
Rättshjälp till brottsoffer
Rättshjälp betyder att du kan få en advokat helt eller delvis för statliga medel.
Du hittar mer information om juridisk hjälp på InfoFinlands sida Behöver du en jurist?
linkkiStatens rättshjälpsbyrå:
Information om rättshjälpfinska _ svenska _ engelska
Om du misstänks för ett brott
Om polisen misstänker att du är skyldig till ett brott, kallar den dig för förhör till polisstationen.
Om det är fråga om ett allvarligt brott, kan polisen gripa eller anhålla den brottsmisstänkta.
Även en brottsmisstänkt har rätt till juridisk hjälp.
Du hittar mer information om juridisk hjälp på InfoFinlands sida Behöver du en jurist?
Behandling av brottmål i Finland
Om polisen misstänker ett brott, inleder den en förundersökning.
När polisen är klar med förundersökningen, övergår brottmålet till åklagaren.
Åklagaren överväger om hen väcker åtal.
Om åklagaren beslutar att väcka åtal, övergår brottmålet till domstolen för behandling.
Åklagaren kan även besluta att inte väcka åtal.
När brottmålet övergår till domstolen, hålls en rättegång i tingsrätten.
Dit kallas brottsoffret, den brottsmisstänkta och vittnen.
Man måste delta i rättegången.
Vissa brottmål kan behandlas skriftligt i domstolen, och då behöver man inte delta i rättegången.
I slutet av rättegången fäller domstolen sin dom.
Inte alla brottmål behandlas i domstolen.
Ett brottmål kan även medlas, om offret och den brottsmisstänkta samtycker till detta.
Syftet med medlingen är att komma överens om hur skadan som uppstått ska ersättas.
Handläggning av brottsmål i tingsrättenfinska _ svenska _ ryska _ arabiska
Enligt Finlands lag ska alla människor behandlas likvärdigt oberoende av deras bakgrund och kön.
Diskriminering (syrjintä) är ett brott.
Vad är diskriminering?
Med diskriminering avses olikvärdig behandling, varvid personen behandlas sämre än en annan person i samma situation.
Grunden för diskriminering kan vara till exempel etniskt ursprung, nationalitet eller religion.
Det är även diskriminering att skapa en hotfull, fientlig, nedsättande eller förödmjukande atmosfär.
Ett exempel på diskriminering är om du inte får betjäning på grund av ditt etniska ursprung eller om man vid en arbetsintervju kräver att du ska behärska finska språket fullständigt trots att det inte är nödvändigt i arbetet.
Att människor behandlas på olika sätt innebär inte alltid att det är fråga om diskriminering.
Människor kan behandlas på olika sätt om det finns en godtagbar grund för detta.
Diskrimineringslagen definierar vad som är diskriminering.
Diskrimineringslagen förbjuder diskriminering på grund av ålder, ursprung, nationalitet, språk, religion, övertygelse, åsikt, politisk verksamhet, fackföreningsverksamhet, familjeförhållanden, hälsotillstånd, funktionsnedsättning, sexuell läggning eller någon annan omständighet som gäller den enskilde som person.
Ingen får missgynnas på grund av dessa omständigheter.
Jämställdhetslagen förbjuder diskriminering på grund av kön.
Information om diskrimineringfinska _ svenska _ engelska
Rasism och rasistiska brott
Rasism (rasismi) innebär att man betraktar någon människogrupp eller en person som hör till gruppen som sämre än andra till exempel på grund av etniskt ursprung, hudfärg, nationalitet, kultur, modersmål eller religion.
Med ett rasistiskt brott avses ett brott som förövaren begår av rasistiska orsaker.
Ett rasistiskt brott kan vara till exempel våld, ärekränkning, diskriminering, hot, trakasserier eller skadegörelse.
Om du blir offer för ett rasistiskt brott ska du anmäla det till polisen.
linkkiBrottsofferjouren:
Hjälp för brottsofferfinska _ svenska _ engelska
Kontaktuppgifter till polisstationernafinska _ svenska _ engelska
Hjälp till offer för diskriminering
Diskriminering på arbetsplatsen
Om du upplever diskriminering på arbetsplatsen ska du först ta kontakt med din förman.
Om du inte får hjälp av din förman ska du ta kontakt med arbetsplatsens arbetarskyddsfullmäktige (työsuojeluvaltuutettuu) eller förtroendeman (luottamusmies).
Om problemet inte blir löst på arbetsplatsen ska du ta kontakt med arbetarskyddsdistriktet (työsuojelupiirii) för ditt eget område eller ditt eget fackförbund.
linkkiArbetarskyddsförvaltningen:
Arbetarskyddfinska _ svenska _ engelska
Rådgivning för att motarbeta diskriminering
Om du misstänker att du har blivit utsatt för diskriminering, kan du kontakta Brottsofferjourens rådgivning för att motarbeta diskriminering.
Rådgivningen för att motarbeta diskriminering betjänar per telefon.
Du hittar kontaktuppgifterna till rådgivningen på Brottsofferjourens webbplats.
linkkiBrottsofferjouren:
Rådgivning för att motarbeta diskrimineringfinska _ svenska _ engelska
Diskrimineringsombudsmannen
Om du upplever diskriminering någon annanstans än på jobbet eller om du har upptäckt diskriminering någonstans kan du ta kontakt med diskrimineringsombudsmannen (yhdenvertaisuusvaltuutettu).
Du kan även ta kontakt på en annan persons eller på någon grupps vägnar.
Diskrimineringsombudsmannen är en självständig och oberoende myndighet, vars uppgift är att främja likvärdighet och ingripa i diskriminering.
Diskrimineringsombudsmannen kan ge anvisningar, råd och rekommendationer samt hjälpa med att åstadkomma förlikning i fall som gäller diskriminering.
Ombudsmannen kan även vid behov be den som misstänks för diskriminering om en redogörelse för det skedda.
Dessutom kan diskrimineringsombudsmannen föra eller hjälpa med att föra ärendet till Diskriminerings- och jämställdhetsnämnden eller inför rätten.
Möten måste avtalas på förhand.
Byråns tjänster är avgiftsfria.
Om du inte kan finska, svenska eller engelska kan du skriva e-post eller brev även på andra språk.
Du hittar kontaktuppgifterna på diskrimineringsombudsmannens webbplats.
Anmäl diskrimineringfinska _ svenska _ engelska
Diskriminerings- och jämställdhetsnämnden
Om du har blivit utsatt för diskriminering kan du även ta kontakt med diskriminerings- och jämställdhetsnämnden (yhdenvertaisuus- ja tasa-arvolautakunta.
Nämnden behandlar ansökningar som berör diskriminering och den kan förbjuda diskrimineringen.
Dessutom kan nämnden utsätta vite, vilket inskärper förbudet för diskriminering.
Nämnden kan även stöda en förlikning mellan parterna.
Nämnden behandlar inte diskrimineringsfall förknippade med arbetsförhållanden.
linkkiDiskriminerings- och jämställdhetsnämnden:
Hjälp vid diskrimineringfinska _ svenska _ engelska
Invandrarorganisationer
Om du utsätts för diskriminering eller rasism kan du få rådgivning och hjälp även av invandrarorganisationerna.
Du hittar organisationernas kontaktuppgifter på InfoFinlands sida Föreningar.
Enligt Finlands lag ska alla människor behandlas likvärdigt oberoende av deras bakgrund och kön.
Diskriminering (syrjintä) är ett brott.
Vad är diskriminering?
Med diskriminering avses olikvärdig behandling, varvid personen behandlas sämre än en annan person i samma situation.
Grunden för diskriminering kan vara till exempel etniskt ursprung, nationalitet eller religion.
Det är även diskriminering att skapa en hotfull, fientlig, nedsättande eller förödmjukande atmosfär.
Ett exempel på diskriminering är om du inte får betjäning på grund av ditt etniska ursprung eller om man vid en arbetsintervju kräver att du ska behärska finska språket fullständigt trots att det inte är nödvändigt i arbetet.
Att människor behandlas på olika sätt innebär inte alltid att det är fråga om diskriminering.
Människor kan behandlas på olika sätt om det finns en godtagbar grund för detta.
Diskrimineringslagen definierar vad som är diskriminering.
Diskrimineringslagen förbjuder diskriminering på grund av ålder, ursprung, nationalitet, språk, religion, övertygelse, åsikt, politisk verksamhet, fackföreningsverksamhet, familjeförhållanden, hälsotillstånd, funktionsnedsättning, sexuell läggning eller någon annan omständighet som gäller den enskilde som person.
Ingen får missgynnas på grund av dessa omständigheter.
Jämställdhetslagen förbjuder diskriminering på grund av kön.
Information om diskrimineringfinska _ svenska _ engelska
Rasism och rasistiska brott
Rasism (rasismi) innebär att man betraktar någon människogrupp eller en person som hör till gruppen som sämre än andra till exempel på grund av etniskt ursprung, hudfärg, nationalitet, kultur, modersmål eller religion.
Med ett rasistiskt brott avses ett brott som förövaren begår av rasistiska orsaker.
Ett rasistiskt brott kan vara till exempel våld, ärekränkning, diskriminering, hot, trakasserier eller skadegörelse.
Om du blir offer för ett rasistiskt brott ska du anmäla det till polisen.
linkkiBrottsofferjouren:
Hjälp för brottsofferfinska _ svenska _ engelska
Kontaktuppgifter till polisstationernafinska _ svenska _ engelska
Hjälp till offer för diskriminering
Diskriminering på arbetsplatsen
Om du upplever diskriminering på arbetsplatsen ska du först ta kontakt med din förman.
Om du inte får hjälp av din förman ska du ta kontakt med arbetsplatsens arbetarskyddsfullmäktige (työsuojeluvaltuutettuu) eller förtroendeman (luottamusmies).
Om problemet inte blir löst på arbetsplatsen ska du ta kontakt med arbetarskyddsdistriktet (työsuojelupiirii) för ditt eget område eller ditt eget fackförbund.
linkkiArbetarskyddsförvaltningen:
Arbetarskyddfinska _ svenska _ engelska
Rådgivning för att motarbeta diskriminering
Om du misstänker att du har blivit utsatt för diskriminering, kan du kontakta Brottsofferjourens rådgivning för att motarbeta diskriminering.
Rådgivningen för att motarbeta diskriminering betjänar per telefon.
Du hittar kontaktuppgifterna till rådgivningen på Brottsofferjourens webbplats.
linkkiBrottsofferjouren:
Rådgivning för att motarbeta diskrimineringfinska _ svenska _ engelska
Diskrimineringsombudsmannen
Om du upplever diskriminering någon annanstans än på jobbet eller om du har upptäckt diskriminering någonstans kan du ta kontakt med diskrimineringsombudsmannen (yhdenvertaisuusvaltuutettu).
Du kan även ta kontakt på en annan persons eller på någon grupps vägnar.
Diskrimineringsombudsmannen är en självständig och oberoende myndighet, vars uppgift är att främja likvärdighet och ingripa i diskriminering.
Diskrimineringsombudsmannen kan ge anvisningar, råd och rekommendationer samt hjälpa med att åstadkomma förlikning i fall som gäller diskriminering.
Ombudsmannen kan även vid behov be den som misstänks för diskriminering om en redogörelse för det skedda.
Dessutom kan diskrimineringsombudsmannen föra eller hjälpa med att föra ärendet till Diskriminerings- och jämställdhetsnämnden eller inför rätten.
Möten måste avtalas på förhand.
Byråns tjänster är avgiftsfria.
Om du inte kan finska, svenska eller engelska kan du skriva e-post eller brev även på andra språk.
Du hittar kontaktuppgifterna på diskrimineringsombudsmannens webbplats.
Anmäl diskrimineringfinska _ svenska _ engelska
Diskriminerings- och jämställdhetsnämnden
Om du har blivit utsatt för diskriminering kan du även ta kontakt med diskriminerings- och jämställdhetsnämnden (yhdenvertaisuus- ja tasa-arvolautakunta.
Nämnden behandlar ansökningar som berör diskriminering och den kan förbjuda diskrimineringen.
Dessutom kan nämnden utsätta vite, vilket inskärper förbudet för diskriminering.
Nämnden kan även stöda en förlikning mellan parterna.
Nämnden behandlar inte diskrimineringsfall förknippade med arbetsförhållanden.
linkkiDiskriminerings- och jämställdhetsnämnden:
Hjälp vid diskrimineringfinska _ svenska _ engelska
Invandrarorganisationer
Om du utsätts för diskriminering eller rasism kan du få rådgivning och hjälp även av invandrarorganisationerna.
Du hittar organisationernas kontaktuppgifter på InfoFinlands sida Föreningar.
Enligt Finlands lag ska alla människor behandlas likvärdigt oberoende av deras bakgrund och kön.
Diskriminering (syrjintä) är ett brott.
Vad är diskriminering?
Med diskriminering avses olikvärdig behandling, varvid personen behandlas sämre än en annan person i samma situation.
Grunden för diskriminering kan vara till exempel etniskt ursprung, nationalitet eller religion.
Det är även diskriminering att skapa en hotfull, fientlig, nedsättande eller förödmjukande atmosfär.
Ett exempel på diskriminering är om du inte får betjäning på grund av ditt etniska ursprung eller om man vid en arbetsintervju kräver att du ska behärska finska språket fullständigt trots att det inte är nödvändigt i arbetet.
Att människor behandlas på olika sätt innebär inte alltid att det är fråga om diskriminering.
Människor kan behandlas på olika sätt om det finns en godtagbar grund för detta.
Diskrimineringslagen definierar vad som är diskriminering.
Diskrimineringslagen förbjuder diskriminering på grund av ålder, ursprung, nationalitet, språk, religion, övertygelse, åsikt, politisk verksamhet, fackföreningsverksamhet, familjeförhållanden, hälsotillstånd, funktionsnedsättning, sexuell läggning eller någon annan omständighet som gäller den enskilde som person.
Ingen får missgynnas på grund av dessa omständigheter.
Jämställdhetslagen förbjuder diskriminering på grund av kön.
Information om diskrimineringfinska _ svenska _ engelska
Rasism och rasistiska brott
Rasism (rasismi) innebär att man betraktar någon människogrupp eller en person som hör till gruppen som sämre än andra till exempel på grund av etniskt ursprung, hudfärg, nationalitet, kultur, modersmål eller religion.
Med ett rasistiskt brott avses ett brott som förövaren begår av rasistiska orsaker.
Ett rasistiskt brott kan vara till exempel våld, ärekränkning, diskriminering, hot, trakasserier eller skadegörelse.
Om du blir offer för ett rasistiskt brott ska du anmäla det till polisen.
linkkiBrottsofferjouren:
Hjälp för brottsofferfinska _ svenska _ engelska
Kontaktuppgifter till polisstationernafinska _ svenska _ engelska
Hjälp till offer för diskriminering
Diskriminering på arbetsplatsen
Om du upplever diskriminering på arbetsplatsen ska du först ta kontakt med din förman.
Om du inte får hjälp av din förman ska du ta kontakt med arbetsplatsens arbetarskyddsfullmäktige (työsuojeluvaltuutettuu) eller förtroendeman (luottamusmies).
Om problemet inte blir löst på arbetsplatsen ska du ta kontakt med arbetarskyddsdistriktet (työsuojelupiirii) för ditt eget område eller ditt eget fackförbund.
linkkiArbetarskyddsförvaltningen:
Arbetarskyddfinska _ svenska _ engelska
Rådgivning för att motarbeta diskriminering
Om du misstänker att du har blivit utsatt för diskriminering, kan du kontakta Brottsofferjourens rådgivning för att motarbeta diskriminering.
Rådgivningen för att motarbeta diskriminering betjänar per telefon.
Du hittar kontaktuppgifterna till rådgivningen på Brottsofferjourens webbplats.
linkkiBrottsofferjouren:
Rådgivning för att motarbeta diskrimineringfinska _ svenska _ engelska
Diskrimineringsombudsmannen
Om du upplever diskriminering någon annanstans än på jobbet eller om du har upptäckt diskriminering någonstans kan du ta kontakt med diskrimineringsombudsmannen (yhdenvertaisuusvaltuutettu).
Du kan även ta kontakt på en annan persons eller på någon grupps vägnar.
Diskrimineringsombudsmannen är en självständig och oberoende myndighet, vars uppgift är att främja likvärdighet och ingripa i diskriminering.
Diskrimineringsombudsmannen kan ge anvisningar, råd och rekommendationer samt hjälpa med att åstadkomma förlikning i fall som gäller diskriminering.
Ombudsmannen kan även vid behov be den som misstänks för diskriminering om en redogörelse för det skedda.
Dessutom kan diskrimineringsombudsmannen föra eller hjälpa med att föra ärendet till Diskriminerings- och jämställdhetsnämnden eller inför rätten.
Möten måste avtalas på förhand.
Byråns tjänster är avgiftsfria.
Om du inte kan finska, svenska eller engelska kan du skriva e-post eller brev även på andra språk.
Du hittar kontaktuppgifterna på diskrimineringsombudsmannens webbplats.
Anmäl diskrimineringfinska _ svenska _ engelska
Diskriminerings- och jämställdhetsnämnden
Om du har blivit utsatt för diskriminering kan du även ta kontakt med diskriminerings- och jämställdhetsnämnden (yhdenvertaisuus- ja tasa-arvolautakunta.
Nämnden behandlar ansökningar som berör diskriminering och den kan förbjuda diskrimineringen.
Dessutom kan nämnden utsätta vite, vilket inskärper förbudet för diskriminering.
Nämnden kan även stöda en förlikning mellan parterna.
Nämnden behandlar inte diskrimineringsfall förknippade med arbetsförhållanden.
linkkiDiskriminerings- och jämställdhetsnämnden:
Hjälp vid diskrimineringfinska _ svenska _ engelska
Invandrarorganisationer
Om du utsätts för diskriminering eller rasism kan du få rådgivning och hjälp även av invandrarorganisationerna.
Du hittar organisationernas kontaktuppgifter på InfoFinlands sida Föreningar.
Om du inte kan betala dina räkningar
Om du har en räkning som du inte kan betala, kontakta avsändaren direkt.
Ofta kan du få betalningstiden förlängd.
Då läggs vanligtvis en liten förseningsavgift på räkningen.
Om du inte betalar räkningen senast på förfallodagen eller inte har kommit överens om att förlänga betalningstiden, måste du betala påminnelse- och inkassokostnader samt dröjsmålsränta.
Inkasso
Om du inte har betalat en räkning senast på förfallodagen får du en betalningspåminnelse.
Efter en eller två påminnelser kan räkningen övergå till en inkassobyrå.
Inkassobyrån skickar dig genast ett betalningskrav.
Om du inte kan betala räkningen på en gång, ska du kontakta inkassobyrån och komma överens om en betalningsplan för räkningen.
Om du inte betalar räkningen eller kommer överens om en betalningsplan kan skulden slutligen gå till utmätning (ulosotto).
Utmätning betyder att myndigheten har rätt att ta en del av dina inkomster för betalning av skulder.
Utmätningsmyndigheten kan även sälja värdefull egendom som du har för att betala skulden.
Ofta behövs ett domstolsbeslut för utmätning.
Vissa betalningar går emellertid direkt till utmätning.
Sådana betalningar är till exempel skatter, hälscentralsavgifter och dagvårdsavgifter.
Betalningsanmärkning
Om du inte betalar en räkning eller en skuld, kan du få en betalningsanmärkning (maksuhäiriömerkintä) i kreditupplysningsregistret.
Detta orsakar många svårigheter för dig.
Hyresvärdar och banker kontrollerar ofta kredituppgifterna i kreditupplysningsregistret.
Om du har en betalningsanmärkning, får du inte nödvändigtvis en hyresbostad, ett banklån eller ett kreditkort.
Även arbetsgivaren kan förutsätta att arbetstagaren inte har betalningsanmärkningar.
linkkiKonkurrens- och konsumentverket:
Information om anmärkning om betalningsstörningfinska _ svenska _ engelska
linkkiRättsväsendet:
Information om utsökningfinska _ svenska _ engelska
Om du inte kan betala din hyra
Hyresvärden har rätt att häva hyresavtalet om du inte betalar din hyra.
Hyresvärden ska meddela hyresgästen om hävandet.
I detta skede finns det vanligtvis ännu en möjlighet att komma överens om hyresbetalningen med hyresvärden.
Om du inte betalar din hyra kan hyresvärden söka ett avhysningsbeslut i domstol.
Det innebär att du måste flytta ut ur bostaden och betala de obetalda hyrorna.
Om du har svårigheter att betala hyran för din bostad ska du ta kontakt med hyresvärden.
Försök att komma överens om att få mer tid på dig att betala.
Du kan även fråga om råd på socialbyrån i din hemkommun.
Kontrollera också om du till exempel har rätt till bostadsbidrag eller utkomststöd.
Din rätt till bostadsbidrag och utkomststöd kan du få reda på hos FPA.
Information om bostadsbidrag finns på InfoFinlands sida Bostadsbidrag.
Hjälp vid ekonomiska problem
Sociala förmåner
Kontrollera att du har ansökt om alla sociala förmåner som du har rätt att få.
Dessa kan vara till exempel arbetslöshetsförsäkring, bostadsbidrag, studiestöd och ekonomiska understöd för barnfamiljer.
Utkomststöd
Om du eller din familj inte har tillräckliga inkomster eller tillgångar för den nödvändiga dagliga försörjningen kan du söka grundläggande utkomststöd (perustoimeentulotuki) hos FPA.
Med den nödvändiga dagliga försörjningen avses skäliga utgifter till exempel för mat, kläder, hälsovård och boende.
Det grundläggande utkomststödet täcker även utgifter för hobby- och rekreationsverksamhet, avgifterna för barndagvård och för skolbarns morgon- och eftermiddagsverksamhet samt nödvändiga kostnader för flytt.
Betalningen av utkomststöd påverkas av alla dina inkomster och tillgångar.
I kalkylen beaktas även de sociala förmåner som du får till exempel av FPA, en arbetspensionsförsäkring eller arbetslöshetskassan.
Innan du ansöker om utkomststöd ska du ansöka om de andra bidragen som du har rätt till (till exempel arbetslöshetsförsäkring, bostadsbidrag, pension, studiestöd, föräldradagpenning, sjukdagpenning, hemvårdsstöd eller underhållsstöd).
Utkomststödet är avsett som en tillfällig hjälp.
Utkomststöd betalas endast om du inte kan få några andra inkomster och bidrag eller om dina övriga inkomster inte räcker till för de nödvändiga utgifterna.
Om du eller din familj har utgifter på grund av särskilda behov, för vilka du inte kan få grundläggande utkomststöd, kan socialbyrån i din hemkommun bevilja kompletterande och förebyggande utkomststöd (täydentävä ja ehkäisevä toimeentulotuki).
Du kan få kompletterande utkomststöd till exempel för att trygga ditt boende eller om din ekonomiska situation oväntat försämrats.
Syftet med det kompletterande och förebyggande utkomststödet är att hjälpa personen att klara sig självständigt och att förebygga utslagning.
Du ska alltid först ansöka om grundläggande utkomststöd hos FPA.
I samma ansökan kan du ange om du också behöver kompletterande eller förebyggande utkomststöd.
FPA kan på din begäran föra över din ansökan om kompletterande och förebyggande utkomststöd till kommunen för behandling.
Vid behov får du rådgivning om hur du ansöker om utkomststödet hos FPA, socialbyrån i din hemkommun eller en rådgivning för invandrare.
Information om utkomststödfinska _ svenska _ engelska _ ryska _ estniska
Rådgivning och hjälp med ekonomin
Om du har problem med att betala räkningar och skulder, kontakta ekonomi- och skuldrådgivningen (talous- ja velkaneuvonta).
Ekonomi- och skuldrådgivning ordnas av kommuner.
Rådgivningen år kostnadsfri.
Hos Takuusäätiö kan du få hjälp och råd med betalningen av skulder.
Stiftelsen kan hjälpa dig att slå ihop dina skulder till ett lån.
Du kan ansöka om lånegaranti vid Takuusäätiö om du behöver ett banklån för att betala dina skulder.
Vid Takuusäätiö kan du även ansöka om ett litet lån, om du behöver pengar för en utgift av engångskaraktär, såsom en hushållsmaskin, möbler, hyresdeposition, reparation av bilen eller glasögon.
Velkalinja är Takuusäätiös kostnadsfria rådgivningstelefon.
Rådgivningsnumret 0800 9 8009 betjänar på finska och vid behov även på engelska eller svenska.
I nödfall, om du till exempel inte har pengar för mat, kan du även kontakta diakoniarbetaren i din församling.
Du hittar kontaktuppgifterna vid din församling.
linkkiKonkurrens- och konsumentverket:
Ekonomi- och skuldrådgivarefinska _ svenska _ engelska
linkkiGaranti-Stiftelsen:
Hjälp med ekonomiska problemfinska _ svenska _ engelska
linkkiKonkurrens- och konsumentverket:
Information om ekonominfinska _ svenska _ engelska
Spelberoende
Om dina ekonomiska problem beror på spelproblem är det bäst att söka hjälp.
Du får hjälp med spelproblem vid A-kliniker (A-klinikka), mentalvårdsbyråer (mielenterveystoimisto) och hälsovårdscentralen (terveyskeskus).
På vissa orter kan även socialbyrån (sosiaalitoimisto) eller församlingarna hjälpa.
Även de anhöriga till en spelberoende person kan få hjälp.
Du kan också söka hjälp för ditt spelproblem vid olika organisationer.
I webbtjänsten Droglänken (Päihdelinkki) finns mycket information om spelproblem på flera språk.
Peluuri är en hjälptelefon för personer med spelproblem, deras närstående och andra som möter spelproblem.
Hjälptelefonen nås på numret 0800 100 101.
Betjäning ges på finska och svenska samt i mån av möjlighet även på engelska.
Peluuri finns även på internet.
linkkiDroglänken:
Information om spelproblemfinska _ svenska _ engelska _ ryska
Hjälp och information till spelberoende och deras anhörigafinska _ svenska _ engelska
Om du inte kan betala dina räkningar
Om du har en räkning som du inte kan betala, kontakta avsändaren direkt.
Ofta kan du få betalningstiden förlängd.
Då läggs vanligtvis en liten förseningsavgift på räkningen.
Om du inte betalar räkningen senast på förfallodagen eller inte har kommit överens om att förlänga betalningstiden, måste du betala påminnelse- och inkassokostnader samt dröjsmålsränta.
Inkasso
Om du inte har betalat en räkning senast på förfallodagen får du en betalningspåminnelse.
Efter en eller två påminnelser kan räkningen övergå till en inkassobyrå.
Inkassobyrån skickar dig genast ett betalningskrav.
Om du inte kan betala räkningen på en gång, ska du kontakta inkassobyrån och komma överens om en betalningsplan för räkningen.
Om du inte betalar räkningen eller kommer överens om en betalningsplan kan skulden slutligen gå till utmätning (ulosotto).
Utmätning betyder att myndigheten har rätt att ta en del av dina inkomster för betalning av skulder.
Utmätningsmyndigheten kan även sälja värdefull egendom som du har för att betala skulden.
Ofta behövs ett domstolsbeslut för utmätning.
Vissa betalningar går emellertid direkt till utmätning.
Sådana betalningar är till exempel skatter, hälscentralsavgifter och dagvårdsavgifter.
Betalningsanmärkning
Om du inte betalar en räkning eller en skuld, kan du få en betalningsanmärkning (maksuhäiriömerkintä) i kreditupplysningsregistret.
Detta orsakar många svårigheter för dig.
Hyresvärdar och banker kontrollerar ofta kredituppgifterna i kreditupplysningsregistret.
Om du har en betalningsanmärkning, får du inte nödvändigtvis en hyresbostad, ett banklån eller ett kreditkort.
Även arbetsgivaren kan förutsätta att arbetstagaren inte har betalningsanmärkningar.
linkkiKonkurrens- och konsumentverket:
Information om anmärkning om betalningsstörningfinska _ svenska _ engelska
linkkiRättsväsendet:
Information om utsökningfinska _ svenska _ engelska
Om du inte kan betala din hyra
Hyresvärden har rätt att häva hyresavtalet om du inte betalar din hyra.
Hyresvärden ska meddela hyresgästen om hävandet.
I detta skede finns det vanligtvis ännu en möjlighet att komma överens om hyresbetalningen med hyresvärden.
Om du inte betalar din hyra kan hyresvärden söka ett avhysningsbeslut i domstol.
Det innebär att du måste flytta ut ur bostaden och betala de obetalda hyrorna.
Om du har svårigheter att betala hyran för din bostad ska du ta kontakt med hyresvärden.
Försök att komma överens om att få mer tid på dig att betala.
Du kan även fråga om råd på socialbyrån i din hemkommun.
Kontrollera också om du till exempel har rätt till bostadsbidrag eller utkomststöd.
Din rätt till bostadsbidrag och utkomststöd kan du få reda på hos FPA.
Information om bostadsbidrag finns på InfoFinlands sida Bostadsbidrag.
Hjälp vid ekonomiska problem
Sociala förmåner
Kontrollera att du har ansökt om alla sociala förmåner som du har rätt att få.
Dessa kan vara till exempel arbetslöshetsförsäkring, bostadsbidrag, studiestöd och ekonomiska understöd för barnfamiljer.
Utkomststöd
Om du eller din familj inte har tillräckliga inkomster eller tillgångar för den nödvändiga dagliga försörjningen kan du söka grundläggande utkomststöd (perustoimeentulotuki) hos FPA.
Med den nödvändiga dagliga försörjningen avses skäliga utgifter till exempel för mat, kläder, hälsovård och boende.
Det grundläggande utkomststödet täcker även utgifter för hobby- och rekreationsverksamhet, avgifterna för barndagvård och för skolbarns morgon- och eftermiddagsverksamhet samt nödvändiga kostnader för flytt.
Betalningen av utkomststöd påverkas av alla dina inkomster och tillgångar.
I kalkylen beaktas även de sociala förmåner som du får till exempel av FPA, en arbetspensionsförsäkring eller arbetslöshetskassan.
Innan du ansöker om utkomststöd ska du ansöka om de andra bidragen som du har rätt till (till exempel arbetslöshetsförsäkring, bostadsbidrag, pension, studiestöd, föräldradagpenning, sjukdagpenning, hemvårdsstöd eller underhållsstöd).
Utkomststödet är avsett som en tillfällig hjälp.
Utkomststöd betalas endast om du inte kan få några andra inkomster och bidrag eller om dina övriga inkomster inte räcker till för de nödvändiga utgifterna.
Om du eller din familj har utgifter på grund av särskilda behov, för vilka du inte kan få grundläggande utkomststöd, kan socialbyrån i din hemkommun bevilja kompletterande och förebyggande utkomststöd (täydentävä ja ehkäisevä toimeentulotuki).
Du kan få kompletterande utkomststöd till exempel för att trygga ditt boende eller om din ekonomiska situation oväntat försämrats.
Syftet med det kompletterande och förebyggande utkomststödet är att hjälpa personen att klara sig självständigt och att förebygga utslagning.
Du ska alltid först ansöka om grundläggande utkomststöd hos FPA.
I samma ansökan kan du ange om du också behöver kompletterande eller förebyggande utkomststöd.
FPA kan på din begäran föra över din ansökan om kompletterande och förebyggande utkomststöd till kommunen för behandling.
Vid behov får du rådgivning om hur du ansöker om utkomststödet hos FPA, socialbyrån i din hemkommun eller en rådgivning för invandrare.
Information om utkomststödfinska _ svenska _ engelska _ ryska _ estniska
Rådgivning och hjälp med ekonomin
Om du har problem med att betala räkningar och skulder, kontakta ekonomi- och skuldrådgivningen (talous- ja velkaneuvonta).
Ekonomi- och skuldrådgivning ordnas av kommuner.
Rådgivningen år kostnadsfri.
Hos Takuusäätiö kan du få hjälp och råd med betalningen av skulder.
Stiftelsen kan hjälpa dig att slå ihop dina skulder till ett lån.
Du kan ansöka om lånegaranti vid Takuusäätiö om du behöver ett banklån för att betala dina skulder.
Vid Takuusäätiö kan du även ansöka om ett litet lån, om du behöver pengar för en utgift av engångskaraktär, såsom en hushållsmaskin, möbler, hyresdeposition, reparation av bilen eller glasögon.
Velkalinja är Takuusäätiös kostnadsfria rådgivningstelefon.
Rådgivningsnumret 0800 9 8009 betjänar på finska och vid behov även på engelska eller svenska.
I nödfall, om du till exempel inte har pengar för mat, kan du även kontakta diakoniarbetaren i din församling.
Du hittar kontaktuppgifterna vid din församling.
linkkiKonkurrens- och konsumentverket:
Ekonomi- och skuldrådgivarefinska _ svenska _ engelska
linkkiGaranti-Stiftelsen:
Hjälp med ekonomiska problemfinska _ svenska _ engelska
linkkiKonkurrens- och konsumentverket:
Information om ekonominfinska _ svenska _ engelska
Spelberoende
Om dina ekonomiska problem beror på spelproblem är det bäst att söka hjälp.
Du får hjälp med spelproblem vid A-kliniker (A-klinikka), mentalvårdsbyråer (mielenterveystoimisto) och hälsovårdscentralen (terveyskeskus).
På vissa orter kan även socialbyrån (sosiaalitoimisto) eller församlingarna hjälpa.
Även de anhöriga till en spelberoende person kan få hjälp.
Du kan också söka hjälp för ditt spelproblem vid olika organisationer.
I webbtjänsten Droglänken (Päihdelinkki) finns mycket information om spelproblem på flera språk.
Peluuri är en hjälptelefon för personer med spelproblem, deras närstående och andra som möter spelproblem.
Hjälptelefonen nås på numret 0800 100 101.
Betjäning ges på finska och svenska samt i mån av möjlighet även på engelska.
Peluuri finns även på internet.
linkkiDroglänken:
Information om spelproblemfinska _ svenska _ engelska _ ryska
Hjälp och information till spelberoende och deras anhörigafinska _ svenska _ engelska
Om du inte kan betala dina räkningar
Om du har en räkning som du inte kan betala, kontakta avsändaren direkt.
Ofta kan du få betalningstiden förlängd.
Då läggs vanligtvis en liten förseningsavgift på räkningen.
Om du inte betalar räkningen senast på förfallodagen eller inte har kommit överens om att förlänga betalningstiden, måste du betala påminnelse- och inkassokostnader samt dröjsmålsränta.
Inkasso
Om du inte har betalat en räkning senast på förfallodagen får du en betalningspåminnelse.
Efter en eller två påminnelser kan räkningen övergå till en inkassobyrå.
Inkassobyrån skickar dig genast ett betalningskrav.
Om du inte kan betala räkningen på en gång, ska du kontakta inkassobyrån och komma överens om en betalningsplan för räkningen.
Om du inte betalar räkningen eller kommer överens om en betalningsplan kan skulden slutligen gå till utmätning (ulosotto).
Utmätning betyder att myndigheten har rätt att ta en del av dina inkomster för betalning av skulder.
Utmätningsmyndigheten kan även sälja värdefull egendom som du har för att betala skulden.
Ofta behövs ett domstolsbeslut för utmätning.
Vissa betalningar går emellertid direkt till utmätning.
Sådana betalningar är till exempel skatter, hälscentralsavgifter och dagvårdsavgifter.
Betalningsanmärkning
Om du inte betalar en räkning eller en skuld, kan du få en betalningsanmärkning (maksuhäiriömerkintä) i kreditupplysningsregistret.
Detta orsakar många svårigheter för dig.
Hyresvärdar och banker kontrollerar ofta kredituppgifterna i kreditupplysningsregistret.
Om du har en betalningsanmärkning, får du inte nödvändigtvis en hyresbostad, ett banklån eller ett kreditkort.
Även arbetsgivaren kan förutsätta att arbetstagaren inte har betalningsanmärkningar.
linkkiKonkurrens- och konsumentverket:
Information om anmärkning om betalningsstörningfinska _ svenska _ engelska
linkkiRättsväsendet:
Information om utsökningfinska _ svenska _ engelska
Om du inte kan betala din hyra
Hyresvärden har rätt att häva hyresavtalet om du inte betalar din hyra.
Hyresvärden ska meddela hyresgästen om hävandet.
I detta skede finns det vanligtvis ännu en möjlighet att komma överens om hyresbetalningen med hyresvärden.
Om du inte betalar din hyra kan hyresvärden söka ett avhysningsbeslut i domstol.
Det innebär att du måste flytta ut ur bostaden och betala de obetalda hyrorna.
Om du har svårigheter att betala hyran för din bostad ska du ta kontakt med hyresvärden.
Försök att komma överens om att få mer tid på dig att betala.
Du kan även fråga om råd på socialbyrån i din hemkommun.
Kontrollera också om du till exempel har rätt till bostadsbidrag eller utkomststöd.
Din rätt till bostadsbidrag och utkomststöd kan du få reda på hos FPA.
Information om bostadsbidrag finns på InfoFinlands sida Bostadsbidrag.
Hjälp vid ekonomiska problem
Sociala förmåner
Kontrollera att du har ansökt om alla sociala förmåner som du har rätt att få.
Dessa kan vara till exempel arbetslöshetsförsäkring, bostadsbidrag, studiestöd och ekonomiska understöd för barnfamiljer.
Utkomststöd
Om du eller din familj inte har tillräckliga inkomster eller tillgångar för den nödvändiga dagliga försörjningen kan du söka grundläggande utkomststöd (perustoimeentulotuki) hos FPA.
Med den nödvändiga dagliga försörjningen avses skäliga utgifter till exempel för mat, kläder, hälsovård och boende.
Det grundläggande utkomststödet täcker även utgifter för hobby- och rekreationsverksamhet, avgifterna för barndagvård och för skolbarns morgon- och eftermiddagsverksamhet samt nödvändiga kostnader för flytt.
Betalningen av utkomststöd påverkas av alla dina inkomster och tillgångar.
I kalkylen beaktas även de sociala förmåner som du får till exempel av FPA, en arbetspensionsförsäkring eller arbetslöshetskassan.
Innan du ansöker om utkomststöd ska du ansöka om de andra bidragen som du har rätt till (till exempel arbetslöshetsförsäkring, bostadsbidrag, pension, studiestöd, föräldradagpenning, sjukdagpenning, hemvårdsstöd eller underhållsstöd).
Utkomststödet är avsett som en tillfällig hjälp.
Utkomststöd betalas endast om du inte kan få några andra inkomster och bidrag eller om dina övriga inkomster inte räcker till för de nödvändiga utgifterna.
Om du eller din familj har utgifter på grund av särskilda behov, för vilka du inte kan få grundläggande utkomststöd, kan socialbyrån i din hemkommun bevilja kompletterande och förebyggande utkomststöd (täydentävä ja ehkäisevä toimeentulotuki).
Du kan få kompletterande utkomststöd till exempel för att trygga ditt boende eller om din ekonomiska situation oväntat försämrats.
Syftet med det kompletterande och förebyggande utkomststödet är att hjälpa personen att klara sig självständigt och att förebygga utslagning.
Du ska alltid först ansöka om grundläggande utkomststöd hos FPA.
I samma ansökan kan du ange om du också behöver kompletterande eller förebyggande utkomststöd.
FPA kan på din begäran föra över din ansökan om kompletterande och förebyggande utkomststöd till kommunen för behandling.
Vid behov får du rådgivning om hur du ansöker om utkomststödet hos FPA, socialbyrån i din hemkommun eller en rådgivning för invandrare.
Information om utkomststödfinska _ svenska _ engelska _ ryska _ estniska
Rådgivning och hjälp med ekonomin
Om du har problem med att betala räkningar och skulder, kontakta ekonomi- och skuldrådgivningen (talous- ja velkaneuvonta).
Ekonomi- och skuldrådgivning ordnas av kommuner.
Rådgivningen år kostnadsfri.
Hos Takuusäätiö kan du få hjälp och råd med betalningen av skulder.
Stiftelsen kan hjälpa dig att slå ihop dina skulder till ett lån.
Du kan ansöka om lånegaranti vid Takuusäätiö om du behöver ett banklån för att betala dina skulder.
Vid Takuusäätiö kan du även ansöka om ett litet lån, om du behöver pengar för en utgift av engångskaraktär, såsom en hushållsmaskin, möbler, hyresdeposition, reparation av bilen eller glasögon.
Velkalinja är Takuusäätiös kostnadsfria rådgivningstelefon.
Rådgivningsnumret 0800 9 8009 betjänar på finska och vid behov även på engelska eller svenska.
I nödfall, om du till exempel inte har pengar för mat, kan du även kontakta diakoniarbetaren i din församling.
Du hittar kontaktuppgifterna vid din församling.
linkkiKonkurrens- och konsumentverket:
Ekonomi- och skuldrådgivarefinska _ svenska _ engelska
linkkiGaranti-Stiftelsen:
Hjälp med ekonomiska problemfinska _ svenska _ engelska
linkkiKonkurrens- och konsumentverket:
Information om ekonominfinska _ svenska _ engelska
Spelberoende
Om dina ekonomiska problem beror på spelproblem är det bäst att söka hjälp.
Du får hjälp med spelproblem vid A-kliniker (A-klinikka), mentalvårdsbyråer (mielenterveystoimisto) och hälsovårdscentralen (terveyskeskus).
På vissa orter kan även socialbyrån (sosiaalitoimisto) eller församlingarna hjälpa.
Även de anhöriga till en spelberoende person kan få hjälp.
Du kan också söka hjälp för ditt spelproblem vid olika organisationer.
I webbtjänsten Droglänken (Päihdelinkki) finns mycket information om spelproblem på flera språk.
Peluuri är en hjälptelefon för personer med spelproblem, deras närstående och andra som möter spelproblem.
Hjälptelefonen nås på numret 0800 100 101.
Betjäning ges på finska och svenska samt i mån av möjlighet även på engelska.
Peluuri finns även på internet.
linkkiDroglänken:
Information om spelproblemfinska _ svenska _ engelska _ ryska
Hjälp och information till spelberoende och deras anhörigafinska _ svenska _ engelska
Om du behöver visum eller uppehållstillstånd för att vistas i Finland, men inte har det, vistas du illegalt i Finland.
Asylsökande har rätt att uppehålla dig i Finland även utan visum eller uppehållstillstånd under den tid som det tar att handlägga asylansökan.
Även om du har kommit lagligt till Finland kan din vistelse i landet bli illegal till exempel om du stannar kvar i landet fastän du inte beviljas ett uppehållstillstånd eller om ditt visum eller uppehållstillstånd har gått ut.
Information om hur du kan få ett uppehållstillstånd i Finland finns på InfoFinlands sida Flytta till Finland.
Hjälp och rådgivning
Mathjälp och inkvartering
Du har rätt till nödinkvartering och mathjälp om du inte har pengar till mat eller någonstans att övernatta.
Kommuner, församlingar och vissa organisationer ordnar nödinkvartering.
Juridisk rådgivning
Flyktingrådgivningen r.f. ger kostnadsfri juridisk rådgivning för papperslösa invandrare.
Rådgivningen betjänar telefonledes på numret 045-237 7104 (måndagar kl. 14–16).
Rådgivningen ges av en jurist.
Fler kontaktuppgifter hittar du på Flyktingrådgivningens webbplats.
Sjukvård
Om du blir sjuk eller skadas, har du rätt till brådskande vård inom den offentliga hälso- och sjukvården, till exempel på en hälsostation eller ett sjukhus.
Du måste i regel själv betala kostnaderna för vården.
I Helsingfors, Åbo, Tammerfors och Esbo får barn och gravida kvinnor samma hälso- och sjukvårdstjänster som övriga invånare.
De måste betala samma avgifter för vården som övriga invånare.
Global Clinic är en klinik där du kan få hjälp eller råd av en läkare eller sjukskötare om du vistas i Finland utan uppehållstillstånd.
Du kan besöka Global Clinic även om du inte behöver brådskande sjukvård.
Global Clinic bedriver verksamhet i följande städer:
Åbo
Tammerfors
Uleåborg
Joensuu
Du kan ringa eller skicka e-post.
En sjukskötare eller läkare besvarar ditt samtal.
Du hittar kontaktinformation på Global Clinic:s hemsidor.
Global Clinic:s tjänster är avgiftsfria för kunderna.
Global Clinic anmäler inte sina kunder till polisen eller andra myndigheter.
Klinikens adress eller öppettider meddelas inte offentligt.
linkkiFlyktingrådgivningen rf:
Juridisk rådgivningfinska _ engelska _ franska _ arabiska
Kontaktuppgifterfinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Om du behöver visum eller uppehållstillstånd för att vistas i Finland, men inte har det, vistas du illegalt i Finland.
Asylsökande har rätt att uppehålla dig i Finland även utan visum eller uppehållstillstånd under den tid som det tar att handlägga asylansökan.
Även om du har kommit lagligt till Finland kan din vistelse i landet bli illegal till exempel om du stannar kvar i landet fastän du inte beviljas ett uppehållstillstånd eller om ditt visum eller uppehållstillstånd har gått ut.
Information om hur du kan få ett uppehållstillstånd i Finland finns på InfoFinlands sida Flytta till Finland.
Hjälp och rådgivning
Mathjälp och inkvartering
Du har rätt till nödinkvartering och mathjälp om du inte har pengar till mat eller någonstans att övernatta.
Kommuner, församlingar och vissa organisationer ordnar nödinkvartering.
Juridisk rådgivning
Flyktingrådgivningen r.f. ger kostnadsfri juridisk rådgivning för papperslösa invandrare.
Rådgivningen betjänar telefonledes på numret 045-237 7104 (måndagar kl. 14–16).
Rådgivningen ges av en jurist.
Fler kontaktuppgifter hittar du på Flyktingrådgivningens webbplats.
Sjukvård
Om du blir sjuk eller skadas, har du rätt till brådskande vård inom den offentliga hälso- och sjukvården, till exempel på en hälsostation eller ett sjukhus.
Du måste i regel själv betala kostnaderna för vården.
I Helsingfors, Åbo, Tammerfors och Esbo får barn och gravida kvinnor samma hälso- och sjukvårdstjänster som övriga invånare.
De måste betala samma avgifter för vården som övriga invånare.
Global Clinic är en klinik där du kan få hjälp eller råd av en läkare eller sjukskötare om du vistas i Finland utan uppehållstillstånd.
Du kan besöka Global Clinic även om du inte behöver brådskande sjukvård.
Global Clinic bedriver verksamhet i följande städer:
Åbo
Tammerfors
Uleåborg
Joensuu
Du kan ringa eller skicka e-post.
En sjukskötare eller läkare besvarar ditt samtal.
Du hittar kontaktinformation på Global Clinic:s hemsidor.
Global Clinic:s tjänster är avgiftsfria för kunderna.
Global Clinic anmäler inte sina kunder till polisen eller andra myndigheter.
Klinikens adress eller öppettider meddelas inte offentligt.
linkkiFlyktingrådgivningen rf:
Juridisk rådgivningfinska _ engelska _ franska _ arabiska
Kontaktuppgifterfinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Om du behöver visum eller uppehållstillstånd för att vistas i Finland, men inte har det, vistas du illegalt i Finland.
Asylsökande har rätt att uppehålla dig i Finland även utan visum eller uppehållstillstånd under den tid som det tar att handlägga asylansökan.
Även om du har kommit lagligt till Finland kan din vistelse i landet bli illegal till exempel om du stannar kvar i landet fastän du inte beviljas ett uppehållstillstånd eller om ditt visum eller uppehållstillstånd har gått ut.
Information om hur du kan få ett uppehållstillstånd i Finland finns på InfoFinlands sida Flytta till Finland.
Hjälp och rådgivning
Mathjälp och inkvartering
Du har rätt till nödinkvartering och mathjälp om du inte har pengar till mat eller någonstans att övernatta.
Kommuner, församlingar och vissa organisationer ordnar nödinkvartering.
Juridisk rådgivning
Flyktingrådgivningen r.f. ger kostnadsfri juridisk rådgivning för papperslösa invandrare.
Rådgivningen betjänar telefonledes på numret 045-237 7104 (måndagar kl. 14–16).
Rådgivningen ges av en jurist.
Fler kontaktuppgifter hittar du på Flyktingrådgivningens webbplats.
Sjukvård
Om du blir sjuk eller skadas, har du rätt till brådskande vård inom den offentliga hälso- och sjukvården, till exempel på en hälsostation eller ett sjukhus.
Du måste i regel själv betala kostnaderna för vården.
I Helsingfors, Åbo, Tammerfors och Esbo får barn och gravida kvinnor samma hälso- och sjukvårdstjänster som övriga invånare.
De måste betala samma avgifter för vården som övriga invånare.
Global Clinic är en klinik där du kan få hjälp eller råd av en läkare eller sjukskötare om du vistas i Finland utan uppehållstillstånd.
Du kan besöka Global Clinic även om du inte behöver brådskande sjukvård.
Global Clinic bedriver verksamhet i följande städer:
Åbo
Tammerfors
Uleåborg
Joensuu
Du kan ringa eller skicka e-post.
En sjukskötare eller läkare besvarar ditt samtal.
Du hittar kontaktinformation på Global Clinic:s hemsidor.
Global Clinic:s tjänster är avgiftsfria för kunderna.
Global Clinic anmäler inte sina kunder till polisen eller andra myndigheter.
Klinikens adress eller öppettider meddelas inte offentligt.
linkkiFlyktingrådgivningen rf:
Juridisk rådgivningfinska _ engelska _ franska _ arabiska
Kontaktuppgifterfinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Återkallande av uppehållstillstånd
Om du flyttar utomlands
Om ditt äktenskap eller registrerade parförhållande upphör
Om du förlorar ditt jobb
Återkallande av uppehållstillstånd
Ditt permanenta eller tidsbegränsade uppehållstillstånd återkallas om
du flyttar permanent från Finland
du har vistats två år utomlands utan avbrott.
Ditt permanenta eller tidsbegränsade uppehållstillstånd kan också återkallas om
du har uppgett felaktiga uppgifter i din ansökan om tillstånd
du har hemlighållit information som hade kunnat förhindra att tillståndet beviljas
ett annat Schengen-land begär att Finland återkallar ditt uppehållstillstånd.
Ett tidsbegränsat uppehållstillstånd kan också återkallas om de grunder på vilka tillståndet beviljades inte längre gäller.
Beslut om återkallelse av uppehållstillstånd fattas av Migrationsverket.
Om du flyttar utomlands
Om du ämnar flytta utomlands från Finland för två år, till exempel på grund av arbete eller studier, kan du ansöka hos Migrationsverket om att ditt uppehållstillstånd inte återkallas.
Ansökan är fritt formulerad men datum, underskrift och dina personuppgifter ska finnas med.
Ur ansökan bör även framgå hur länge och varför du studerar utomlands.
I din ansökning ska du motivera varför ditt uppehållstillstånd inte bör återkallas.
Ansökan ska göras innan du har vistats utomlands två år.
Om din finländska arbetsgivare har sänt dig utomlands för att arbeta förlorar du inte ditt uppehållstillstånd i Finland även om du vistas utomlands på grund av arbetet i över två år.
Om ditt äktenskap eller registrerade parförhållande upphör
Om du har ett tidsbestämt uppehållstillstånd med familjeband som grund kan det faktum att äktenskapet eller det registrerade parförhållandet upphör påverka uppehållstillståndet.
Om familjebandet inte längre existerar kan det hända att uppehållstillståndet inte förlängs.
Det är även möjligt att ett existerande tillstånd upphävs.
Uppehållstillståndet kan dock förlängas om du fortsättningsvis har starka band till Finland.
Exempel på sådana är:
barn eller andra familjemedlemmar i Finland
arbetsplats eller eget företag i Finland
studieplats i Finland
Om du skiljer dig på grund av att din make/maka varit våldsam mot dig kan ditt uppehållstillstånd förlängas trots skilsmässan.
Du ska lämna in en redovisning, exempelvis läkarintyg eller utlåtande från familjerådgivning.
Bifoga även till ansökan om uppehållstillstånd din egen redovisning av situationen.
Mer information om skilsmässa och upplösande av ett registrerat parförhållande hittar du på InfoFinlands sidor Skilsmässa.
Om du förlorar ditt jobb
Om du har ett uppehållstillstånd för arbetstagare som endast gäller arbete för en viss arbetsgivare och du förlorar din arbetsplats, ska du ansöka om ett nytt uppehållstillstånd för arbetstagare eller ett uppehållstillstånd på andra grunder.
Om Migrationsverket har beviljat dig ett uppehållstillstånd för arbetstagare och din anställning upphör tidigare än uppehållstillståndet, måste du eller din arbetsgivare skriftligt meddela Migrationsverket att din anställning upphör.
Om ditt uppehållstillstånd för arbetstagare inte har begränsats att gälla arbete för en viss arbetsgivare, utan för en viss bransch och tillståndet är fortfarande giltigt, kan du byta jobb inom samma bransch.
Mer information om arbete och företagande i Finland hittar du på InfoFinlands sida Arbete och entreprenörskap.
Mer information om uppehållstillstånd för arbetstagare och företagare hittar du på sidan Arbeta i Finland och Till Finland som företagare.
Om du redan har haft ett uppehållstillstånd i Finland, men tillståndet inte förlängs, fattar Migrationsverket beslut om utvisning.
Om du begår brott i Finland, kan du även utvisas på grund av brotten.
Om du blir utvisad, förfaller ditt eventuella giltiga uppehållstillstånd och du måste lämna landet.
Vanligtvis får du en tidsfrist inom vilken du måste lämna Finland.
Om du inte lämnar Finland inom tidsfristen avlägsnar polisen eller gränsbevakningsväsendet dig ur landet.
Enligt lag kan du inte utvisas om du hotas av dödsstraff, tortyr, förföljelse eller någon annan behandling som är omänsklig eller kränker människovärdet i ditt hemland.
Återkallelse av uppehållstillståndfinska _ svenska _ engelska
Avvisning och utvisningfinska _ svenska _ engelska
Återkallande av uppehållstillstånd
Om du flyttar utomlands
Om ditt äktenskap eller registrerade parförhållande upphör
Om du förlorar ditt jobb
Återkallande av uppehållstillstånd
Ditt permanenta eller tidsbegränsade uppehållstillstånd återkallas om
du flyttar permanent från Finland
du har vistats två år utomlands utan avbrott.
Ditt permanenta eller tidsbegränsade uppehållstillstånd kan också återkallas om
du har uppgett felaktiga uppgifter i din ansökan om tillstånd
du har hemlighållit information som hade kunnat förhindra att tillståndet beviljas
ett annat Schengen-land begär att Finland återkallar ditt uppehållstillstånd.
Ett tidsbegränsat uppehållstillstånd kan också återkallas om de grunder på vilka tillståndet beviljades inte längre gäller.
Beslut om återkallelse av uppehållstillstånd fattas av Migrationsverket.
Om du flyttar utomlands
Om du ämnar flytta utomlands från Finland för två år, till exempel på grund av arbete eller studier, kan du ansöka hos Migrationsverket om att ditt uppehållstillstånd inte återkallas.
Ansökan är fritt formulerad men datum, underskrift och dina personuppgifter ska finnas med.
Ur ansökan bör även framgå hur länge och varför du studerar utomlands.
I din ansökning ska du motivera varför ditt uppehållstillstånd inte bör återkallas.
Ansökan ska göras innan du har vistats utomlands två år.
Om din finländska arbetsgivare har sänt dig utomlands för att arbeta förlorar du inte ditt uppehållstillstånd i Finland även om du vistas utomlands på grund av arbetet i över två år.
Om ditt äktenskap eller registrerade parförhållande upphör
Om du har ett tidsbestämt uppehållstillstånd med familjeband som grund kan det faktum att äktenskapet eller det registrerade parförhållandet upphör påverka uppehållstillståndet.
Om familjebandet inte längre existerar kan det hända att uppehållstillståndet inte förlängs.
Det är även möjligt att ett existerande tillstånd upphävs.
Uppehållstillståndet kan dock förlängas om du fortsättningsvis har starka band till Finland.
Exempel på sådana är:
barn eller andra familjemedlemmar i Finland
arbetsplats eller eget företag i Finland
studieplats i Finland
Om du skiljer dig på grund av att din make/maka varit våldsam mot dig kan ditt uppehållstillstånd förlängas trots skilsmässan.
Du ska lämna in en redovisning, exempelvis läkarintyg eller utlåtande från familjerådgivning.
Bifoga även till ansökan om uppehållstillstånd din egen redovisning av situationen.
Mer information om skilsmässa och upplösande av ett registrerat parförhållande hittar du på InfoFinlands sidor Skilsmässa.
Om du förlorar ditt jobb
Om du har ett uppehållstillstånd för arbetstagare som endast gäller arbete för en viss arbetsgivare och du förlorar din arbetsplats, ska du ansöka om ett nytt uppehållstillstånd för arbetstagare eller ett uppehållstillstånd på andra grunder.
Om Migrationsverket har beviljat dig ett uppehållstillstånd för arbetstagare och din anställning upphör tidigare än uppehållstillståndet, måste du eller din arbetsgivare skriftligt meddela Migrationsverket att din anställning upphör.
Om ditt uppehållstillstånd för arbetstagare inte har begränsats att gälla arbete för en viss arbetsgivare, utan för en viss bransch och tillståndet är fortfarande giltigt, kan du byta jobb inom samma bransch.
Mer information om arbete och företagande i Finland hittar du på InfoFinlands sida Arbete och entreprenörskap.
Mer information om uppehållstillstånd för arbetstagare och företagare hittar du på sidan Arbeta i Finland och Till Finland som företagare.
Om du redan har haft ett uppehållstillstånd i Finland, men tillståndet inte förlängs, fattar Migrationsverket beslut om utvisning.
Om du begår brott i Finland, kan du även utvisas på grund av brotten.
Om du blir utvisad, förfaller ditt eventuella giltiga uppehållstillstånd och du måste lämna landet.
Vanligtvis får du en tidsfrist inom vilken du måste lämna Finland.
Om du inte lämnar Finland inom tidsfristen avlägsnar polisen eller gränsbevakningsväsendet dig ur landet.
Enligt lag kan du inte utvisas om du hotas av dödsstraff, tortyr, förföljelse eller någon annan behandling som är omänsklig eller kränker människovärdet i ditt hemland.
Återkallelse av uppehållstillståndfinska _ svenska _ engelska
Avvisning och utvisningfinska _ svenska _ engelska
Återkallande av uppehållstillstånd
Om du flyttar utomlands
Om ditt äktenskap eller registrerade parförhållande upphör
Om du förlorar ditt jobb
Återkallande av uppehållstillstånd
Ditt permanenta eller tidsbegränsade uppehållstillstånd återkallas om
du flyttar permanent från Finland
du har vistats två år utomlands utan avbrott.
Ditt permanenta eller tidsbegränsade uppehållstillstånd kan också återkallas om
du har uppgett felaktiga uppgifter i din ansökan om tillstånd
du har hemlighållit information som hade kunnat förhindra att tillståndet beviljas
ett annat Schengen-land begär att Finland återkallar ditt uppehållstillstånd.
Ett tidsbegränsat uppehållstillstånd kan också återkallas om de grunder på vilka tillståndet beviljades inte längre gäller.
Beslut om återkallelse av uppehållstillstånd fattas av Migrationsverket.
Om du flyttar utomlands
Om du ämnar flytta utomlands från Finland för två år, till exempel på grund av arbete eller studier, kan du ansöka hos Migrationsverket om att ditt uppehållstillstånd inte återkallas.
Ansökan är fritt formulerad men datum, underskrift och dina personuppgifter ska finnas med.
Ur ansökan bör även framgå hur länge och varför du studerar utomlands.
I din ansökning ska du motivera varför ditt uppehållstillstånd inte bör återkallas.
Ansökan ska göras innan du har vistats utomlands två år.
Om din finländska arbetsgivare har sänt dig utomlands för att arbeta förlorar du inte ditt uppehållstillstånd i Finland även om du vistas utomlands på grund av arbetet i över två år.
Om ditt äktenskap eller registrerade parförhållande upphör
Om du har ett tidsbestämt uppehållstillstånd med familjeband som grund kan det faktum att äktenskapet eller det registrerade parförhållandet upphör påverka uppehållstillståndet.
Om familjebandet inte längre existerar kan det hända att uppehållstillståndet inte förlängs.
Det är även möjligt att ett existerande tillstånd upphävs.
Uppehållstillståndet kan dock förlängas om du fortsättningsvis har starka band till Finland.
Exempel på sådana är:
barn eller andra familjemedlemmar i Finland
arbetsplats eller eget företag i Finland
studieplats i Finland
Om du skiljer dig på grund av att din make/maka varit våldsam mot dig kan ditt uppehållstillstånd förlängas trots skilsmässan.
Du ska lämna in en redovisning, exempelvis läkarintyg eller utlåtande från familjerådgivning.
Bifoga även till ansökan om uppehållstillstånd din egen redovisning av situationen.
Mer information om skilsmässa och upplösande av ett registrerat parförhållande hittar du på InfoFinlands sidor Skilsmässa.
Om du förlorar ditt jobb
Om du har ett uppehållstillstånd för arbetstagare som endast gäller arbete för en viss arbetsgivare och du förlorar din arbetsplats, ska du ansöka om ett nytt uppehållstillstånd för arbetstagare eller ett uppehållstillstånd på andra grunder.
Om Migrationsverket har beviljat dig ett uppehållstillstånd för arbetstagare och din anställning upphör tidigare än uppehållstillståndet, måste du eller din arbetsgivare skriftligt meddela Migrationsverket att din anställning upphör.
Om ditt uppehållstillstånd för arbetstagare inte har begränsats att gälla arbete för en viss arbetsgivare, utan för en viss bransch och tillståndet är fortfarande giltigt, kan du byta jobb inom samma bransch.
Mer information om arbete och företagande i Finland hittar du på InfoFinlands sida Arbete och entreprenörskap.
Mer information om uppehållstillstånd för arbetstagare och företagare hittar du på sidan Arbeta i Finland och Till Finland som företagare.
Om du redan har haft ett uppehållstillstånd i Finland, men tillståndet inte förlängs, fattar Migrationsverket beslut om utvisning.
Om du begår brott i Finland, kan du även utvisas på grund av brotten.
Om du blir utvisad, förfaller ditt eventuella giltiga uppehållstillstånd och du måste lämna landet.
Vanligtvis får du en tidsfrist inom vilken du måste lämna Finland.
Om du inte lämnar Finland inom tidsfristen avlägsnar polisen eller gränsbevakningsväsendet dig ur landet.
Enligt lag kan du inte utvisas om du hotas av dödsstraff, tortyr, förföljelse eller någon annan behandling som är omänsklig eller kränker människovärdet i ditt hemland.
Återkallelse av uppehållstillståndfinska _ svenska _ engelska
Avvisning och utvisningfinska _ svenska _ engelska
Om du redan är i Finland och får ett negativt beslut om uppehållstillstånd från Migrationsverket (Maahanmuuttovirasto), måste du antingen lämna Finland eller överklaga beslutet.
Du får vistas i Finland så länge som behandlingen av besvären pågår.
Du kan överklaga också om du har ansökt om uppehållstillstånd utomlands.
Då måste du vänta på behandlingen av besvären utomlands.
Om du är asylsökande i Finland eller offer för människohandel, har du rätt att få stöd för frivillig återresa (vapaaehtoisen paluun tuki), om du beslutar att återvända till ditt hemland.
Läs mer under rubriken Stöd för frivillig återresa.
Att överklaga ett beslut om uppehållstillstånd
En besvärsanvisning om hur beslutet får överklagas bifogas alltid beslutet.
Besvären behandlas av förvaltningsdomstolen (hallinto-oikeus).
Förvaltningsdomstolen kan antingen avslå besvären eller sända ärendet till Migrationsverket för ny behandling.
Avslag innebär att Migrationsverkets beslut förblir gällande.
Om förvaltningsdomstolen avslår besvären kan du i vissa fall ansöka om besvärstillstånd hos högsta förvaltningsdomstolen (korkein hallinto-oikeus).
Om högsta förvaltningsdomstolen beviljar besvärstillstånd, behandlar den besvären.
Du kan få hjälp med att överklaga av antingen en privat jurist, en statlig rättshjälpsbyrå (valtion oikeusaputoimisto) eller Flyktingrådgivningen rf (Pakolaisneuvonta) (endast asylsökande).
På InfoFinlands sida Behöver du en jurist? finns mer information om hur du kan få hjälp i juridiska ärenden.
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Att lämna Finland
Om du får avslag på din ansökan om uppehållstillstånd eller om förvaltningsrätten avslår ditt överklagande, måste du lämna Finland.
Du ges möjlighet att lämna landet frivilligt.
Tidsfristen är vanligtvis 30 dagar.
Om du inte lämnar landet inom tidsfristen, avlägsnar polisen eller gränsbevakningsväsendet dig ur landet.
Du får inreseförbud till Schengenområdet om:
Du har brutit mot inresereglerna och din ansökan har avslagits, till exempel på grund av skenäktenskap.
Du har begått brott och du anses utgöra ett hot mot den allmänna ordningen och säkerheten.
Din asylansökan avslås i ett påskyndat förfarande.
Du inte lämnar landet frivilligt inom den tidsfrist som meddelats för dig.
När du har inreseförbud kan du inte besöka Finland eller något annat Schengenland.
Avvisning och utvisningfinska _ svenska _ engelska
Stöd för frivillig återresa
Om du vill återvända till ditt hemland kan du i vissa fall få stöd för frivilligt återvändande.
Stödet består antingen av pengar eller tjänster.
Penningsummans storlek beror på vilket land du återvänder till.
Tjänsten kan till exempel vara att du får hjälp med att leta efter en bostad eller arbetsplats i det land dit du återvänder.
Du kan få stöd om:
du har fått ett negativt beslut på din asylansökan
du återkallar din asylansökan
du är ett offer för människohandel och du inte har en hemkommun i Finland
du har ett tillfälligt uppehållstillstånd på grund av hinder för avlägsnande ur landet
du har fått tillfälligt skydd
din flyktingstatus i Finland har upphört eller återkallats eller det har fattats beslut om att avvisa dig
du har fått humanitärt skydd, men ditt uppehållstillstånd löper ut eller har redan löpt ut.
Om du är kund hos en mottagningscentral kan du ansöka om stöd för frivilligt återvändande vid din egen mottagningscentral.
Om du inte är kund hos en mottagningscentral kan du ansöka om stöd hos Migrationsverket.
Frivillig återflyttningfinska _ svenska _ engelska
Om du redan är i Finland och får ett negativt beslut om uppehållstillstånd från Migrationsverket (Maahanmuuttovirasto), måste du antingen lämna Finland eller överklaga beslutet.
Du får vistas i Finland så länge som behandlingen av besvären pågår.
Du kan överklaga också om du har ansökt om uppehållstillstånd utomlands.
Då måste du vänta på behandlingen av besvären utomlands.
Om du är asylsökande i Finland eller offer för människohandel, har du rätt att få stöd för frivillig återresa (vapaaehtoisen paluun tuki), om du beslutar att återvända till ditt hemland.
Läs mer under rubriken Stöd för frivillig återresa.
Att överklaga ett beslut om uppehållstillstånd
En besvärsanvisning om hur beslutet får överklagas bifogas alltid beslutet.
Besvären behandlas av förvaltningsdomstolen (hallinto-oikeus).
Förvaltningsdomstolen kan antingen avslå besvären eller sända ärendet till Migrationsverket för ny behandling.
Avslag innebär att Migrationsverkets beslut förblir gällande.
Om förvaltningsdomstolen avslår besvären kan du i vissa fall ansöka om besvärstillstånd hos högsta förvaltningsdomstolen (korkein hallinto-oikeus).
Om högsta förvaltningsdomstolen beviljar besvärstillstånd, behandlar den besvären.
Du kan få hjälp med att överklaga av antingen en privat jurist, en statlig rättshjälpsbyrå (valtion oikeusaputoimisto) eller Flyktingrådgivningen rf (Pakolaisneuvonta) (endast asylsökande).
På InfoFinlands sida Behöver du en jurist? finns mer information om hur du kan få hjälp i juridiska ärenden.
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Att lämna Finland
Om du får avslag på din ansökan om uppehållstillstånd eller om förvaltningsrätten avslår ditt överklagande, måste du lämna Finland.
Du ges möjlighet att lämna landet frivilligt.
Tidsfristen är vanligtvis 30 dagar.
Om du inte lämnar landet inom tidsfristen, avlägsnar polisen eller gränsbevakningsväsendet dig ur landet.
Du får inreseförbud till Schengenområdet om:
Du har brutit mot inresereglerna och din ansökan har avslagits, till exempel på grund av skenäktenskap.
Du har begått brott och du anses utgöra ett hot mot den allmänna ordningen och säkerheten.
Din asylansökan avslås i ett påskyndat förfarande.
Du inte lämnar landet frivilligt inom den tidsfrist som meddelats för dig.
När du har inreseförbud kan du inte besöka Finland eller något annat Schengenland.
Avvisning och utvisningfinska _ svenska _ engelska
Stöd för frivillig återresa
Om du vill återvända till ditt hemland kan du i vissa fall få stöd för frivilligt återvändande.
Stödet består antingen av pengar eller tjänster.
Penningsummans storlek beror på vilket land du återvänder till.
Tjänsten kan till exempel vara att du får hjälp med att leta efter en bostad eller arbetsplats i det land dit du återvänder.
Du kan få stöd om:
du har fått ett negativt beslut på din asylansökan
du återkallar din asylansökan
du är ett offer för människohandel och du inte har en hemkommun i Finland
du har ett tillfälligt uppehållstillstånd på grund av hinder för avlägsnande ur landet
du har fått tillfälligt skydd
din flyktingstatus i Finland har upphört eller återkallats eller det har fattats beslut om att avvisa dig
du har fått humanitärt skydd, men ditt uppehållstillstånd löper ut eller har redan löpt ut.
Om du är kund hos en mottagningscentral kan du ansöka om stöd för frivilligt återvändande vid din egen mottagningscentral.
Om du inte är kund hos en mottagningscentral kan du ansöka om stöd hos Migrationsverket.
Frivillig återflyttningfinska _ svenska _ engelska
Stöd för frivilligt återvändandefinska _ svenska _ engelska _ persiska _ arabiska
Om du redan är i Finland och får ett negativt beslut om uppehållstillstånd från Migrationsverket (Maahanmuuttovirasto), måste du antingen lämna Finland eller överklaga beslutet.
Du får vistas i Finland så länge som behandlingen av besvären pågår.
Du kan överklaga också om du har ansökt om uppehållstillstånd utomlands.
Då måste du vänta på behandlingen av besvären utomlands.
Om du är asylsökande i Finland eller offer för människohandel, har du rätt att få stöd för frivillig återresa (vapaaehtoisen paluun tuki), om du beslutar att återvända till ditt hemland.
Läs mer under rubriken Stöd för frivillig återresa.
Att överklaga ett beslut om uppehållstillstånd
En besvärsanvisning om hur beslutet får överklagas bifogas alltid beslutet.
Besvären behandlas av förvaltningsdomstolen (hallinto-oikeus).
Förvaltningsdomstolen kan antingen avslå besvären eller sända ärendet till Migrationsverket för ny behandling.
Avslag innebär att Migrationsverkets beslut förblir gällande.
Om förvaltningsdomstolen avslår besvären kan du i vissa fall ansöka om besvärstillstånd hos högsta förvaltningsdomstolen (korkein hallinto-oikeus).
Om högsta förvaltningsdomstolen beviljar besvärstillstånd, behandlar den besvären.
Du kan få hjälp med att överklaga av antingen en privat jurist, en statlig rättshjälpsbyrå (valtion oikeusaputoimisto) eller Flyktingrådgivningen rf (Pakolaisneuvonta) (endast asylsökande).
På InfoFinlands sida Behöver du en jurist? finns mer information om hur du kan få hjälp i juridiska ärenden.
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Att lämna Finland
Om du får avslag på din ansökan om uppehållstillstånd eller om förvaltningsrätten avslår ditt överklagande, måste du lämna Finland.
Du ges möjlighet att lämna landet frivilligt.
Tidsfristen är vanligtvis 30 dagar.
Om du inte lämnar landet inom tidsfristen, avlägsnar polisen eller gränsbevakningsväsendet dig ur landet.
Du får inreseförbud till Schengenområdet om:
Du har brutit mot inresereglerna och din ansökan har avslagits, till exempel på grund av skenäktenskap.
Du har begått brott och du anses utgöra ett hot mot den allmänna ordningen och säkerheten.
Din asylansökan avslås i ett påskyndat förfarande.
Du inte lämnar landet frivilligt inom den tidsfrist som meddelats för dig.
När du har inreseförbud kan du inte besöka Finland eller något annat Schengenland.
Avvisning och utvisningfinska _ svenska _ engelska
Stöd för frivillig återresa
Om du vill återvända till ditt hemland kan du i vissa fall få stöd för frivilligt återvändande.
Stödet består antingen av pengar eller tjänster.
Penningsummans storlek beror på vilket land du återvänder till.
Tjänsten kan till exempel vara att du får hjälp med att leta efter en bostad eller arbetsplats i det land dit du återvänder.
Du kan få stöd om:
du har fått ett negativt beslut på din asylansökan
du återkallar din asylansökan
du är ett offer för människohandel och du inte har en hemkommun i Finland
du har ett tillfälligt uppehållstillstånd på grund av hinder för avlägsnande ur landet
du har fått tillfälligt skydd
din flyktingstatus i Finland har upphört eller återkallats eller det har fattats beslut om att avvisa dig
du har fått humanitärt skydd, men ditt uppehållstillstånd löper ut eller har redan löpt ut.
Om du är kund hos en mottagningscentral kan du ansöka om stöd för frivilligt återvändande vid din egen mottagningscentral.
Om du inte är kund hos en mottagningscentral kan du ansöka om stöd hos Migrationsverket.
Frivillig återflyttningfinska _ svenska _ engelska
Stöd för frivilligt återvändandefinska _ svenska _ engelska _ persiska _ arabiska
Rådgivning i uppehållstillståndsärenden
Om du har problem eller oklarheter med uppehållstillståndet, kan du ta kontakt med följande instanser för att be om råd:
Finlands beskickningar utomlands
Invandrarrådgivarna i din kommun i Finland
På Migrationsverkets webbplats finns mycket information om uppehållstillstånd.
Migrationsverket ger rådgivning angående tillstånd också per telefon.
Finlands beskickningar utomlands betjänar personer som ansöker om uppehållstillstånd i utlandet.
Många städer har rådgivningstjänster för invandrare med rådgivare som specialiserat sig på invandringsfrågor.
Flyktingsrådgivningen bistår asylsökande juridiskt i asylprocessen.
Dessutom tillhandahåller Flyktingrådgivningen allmän juridisk rådgivning för andra utlänningar.
Vänligen observera att endast Migrationsverket kan fatta beslut om uppehållstillstånd.
Information om uppehållstillståndfinska _ svenska _ engelska
linkkiFlyktingrådgivningen rf:
Juridisk rådgivningfinska _ engelska _ franska _ arabiska
Rådgivning i uppehållstillståndsärenden
Om du har problem eller oklarheter med uppehållstillståndet, kan du ta kontakt med följande instanser för att be om råd:
Finlands beskickningar utomlands
Invandrarrådgivarna i din kommun i Finland
På Migrationsverkets webbplats finns mycket information om uppehållstillstånd.
Migrationsverket ger rådgivning angående tillstånd också per telefon.
Finlands beskickningar utomlands betjänar personer som ansöker om uppehållstillstånd i utlandet.
Många städer har rådgivningstjänster för invandrare med rådgivare som specialiserat sig på invandringsfrågor.
Flyktingsrådgivningen bistår asylsökande juridiskt i asylprocessen.
Dessutom tillhandahåller Flyktingrådgivningen allmän juridisk rådgivning för andra utlänningar.
Vänligen observera att endast Migrationsverket kan fatta beslut om uppehållstillstånd.
Information om uppehållstillståndfinska _ svenska _ engelska
linkkiFlyktingrådgivningen rf:
Juridisk rådgivningfinska _ engelska _ franska _ arabiska
Rådgivning i uppehållstillståndsärenden
Om du har problem eller oklarheter med uppehållstillståndet, kan du ta kontakt med följande instanser för att be om råd:
Finlands beskickningar utomlands
Invandrarrådgivarna i din kommun i Finland
På Migrationsverkets webbplats finns mycket information om uppehållstillstånd.
Migrationsverket ger rådgivning angående tillstånd också per telefon.
Finlands beskickningar utomlands betjänar personer som ansöker om uppehållstillstånd i utlandet.
Många städer har rådgivningstjänster för invandrare med rådgivare som specialiserat sig på invandringsfrågor.
Flyktingsrådgivningen bistår asylsökande juridiskt i asylprocessen.
Dessutom tillhandahåller Flyktingrådgivningen allmän juridisk rådgivning för andra utlänningar.
Vänligen observera att endast Migrationsverket kan fatta beslut om uppehållstillstånd.
Information om uppehållstillståndfinska _ svenska _ engelska
linkkiFlyktingrådgivningen rf:
Juridisk rådgivningfinska _ engelska _ franska _ arabiska
Nödnumret (hätänumero) i Finland är 112.
Du får ringa nödnumret endast i brådskande nödfall där liv, hälsa, egendom eller miljö är i fara.
I nödsituationer får du vård även om du inte har en hemkommun i Finland.
Vårdavgifter kan komma att debiteras av dig i efterhand.
Ring 112 till exempel i följande situationer:
du har råkat ut för en bilolycka (auto-onnettomuus) eller är vittne till en olycka
någon är i livsfara (hengenvaara)
du upptäcker en brand (tulipalo)
du upptäcker ett inbrott (murto)
Ring inte nödnumret om ärendet inte är brådskande.
Du ska inte ringa nödnumret vid vanliga sjukdomsfall.
Du ska inte heller ringa nödnumret om du vill fråga polisen (poliisi) till exempel om ett tillståndsärende.
Onödiga samtal kan orsaka att hjälpen kommer för sent i verkliga nödsituationer.
Du kan straffas för att ha missbrukat nödnumret.
Samtalet besvaras av en utbildad nödcentraloperatör.
Han eller hon ställer dig frågor och bedömer hjälpbehovet.
Därefter larmar han eller hon hjälp.
Operatören berättar också vad du ska göra.
Operatören kopplar inte samtalet vidare, så besvara frågorna noga.
Du kan tala finska eller svenska när du ringer nödnumret.
Du kan också fråga om nödcentraloperatören förstår engelska, med det är inte säkert.
Vid behov bistås nödcentralen av en tolktjänst.
Du kan ringa nödnumret gratis från alla telefoner.
Du behöver inget riktnummer.
Du kan ringa nödnumret utan riktnummer även om du har ett utländskt mobilabonnemang.
Nödnumret 112 fungerar i alla EU-länder.
Om du har installerat den kostnadsfria mobilappen 112 Suomi i din telefon, behöver du inte nödvändigtvis kunna berätta var du befinner dig.
Nödcentraloperatören ser var du är, när du ringer ett nödsamtal via appen.
Du kan ladda ned appen i applikationsbutiken.
När du ringer nödnumret 112:
uppge ditt namn
berätta vad som har hänt
ange exakt adress och kommun
svara på nödcentraloperatörens frågor
följ instruktionerna
avsluta inte samtalet förrän du får lov.
Mer information om nödnumret får du på Nödcentralsverkets (Hätäkeskuslaitos) webbplats.
Om du behöver information om tillståndsärenden som sköts av polisen, fordonsföreskrifter eller hur undersökningen i ett brott som skett tidigare framskrider ska du ringa polisens egna nummer under tjänstetid.
Om du misstänker att någon har förgiftats kan du fråga råd vid Giftinformationscentralen (Myrkytystietokeskus).
Giftinformationscentralens telefontjänst är öppen 24 timmar om dygnet.
Telefonnumret är (09) 471 977.
linkkiNödcentralsverket:
Nödsituationfinska _ svenska _ engelska
linkkiNödcentralsverket:
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
linkkiRöda Kors:
Första hjälpen-anvisningar för olika situationerfinska _ svenska _ engelska
Första hjälpen-anvisningar vid förgiftningfinska _ svenska _ engelska
Nödnumret (hätänumero) i Finland är 112.
Du får ringa nödnumret endast i brådskande nödfall där liv, hälsa, egendom eller miljö är i fara.
I nödsituationer får du vård även om du inte har en hemkommun i Finland.
Vårdavgifter kan komma att debiteras av dig i efterhand.
Ring 112 till exempel i följande situationer:
du har råkat ut för en bilolycka (auto-onnettomuus) eller är vittne till en olycka
någon är i livsfara (hengenvaara)
du upptäcker en brand (tulipalo)
du upptäcker ett inbrott (murto)
Ring inte nödnumret om ärendet inte är brådskande.
Du ska inte ringa nödnumret vid vanliga sjukdomsfall.
Du ska inte heller ringa nödnumret om du vill fråga polisen (poliisi) till exempel om ett tillståndsärende.
Onödiga samtal kan orsaka att hjälpen kommer för sent i verkliga nödsituationer.
Du kan straffas för att ha missbrukat nödnumret.
Samtalet besvaras av en utbildad nödcentraloperatör.
Han eller hon ställer dig frågor och bedömer hjälpbehovet.
Därefter larmar han eller hon hjälp.
Operatören berättar också vad du ska göra.
Operatören kopplar inte samtalet vidare, så besvara frågorna noga.
Du kan tala finska eller svenska när du ringer nödnumret.
Du kan också fråga om nödcentraloperatören förstår engelska, med det är inte säkert.
Vid behov bistås nödcentralen av en tolktjänst.
Du kan ringa nödnumret gratis från alla telefoner.
Du behöver inget riktnummer.
Du kan ringa nödnumret utan riktnummer även om du har ett utländskt mobilabonnemang.
Nödnumret 112 fungerar i alla EU-länder.
Om du har installerat den kostnadsfria mobilappen 112 Suomi i din telefon, behöver du inte nödvändigtvis kunna berätta var du befinner dig.
Nödcentraloperatören ser var du är, när du ringer ett nödsamtal via appen.
Du kan ladda ned appen i applikationsbutiken.
När du ringer nödnumret 112:
uppge ditt namn
berätta vad som har hänt
ange exakt adress och kommun
svara på nödcentraloperatörens frågor
följ instruktionerna
avsluta inte samtalet förrän du får lov.
Mer information om nödnumret får du på Nödcentralsverkets (Hätäkeskuslaitos) webbplats.
Om du behöver information om tillståndsärenden som sköts av polisen, fordonsföreskrifter eller hur undersökningen i ett brott som skett tidigare framskrider ska du ringa polisens egna nummer under tjänstetid.
Om du misstänker att någon har förgiftats kan du fråga råd vid Giftinformationscentralen (Myrkytystietokeskus).
Giftinformationscentralens telefontjänst är öppen 24 timmar om dygnet.
Telefonnumret är (09) 471 977.
linkkiNödcentralsverket:
Nödsituationfinska _ svenska _ engelska
linkkiNödcentralsverket:
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
linkkiRöda Kors:
Första hjälpen-anvisningar för olika situationerfinska _ svenska _ engelska
Första hjälpen-anvisningar vid förgiftningfinska _ svenska _ engelska
Nödnumret (hätänumero) i Finland är 112.
Du får ringa nödnumret endast i brådskande nödfall där liv, hälsa, egendom eller miljö är i fara.
I nödsituationer får du vård även om du inte har en hemkommun i Finland.
Vårdavgifter kan komma att debiteras av dig i efterhand.
Ring 112 till exempel i följande situationer:
du har råkat ut för en bilolycka (auto-onnettomuus) eller är vittne till en olycka
någon är i livsfara (hengenvaara)
du upptäcker en brand (tulipalo)
du upptäcker ett inbrott (murto)
Ring inte nödnumret om ärendet inte är brådskande.
Du ska inte ringa nödnumret vid vanliga sjukdomsfall.
Du ska inte heller ringa nödnumret om du vill fråga polisen (poliisi) till exempel om ett tillståndsärende.
Onödiga samtal kan orsaka att hjälpen kommer för sent i verkliga nödsituationer.
Du kan straffas för att ha missbrukat nödnumret.
Samtalet besvaras av en utbildad nödcentraloperatör.
Han eller hon ställer dig frågor och bedömer hjälpbehovet.
Därefter larmar han eller hon hjälp.
Operatören berättar också vad du ska göra.
Operatören kopplar inte samtalet vidare, så besvara frågorna noga.
Du kan tala finska eller svenska när du ringer nödnumret.
Du kan också fråga om nödcentraloperatören förstår engelska, med det är inte säkert.
Vid behov bistås nödcentralen av en tolktjänst.
Du kan ringa nödnumret gratis från alla telefoner.
Du behöver inget riktnummer.
Du kan ringa nödnumret utan riktnummer även om du har ett utländskt mobilabonnemang.
Nödnumret 112 fungerar i alla EU-länder.
Om du har installerat den kostnadsfria mobilappen 112 Suomi i din telefon, behöver du inte nödvändigtvis kunna berätta var du befinner dig.
Nödcentraloperatören ser var du är, när du ringer ett nödsamtal via appen.
Du kan ladda ned appen i applikationsbutiken.
När du ringer nödnumret 112:
uppge ditt namn
berätta vad som har hänt
ange exakt adress och kommun
svara på nödcentraloperatörens frågor
följ instruktionerna
avsluta inte samtalet förrän du får lov.
Mer information om nödnumret får du på Nödcentralsverkets (Hätäkeskuslaitos) webbplats.
Om du behöver information om tillståndsärenden som sköts av polisen, fordonsföreskrifter eller hur undersökningen i ett brott som skett tidigare framskrider ska du ringa polisens egna nummer under tjänstetid.
Om du misstänker att någon har förgiftats kan du fråga råd vid Giftinformationscentralen (Myrkytystietokeskus).
Giftinformationscentralens telefontjänst är öppen 24 timmar om dygnet.
Telefonnumret är (09) 471 977.
linkkiNödcentralsverket:
Nödsituationfinska _ svenska _ engelska
linkkiNödcentralsverket:
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
linkkiRöda Kors:
Första hjälpen-anvisningar för olika situationerfinska _ svenska _ engelska
Första hjälpen-anvisningar vid förgiftningfinska _ svenska _ engelska
I Finland ordnar kommunerna tjänster för äldre för att underlätta deras vardag och för att de ska kunna bo hemma så länge som möjligt.
Om du har hemkommun i Finland har du rätt att använda de tjänster som kommunen tillhandahåller.
Boende
Om ditt hem är funktionellt kan du bo hemma även om du har lite svag hälsa.
Du kan låta utföra ändringsarbeten i ditt hem som underlättar boendet.
Det åligger kommunerna att ordna serviceboende och stödboende för personer som behöver det.
Läs mer på InfoFinlands sida Stöd- och serviceboende.
Invandrare som har bott tillräckligt länge i Finland får ålders- eller invalidpension på samma grunder som alla andra som är bosatta i Finland.
Pensionsbeloppet beror på hur länge personen har bott eller arbetat i Finland.
Efter tre års boende tryggar dock garantipensionen ett existensminimum.
Stöden för pensionärerfinska _ svenska _ engelska
Att röra sig
Du kan få låna olika hjälpmedel för att lättare kunna röra på dig, till exempel en käpp eller en rullator.
Om du behöver hjälpmedel ska du först kontakta din egen hälsostation.
Vid hälsostationen får du mer information om hjälpmedlen.
På vintern är det ofta halt ute.
Skomakare och en del stora varuhus säljer halkskydd (liukueste) som kan fästas under sulan på vanliga skor.
Du kan också köpa skor med dubbar (nastakengät) på en skoaffär. Med dem är det lättare att gå på hala gator.
Hemvård
För äldre personer ordnar kommunerna hemvård (kotihoito) som omfattar hjälp med vardagssysslor och sjukvård i hemmet.
Hemvården omfattar hemtjänster, hemsjukvård och stödtjänster.
Hemtjänsterna är hjälp med vardagssysslor, till exempel med att tvätta sig, klä på sig och måltider.
Hemsjukvård är sjukvård och rehabilitering som ges i hemmet.
Remiss för hemsjukvården skrivs av läkare.
Utöver dessa finns det stödtjänster, som är till exempel måltids-, städ-, inköps-, säkerhets- och transporthjälp.
Kontakta hemvårdsenheten i din hemkommun när du behöver hemvård.
Kommunens hemvård är avgiftsbelagd.
När hemvården är regelbunden påverkar dina egna och din makas eller makes inkomster hemvårdsavgiften.
Tillfällig hemvård kostar lika mycket för alla.
Kommunen kan även ge dig servicesedlar med vilka du kan köpa tjänsten av en serviceproducent som kommunen godkänt.
Hälsa
Om du har hemkommun i Finland kan du utnyttja de offentliga hälsovårdstjänsterna.
När du blir sjuk ska du kontakta hälsostationen i ditt område.
Du får mer information på InfoFinlands sida Hälsotjänsterna i Finland och Äldre människors hälsa.
När du vårdar en närstående i hemmet
När din familjemedlem kontinuerligt behöver hjälp och vården är bindande och krävande kan det vara möjligt att få stöd för närståendevård.
Stödet är avsett för dem som har en hemkommun i Finland.
Stödets storlek och villkoren för att erhålla stödet kan variera mellan olika kommuner.
Man kan ansöka om stödet vid socialbyrån i den egna kommunen.
För att få stöd måste du göra ett avtal om närståendevård med din kommun.
Du får mer information om stöd för närståendevård vid socialbyrån på din egen ort.
Utöver en ersättning kan kommunen ordna även andra tjänster genom vilka vården i hemmet stöds.
Kommunerna ordnar även dagverksamhet för åldringar.
Dagverksamheten innefattar transport, en måltid, motion eller annan verksamhet.
Fråga mer vid socialbyrån på din egen ort.
linkkiPolli.fi:
Information för närståendevårdare(pdf, MB)finska _ engelska _ ryska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska
linkkiNärståendevårdare och Vänner -Förbundet rf:
linkkiNärståendevårdare och Vänner -Förbundet rf:
Stöd för närståendevårdfinska
linkkiSocial- och hälsovårdsministeriet:
Stöd för närståendevårdfinska _ svenska
I Finland ordnar kommunerna tjänster för äldre för att underlätta deras vardag och för att de ska kunna bo hemma så länge som möjligt.
Om du har hemkommun i Finland har du rätt att använda de tjänster som kommunen tillhandahåller.
Boende
Om ditt hem är funktionellt kan du bo hemma även om du har lite svag hälsa.
Du kan låta utföra ändringsarbeten i ditt hem som underlättar boendet.
Det åligger kommunerna att ordna serviceboende och stödboende för personer som behöver det.
Läs mer på InfoFinlands sida Stöd- och serviceboende.
Invandrare som har bott tillräckligt länge i Finland får ålders- eller invalidpension på samma grunder som alla andra som är bosatta i Finland.
Pensionsbeloppet beror på hur länge personen har bott eller arbetat i Finland.
Efter tre års boende tryggar dock garantipensionen ett existensminimum.
Stöden för pensionärerfinska _ svenska _ engelska
Att röra sig
Du kan få låna olika hjälpmedel för att lättare kunna röra på dig, till exempel en käpp eller en rullator.
Om du behöver hjälpmedel ska du först kontakta din egen hälsostation.
Vid hälsostationen får du mer information om hjälpmedlen.
På vintern är det ofta halt ute.
Skomakare och en del stora varuhus säljer halkskydd (liukueste) som kan fästas under sulan på vanliga skor.
Du kan också köpa skor med dubbar (nastakengät) på en skoaffär. Med dem är det lättare att gå på hala gator.
Hemvård
För äldre personer ordnar kommunerna hemvård (kotihoito) som omfattar hjälp med vardagssysslor och sjukvård i hemmet.
Hemvården omfattar hemtjänster, hemsjukvård och stödtjänster.
Hemtjänsterna är hjälp med vardagssysslor, till exempel med att tvätta sig, klä på sig och måltider.
Hemsjukvård är sjukvård och rehabilitering som ges i hemmet.
Remiss för hemsjukvården skrivs av läkare.
Utöver dessa finns det stödtjänster, som är till exempel måltids-, städ-, inköps-, säkerhets- och transporthjälp.
Kontakta hemvårdsenheten i din hemkommun när du behöver hemvård.
Kommunens hemvård är avgiftsbelagd.
När hemvården är regelbunden påverkar dina egna och din makas eller makes inkomster hemvårdsavgiften.
Tillfällig hemvård kostar lika mycket för alla.
Kommunen kan även ge dig servicesedlar med vilka du kan köpa tjänsten av en serviceproducent som kommunen godkänt.
Hälsa
Om du har hemkommun i Finland kan du utnyttja de offentliga hälsovårdstjänsterna.
När du blir sjuk ska du kontakta hälsostationen i ditt område.
Du får mer information på InfoFinlands sida Hälsotjänsterna i Finland.
När du vårdar en närstående i hemmet
När din familjemedlem kontinuerligt behöver hjälp och vården är bindande och krävande kan det vara möjligt att få stöd för närståendevård.
Stödet är avsett för dem som har en hemkommun i Finland.
Stödets storlek och villkoren för att erhålla stödet kan variera mellan olika kommuner.
Man kan ansöka om stödet vid socialbyrån i den egna kommunen.
För att få stöd måste du göra ett avtal om närståendevård med din kommun.
Du får mer information om stöd för närståendevård vid socialbyrån på din egen ort.
Utöver en ersättning kan kommunen ordna även andra tjänster genom vilka vården i hemmet stöds.
Kommunerna ordnar även dagverksamhet för åldringar.
Dagverksamheten innefattar transport, en måltid, motion eller annan verksamhet.
Fråga mer vid socialbyrån på din egen ort.
linkkiPolli.fi:
Information för närståendevårdare(pdf, MB)finska _ engelska _ ryska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska
linkkiNärståendevårdare och Vänner -Förbundet rf:
linkkiNärståendevårdare och Vänner -Förbundet rf:
Stöd för närståendevårdfinska
linkkiSocial- och hälsovårdsministeriet:
Stöd för närståendevårdfinska _ svenska
I Finland ordnar kommunerna tjänster för äldre för att underlätta deras vardag och för att de ska kunna bo hemma så länge som möjligt.
Om du har hemkommun i Finland har du rätt att använda de tjänster som kommunen tillhandahåller.
Boende
Om ditt hem är funktionellt kan du bo hemma även om du har lite svag hälsa.
Du kan låta utföra ändringsarbeten i ditt hem som underlättar boendet.
Det åligger kommunerna att ordna serviceboende och stödboende för personer som behöver det.
Läs mer på InfoFinlands sida Stöd- och serviceboende.
Invandrare som har bott tillräckligt länge i Finland får ålders- eller invalidpension på samma grunder som alla andra som är bosatta i Finland.
Pensionsbeloppet beror på hur länge personen har bott eller arbetat i Finland.
Efter tre års boende tryggar dock garantipensionen ett existensminimum.
Stöden för pensionärerfinska _ svenska _ engelska
Att röra sig
Du kan få låna olika hjälpmedel för att lättare kunna röra på dig, till exempel en käpp eller en rullator.
Om du behöver hjälpmedel ska du först kontakta din egen hälsostation.
Vid hälsostationen får du mer information om hjälpmedlen.
På vintern är det ofta halt ute.
Skomakare och en del stora varuhus säljer halkskydd (liukueste) som kan fästas under sulan på vanliga skor.
Du kan också köpa skor med dubbar (nastakengät) på en skoaffär. Med dem är det lättare att gå på hala gator.
Hemvård
För äldre personer ordnar kommunerna hemvård (kotihoito) som omfattar hjälp med vardagssysslor och sjukvård i hemmet.
Hemvården omfattar hemtjänster, hemsjukvård och stödtjänster.
Hemtjänsterna är hjälp med vardagssysslor, till exempel med att tvätta sig, klä på sig och måltider.
Hemsjukvård är sjukvård och rehabilitering som ges i hemmet.
Remiss för hemsjukvården skrivs av läkare.
Utöver dessa finns det stödtjänster, som är till exempel måltids-, städ-, inköps-, säkerhets- och transporthjälp.
Kontakta hemvårdsenheten i din hemkommun när du behöver hemvård.
Kommunens hemvård är avgiftsbelagd.
När hemvården är regelbunden påverkar dina egna och din makas eller makes inkomster hemvårdsavgiften.
Tillfällig hemvård kostar lika mycket för alla.
Kommunen kan även ge dig servicesedlar med vilka du kan köpa tjänsten av en serviceproducent som kommunen godkänt.
Hälsa
Om du har hemkommun i Finland kan du utnyttja de offentliga hälsovårdstjänsterna.
När du blir sjuk ska du kontakta hälsostationen i ditt område.
Du får mer information på InfoFinlands sida Hälsotjänsterna i Finland.
När du vårdar en närstående i hemmet
När din familjemedlem kontinuerligt behöver hjälp och vården är bindande och krävande kan det vara möjligt att få stöd för närståendevård.
Stödet är avsett för dem som har en hemkommun i Finland.
Stödets storlek och villkoren för att erhålla stödet kan variera mellan olika kommuner.
Man kan ansöka om stödet vid socialbyrån i den egna kommunen.
För att få stöd måste du göra ett avtal om närståendevård med din kommun.
Du får mer information om stöd för närståendevård vid socialbyrån på din egen ort.
Utöver en ersättning kan kommunen ordna även andra tjänster genom vilka vården i hemmet stöds.
Kommunerna ordnar även dagverksamhet för åldringar.
Dagverksamheten innefattar transport, en måltid, motion eller annan verksamhet.
Fråga mer vid socialbyrån på din egen ort.
linkkiPolli.fi:
Information för närståendevårdare(pdf, MB)finska _ engelska _ ryska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska
linkkiNärståendevårdare och Vänner -Förbundet rf:
linkkiNärståendevårdare och Vänner -Förbundet rf:
Stöd för närståendevårdfinska
linkkiSocial- och hälsovårdsministeriet:
Stöd för närståendevårdfinska _ svenska
Småbarnspedagogik är avsedd för barn under skolåldern.
I Finland tillhandahåller kommunerna kommunal småbarnspedagogik bland annat i daghem.
Dessutom finns det privata daghem.
Småbarnspedagogik är fostran, undervisning och omsorg som är pedagogiskt planerad och som har noga genomtänkta mål.
Inom småbarnspedagogiken arbetar utbildade lärare i småbarnspedagogik och barnskötare.
Vanligen vårdar någondera av föräldrarna barnet hemma åtminstone under föräldraledigheten (vanhempainvapaa), det vill säga tills barnet är ungefär 9 månader gammalt.
Om du vårdar ditt barn hemma även efter detta har du rätt att vara ledig från ditt arbete för vård av barn tills barnet fyller tre år.
Mer information om ledigheterna får du på InfoFinlands sida Familjeledighet.
Du kan ansöka från Kela om ekonomiskt stöd för hemvård av barn.
Läs mer på InfoFinlands sida Stöd för vård av barn i hemmet.
Kommunal småbarnspedagogik
Om du har din hemkommun i Finland, kan du ansöka om en plats inom den kommunala småbarnspedagogiken för barnet efter föräldraledigheten.
Då är barnet ca nio månader gammalt.
Om du inte har en hemkommun i Finland, räknas du som invånare i den kommun där du vistas.
Om båda föräldrarna arbetar, har barnet rätt till småbarnspedagogik på heltid.
Om den ena föräldern är hemma, beror rätten till småbarnspedagogik på hemkommunen.
I vissa kommuner har barnet rätt till småbarnspedagogik på heltid även då den ena föräldern är hemma.
I vissa kommuner har barnet rätt till 20 timmar småbarnspedagogik per vecka om den ena föräldern är hemma.
Familjen kan ändå söka rätt till småbarnspedagogik på heltid om barnet behöver särskilt stöd till exempel i att lära sig det finska språket eller på grund av att familjen befinner sig i en svår situation.
Du kan ansöka om en plats
på ett daghem (päiväkoti)
På daghemmet är barnen i större gruppen är i gruppfamiljedagvården.
Familjedagvård innebär att skötaren vårdar barnen i sitt eget hem.
Vissa familjedagvårdare vårdar barnen hemma hos de barn som ingår i gruppen.
Ansök om en plats inom den kommunala småbarnspedagogiken från din egen kommun senast fyra månader innan du behöver den.
Man kan få en plats inom två veckor, om föräldrarna får ett arbete eller en studieplats.
Avgiften för småbarnspedagogik (varhaiskasvatusmaksu) beror på
familjens inkomster
familjens storlek och
på hur många timmar per vecka barnet deltar i småbarnspedagogik.
Man får syskonrabatt.
Om familjen inkomster är mycket låga, kan småbarnspedagogiken vara kostnadsfri för familjen.
Fråga mer i din kommuns rådgivningstjänster.
Privat småbarnspedagogik
En plats inom den privata småbarnspedagogiken kan finnas
i ett privat daghem eller i ett gruppfamiljedaghem
i familjedagvård eller
hemma, då familjen anställer en skötare i hemmet
Du kan ansöka om en plats inom småbarnspedagogiken direkt från det privata daghemmet eller gruppfamiljedaghemmet.
Du kan också leta upp en privat familjedagvårdare som vårdar barnen hemma hos sig, eller anställa en skötare i ditt eget hem.
Om du anställer en skötare i ditt hem blir du en arbetsgivare, och du måste uppfylla en arbetsgivares skyldigheter.
Läs mera på InfoFinlands sida Arbetsgivarens rättigheter och skyldigheter.
Familjen kan anställa en skötare i sitt hem även tillsammans med en annan familj.
Kommunen övervakar den privata småbarnspedagogiken.
Priserna för den privata småbarnspedagogiken varierar.
Du kan ändå få stöd för den från FPA.
Då är den inte nödvändigtvis mycket dyrare än den kommunala småbarnspedagogiken.
Stöd för privat dagvård
Om barnet har en hemkommun i Finland, kan du ansöka om Fpa-stöd för privat vård.
Dagvårdsproducenten måste ha kommunens godkännande.
Du kan ansöka om privatvårdsstöd (yksityisen hoidon tuki), om
ditt barn som är under skolåldern är i privat dagvård; eller
barnet har någon annan privat skötare.
Du kan inte ansöka om privatvårdsstöd om skötaren är en medlem i barnets familj eller om barnet och skötaren bor i samma hushåll.
Du kan inte heller ansöka om privatvårdsstöd för den kommunala småbarnspedagogiken.
Stödets storlek beror bland annat på familjens inkomster och kommunen som familjen bor i.
Kela betalar stödet direkt till skötaren eller dagvårdsproducenten.
Man måste betala skatt för privatvårdsstödet.
Stödet betalas inte till utlandet.
Läs mera om privatvårdsstöd på Fpa:s sidor.
Fpa har en telefontjänst för barnfamiljer.
på finska tfn +358 (0)20 692 206
på svenska och engelska tfn +358 (0)20 692 226
På Fpas byråer får du betjäning även på andra språk med hjälp av en tolk.
Stöd för privat vårdfinska _ svenska _ engelska
Vad händer i småbarnspedagogiken?
Till småbarnspedagogiken hör mångsidig verksamhet, till exempel lekar, motion, utevistelse, musik, pyssel och utfärder.
I dagen ingår också en vilostund.
Målsättningen med verksamheten är att främja barnets utveckling och lärande.
Barnet lär sig även sociala färdigheter.
Barnet får stöd i att lära sig det finska eller svenska språket, om hans/hennes modersmål är ett annat språk.
Om barnet behöver, kan hen även få specialundervisning.
Daghemmet är ändå inte en skola.
Barnen studerar inte skolämnen och har inte lektioner.
Barnen äter tre måltider under dagen: frukost, lunch och mellanmål.
Om ditt barn har en specialdiet ska du berätta om det för lärarna i småbarnspedagogiken.
I småbarnspedagogiken beaktas familjens religion eller livsåskådning.
På vissa orter finns det daghem, som fungerar på andra språk än finska eller svenska.
Vanligen börjar daghemsdagen på morgonen och tar slut på eftermiddagen.
Vissa daghem och familjedagvårdare har öppet dygnet runt med anledning av föräldrarnas arbete eller studier.
linkkiFinlands Flyktinghjälp:
Klubbar
Kommunerna, föreningar och församlingar ordnar dagklubbar för barn.
Klubbarna räcker vanligen ett par timmar.
I klubbarna ordnas handledda lekar, sång, pyssel och annat program.
linkkiUndervisnings- och kulturministeriet:
Information om småbarnspedagogikfinska _ svenska _ engelska
Småbarnspedagogik är avsedd för barn under skolåldern.
I Finland tillhandahåller kommunerna kommunal småbarnspedagogik bland annat i daghem.
Dessutom finns det privata daghem.
Småbarnspedagogik är fostran, undervisning och omsorg som är pedagogiskt planerad och som har noga genomtänkta mål.
Inom småbarnspedagogiken arbetar utbildade lärare i småbarnspedagogik och barnskötare.
Vanligen vårdar någondera av föräldrarna barnet hemma åtminstone under föräldraledigheten (vanhempainvapaa), det vill säga tills barnet är ungefär 9 månader gammalt.
Om du vårdar ditt barn hemma även efter detta har du rätt att vara ledig från ditt arbete för vård av barn tills barnet fyller tre år.
Mer information om ledigheterna får du på InfoFinlands sida Familjeledighet.
Du kan ansöka från Kela om ekonomiskt stöd för hemvård av barn.
Läs mer på InfoFinlands sida Stöd för vård av barn i hemmet.
Kommunal småbarnspedagogik
Om du har din hemkommun i Finland, kan du ansöka om en plats inom den kommunala småbarnspedagogiken för barnet efter föräldraledigheten.
Då är barnet ca nio månader gammalt.
Om du inte har en hemkommun i Finland, räknas du som invånare i den kommun där du vistas.
Om båda föräldrarna arbetar, har barnet rätt till småbarnspedagogik på heltid.
Om den ena föräldern är hemma, beror rätten till småbarnspedagogik på hemkommunen.
I vissa kommuner har barnet rätt till småbarnspedagogik på heltid även då den ena föräldern är hemma.
I vissa kommuner har barnet rätt till 20 timmar småbarnspedagogik per vecka om den ena föräldern är hemma.
Familjen kan ändå söka rätt till småbarnspedagogik på heltid om barnet behöver särskilt stöd till exempel i att lära sig det finska språket eller på grund av att familjen befinner sig i en svår situation.
Du kan ansöka om en plats
på ett daghem (päiväkoti)
På daghemmet är barnen i större gruppen är i gruppfamiljedagvården.
Familjedagvård innebär att skötaren vårdar barnen i sitt eget hem.
Vissa familjedagvårdare vårdar barnen hemma hos de barn som ingår i gruppen.
Ansök om en plats inom den kommunala småbarnspedagogiken från din egen kommun senast fyra månader innan du behöver den.
Man kan få en plats inom två veckor, om föräldrarna får ett arbete eller en studieplats.
Avgiften för småbarnspedagogik (varhaiskasvatusmaksu) beror på
familjens inkomster
familjens storlek och
på hur många timmar per vecka barnet deltar i småbarnspedagogik.
Man får syskonrabatt.
Om familjen inkomster är mycket låga, kan småbarnspedagogiken vara kostnadsfri för familjen.
Fråga mer i din kommuns rådgivningstjänster.
Privat småbarnspedagogik
En plats inom den privata småbarnspedagogiken kan finnas
i ett privat daghem eller i ett gruppfamiljedaghem
i familjedagvård eller
hemma, då familjen anställer en skötare i hemmet
Du kan ansöka om en plats inom småbarnspedagogiken direkt från det privata daghemmet eller gruppfamiljedaghemmet.
Du kan också leta upp en privat familjedagvårdare som vårdar barnen hemma hos sig, eller anställa en skötare i ditt eget hem.
Om du anställer en skötare i ditt hem blir du en arbetsgivare, och du måste uppfylla en arbetsgivares skyldigheter.
Läs mera på InfoFinlands sida Arbetsgivarens rättigheter och skyldigheter.
Familjen kan anställa en skötare i sitt hem även tillsammans med en annan familj.
Kommunen övervakar den privata småbarnspedagogiken.
Priserna för den privata småbarnspedagogiken varierar.
Du kan ändå få stöd för den från FPA.
Då är den inte nödvändigtvis mycket dyrare än den kommunala småbarnspedagogiken.
Stöd för privat dagvård
Om barnet har en hemkommun i Finland, kan du ansöka om Fpa-stöd för privat vård.
Dagvårdsproducenten måste ha kommunens godkännande.
Du kan ansöka om privatvårdsstöd (yksityisen hoidon tuki), om
ditt barn som är under skolåldern är i privat dagvård; eller
barnet har någon annan privat skötare.
Du kan inte ansöka om privatvårdsstöd om skötaren är en medlem i barnets familj eller om barnet och skötaren bor i samma hushåll.
Du kan inte heller ansöka om privatvårdsstöd för den kommunala småbarnspedagogiken.
Stödets storlek beror bland annat på familjens inkomster och kommunen som familjen bor i.
Kela betalar stödet direkt till skötaren eller dagvårdsproducenten.
Man måste betala skatt för privatvårdsstödet.
Stödet betalas inte till utlandet.
Läs mera om privatvårdsstöd på Fpa:s sidor.
Fpa har en telefontjänst för barnfamiljer.
på finska tfn +358 (0)20 692 206
på svenska och engelska tfn +358 (0)20 692 226
På Fpas byråer får du betjäning även på andra språk med hjälp av en tolk.
Stöd för privat vårdfinska _ svenska _ engelska
Vad händer i småbarnspedagogiken?
Till småbarnspedagogiken hör mångsidig verksamhet, till exempel lekar, motion, utevistelse, musik, pyssel och utfärder.
I dagen ingår också en vilostund.
Målsättningen med verksamheten är att främja barnets utveckling och lärande.
Barnet lär sig även sociala färdigheter.
Barnet får stöd i att lära sig det finska eller svenska språket, om hans/hennes modersmål är ett annat språk.
Om barnet behöver, kan hen även få specialundervisning.
Daghemmet är ändå inte en skola.
Barnen studerar inte skolämnen och har inte lektioner.
Barnen äter tre måltider under dagen: frukost, lunch och mellanmål.
Om ditt barn har en specialdiet ska du berätta om det för lärarna i småbarnspedagogiken.
I småbarnspedagogiken beaktas familjens religion eller livsåskådning.
På vissa orter finns det daghem, som fungerar på andra språk än finska eller svenska.
Vanligen börjar daghemsdagen på morgonen och tar slut på eftermiddagen.
Vissa daghem och familjedagvårdare har öppet dygnet runt med anledning av föräldrarnas arbete eller studier.
linkkiFinlands Flyktinghjälp:
Klubbar
Kommunerna, föreningar och församlingar ordnar dagklubbar för barn.
Klubbarna räcker vanligen ett par timmar.
I klubbarna ordnas handledda lekar, sång, pyssel och annat program.
linkkiUndervisnings- och kulturministeriet:
Information om småbarnspedagogikfinska _ svenska _ engelska
Småbarnspedagogik är avsedd för barn under skolåldern.
I Finland tillhandahåller kommunerna kommunal småbarnspedagogik bland annat i daghem.
Dessutom finns det privata daghem.
Småbarnspedagogik är fostran, undervisning och omsorg som är pedagogiskt planerad och som har noga genomtänkta mål.
Inom småbarnspedagogiken arbetar utbildade lärare i småbarnspedagogik och barnskötare.
Vanligen vårdar någondera av föräldrarna barnet hemma åtminstone under föräldraledigheten (vanhempainvapaa), det vill säga tills barnet är ungefär 9 månader gammalt.
Om du vårdar ditt barn hemma även efter detta har du rätt att vara ledig från ditt arbete för vård av barn tills barnet fyller tre år.
Mer information om ledigheterna får du på InfoFinlands sida Familjeledighet.
Du kan ansöka från Kela om ekonomiskt stöd för hemvård av barn.
Läs mer på InfoFinlands sida Stöd för vård av barn i hemmet.
Kommunal småbarnspedagogik
Om du har din hemkommun i Finland, kan du ansöka om en plats inom den kommunala småbarnspedagogiken för barnet efter föräldraledigheten.
Då är barnet ca nio månader gammalt.
Om du inte har en hemkommun i Finland, räknas du som invånare i den kommun där du vistas.
Om båda föräldrarna arbetar, har barnet rätt till småbarnspedagogik på heltid.
Om den ena föräldern är hemma, beror rätten till småbarnspedagogik på hemkommunen.
I vissa kommuner har barnet rätt till småbarnspedagogik på heltid även då den ena föräldern är hemma.
I vissa kommuner har barnet rätt till 20 timmar småbarnspedagogik per vecka om den ena föräldern är hemma.
Familjen kan ändå söka rätt till småbarnspedagogik på heltid om barnet behöver särskilt stöd till exempel i att lära sig det finska språket eller på grund av att familjen befinner sig i en svår situation.
Du kan ansöka om en plats
på ett daghem (päiväkoti)
På daghemmet är barnen i större gruppen är i gruppfamiljedagvården.
Familjedagvård innebär att skötaren vårdar barnen i sitt eget hem.
Vissa familjedagvårdare vårdar barnen hemma hos de barn som ingår i gruppen.
Ansök om en plats inom den kommunala småbarnspedagogiken från din egen kommun senast fyra månader innan du behöver den.
Man kan få en plats inom två veckor, om föräldrarna får ett arbete eller en studieplats.
Avgiften för småbarnspedagogik (varhaiskasvatusmaksu) beror på
familjens inkomster
familjens storlek och
på hur många timmar per vecka barnet deltar i småbarnspedagogik.
Man får syskonrabatt.
Om familjen inkomster är mycket låga, kan småbarnspedagogiken vara kostnadsfri för familjen.
Fråga mer i din kommuns rådgivningstjänster.
Privat småbarnspedagogik
En plats inom den privata småbarnspedagogiken kan finnas
i ett privat daghem eller i ett gruppfamiljedaghem
i familjedagvård eller
hemma, då familjen anställer en skötare i hemmet
Du kan ansöka om en plats inom småbarnspedagogiken direkt från det privata daghemmet eller gruppfamiljedaghemmet.
Du kan också leta upp en privat familjedagvårdare som vårdar barnen hemma hos sig, eller anställa en skötare i ditt eget hem.
Om du anställer en skötare i ditt hem blir du en arbetsgivare, och du måste uppfylla en arbetsgivares skyldigheter.
Läs mera på InfoFinlands sida Arbetsgivarens rättigheter och skyldigheter.
Familjen kan anställa en skötare i sitt hem även tillsammans med en annan familj.
Kommunen övervakar den privata småbarnspedagogiken.
Priserna för den privata småbarnspedagogiken varierar.
Du kan ändå få stöd för den från FPA.
Då är den inte nödvändigtvis mycket dyrare än den kommunala småbarnspedagogiken.
Stöd för privat dagvård
Om barnet har en hemkommun i Finland, kan du ansöka om Fpa-stöd för privat vård.
Dagvårdsproducenten måste ha kommunens godkännande.
Du kan ansöka om privatvårdsstöd (yksityisen hoidon tuki), om
ditt barn som är under skolåldern är i privat dagvård; eller
barnet har någon annan privat skötare.
Du kan inte ansöka om privatvårdsstöd om skötaren är en medlem i barnets familj eller om barnet och skötaren bor i samma hushåll.
Du kan inte heller ansöka om privatvårdsstöd för den kommunala småbarnspedagogiken.
Stödets storlek beror bland annat på familjens inkomster och kommunen som familjen bor i.
Kela betalar stödet direkt till skötaren eller dagvårdsproducenten.
Man måste betala skatt för privatvårdsstödet.
Stödet betalas inte till utlandet.
Läs mera om privatvårdsstöd på Fpa:s sidor.
Fpa har en telefontjänst för barnfamiljer.
på finska tfn +358 (0)20 692 206
på svenska och engelska tfn +358 (0)20 692 226
På Fpas byråer får du betjäning även på andra språk med hjälp av en tolk.
Stöd för privat vårdfinska _ svenska _ engelska
Vad händer i småbarnspedagogiken?
Till småbarnspedagogiken hör mångsidig verksamhet, till exempel lekar, motion, utevistelse, musik, pyssel och utfärder.
I dagen ingår också en vilostund.
Målsättningen med verksamheten är att främja barnets utveckling och lärande.
Barnet lär sig även sociala färdigheter.
Barnet får stöd i att lära sig det finska eller svenska språket, om hans/hennes modersmål är ett annat språk.
Om barnet behöver, kan hen även få specialundervisning.
Daghemmet är ändå inte en skola.
Barnen studerar inte skolämnen och har inte lektioner.
Barnen äter tre måltider under dagen: frukost, lunch och mellanmål.
Om ditt barn har en specialdiet ska du berätta om det för lärarna i småbarnspedagogiken.
I småbarnspedagogiken beaktas familjens religion eller livsåskådning.
På vissa orter finns det daghem, som fungerar på andra språk än finska eller svenska.
Vanligen börjar daghemsdagen på morgonen och tar slut på eftermiddagen.
Vissa daghem och familjedagvårdare har öppet dygnet runt med anledning av föräldrarnas arbete eller studier.
linkkiFinlands Flyktinghjälp:
Klubbar
Kommunerna, föreningar och församlingar ordnar dagklubbar för barn.
Klubbarna räcker vanligen ett par timmar.
I klubbarna ordnas handledda lekar, sång, pyssel och annat program.
linkkiUndervisnings- och kulturministeriet:
Information om småbarnspedagogikfinska _ svenska _ engelska
På den här sidan finns information om tjänsterna i Rovaniemi.
Nödfall
När du är sjuk
Akutmottagningen
Tandvård
Mental hälsa
Nödfall
Ett nödfall är en verklig och akut farlig situation där ens liv, hälsa, egendom eller miljön är hotad.
I nödsituationer ska du alltid ringa nödnumret 112.
Mer information hittar du på Nödcentralsverkets webbplats.
Nödcentralsverketfinska _ svenska _ engelska
När du är sjuk
I Rovaniemi finns två hälsostationer:
linkkiHälsovårdscentralen:
Hälsostationen på Rinteenkulmafinska
linkkiHälsovårdscentralen:
Hälsostationen på Pulkamontiefinska
I brådskande situationer kan du ringa vårdteamet för ditt eget område.
Du får en tid på mottagningen inom 1–3 dagar.
Brådskande ärenden är till exempel bihåleinflammation, ögoninfektion, ryggvärk, en lindrig urinvägsinfektion, en vaginal infektion eller eksem.
Akutmottagningen
Du kan gå till akutmottagningen vid akuta sjukfall där du inte kan vänta till följande dag på vård. Sådana fall är till exempel blödande sår, bröstsmärtor, brännskador med mera.
dagtid kl. 8–22
Jourmottagningen vid
Lapplands centralsjukhus
Ounasrinteentie 22
tfn 016 328 2140
nattetid kl. 22–8
Akutmottagningen vid Lapplands centralsjukhus
Ounasrinteentie 22
tfn 016 328 2100
På natten vårdas endast nödfall.
Tandvård
Tandvårdens tidsbeställning och värkjouren nås vardagar kl. 8–15 på tfn 016 322 2562 eller 016 356 1750. Kvällstid och på veckoslut kan du ta kontakt med läkarmottagningen om du är i brådskande behov av vård.
Tfn 016 322 4900.
Tandvården vid hälsovårdscentralen är avgiftsfri för barn under 18 år.
Om du har bokat en tid hos tandläkaren, men inte kan komma på avtalad tid ska du komma ihåg att avboka din tid.
Om du inte avbokar debiteras du på en avgift om 27 euro.
Du kan även gå till en privat tandläkarmottagning.
Mental hälsa
Om du behöver hjälp med något som rör den mentala hälsan, kan du kontakta mentalvårdsenheten.
Mentalvårdsenheterna har verksamhet på två adresser:
tfn 016 322 2269
Pulkamontie 6, vån. 2
tfn 016 322 4600
På den här sidan finns information om tjänsterna i Rovaniemi.
Nödfall
När du är sjuk
Akutmottagningen
Tandvård
Mental hälsa
Nödfall
Ett nödfall är en verklig och akut farlig situation där ens liv, hälsa, egendom eller miljön är hotad.
I nödsituationer ska du alltid ringa nödnumret 112.
Mer information hittar du på Nödcentralsverkets webbplats.
Nödcentralsverketfinska _ svenska _ engelska
När du är sjuk
I Rovaniemi finns två hälsostationer:
linkkiHälsovårdscentralen:
Hälsostationen på Rinteenkulmafinska
linkkiHälsovårdscentralen:
Hälsostationen på Pulkamontiefinska
I brådskande situationer kan du ringa vårdteamet för ditt eget område.
Du får en tid på mottagningen inom 1–3 dagar.
Brådskande ärenden är till exempel bihåleinflammation, ögoninfektion, ryggvärk, en lindrig urinvägsinfektion, en vaginal infektion eller eksem.
Akutmottagningen
Du kan gå till akutmottagningen vid akuta sjukfall där du inte kan vänta till följande dag på vård. Sådana fall är till exempel blödande sår, bröstsmärtor, brännskador med mera.
dagtid kl. 8–22
Jourmottagningen vid
Lapplands centralsjukhus
Ounasrinteentie 22
tfn 016 328 2140
nattetid kl. 22–8
Akutmottagningen vid Lapplands centralsjukhus
Ounasrinteentie 22
tfn 016 328 2100
På natten vårdas endast nödfall.
Tandvård
Tandvårdens tidsbeställning och värkjouren nås vardagar kl. 8–15 på tfn 016 322 2562 eller 016 356 1750. Kvällstid och på veckoslut kan du ta kontakt med läkarmottagningen om du är i brådskande behov av vård.
Tfn 016 322 4900.
Tandvården vid hälsovårdscentralen är avgiftsfri för barn under 18 år.
Om du har bokat en tid hos tandläkaren, men inte kan komma på avtalad tid ska du komma ihåg att avboka din tid.
Om du inte avbokar debiteras du på en avgift om 27 euro.
Du kan även gå till en privat tandläkarmottagning.
Mental hälsa
Om du behöver hjälp med något som rör den mentala hälsan, kan du kontakta mentalvårdsenheten.
Mentalvårdsenheterna har verksamhet på två adresser:
tfn 016 322 2269
Pulkamontie 6, vån. 2
tfn 016 322 4600
På den här sidan finns information om tjänsterna i Rovaniemi.
Nödfall
När du är sjuk
Akutmottagningen
Tandvård
Mental hälsa
Nödfall
Ett nödfall är en verklig och akut farlig situation där ens liv, hälsa, egendom eller miljön är hotad.
I nödsituationer ska du alltid ringa nödnumret 112.
Mer information hittar du på Nödcentralsverkets webbplats.
Nödcentralsverketfinska _ svenska _ engelska
När du är sjuk
I Rovaniemi finns två hälsostationer:
linkkiHälsovårdscentralen:
Hälsostationen på Rinteenkulmafinska
linkkiHälsovårdscentralen:
Hälsostationen på Pulkamontiefinska
I brådskande situationer kan du ringa vårdteamet för ditt eget område.
Du får en tid på mottagningen inom 1–3 dagar.
Brådskande ärenden är till exempel bihåleinflammation, ögoninfektion, ryggvärk, en lindrig urinvägsinfektion, en vaginal infektion eller eksem.
Akutmottagningen
Du kan gå till akutmottagningen vid akuta sjukfall där du inte kan vänta till följande dag på vård. Sådana fall är till exempel blödande sår, bröstsmärtor, brännskador med mera.
dagtid kl. 8–22
Jourmottagningen vid
Lapplands centralsjukhus
Ounasrinteentie 22
tfn 016 328 2140
nattetid kl. 22–8
Akutmottagningen vid Lapplands centralsjukhus
Ounasrinteentie 22
tfn 016 328 2100
På natten vårdas endast nödfall.
Tandvård
Tandvårdens tidsbeställning och värkjouren nås vardagar kl. 8–15 på tfn 016 322 2562 eller 016 356 1750. Kvällstid och på veckoslut kan du ta kontakt med läkarmottagningen om du är i brådskande behov av vård.
Tfn 016 322 4900.
Tandvården vid hälsovårdscentralen är avgiftsfri för barn under 18 år.
Om du har bokat en tid hos tandläkaren, men inte kan komma på avtalad tid ska du komma ihåg att avboka din tid.
Om du inte avbokar debiteras du på en avgift om 27 euro.
Du kan även gå till en privat tandläkarmottagning.
Mental hälsa
Om du behöver hjälp med något som rör den mentala hälsan, kan du kontakta mentalvårdsenheten.
Mentalvårdsenheterna har verksamhet på två adresser:
tfn 016 322 2269
Pulkamontie 6, vån. 2
tfn 016 322 4600
Familjer kan få olika slags understöd för sina levnadskostnader.
Förutsättningen för att få de flesta understöden är att du omfattas av den sociala tryggheten i Finland eller att du har hemkommun i Finland.
Om familjens pengar inte räcker till att betala hyran för bostaden eller kostnaderna för en ägarbostad kan familjen ansöka om allmänt bostadsbidrag vid Fpa.
Om barnets vårdnadshavare är pensionerad kan han eller hon ansöka om en barnförhöjning på sin pension från Fpa.
Fpa betalar barnförhöjningen tills barnet fyller 16 år.
Familjen kan ansöka om utkomststöd om den har ekonomiska problem som den inte klarar av annars.
Utkomststöd söks hos FPA.
Om du hemma vårdar en långtidssjuk, handikappad eller äldre familjemedlem kan din hemkommun betala stöd för närståendevård (omaishoidontuki) till dig.
Du kan ansöka om stöd för närståendevård hos socialbyrån i din hemkommun.
Läs mer på InfoFinlands sida Ekonomiskt stöd och under rubriken När du vårdar en närstående i hemmet på sidan Äldre människor.
På InfoFinlands sida Familjer med en förälder finns information om hurdant understöd den vårdnadshavare som bor med sitt barn kan få om föräldrarna inte bor tillsammans.
Underhållsbidraget är ett bidrag som den förälder som inte bor med barnet betalar för att delta i barnets levnadskostnader.
Den förälder som inte bor med barnet betalar underhållsbidrag till den förälder hos vilken barnet bor officiellt.
Barnförhöjningfinska _ svenska _ engelska
Familjer kan få olika slags understöd för sina levnadskostnader.
Förutsättningen för att få de flesta understöden är att du omfattas av den sociala tryggheten i Finland eller att du har hemkommun i Finland.
Om familjens pengar inte räcker till att betala hyran för bostaden eller kostnaderna för en ägarbostad kan familjen ansöka om allmänt bostadsbidrag vid Fpa.
Om barnets vårdnadshavare är pensionerad kan han eller hon ansöka om en barnförhöjning på sin pension från Fpa.
Fpa betalar barnförhöjningen tills barnet fyller 16 år.
Familjen kan ansöka om utkomststöd om den har ekonomiska problem som den inte klarar av annars.
Utkomststöd söks hos FPA.
Om du hemma vårdar en långtidssjuk, handikappad eller äldre familjemedlem kan din hemkommun betala stöd för närståendevård (omaishoidontuki) till dig.
Du kan ansöka om stöd för närståendevård hos socialbyrån i din hemkommun.
Läs mer på InfoFinlands sida Ekonomiskt stöd och under rubriken När du vårdar en närstående i hemmet på sidan Äldre människor.
På InfoFinlands sida Familjer med en förälder finns information om hurdant understöd den vårdnadshavare som bor med sitt barn kan få om föräldrarna inte bor tillsammans.
Underhållsbidraget är ett bidrag som den förälder som inte bor med barnet betalar för att delta i barnets levnadskostnader.
Den förälder som inte bor med barnet betalar underhållsbidrag till den förälder hos vilken barnet bor officiellt.
Barnförhöjningfinska _ svenska _ engelska
Familjer kan få olika slags understöd för sina levnadskostnader.
Förutsättningen för att få de flesta understöden är att du omfattas av den sociala tryggheten i Finland eller att du har hemkommun i Finland.
Om familjens pengar inte räcker till att betala hyran för bostaden eller kostnaderna för en ägarbostad kan familjen ansöka om allmänt bostadsbidrag vid Fpa.
Om barnets vårdnadshavare är pensionerad kan han eller hon ansöka om en barnförhöjning på sin pension från Fpa.
Fpa betalar barnförhöjningen tills barnet fyller 16 år.
Familjen kan ansöka om utkomststöd om den har ekonomiska problem som den inte klarar av annars.
Utkomststöd söks hos FPA.
Om du hemma vårdar en långtidssjuk, handikappad eller äldre familjemedlem kan din hemkommun betala stöd för närståendevård (omaishoidontuki) till dig.
Du kan ansöka om stöd för närståendevård hos socialbyrån i din hemkommun.
Läs mer på InfoFinlands sida Ekonomiskt stöd och under rubriken När du vårdar en närstående i hemmet på sidan Äldre människor.
På InfoFinlands sida Familjer med en förälder finns information om hurdant understöd den vårdnadshavare som bor med sitt barn kan få om föräldrarna inte bor tillsammans.
Underhållsbidraget är ett bidrag som den förälder som inte bor med barnet betalar för att delta i barnets levnadskostnader.
Den förälder som inte bor med barnet betalar underhållsbidrag till den förälder hos vilken barnet bor officiellt.
Barnförhöjningfinska _ svenska _ engelska
FPA betalar ut barnbidrag för varje barn som bor i Finland och omfattas av den sociala tryggheten i Finland.
Barnbidrag betalas ut fram till dess att barnet fyller 17 år.
Du kan ansöka om barnbidrag från FPA antingen via FPA:s webbsidor eller med en pappersblankett.
Webbtjänsten är på finska och svenska.
Du kan ansöka om barnbidrag på samma gång som du ansöker om moderskapspenning.
Ansök om barnbidrag i tid, du kan få barnbidrag retroaktivt för en period på högst sex månader.
Barnbidraget för det första barnet uppgår till cirka 100 euro per månad.
Barnbidragsbeloppet är en aning högre för varje följande barn.
En förälder som bor ensam med ett eller flera barn kan få förhöjt barnbidrag.
Barnbidrag betalas ut månatligen antingen till moderns, faderns eller en annan vårdnadshavares bankkonto.
Ingen skatt tas ut på barnbidrag.
I vissa situationer kan barnbidrag också betalas ut till utlandet, om du eller din make/maka omfattas av den sociala tryggheten i Finland.
Läs på FPA:s webbsidor när familjeförmåner betalas ut till utlandet.
Sköta ärenden på Internetfinska _ svenska _ engelska
Kontaktuppgifter till FPAfinska _ svenska _ engelska
Elektronisk tidsbeställningfinska _ svenska _ engelska
FPA betalar ut barnbidrag för varje barn som bor i Finland och omfattas av den sociala tryggheten i Finland.
Barnbidrag betalas ut fram till dess att barnet fyller 17 år.
Du kan ansöka om barnbidrag från FPA antingen via FPA:s webbsidor eller med en pappersblankett.
Webbtjänsten är på finska och svenska.
Du kan ansöka om barnbidrag på samma gång som du ansöker om moderskapspenning.
Ansök om barnbidrag i tid, du kan få barnbidrag retroaktivt för en period på högst sex månader.
Barnbidraget för det första barnet uppgår till cirka 100 euro per månad.
Barnbidragsbeloppet är en aning högre för varje följande barn.
En förälder som bor ensam med ett eller flera barn kan få förhöjt barnbidrag.
Barnbidrag betalas ut månatligen antingen till moderns, faderns eller en annan vårdnadshavares bankkonto.
Ingen skatt tas ut på barnbidrag.
I vissa situationer kan barnbidrag också betalas ut till utlandet, om du eller din make/maka omfattas av den sociala tryggheten i Finland.
Läs på FPA:s webbsidor när familjeförmåner betalas ut till utlandet.
Sköta ärenden på Internetfinska _ svenska _ engelska
Kontaktuppgifter till FPAfinska _ svenska _ engelska
Elektronisk tidsbeställningfinska _ svenska _ engelska
FPA betalar ut barnbidrag för varje barn som bor i Finland och omfattas av den sociala tryggheten i Finland.
Barnbidrag betalas ut fram till dess att barnet fyller 17 år.
Du kan ansöka om barnbidrag från FPA antingen via FPA:s webbsidor eller med en pappersblankett.
Webbtjänsten är på finska och svenska.
Du kan ansöka om barnbidrag på samma gång som du ansöker om moderskapspenning.
Ansök om barnbidrag i tid, du kan få barnbidrag retroaktivt för en period på högst sex månader.
Barnbidraget för det första barnet uppgår till cirka 100 euro per månad.
Barnbidragsbeloppet är en aning högre för varje följande barn.
En förälder som bor ensam med ett eller flera barn kan få förhöjt barnbidrag.
Barnbidrag betalas ut månatligen antingen till moderns, faderns eller en annan vårdnadshavares bankkonto.
Ingen skatt tas ut på barnbidrag.
I vissa situationer kan barnbidrag också betalas ut till utlandet, om du eller din make/maka omfattas av den sociala tryggheten i Finland.
Läs på FPA:s webbsidor när familjeförmåner betalas ut till utlandet.
Sköta ärenden på Internetfinska _ svenska _ engelska
Kontaktuppgifter till FPAfinska _ svenska _ engelska
Elektronisk tidsbeställningfinska _ svenska _ engelska
Vanligen vårdar någondera av föräldrarna barnet i hemmet åtminstone under föräldraledigheten, det vill säga tills barnet är ca 9 månader gammalt.
Efter föräldraledigheten kan barnet börja i dagvård eller någondera av föräldrarna kan vårda barnet hemma.
Läs mer om dagvård på InfoFinlands sida Dagvård.
Hemvårdsstöd
Om du vårdar ett barn som är yngre än tre år hemma kan du ansöka om hemvårdsstöd från Fpa. Skötaren kan till exempel vara barnets vårdnadshavare eller annan släkting.
Du kan inte få hemvårdsstöd om barnet går i den kommunala dagvården.
Hemvårdsstöd betalas vanligen inte till utlandet.
Be Fpa om mera information.
FPA betalar hemvårdsstöd om
den ena föräldern eller båda föräldrarna har hemkommun i Finland eller
minst en av föräldrarna arbetar i Finland och därmed omfattas av den sociala tryggheten i Finland.
Hemvårdsstödet består av en vårdpenning och ett vårdtillägg som är beroende av familjens inkomster samt ett eventuellt kommuntillägg.
Fråga vid socialbyrån om kommuntillägg betalas i din kommun.
Hemvårdsstödets vårdpenning är lika stor för alla; beloppet påverkas inte av familjens inkomster.
Hemvårdsstödet är skattepliktig inkomst.
Hemvårdsstöd kan i vissa fall även betalas till familjemedlemmar som vistas i ett annat EU- eller EES-land.
Fråga mer på FPA.
Information om hemvårdsstödfinska _ svenska _ engelska
Vårdledighet
Om du vårdar barnet i hemmet har du rätt att ta ut oavlönad vårdledighet från ditt arbete ända tills barnet fyller tre år.
Under vårdledigheten kan du ansöka om hemvårdsstöd av Fpa.
Du kan ta ut vårdledighet om du har befunnit dig i samma arbetsgivares tjänst under minst 6 månader under det senaste året.
Meddela arbetsgivaren om vårdledigheten senast 2 månader innan den börjar.
Flexibel och partiell vårdpenning
Du kan också vara partiellt vårdledig.
Då arbetar du kortare dagar och får på motsvarande sätt mindre lön.
Om du har hemkommun i Finland kan du ansöka om flexibel vårdpenning (joustava hoitoraha) för vård av barn under tre år och partiell vårdpenning (osittainen hoitoraha) för vård av skolbarn i årskurserna 1 eller 2 hos FPA.
Flexibel eller partiell vårdpenning betalas inte för vård av ett barn som fyllt tre, men som ännu inte går i skolan.
Ett barn under tre år kan vara i kommunal dagvård på deltid under tiden för flexibel vårdledighet.
Du kan ansöka om flexibel eller partiell vårdpenning om du förkortar din normala arbetstid så att du arbetar högst 30 timmar i veckan för att ta hand om barnet.
Modern och fadern kan få flexibel eller partiell vårdpenning samtidigt om båda har förkortat sin arbetstid och tar hand om barnet under olika tider.
Vårdpenning betalas bara för ett barn i taget och är skattepliktig inkomst.
Du kan inte få flexibel eller partiell vårdpenning om du får föräldradagpenning och/eller hemvårdsstöd och själv tar hand om dina barn.
Information om stöd till barnfamiljerfinska _ svenska _ engelska
linkkiSkattemyndigheten:
Skattekortfinska _ svenska _ engelska
Vanligen vårdar någondera av föräldrarna barnet i hemmet åtminstone under föräldraledigheten, det vill säga tills barnet är ca 9 månader gammalt.
Efter föräldraledigheten kan barnet börja i dagvård eller någondera av föräldrarna kan vårda barnet hemma.
Läs mer om dagvård på InfoFinlands sida Dagvård.
Hemvårdsstöd
Om du vårdar ett barn som är yngre än tre år hemma kan du ansöka om hemvårdsstöd från Fpa. Skötaren kan till exempel vara barnets vårdnadshavare eller annan släkting.
Du kan inte få hemvårdsstöd om barnet går i den kommunala dagvården.
Hemvårdsstöd betalas vanligen inte till utlandet.
Be Fpa om mera information.
FPA betalar hemvårdsstöd om
den ena föräldern eller båda föräldrarna har hemkommun i Finland eller
minst en av föräldrarna arbetar i Finland och därmed omfattas av den sociala tryggheten i Finland.
Hemvårdsstödet består av en vårdpenning och ett vårdtillägg som är beroende av familjens inkomster samt ett eventuellt kommuntillägg.
Fråga vid socialbyrån om kommuntillägg betalas i din kommun.
Hemvårdsstödets vårdpenning är lika stor för alla; beloppet påverkas inte av familjens inkomster.
Hemvårdsstödet är skattepliktig inkomst.
Hemvårdsstöd kan i vissa fall även betalas till familjemedlemmar som vistas i ett annat EU- eller EES-land.
Fråga mer på FPA.
Information om hemvårdsstödfinska _ svenska _ engelska
Vårdledighet
Om du vårdar barnet i hemmet har du rätt att ta ut oavlönad vårdledighet från ditt arbete ända tills barnet fyller tre år.
Under vårdledigheten kan du ansöka om hemvårdsstöd av Fpa.
Du kan ta ut vårdledighet om du har befunnit dig i samma arbetsgivares tjänst under minst 6 månader under det senaste året.
Meddela arbetsgivaren om vårdledigheten senast 2 månader innan den börjar.
Flexibel och partiell vårdpenning
Du kan också vara partiellt vårdledig.
Då arbetar du kortare dagar och får på motsvarande sätt mindre lön.
Om du har hemkommun i Finland kan du ansöka om flexibel vårdpenning (joustava hoitoraha) för vård av barn under tre år och partiell vårdpenning (osittainen hoitoraha) för vård av skolbarn i årskurserna 1 eller 2 hos FPA.
Flexibel eller partiell vårdpenning betalas inte för vård av ett barn som fyllt tre, men som ännu inte går i skolan.
Ett barn under tre år kan vara i kommunal dagvård på deltid under tiden för flexibel vårdledighet.
Du kan ansöka om flexibel eller partiell vårdpenning om du förkortar din normala arbetstid så att du arbetar högst 30 timmar i veckan för att ta hand om barnet.
Modern och fadern kan få flexibel eller partiell vårdpenning samtidigt om båda har förkortat sin arbetstid och tar hand om barnet under olika tider.
Vårdpenning betalas bara för ett barn i taget och är skattepliktig inkomst.
Du kan inte få flexibel eller partiell vårdpenning om du får föräldradagpenning och/eller hemvårdsstöd och själv tar hand om dina barn.
Information om stöd till barnfamiljerfinska _ svenska _ engelska
linkkiSkattemyndigheten:
Skattekortfinska _ svenska _ engelska
Vanligen vårdar någondera av föräldrarna barnet i hemmet åtminstone under föräldraledigheten, det vill säga tills barnet är ca 9 månader gammalt.
Efter föräldraledigheten kan barnet börja i dagvård eller någondera av föräldrarna kan vårda barnet hemma.
Läs mer om dagvård på InfoFinlands sida Dagvård.
Hemvårdsstöd
Om du vårdar ett barn som är yngre än tre år hemma kan du ansöka om hemvårdsstöd från Fpa. Skötaren kan till exempel vara barnets vårdnadshavare eller annan släkting.
Du kan inte få hemvårdsstöd om barnet går i den kommunala dagvården.
Hemvårdsstöd betalas vanligen inte till utlandet.
Be Fpa om mera information.
FPA betalar hemvårdsstöd om
den ena föräldern eller båda föräldrarna har hemkommun i Finland eller
minst en av föräldrarna arbetar i Finland och därmed omfattas av den sociala tryggheten i Finland.
Hemvårdsstödet består av en vårdpenning och ett vårdtillägg som är beroende av familjens inkomster samt ett eventuellt kommuntillägg.
Fråga vid socialbyrån om kommuntillägg betalas i din kommun.
Hemvårdsstödets vårdpenning är lika stor för alla; beloppet påverkas inte av familjens inkomster.
Hemvårdsstödet är skattepliktig inkomst.
Hemvårdsstöd kan i vissa fall även betalas till familjemedlemmar som vistas i ett annat EU- eller EES-land.
Fråga mer på FPA.
Information om hemvårdsstödfinska _ svenska _ engelska
Vårdledighet
Om du vårdar barnet i hemmet har du rätt att ta ut oavlönad vårdledighet från ditt arbete ända tills barnet fyller tre år.
Under vårdledigheten kan du ansöka om hemvårdsstöd av Fpa.
Du kan ta ut vårdledighet om du har befunnit dig i samma arbetsgivares tjänst under minst 6 månader under det senaste året.
Meddela arbetsgivaren om vårdledigheten senast 2 månader innan den börjar.
Flexibel och partiell vårdpenning
Du kan också vara partiellt vårdledig.
Då arbetar du kortare dagar och får på motsvarande sätt mindre lön.
Om du har hemkommun i Finland kan du ansöka om flexibel vårdpenning (joustava hoitoraha) för vård av barn under tre år och partiell vårdpenning (osittainen hoitoraha) för vård av skolbarn i årskurserna 1 eller 2 hos FPA.
Flexibel eller partiell vårdpenning betalas inte för vård av ett barn som fyllt tre, men som ännu inte går i skolan.
Ett barn under tre år kan vara i kommunal dagvård på deltid under tiden för flexibel vårdledighet.
Du kan ansöka om flexibel eller partiell vårdpenning om du förkortar din normala arbetstid så att du arbetar högst 30 timmar i veckan för att ta hand om barnet.
Modern och fadern kan få flexibel eller partiell vårdpenning samtidigt om båda har förkortat sin arbetstid och tar hand om barnet under olika tider.
Vårdpenning betalas bara för ett barn i taget och är skattepliktig inkomst.
Du kan inte få flexibel eller partiell vårdpenning om du får föräldradagpenning och/eller hemvårdsstöd och själv tar hand om dina barn.
Information om stöd till barnfamiljerfinska _ svenska _ engelska
linkkiSkattemyndigheten:
Skattekortfinska _ svenska _ engelska
Efter att barnet fötts sköter vanligtvis en av föräldrarna barnet hemma i en viss tid.
Under denna tid betalar FPA ut olika föräldradagpenningar (vanhempainpäiväraha).
Föräldradagpenningarna omfattar
moderskapspenning och särskild moderskapspenning
föräldrapenning
faderskapspenning.
Därtill utbetalas barnbidrag (lapsilisä) till barnets vårdnadshavare fram till dess att barnet fyller 17 år.
Läs mer på InfoFinlands sida Barnbidrag.
Ansökan om föräldradagpenningar
Du kan ansöka om föräldradagpenningar om du omfattas av den sociala tryggheten i Finland och varit sjukförsäkrad i Finland, ett annat EU- eller EES-land eller Schweiz oavbrutet i 180 dagar före det beräknade förslossningsdatumet.
Du kan göra en ansökan om föräldradagpenning på FPA:s webbsidor.
Logga in med nätbankskoder eller ett mobilcertifikat.
Tjänsten innehåller anvisningar för att fylla i ansökan.
På samma adress ser du också hur behandlingen av din ansökan framskrider.
När ansökan avgjorts, ser du beloppet på ditt stöd och tidpunkten för utbetalningen.
Tjänsten är på finska och svenska.
Du kan ansöka om föräldradagpenningar också genom att fylla i en pappersblankett och skicka den jämte nödvändiga bilagor till vilken FPA-byrå som helst.
Rådgivningen hjälper dig att fylla i ansökan.
Beloppet på din föräldradagpenning beror på hur höga inkomster du har.
Dagpenningen är alltid lägre än lönen, vanligen cirka 70 procent av inkomsterna.
Om du inte har några inkomster, får du föräldradagpenningens minimibelopp.
Också en arbetslös förälder har rätt till föräldradagpenning.
Om din arbetsgivare betalar ut lön till dig under föräldradagpenningperioden, betalar FPA dagpenningen till din arbetsgivare.
Meddela din arbetsgivare om din föräldraledighet två månader innan den börjar.
Om din ledighet varar i 12 vardagar eller mindre, ska du meddela om ledigheten till din arbetsgivare en månad på förhand.
Läs mer på InfoFinlands sida Familjeledighet.
Föräldradagpenningar är skattepliktiga inkomster och följaktligen behöver du ett skattekort (verokortti).
Läs mer på InfoFinlands sida Beskattning.
linkkiSkattemyndigheten:
Skattekortfinska _ svenska _ engelska
Moderskapspenningperioden varar i cirka tre månader.
Den börjar vanligen 30 vardagar för det beräknade förlossningsdatumet.
Läs mer på InfoFinlands sidor Stöd till gravida.
Föräldrapenning
Efter utgången av moderskapspenningperioden kan en av vårdnadshavarna ta ut föräldraledighet.
I så fall sköter en av föräldrarna barnet hemma och får en föräldrapenning.
Ansökan ska lämnas in till FPA senast en månad innan moderskapspenningperiodens utgång och föräldrapenningperiodens början.
Föräldrapenningperioden varar i cirka sex månader.
Om familjen får tvillingar är föräldrapenningperioden 60 vardagar längre.
Modern ska genomgå en läkarundersökning 5–12 veckor efter förlossningen och skicka läkarintyget till FPA.
Annars utbetalas inte föräldradagpenning.
Vilken som helst av vårdnadshavarna kan vara föräldraledig.
De kan också vara lediga turvis.
Föräldrarna kan också arbeta deltid och tillsammans sköta barnet på deltid.
Under denna tid betalar FPA partiell föräldrapenning till bägge föräldrar.
Om en av föräldrarna vill sköta barnet hemma efter föräldrapenningperioden, kan han eller hon få hemvårdsstöd.
Läs mer på InfoFinlands sida Stöd för vård av barn i hemmet.
Föräldrapenning till modern eller fadernfinska _ svenska _ engelska
Faderskapspenning
Faderskapspenningen (Isyysraha) är avsedd för fadern då han tar hand om barnet.
FPA (Kela) betalar ut faderskapspenning under faderskapsledigheten.
Du kan ansöka om faderskapspenning även om du är till exempel företagare, arbetslös eller studerande.
Faderskapspenning betalas ut för 54 vardagar, alltså ungefär nio veckor.
Dessa dagar kan inte överföras till modern.
Du får själv bestämma om du tar ut alla faderskapspenningdagar eller bara en del av dem.
Du får faderskapspenning även om du inte bor tillsammans med barnets mor.
Du kan vara pappaledig samtidigt som barnets mor är mamma- eller föräldraledig.
Då kan du ta ut högst 18 faderskapspenningdagar.
Du kan också ta ut alla 54 faderskapspenningdagar separat, till exempel efter föräldraledigheten.
De 1–18 vardagar av faderskapsledigheten som du kan ta ut samtidigt med barnets mor kan delas upp i högst fyra perioder.
Faderskapsledighet som tas ut efter föräldrapenningperioden kan delas upp i högst två perioder.
Du kan endast använda faderskapspenningdagar för vård av ett barn under två år.
När barnet fyller två år kan du inte längre använda dina faderskapspenningdagar även om sådana finns kvar.
Efter att barnet fötts sköter vanligtvis en av föräldrarna barnet hemma i en viss tid.
Under denna tid betalar FPA ut olika föräldradagpenningar (vanhempainpäiväraha).
Föräldradagpenningarna omfattar
moderskapspenning och särskild moderskapspenning
föräldrapenning
faderskapspenning.
Därtill utbetalas barnbidrag (lapsilisä) till barnets vårdnadshavare fram till dess att barnet fyller 17 år.
Läs mer på InfoFinlands sida Barnbidrag.
Ansökan om föräldradagpenningar
Du kan ansöka om föräldradagpenningar om du omfattas av den sociala tryggheten i Finland och varit sjukförsäkrad i Finland, ett annat EU- eller EES-land eller Schweiz oavbrutet i 180 dagar före det beräknade förslossningsdatumet.
Du kan göra en ansökan om föräldradagpenning på FPA:s webbsidor.
Logga in med nätbankskoder eller ett mobilcertifikat.
Tjänsten innehåller anvisningar för att fylla i ansökan.
På samma adress ser du också hur behandlingen av din ansökan framskrider.
När ansökan avgjorts, ser du beloppet på ditt stöd och tidpunkten för utbetalningen.
Tjänsten är på finska och svenska.
Du kan ansöka om föräldradagpenningar också genom att fylla i en pappersblankett och skicka den jämte nödvändiga bilagor till vilken FPA-byrå som helst.
Rådgivningen hjälper dig att fylla i ansökan.
Beloppet på din föräldradagpenning beror på hur höga inkomster du har.
Dagpenningen är alltid lägre än lönen, vanligen cirka 70 procent av inkomsterna.
Om du inte har några inkomster, får du föräldradagpenningens minimibelopp.
Också en arbetslös förälder har rätt till föräldradagpenning.
Om din arbetsgivare betalar ut lön till dig under föräldradagpenningperioden, betalar FPA dagpenningen till din arbetsgivare.
Meddela din arbetsgivare om din föräldraledighet två månader innan den börjar.
Om din ledighet varar i 12 vardagar eller mindre, ska du meddela om ledigheten till din arbetsgivare en månad på förhand.
Läs mer på InfoFinlands sida Familjeledighet.
Föräldradagpenningar är skattepliktiga inkomster och följaktligen behöver du ett skattekort (verokortti).
Läs mer på InfoFinlands sida Beskattning.
linkkiSkattemyndigheten:
Skattekortfinska _ svenska _ engelska
Moderskapspenningperioden varar i cirka tre månader.
Den börjar vanligen 30 vardagar för det beräknade förlossningsdatumet.
Läs mer på InfoFinlands sidor Stöd till gravida.
Föräldrapenning
Efter utgången av moderskapspenningperioden kan en av vårdnadshavarna ta ut föräldraledighet.
I så fall sköter en av föräldrarna barnet hemma och får en föräldrapenning.
Ansökan ska lämnas in till FPA senast en månad innan moderskapspenningperiodens utgång och föräldrapenningperiodens början.
Föräldrapenningperioden varar i cirka sex månader.
Om familjen får tvillingar är föräldrapenningperioden 60 vardagar längre.
Modern ska genomgå en läkarundersökning 5–12 veckor efter förlossningen och skicka läkarintyget till FPA.
Annars utbetalas inte föräldradagpenning.
Vilken som helst av vårdnadshavarna kan vara föräldraledig.
De kan också vara lediga turvis.
Föräldrarna kan också arbeta deltid och tillsammans sköta barnet på deltid.
Under denna tid betalar FPA partiell föräldrapenning till bägge föräldrar.
Om en av föräldrarna vill sköta barnet hemma efter föräldrapenningperioden, kan han eller hon få hemvårdsstöd.
Läs mer på InfoFinlands sida Stöd för vård av barn i hemmet.
Föräldrapenning till modern eller fadernfinska _ svenska _ engelska
Faderskapspenning
Faderskapspenningen (Isyysraha) är avsedd för fadern då han tar hand om barnet.
FPA (Kela) betalar ut faderskapspenning under faderskapsledigheten.
Du kan ansöka om faderskapspenning även om du är till exempel företagare, arbetslös eller studerande.
Faderskapspenning betalas ut för 54 vardagar, alltså ungefär nio veckor.
Dessa dagar kan inte överföras till modern.
Du får själv bestämma om du tar ut alla faderskapspenningdagar eller bara en del av dem.
Du får faderskapspenning även om du inte bor tillsammans med barnets mor.
Du kan vara pappaledig samtidigt som barnets mor är mamma- eller föräldraledig.
Då kan du ta ut högst 18 faderskapspenningdagar.
Du kan också ta ut alla 54 faderskapspenningdagar separat, till exempel efter föräldraledigheten.
De 1–18 vardagar av faderskapsledigheten som du kan ta ut samtidigt med barnets mor kan delas upp i högst fyra perioder.
Faderskapsledighet som tas ut efter föräldrapenningperioden kan delas upp i högst två perioder.
Du kan endast använda faderskapspenningdagar för vård av ett barn under två år.
När barnet fyller två år kan du inte längre använda dina faderskapspenningdagar även om sådana finns kvar.
Efter att barnet fötts sköter vanligtvis en av föräldrarna barnet hemma i en viss tid.
Under denna tid betalar FPA ut olika föräldradagpenningar (vanhempainpäiväraha).
Föräldradagpenningarna omfattar
moderskapspenning och särskild moderskapspenning
föräldrapenning
faderskapspenning.
Därtill utbetalas barnbidrag (lapsilisä) till barnets vårdnadshavare fram till dess att barnet fyller 17 år.
Läs mer på InfoFinlands sida Barnbidrag.
Ansökan om föräldradagpenningar
Du kan ansöka om föräldradagpenningar om du omfattas av den sociala tryggheten i Finland och varit sjukförsäkrad i Finland, ett annat EU- eller EES-land eller Schweiz oavbrutet i 180 dagar före det beräknade förslossningsdatumet.
Du kan göra en ansökan om föräldradagpenning på FPA:s webbsidor.
Logga in med nätbankskoder eller ett mobilcertifikat.
Tjänsten innehåller anvisningar för att fylla i ansökan.
På samma adress ser du också hur behandlingen av din ansökan framskrider.
När ansökan avgjorts, ser du beloppet på ditt stöd och tidpunkten för utbetalningen.
Tjänsten är på finska och svenska.
Du kan ansöka om föräldradagpenningar också genom att fylla i en pappersblankett och skicka den jämte nödvändiga bilagor till vilken FPA-byrå som helst.
Rådgivningen hjälper dig att fylla i ansökan.
Beloppet på din föräldradagpenning beror på hur höga inkomster du har.
Dagpenningen är alltid lägre än lönen, vanligen cirka 70 procent av inkomsterna.
Om du inte har några inkomster, får du föräldradagpenningens minimibelopp.
Också en arbetslös förälder har rätt till föräldradagpenning.
Om din arbetsgivare betalar ut lön till dig under föräldradagpenningperioden, betalar FPA dagpenningen till din arbetsgivare.
Meddela din arbetsgivare om din föräldraledighet två månader innan den börjar.
Om din ledighet varar i 12 vardagar eller mindre, ska du meddela om ledigheten till din arbetsgivare en månad på förhand.
Läs mer på InfoFinlands sida Familjeledighet.
Föräldradagpenningar är skattepliktiga inkomster och följaktligen behöver du ett skattekort (verokortti).
Läs mer på InfoFinlands sida Beskattning.
linkkiSkattemyndigheten:
Skattekortfinska _ svenska _ engelska
Moderskapspenningperioden varar i cirka tre månader.
Den börjar vanligen 30 vardagar för det beräknade förlossningsdatumet.
Läs mer på InfoFinlands sidor Stöd till gravida.
Föräldrapenning
Efter utgången av moderskapspenningperioden kan en av vårdnadshavarna ta ut föräldraledighet.
I så fall sköter en av föräldrarna barnet hemma och får en föräldrapenning.
Ansökan ska lämnas in till FPA senast en månad innan moderskapspenningperiodens utgång och föräldrapenningperiodens början.
Föräldrapenningperioden varar i cirka sex månader.
Om familjen får tvillingar är föräldrapenningperioden 60 vardagar längre.
Modern ska genomgå en läkarundersökning 5–12 veckor efter förlossningen och skicka läkarintyget till FPA.
Annars utbetalas inte föräldradagpenning.
Vilken som helst av vårdnadshavarna kan vara föräldraledig.
De kan också vara lediga turvis.
Föräldrarna kan också arbeta deltid och tillsammans sköta barnet på deltid.
Under denna tid betalar FPA partiell föräldrapenning till bägge föräldrar.
Om en av föräldrarna vill sköta barnet hemma efter föräldrapenningperioden, kan han eller hon få hemvårdsstöd.
Läs mer på InfoFinlands sida Stöd för vård av barn i hemmet.
Föräldrapenning till modern eller fadernfinska _ svenska _ engelska
Faderskapspenning
Faderskapspenningen (Isyysraha) är avsedd för fadern då han tar hand om barnet.
FPA (Kela) betalar ut faderskapspenning under faderskapsledigheten.
Du kan ansöka om faderskapspenning även om du är till exempel företagare, arbetslös eller studerande.
Faderskapspenning betalas ut för 54 vardagar, alltså ungefär nio veckor.
Dessa dagar kan inte överföras till modern.
Du får själv bestämma om du tar ut alla faderskapspenningdagar eller bara en del av dem.
Du får faderskapspenning även om du inte bor tillsammans med barnets mor.
Du kan vara pappaledig samtidigt som barnets mor är mamma- eller föräldraledig.
Då kan du ta ut högst 18 faderskapspenningdagar.
Du kan också ta ut alla 54 faderskapspenningdagar separat, till exempel efter föräldraledigheten.
De 1–18 vardagar av faderskapsledigheten som du kan ta ut samtidigt med barnets mor kan delas upp i högst fyra perioder.
Faderskapsledighet som tas ut efter föräldrapenningperioden kan delas upp i högst två perioder.
Du kan endast använda faderskapspenningdagar för vård av ett barn under två år.
När barnet fyller två år kan du inte längre använda dina faderskapspenningdagar även om sådana finns kvar.
Moderskapsförpackning
Om du bor i Finland kan du ha rätt till moderskapsunderstöd (äitiysavustus).
Moderskapsunderstödet är antingen en moderskapsförpackning (äitiyspakkaus) eller ett fast skattefritt belopp, du väljer vilket alternativ du vill ha.
Moderskapsförpackningen innehåller bebiskläder och vårdartiklar.
Största delen av mödrarna väljer moderskapsförpackningen, eftersom dess penningvärde är högre.
Du har rätt till moderskapsunderstöd då
graviditeten varat i cirka fem månader
du genomgått läkarundersökning före utgången av fjärde graviditetsmånaden
du omfattas av den sociala tryggheten i Finland.
Moderskapsförpackningfinska _ svenska _ engelska
Moderskapspenning
När du är gravid kan FPA betala ut moderskapspenning (äitiysraha) till dig.
Modern inleder i allmänhet moderskapsledigheten 30 vardagar för det beräknade förlossningsdatumet.
Du kan ansöka om moderskapspenning om du omfattas av den sociala tryggheten i Finland och varit sjukförsäkrad i Finland, ett annat EU- eller EES-land eller Schweiz oavbrutet i 180 dagar före det beräknade förslossningsdatumet.
FPA betalar ut moderskapspenning på samma villkor också till studeranden och arbetslösa.
Ansökan om moderskapsunderstöd och moderskapspenning
Ansök om moderskapsunderstöd och moderskapspenning hos FPA senast två månader före det beräknade förlossningsdatumet.
Du kan göra en ansökan om moderskapsunderstöd och moderskapspenning via FPA:s webbsidor.
Logga in med nätbankskoder eller ett mobilcertifikat.
Tjänsten innehåller anvisningar för att fylla i ansökan.
På samma adress ser du också hur behandlingen av din ansökan framskrider.
När ansökan avgjorts, ser du beloppet på ditt stöd och tidpunkten för utbetalningen.
Tjänsten är på finska och svenska.
Du kan ansöka om moderskapsunderstöd och moderskapspenning också genom att fylla i en pappersblankett och skicka den jämte nödvändiga bilagor till vilken FPA-byrå som helst.
Rådgivningen hjälper dig att fylla i ansökan.
Föräldradagpenningar är skattepliktiga inkomster och följaktligen behöver du ett skattekort (verokortti).
Läs mer på InfoFinlands sida Beskattning.
Kom ihåg att meddela din arbetsgivare om moderskapsledigheten senast två månader innan den börjar.
Tidigarelagd moderskapspenning
En moder kan bli moderskapsledig redan 31–50 vardagar innan det beräknade förlossningsdatumet.
Moderskapspenning utbetalas under sammanlagt fyra månader från moderskapsledighetens början.
Särskild moderskapspenning
Om du är utsatt för strålning, kemiska ämnen eller smittsamma sjukdomar i ditt arbete kan du sluta arbeta genast då graviditeten konstaterats.
Under denna tid får du särskild moderskapspenning (erityisäitiysraha).
Kom ihåg att ansöka om särskild moderskapspenning hos FPA inom fyra månader från den dag du slutar arbeta.
Särskild moderskapspenning betalas inte alls ut till arbetslösa och endast i vissa fall till studeranden.
Fråga närmare av FPA.
På FPA:s webbsidor kan du ta del av alla förmåner som FPA erbjuder till barnfamiljer.
Information om stöd till barnfamiljerfinska _ svenska _ engelska
Moderskapsförpackning
Om du bor i Finland kan du ha rätt till moderskapsunderstöd (äitiysavustus).
Moderskapsunderstödet är antingen en moderskapsförpackning (äitiyspakkaus) eller ett fast skattefritt belopp, du väljer vilket alternativ du vill ha.
Moderskapsförpackningen innehåller bebiskläder och vårdartiklar.
Största delen av mödrarna väljer moderskapsförpackningen, eftersom dess penningvärde är högre.
Du har rätt till moderskapsunderstöd då
graviditeten varat i cirka fem månader
du genomgått läkarundersökning före utgången av fjärde graviditetsmånaden
du omfattas av den sociala tryggheten i Finland.
Moderskapsförpackningfinska _ svenska _ engelska
Moderskapspenning
När du är gravid kan FPA betala ut moderskapspenning (äitiysraha) till dig.
Modern inleder i allmänhet moderskapsledigheten 30 vardagar för det beräknade förlossningsdatumet.
Du kan ansöka om moderskapspenning om du omfattas av den sociala tryggheten i Finland och varit sjukförsäkrad i Finland, ett annat EU- eller EES-land eller Schweiz oavbrutet i 180 dagar före det beräknade förslossningsdatumet.
FPA betalar ut moderskapspenning på samma villkor också till studeranden och arbetslösa.
Ansökan om moderskapsunderstöd och moderskapspenning
Ansök om moderskapsunderstöd och moderskapspenning hos FPA senast två månader före det beräknade förlossningsdatumet.
Du kan göra en ansökan om moderskapsunderstöd och moderskapspenning via FPA:s webbsidor.
Logga in med nätbankskoder eller ett mobilcertifikat.
Tjänsten innehåller anvisningar för att fylla i ansökan.
På samma adress ser du också hur behandlingen av din ansökan framskrider.
När ansökan avgjorts, ser du beloppet på ditt stöd och tidpunkten för utbetalningen.
Tjänsten är på finska och svenska.
Du kan ansöka om moderskapsunderstöd och moderskapspenning också genom att fylla i en pappersblankett och skicka den jämte nödvändiga bilagor till vilken FPA-byrå som helst.
Rådgivningen hjälper dig att fylla i ansökan.
Föräldradagpenningar är skattepliktiga inkomster och följaktligen behöver du ett skattekort (verokortti).
Läs mer på InfoFinlands sida Beskattning.
Kom ihåg att meddela din arbetsgivare om moderskapsledigheten senast två månader innan den börjar.
Tidigarelagd moderskapspenning
En moder kan bli moderskapsledig redan 31–50 vardagar innan det beräknade förlossningsdatumet.
Moderskapspenning utbetalas under sammanlagt fyra månader från moderskapsledighetens början.
Särskild moderskapspenning
Om du är utsatt för strålning, kemiska ämnen eller smittsamma sjukdomar i ditt arbete kan du sluta arbeta genast då graviditeten konstaterats.
Under denna tid får du särskild moderskapspenning (erityisäitiysraha).
Kom ihåg att ansöka om särskild moderskapspenning hos FPA inom fyra månader från den dag du slutar arbeta.
Särskild moderskapspenning betalas inte alls ut till arbetslösa och endast i vissa fall till studeranden.
Fråga närmare av FPA.
På FPA:s webbsidor kan du ta del av alla förmåner som FPA erbjuder till barnfamiljer.
Information om stöd till barnfamiljerfinska _ svenska _ engelska
Moderskapsförpackning
Om du bor i Finland kan du ha rätt till moderskapsunderstöd (äitiysavustus).
Moderskapsunderstödet är antingen en moderskapsförpackning (äitiyspakkaus) eller ett fast skattefritt belopp, du väljer vilket alternativ du vill ha.
Moderskapsförpackningen innehåller bebiskläder och vårdartiklar.
Största delen av mödrarna väljer moderskapsförpackningen, eftersom dess penningvärde är högre.
Du har rätt till moderskapsunderstöd då
graviditeten varat i cirka fem månader
du genomgått läkarundersökning före utgången av fjärde graviditetsmånaden
du omfattas av den sociala tryggheten i Finland.
Moderskapsförpackningfinska _ svenska _ engelska
Moderskapspenning
När du är gravid kan FPA betala ut moderskapspenning (äitiysraha) till dig.
Modern inleder i allmänhet moderskapsledigheten 30 vardagar för det beräknade förlossningsdatumet.
Du kan ansöka om moderskapspenning om du omfattas av den sociala tryggheten i Finland och varit sjukförsäkrad i Finland, ett annat EU- eller EES-land eller Schweiz oavbrutet i 180 dagar före det beräknade förslossningsdatumet.
FPA betalar ut moderskapspenning på samma villkor också till studeranden och arbetslösa.
Ansökan om moderskapsunderstöd och moderskapspenning
Ansök om moderskapsunderstöd och moderskapspenning hos FPA senast två månader före det beräknade förlossningsdatumet.
Du kan göra en ansökan om moderskapsunderstöd och moderskapspenning via FPA:s webbsidor.
Logga in med nätbankskoder eller ett mobilcertifikat.
Tjänsten innehåller anvisningar för att fylla i ansökan.
På samma adress ser du också hur behandlingen av din ansökan framskrider.
När ansökan avgjorts, ser du beloppet på ditt stöd och tidpunkten för utbetalningen.
Tjänsten är på finska och svenska.
Du kan ansöka om moderskapsunderstöd och moderskapspenning också genom att fylla i en pappersblankett och skicka den jämte nödvändiga bilagor till vilken FPA-byrå som helst.
Rådgivningen hjälper dig att fylla i ansökan.
Föräldradagpenningar är skattepliktiga inkomster och följaktligen behöver du ett skattekort (verokortti).
Läs mer på InfoFinlands sida Beskattning.
Kom ihåg att meddela din arbetsgivare om moderskapsledigheten senast två månader innan den börjar.
Tidigarelagd moderskapspenning
En moder kan bli moderskapsledig redan 31–50 vardagar innan det beräknade förlossningsdatumet.
Moderskapspenning utbetalas under sammanlagt fyra månader från moderskapsledighetens början.
Särskild moderskapspenning
Om du är utsatt för strålning, kemiska ämnen eller smittsamma sjukdomar i ditt arbete kan du sluta arbeta genast då graviditeten konstaterats.
Under denna tid får du särskild moderskapspenning (erityisäitiysraha).
Kom ihåg att ansöka om särskild moderskapspenning hos FPA inom fyra månader från den dag du slutar arbeta.
Särskild moderskapspenning betalas inte alls ut till arbetslösa och endast i vissa fall till studeranden.
Fråga närmare av FPA.
På FPA:s webbsidor kan du ta del av alla förmåner som FPA erbjuder till barnfamiljer.
Information om stöd till barnfamiljerfinska _ svenska _ engelska
På dessa sidor redogörs det för hurdant ekonomiskt stöd barnfamiljer kan få i Finland.
De flesta stöd ansöker man om av Fpa.
Läs mer om Fpa på InfoFinlands sida Viktiga myndigheter.
Vanligen måste du omfattas av Den sociala tryggheten i Finland eller ha en hemkommun i Finland för att du ska kunna få stöd.
Barnets medborgarskap påverkar inte huruvida du får stöd eller ej.
Föräldrarnas uppehållstillstånd kan dock påverka vilka stöd familjen kan få.
Du kan ha rätt att få stöd från ditt eget hemland.
Om du omfattas av Den sociala tryggheten i Finland och bor utomlands kan du få vissa av de Fpa-stöd som du skulle få i Finland.
Till exempel barnbidrag, moderskapsunderstöd och föräldrapenning betalas även till utlandet.
Moderskaps- och föräldrapenning kan betalas till exempel till mödrar som mitt under föräldrapenningsperioden flyttar till ett annat EU/EES-land eller Schweiz för mindre än ett år.
Meddela alltid
Fpa om du flyttar utomlands permanent eller vistas utomlands mer än tre månader.
Se Fpas hemsidor för mer information.
Hem och familjsvenska _ engelska _ ryska _ estniska
Familjeförmåner utomlandsfinska _ svenska _ engelska
På dessa sidor redogörs det för hurdant ekonomiskt stöd barnfamiljer kan få i Finland.
De flesta stöd ansöker man om av Fpa.
Läs mer om Fpa på InfoFinlands sida Viktiga myndigheter.
Vanligen måste du omfattas av Den sociala tryggheten i Finland eller ha en hemkommun i Finland för att du ska kunna få stöd.
Barnets medborgarskap påverkar inte huruvida du får stöd eller ej.
Föräldrarnas uppehållstillstånd kan dock påverka vilka stöd familjen kan få.
Du kan ha rätt att få stöd från ditt eget hemland.
Om du omfattas av Den sociala tryggheten i Finland och bor utomlands kan du få vissa av de Fpa-stöd som du skulle få i Finland.
Till exempel barnbidrag, moderskapsunderstöd och föräldrapenning betalas även till utlandet.
Moderskaps- och föräldrapenning kan betalas till exempel till mödrar som mitt under föräldrapenningsperioden flyttar till ett annat EU/EES-land eller Schweiz för mindre än ett år.
Meddela alltid
Fpa om du flyttar utomlands permanent eller vistas utomlands mer än tre månader.
Se Fpas hemsidor för mer information.
Hem och familjsvenska _ engelska _ ryska _ estniska
Familjeförmåner utomlandsfinska _ svenska _ engelska
På dessa sidor redogörs det för hurdant ekonomiskt stöd barnfamiljer kan få i Finland.
De flesta stöd ansöker man om av Fpa.
Läs mer om Fpa på InfoFinlands sida Viktiga myndigheter.
Vanligen måste du omfattas av Den sociala tryggheten i Finland eller ha en hemkommun i Finland för att du ska kunna få stöd.
Barnets medborgarskap påverkar inte huruvida du får stöd eller ej.
Föräldrarnas uppehållstillstånd kan dock påverka vilka stöd familjen kan få.
Du kan ha rätt att få stöd från ditt eget hemland.
Om du omfattas av Den sociala tryggheten i Finland och bor utomlands kan du få vissa av de Fpa-stöd som du skulle få i Finland.
Till exempel barnbidrag, moderskapsunderstöd och föräldrapenning betalas även till utlandet.
Moderskaps- och föräldrapenning kan betalas till exempel till mödrar som mitt under föräldrapenningsperioden flyttar till ett annat EU/EES-land eller Schweiz för mindre än ett år.
Meddela alltid
Fpa om du flyttar utomlands permanent eller vistas utomlands mer än tre månader.
Se Fpas hemsidor för mer information.
Hem och familjfinska _ svenska _ engelska _ ryska _ estniska
Familjeförmåner utomlandsfinska _ svenska _ engelska
Varje barn har rätt till en god och trygg barndom.
Barnskydd innebär att kommunens socialarbetare hjälper barn och familjer i problematiska situationer.
Man försöker alltid ingripa i problem redan innan de blivit alltför stora.
Barnskydd är alltid det sista alternativet.
Det betyder att barnet och familjen får stöd till exempel i skolan eller rådgivningen innan man kontaktar barnskyddet.
Kontakten med barnskyddet inleds med en barnskyddsanmälan.
Familjen kan själv be barnskyddsmyndigheterna om hjälp.
Vem som helst som oroar sig för familjens välbefinnande kan göra en barnskyddsanmälan.
Till exempel kan barnets lärare kontakta barnskyddsmyndigheterna.
Ibland kan föräldrarna inte sörja för barnets välfärd.
Då måste samhället ingripa i familjens situation.
Inom barnskyddet är barnets bästa den högsta prioriteten.
Barnskyddet stöder familjer i problematiska situationer
Man kan själv be om hjälp hos barnskyddet om föräldrarna är utmattade eller familjen genomgår en svår förändring i livet.
Barnskyddet stöder familjen även då ett barn eller en ung till exempel använder mycket rusmedel eller begår brott.
Barnskyddet har många slags medel som de kan använda för att hjälpa familjen.
I första hand försöker man använda öppenvården alltså att barnet bor tillsammans med sin familj.
Socialarbetaren kan ordna familjen till exempel hemhjälp eller en stödperson.
Om det förekommer våld eller missbruk i familjen ingriper barnskyddets socialarbetare i situationen.
Om barnet inte är tryggt i sitt hem eller om situationen med barnet är mycket svårt, kan det fattas ett beslut om vård utom hemmet eller omhändertagande.
Man försöker emellertid alltid först hjälpa barnet så att det kan bo kvar hemma.
Barnskyddet är baserat på lag
Barnskyddet är baserat på barnskyddslagen och internationella konventioner.
Barnskyddslagen gäller alla barn som bor i Finland oavsett deras nationalitet, religion eller kultur.
Information om barnskyddfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
Barnskyddslagenfinska _ svenska _ engelska
Varje barn har rätt till en god och trygg barndom.
Barnskydd innebär att kommunens socialarbetare hjälper barn och familjer i problematiska situationer.
Man försöker alltid ingripa i problem redan innan de blivit alltför stora.
Barnskydd är alltid det sista alternativet.
Det betyder att barnet och familjen får stöd till exempel i skolan eller rådgivningen innan man kontaktar barnskyddet.
Kontakten med barnskyddet inleds med en barnskyddsanmälan.
Familjen kan själv be barnskyddsmyndigheterna om hjälp.
Vem som helst som oroar sig för familjens välbefinnande kan göra en barnskyddsanmälan.
Till exempel kan barnets lärare kontakta barnskyddsmyndigheterna.
Ibland kan föräldrarna inte sörja för barnets välfärd.
Då måste samhället ingripa i familjens situation.
Inom barnskyddet är barnets bästa den högsta prioriteten.
Barnskyddet stöder familjer i problematiska situationer
Man kan själv be om hjälp hos barnskyddet om föräldrarna är utmattade eller familjen genomgår en svår förändring i livet.
Barnskyddet stöder familjen även då ett barn eller en ung till exempel använder mycket rusmedel eller begår brott.
Barnskyddet har många slags medel som de kan använda för att hjälpa familjen.
I första hand försöker man använda öppenvården alltså att barnet bor tillsammans med sin familj.
Socialarbetaren kan ordna familjen till exempel hemhjälp eller en stödperson.
Om det förekommer våld eller missbruk i familjen ingriper barnskyddets socialarbetare i situationen.
Om barnet inte är tryggt i sitt hem eller om situationen med barnet är mycket svårt, kan det fattas ett beslut om vård utom hemmet eller omhändertagande.
Man försöker emellertid alltid först hjälpa barnet så att det kan bo kvar hemma.
Barnskyddet är baserat på lag
Barnskyddet är baserat på barnskyddslagen och internationella konventioner.
Barnskyddslagen gäller alla barn som bor i Finland oavsett deras nationalitet, religion eller kultur.
Information om barnskyddfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
Barnskyddslagenfinska _ svenska _ engelska
Varje barn har rätt till en god och trygg barndom.
Barnskydd innebär att kommunens socialarbetare hjälper barn och familjer i problematiska situationer.
Man försöker alltid ingripa i problem redan innan de blivit alltför stora.
Barnskydd är alltid det sista alternativet.
Det betyder att barnet och familjen får stöd till exempel i skolan eller rådgivningen innan man kontaktar barnskyddet.
Kontakten med barnskyddet inleds med en barnskyddsanmälan.
Familjen kan själv be barnskyddsmyndigheterna om hjälp.
Vem som helst som oroar sig för familjens välbefinnande kan göra en barnskyddsanmälan.
Till exempel kan barnets lärare kontakta barnskyddsmyndigheterna.
Ibland kan föräldrarna inte sörja för barnets välfärd.
Då måste samhället ingripa i familjens situation.
Inom barnskyddet är barnets bästa den högsta prioriteten.
Barnskyddet stöder familjer i problematiska situationer
Man kan själv be om hjälp hos barnskyddet om föräldrarna är utmattade eller familjen genomgår en svår förändring i livet.
Barnskyddet stöder familjen även då ett barn eller en ung till exempel använder mycket rusmedel eller begår brott.
Barnskyddet har många slags medel som de kan använda för att hjälpa familjen.
I första hand försöker man använda öppenvården alltså att barnet bor tillsammans med sin familj.
Socialarbetaren kan ordna familjen till exempel hemhjälp eller en stödperson.
Om det förekommer våld eller missbruk i familjen ingriper barnskyddets socialarbetare i situationen.
Om barnet inte är tryggt i sitt hem eller om situationen med barnet är mycket svårt, kan det fattas ett beslut om vård utom hemmet eller omhändertagande.
Man försöker emellertid alltid först hjälpa barnet så att det kan bo kvar hemma.
Barnskyddet är baserat på lag
Barnskyddet är baserat på barnskyddslagen och internationella konventioner.
Barnskyddslagen gäller alla barn som bor i Finland oavsett deras nationalitet, religion eller kultur.
linkkiSocial- och hälsovårdsministeriet:
Barnskyddfinska _ svenska _ engelska _ ryska
Information om barnskyddfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
Barnskyddslagenfinska _ svenska _ engelska
Samhället tryggar barnets rättigheter med hjälp av lagar och författningar.
Enligt lagen har barnets föräldrar eller vårdnadshavare huvudansvaret för barnets välfärd och harmoniska utveckling.
I Finland är kroppsaga på barn (våld i syfte att straffa) förbjuden i lag.
Barn får till exempel inte slås eller luggas.
I Finland framhävs jämställdhet.
Till exempel kan mamman till ett litet barn förvärvsarbeta medan den andra föräldern stannar hemma för att ta hand om barnet.
I Finland sköter och uppfostrar både män och kvinnor barnen.
Barnet uppmuntras till självständigt tänkande.
Barnet får till exempel ha andra åsikter än föräldrarna.
I Finland flyttar ungdomar oftast hemifrån när de är myndiga och börjar studera eller arbeta.
Det är vanligt att de bor antingen ensamma eller med studiekamrater innan de grundar sin egen familj.
Utbildning skattas högt i Finland och det är viktigt att föräldrarna uppmuntrar skolgången.
Visa intresse för barnets skolgång och delta till exempel i föräldramöten som skolan ordnar.
Det är viktigt att sätta upp tydliga gränser och regler för barn och unga.
Man kan till exempel komma överens om gemensamma regler med andra föräldrar.
Det är viktigt att komma ihåg att man inte får ge tobak eller alkohol till barn under 18 år.
När en person fyller 18 år är han eller hon enligt lagen myndig.
Då är den unga en myndig samhällsmedlem som har rätt att besluta om sitt eget liv.
Också barn under 18 har rätt att fatta beslut i vissa ärenden.
Mer information om barnets rättigheter i olika åldrar finns på InfoFinlands sida Barns och ungdomars rättigheter och skyldigheter.
Det finns mycket hjälp och stöd att få när det gäller uppfostring av barn.
Om du behöver stöd eller är orolig för barnet är det bäst att i god tid be om råd till exempel vid den egna kommunens socialtjänst.
Läs mer på InfoFinlands sida Barns och ungas problem.
Uppfostring av barn i Finland(pdf, 8,08 Mt)finska _ engelska _ ryska _ somaliska _ kurdiska _ albanska _ burmesiska
linkkiUnicef:
Konvention om barnets rättigheterfinska _ engelska _ franska _ spanska _ kinesiska
linkkiBarnombudsmannen:
Broschyren Barnets rättigheterfinska _ svenska _ engelska _ ryska
linkkiSocial- och hälsovårdsministeriet:
Lagstiftning som rör barn, unga och familjerfinska _ svenska _ engelska
Samhället tryggar barnets rättigheter med hjälp av lagar och författningar.
Enligt lagen har barnets föräldrar eller vårdnadshavare huvudansvaret för barnets välfärd och harmoniska utveckling.
I Finland är kroppsaga på barn (våld i syfte att straffa) förbjuden i lag.
Barn får till exempel inte slås eller luggas.
I Finland framhävs jämställdhet.
Till exempel kan mamman till ett litet barn förvärvsarbeta medan den andra föräldern stannar hemma för att ta hand om barnet.
I Finland sköter och uppfostrar både män och kvinnor barnen.
Barnet uppmuntras till självständigt tänkande.
Barnet får till exempel ha andra åsikter än föräldrarna.
I Finland flyttar ungdomar oftast hemifrån när de är myndiga och börjar studera eller arbeta.
Det är vanligt att de bor antingen ensamma eller med studiekamrater innan de grundar sin egen familj.
Utbildning skattas högt i Finland och det är viktigt att föräldrarna uppmuntrar skolgången.
Visa intresse för barnets skolgång och delta till exempel i föräldramöten som skolan ordnar.
Det är viktigt att sätta upp tydliga gränser och regler för barn och unga.
Man kan till exempel komma överens om gemensamma regler med andra föräldrar.
Det är viktigt att komma ihåg att man inte får ge tobak eller alkohol till barn under 18 år.
När en person fyller 18 år är han eller hon enligt lagen myndig.
Då är den unga en myndig samhällsmedlem som har rätt att besluta om sitt eget liv.
Också barn under 18 har rätt att fatta beslut i vissa ärenden.
Mer information om barnets rättigheter i olika åldrar finns på InfoFinlands sida Barns och ungdomars rättigheter och skyldigheter.
Det finns mycket hjälp och stöd att få när det gäller uppfostring av barn.
Om du behöver stöd eller är orolig för barnet är det bäst att i god tid be om råd till exempel vid den egna kommunens socialtjänst.
Läs mer på InfoFinlands sida Barns och ungas problem.
Uppfostring av barn i Finland(pdf, 8,08 Mt)finska _ engelska _ ryska _ somaliska _ kurdiska _ albanska _ burmesiska
linkkiUnicef:
Konvention om barnets rättigheterfinska _ engelska _ franska _ spanska _ kinesiska
linkkiBarnombudsmannen:
Broschyren Barnets rättigheterfinska _ svenska _ engelska _ ryska
linkkiSocial- och hälsovårdsministeriet:
Lagstiftning som rör barn, unga och familjerfinska _ svenska _ engelska
Samhället tryggar barnets rättigheter med hjälp av lagar och författningar.
Enligt lagen har barnets föräldrar eller vårdnadshavare huvudansvaret för barnets välfärd och harmoniska utveckling.
I Finland är kroppsaga på barn (våld i syfte att straffa) förbjuden i lag.
Barn får till exempel inte slås eller luggas.
I Finland framhävs jämställdhet.
Till exempel kan mamman till ett litet barn förvärvsarbeta medan den andra föräldern stannar hemma för att ta hand om barnet.
I Finland sköter och uppfostrar både män och kvinnor barnen.
Barnet uppmuntras till självständigt tänkande.
Barnet får till exempel ha andra åsikter än föräldrarna.
I Finland flyttar ungdomar oftast hemifrån när de är myndiga och börjar studera eller arbeta.
Det är vanligt att de bor antingen ensamma eller med studiekamrater innan de grundar sin egen familj.
Utbildning skattas högt i Finland och det är viktigt att föräldrarna uppmuntrar skolgången.
Visa intresse för barnets skolgång och delta till exempel i föräldramöten som skolan ordnar.
Det är viktigt att sätta upp tydliga gränser och regler för barn och unga.
Man kan till exempel komma överens om gemensamma regler med andra föräldrar.
Det är viktigt att komma ihåg att man inte får ge tobak eller alkohol till barn under 18 år.
När en person fyller 18 år är han eller hon enligt lagen myndig.
Då är den unga en myndig samhällsmedlem som har rätt att besluta om sitt eget liv.
Också barn under 18 har rätt att fatta beslut i vissa ärenden.
Mer information om barnets rättigheter i olika åldrar finns på InfoFinlands sida Barns och ungdomars rättigheter och skyldigheter.
Det finns mycket hjälp och stöd att få när det gäller uppfostring av barn.
Om du behöver stöd eller är orolig för barnet är det bäst att i god tid be om råd till exempel vid den egna kommunens socialtjänst.
Läs mer på InfoFinlands sida Barns och ungas problem.
Uppfostring av barn i Finland(pdf, 8,08 Mt)finska _ engelska _ ryska _ somaliska _ kurdiska _ albanska _ burmesiska
linkkiUnicef:
Konvention om barnets rättigheterfinska _ engelska _ franska _ spanska _ kinesiska
linkkiBarnombudsmannen:
Broschyren Barnets rättigheterfinska _ svenska _ engelska _ ryska
linkkiSocial- och hälsovårdsministeriet:
Lagstiftning som rör barn, unga och familjerfinska _ svenska _ engelska
6 år
Rättighet och skyldighet:
Barnet måste delta i förskoleundervisningen.
Barnet kan få dispens för att börja i skolan.
7 år
Rättighet och skyldighet:
Skolan börjar (läroplikt).
I särskilda fall kan barnet börja skolan senare.
12 år
Rättighet:
Barnets för- eller efternamn kan inte bytas utan barnets tillstånd.
Barnet kan inte anslutas till ett trossamfund utan barnets tillstånd.
Barnets tillstånd behövs också för utträde ur ett trossamfund.
Barn, vars föräldrar har skilt sig, har rätt att vägra träffa någon av föräldrarna.
Barnet kan inte adopteras utan barnets medgivande.
Om det finns problem i familjen kan barnet själv be om vård utom hemmet.
Vård utom hemmet betyder att barnet bor någon annanstans än hos sina föräldrar.
Skyldighet:
Barn får inte l ängre cykla på trottoaren.
14 år
Rättighet:
Barnet får utföra lätt arbete några timmar om dagen om det inte skadar hennes hälsa eller skolgång.
Vårdnadshavaren måste underteckna arbetsavtalet.
15 år
Rättighet
Den unga kan själv ingå ett arbetsavtal.
Föräldrarna kan dock häva ett avtal som ingåtts av ett barn under 18 år om barnet inte har berättat för föräldrarna om arbetet.
Den unga har rätt att öppna ett eget bankkonto och förvalta de medel som han eller hon förtjänat med sitt eget arbete.
När den unga har fullgjort sin läroplikt får han eller hon arbeta heltid mellan klockan 6.00 och 22.00.
Den unga kan avlägga körtillstånd som behövs för att köra moped, traktor och motorbåt.
Den unga kan ansluta sig till ett trossamfund eller utträda ur ett trossamfund med föräldrarnas skriftliga tillstånd
Skyldighet
Den unga kan ställas till svars för brott som han eller hon begått.
Om den unga begår ett brott kan han eller hon åtalas och dömas för det.
16 år
Den sexuella skyddsåldersgränsen för barn är 16 år.
Detta betyder att sexuellt umgänge med barn under 16 år är straffbart. (Undantag från detta är en sexuell förbindelse mellan två ungdomar som befinner sig på samma utvecklingsstadium.)
Att köpa sexuella tjänster av ett barn under 18 år är ett brott.
Rättighet
Rätt att avlägga A-körkortet som behövs för att köra lätt motorcykel.
Rätt att få eget sjukförsäkringskort.
Detta betyder att en 16-åring är försäkrad mot ålderdom, arbetslöshet och arbetsoförmåga och att sjukförsäkringsersättningen betalas till den unga själv, inte dennes föräldrar.
17 år
Rättighet
Läroplikten upphör om den inte redan har fullgjorts.
Rätten till barnbidrag upphör.
Den unga kan ansöka om studiestöd hos Fpa.
Vårdnadshavarens inkomster påverkar dock studiestödets storlek och beviljande.
18 år
Myndighet
Rättighet
rösta i nationella val och kommunalval
skaffa sig ett eget pass
inträda i eller utträda ur ett trossamfund
disponera över sin egendom
skaffa sig ett körkort (till exempel för motorcykel, personbil)
få finskt medborgarskap (18–22-åringar), om personen bott länge i Finland.
Skyldighet
värnplikt för män (armé eller civiltjänstgöring)
Läs mer om myndiga medborgares rättigheter och skyldigheter på InfoFinlands sida Dina rättigheter och skyldigheter i Finland.
linkkiBarnombudsmannen:
Broschyren Barnets rättigheterfinska _ svenska _ engelska _ ryska
6 år
Rättighet och skyldighet:
Barnet måste delta i förskoleundervisningen.
Barnet kan få dispens för att börja i skolan.
7 år
Rättighet och skyldighet:
Skolan börjar (läroplikt).
I särskilda fall kan barnet börja skolan senare.
12 år
Rättighet:
Barnets för- eller efternamn kan inte bytas utan barnets tillstånd.
Barnet kan inte anslutas till ett trossamfund utan barnets tillstånd.
Barnets tillstånd behövs också för utträde ur ett trossamfund.
Barn, vars föräldrar har skilt sig, har rätt att vägra träffa någon av föräldrarna.
Barnet kan inte adopteras utan barnets medgivande.
Om det finns problem i familjen kan barnet själv be om vård utom hemmet.
Vård utom hemmet betyder att barnet bor någon annanstans än hos sina föräldrar.
Skyldighet:
Barn får inte l ängre cykla på trottoaren.
14 år
Rättighet:
Barnet får utföra lätt arbete några timmar om dagen om det inte skadar hennes hälsa eller skolgång.
Vårdnadshavaren måste underteckna arbetsavtalet.
15 år
Rättighet
Den unga kan själv ingå ett arbetsavtal.
Föräldrarna kan dock häva ett avtal som ingåtts av ett barn under 18 år om barnet inte har berättat för föräldrarna om arbetet.
Den unga har rätt att öppna ett eget bankkonto och förvalta de medel som han eller hon förtjänat med sitt eget arbete.
När den unga har fullgjort sin läroplikt får han eller hon arbeta heltid mellan klockan 6.00 och 22.00.
Den unga kan avlägga körtillstånd som behövs för att köra moped, traktor och motorbåt.
Den unga kan ansluta sig till ett trossamfund eller utträda ur ett trossamfund med föräldrarnas skriftliga tillstånd
Skyldighet
Den unga kan ställas till svars för brott som han eller hon begått.
Om den unga begår ett brott kan han eller hon åtalas och dömas för det.
16 år
Den sexuella skyddsåldersgränsen för barn är 16 år.
Detta betyder att sexuellt umgänge med barn under 16 år är straffbart. (Undantag från detta är en sexuell förbindelse mellan två ungdomar som befinner sig på samma utvecklingsstadium.)
Att köpa sexuella tjänster av ett barn under 18 år är ett brott.
Rättighet
Rätt att avlägga A-körkortet som behövs för att köra lätt motorcykel.
Rätt att få eget sjukförsäkringskort.
Detta betyder att en 16-åring är försäkrad mot ålderdom, arbetslöshet och arbetsoförmåga och att sjukförsäkringsersättningen betalas till den unga själv, inte dennes föräldrar.
17 år
Rättighet
Läroplikten upphör om den inte redan har fullgjorts.
Rätten till barnbidrag upphör.
Den unga kan ansöka om studiestöd hos Fpa.
Vårdnadshavarens inkomster påverkar dock studiestödets storlek och beviljande.
18 år
Myndighet
Rättighet
rösta i nationella val och kommunalval
skaffa sig ett eget pass
inträda i eller utträda ur ett trossamfund
disponera över sin egendom
skaffa sig ett körkort (till exempel för motorcykel, personbil)
få finskt medborgarskap (18–22-åringar), om personen bott länge i Finland.
Skyldighet
värnplikt för män (armé eller civiltjänstgöring)
Läs mer om myndiga medborgares rättigheter och skyldigheter på InfoFinlands sida Dina rättigheter och skyldigheter i Finland.
linkkiBarnombudsmannen:
Broschyren Barnets rättigheterfinska _ svenska _ engelska _ ryska
6 år
Rättighet och skyldighet:
Barnet måste delta i förskoleundervisningen.
Barnet kan få dispens för att börja i skolan.
7 år
Rättighet och skyldighet:
Skolan börjar (läroplikt).
I särskilda fall kan barnet börja skolan senare.
12 år
Rättighet:
Barnets för- eller efternamn kan inte bytas utan barnets tillstånd.
Barnet kan inte anslutas till ett trossamfund utan barnets tillstånd.
Barnets tillstånd behövs också för utträde ur ett trossamfund.
Barn, vars föräldrar har skilt sig, har rätt att vägra träffa någon av föräldrarna.
Barnet kan inte adopteras utan barnets medgivande.
Om det finns problem i familjen kan barnet själv be om vård utom hemmet.
Vård utom hemmet betyder att barnet bor någon annanstans än hos sina föräldrar.
Skyldighet:
Barn får inte l ängre cykla på trottoaren.
14 år
Rättighet:
Barnet får utföra lätt arbete några timmar om dagen om det inte skadar hennes hälsa eller skolgång.
Vårdnadshavaren måste underteckna arbetsavtalet.
15 år
Rättighet
Den unga kan själv ingå ett arbetsavtal.
Föräldrarna kan dock häva ett avtal som ingåtts av ett barn under 18 år om barnet inte har berättat för föräldrarna om arbetet.
Den unga har rätt att öppna ett eget bankkonto och förvalta de medel som han eller hon förtjänat med sitt eget arbete.
När den unga har fullgjort sin läroplikt får han eller hon arbeta heltid mellan klockan 6.00 och 22.00.
Den unga kan avlägga körtillstånd som behövs för att köra moped, traktor och motorbåt.
Den unga kan ansluta sig till ett trossamfund eller utträda ur ett trossamfund med föräldrarnas skriftliga tillstånd
Skyldighet
Den unga kan ställas till svars för brott som han eller hon begått.
Om den unga begår ett brott kan han eller hon åtalas och dömas för det.
16 år
Den sexuella skyddsåldersgränsen för barn är 16 år.
Detta betyder att sexuellt umgänge med barn under 16 år är straffbart. (Undantag från detta är en sexuell förbindelse mellan två ungdomar som befinner sig på samma utvecklingsstadium.)
Att köpa sexuella tjänster av ett barn under 18 år är ett brott.
Rättighet
Rätt att avlägga A-körkortet som behövs för att köra lätt motorcykel.
Rätt att få eget sjukförsäkringskort.
Detta betyder att en 16-åring är försäkrad mot ålderdom, arbetslöshet och arbetsoförmåga och att sjukförsäkringsersättningen betalas till den unga själv, inte dennes föräldrar.
17 år
Rättighet
Läroplikten upphör om den inte redan har fullgjorts.
Rätten till barnbidrag upphör.
Den unga kan ansöka om studiestöd hos Fpa.
Vårdnadshavarens inkomster påverkar dock studiestödets storlek och beviljande.
18 år
Myndighet
Rättighet
rösta i nationella val och kommunalval
skaffa sig ett eget pass
inträda i eller utträda ur ett trossamfund
disponera över sin egendom
skaffa sig ett körkort (till exempel för motorcykel, personbil)
få finskt medborgarskap (18–22-åringar), om personen bott länge i Finland.
Skyldighet
värnplikt för män (armé eller civiltjänstgöring)
Läs mer om myndiga medborgares rättigheter och skyldigheter på InfoFinlands sida Dina rättigheter och skyldigheter i Finland.
linkkiBarnombudsmannen:
Broschyren Barnets rättigheterfinska _ svenska _ engelska _ ryska
Barnets födelse registreras på sjukhuset
Vilket medborgarskap får barnet?
Om barnet inte får finskt medborgarskap
Barnets sociala trygghet
Erkännande av faderskap
Barnet måste ha en vårdnadshavare
Barnets födelse registreras på sjukhuset
När ett barn har fötts registrerar sjukhuset födelsen i Finlands befolkningsdatasystem, och barnet får en tillfällig personbeteckning.
Detta görs om
barnets mor har uppehållsrätt i Finland,
modern har en hemkommun i Finland och
modern har en finsk personbeteckning.
Om barnets mor inte är registrerad i Finland kan sjukhuset inte registrera födelsen och magistraten skickar ingen blankett till modern.
I detta fall ska du kontakta magistraten och be om anvisningar om hur barnet registreras.
Du kan läsa mer om registreringen av modern på InfoFinlands sida Registrering som invånare.
Kontaktuppgifter till magistratfinska _ svenska _ engelska
Inom två veckor efter att barnets födelse registrerats skickar magistraten en blankett hem till modern.
Med den här blanketten kan du meddela följande information till myndigheterna:
modersmål
religion.
Fyll i blanketten noggrant och underteckna den.
Om föräldrarna är gifta ska båda föräldrarna underteckna blanketten.
Returnera blanketten till magistraten inom två månader efter att barnet fötts.
Du kan skicka blanketten per post eller lämna den personligen till magistraten i ditt område.
Först efter detta registreras ditt barn i befolkningsdatasystemet.
I Finland finns en namnlag. Enligt den ska alla som har en hemort i Finland ha ett efternamn och 1–4 förnamn.
Förnamnen ska vara förenliga med Finlands namnlag.
Till exempel får syskon inte ha samma namn som första namn.
Barnet får efternamn av sina föräldrar.
Om föräldrarna har samma efternamn, blir detta även barnets efternamn.
Om föräldrarna har olika efternamn beror barnets efternamn på situationen.
Om föräldrarna är gifta kan de välja endera makens efternamn till barnet.
Om föräldrarna inte är gifta kan barnet få antingen moderns eller faderns efternamn, om faderskapet har fastställts.
Läs mer om fastställande av faderskap vid punkten Erkännande av faderskap på den här sidan.
Om föräldrarna har ett kombinerat efternamn, blir detta även barnets efternamn.
Om föräldrarna har gemensamma barn sedan tidigare, ska minderåriga syskon ha samma efternamn.
Om föräldrarna har separerat, bestämmer barnets vårdnadshavare vilket namn barnet får.
Om föräldrarna inte kommer överens om barnets efternamn, får barnet moderns efternamn.
Broschyren Makens efternamn och barnets efternamnfinska _ svenska _ engelska
Namnlagenfinska _ svenska
Barnets modersmål
När barnet föds måste man registrera dess modersmål.
Det är obligatoriskt att registrera språket.
Ditt barn kan endast ha ett språk som modersmål.
Du kan ändra språket senare om du vill.
Det är bra att fundera på vilket språk du vill registrera för ditt barn.
Språkvalet kan påverka barnets möjligheter att studera olika språk i skolan.
Barn, vars modersmål inte är finska eller svenska, studerar finska eller svenska som andraspråk i den så kallade S2-undervisningen.
Barnet kan även läsa sitt eget modersmål om man har registrerat något annat språk än finska eller svenska som modersmål för barnet.
Att delta i modersmålsundervisningen är frivilligt.
linkkiUtbildningsstyrelsen:
Eget språk, eget sinnefinska _ engelska _ ryska _ estniska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ burmesiska _ bosniska
Barnets religion
Barnets religion är familjens ensak.
Du får själv bestämma vilket trossamfund ditt barn ska höra till.
Det är inte obligatoriskt att ange barnets religion.
Om den ena föräldern har ensam vårdnad om barnet, kan den föräldern ensam bestämma vilket trossamfund barnet ska höra till.
linkkiUndervisnings- och kulturministeriet:
Religionsfrihetfinska _ svenska _ engelska
linkkiFritänkarförbundet r.f.:
Religionsfriheten för barn och ungafinska
Vilket medborgarskap får barnet?
Barnets medborgarskap beror på föräldrarnas medborgarskap.
När ett barn föds, får barnet finskt medborgarskap om
barnets mor är finsk medborgare,
barnets far är finsk medborgare och föräldrarna är gifta,
barnets far är finsk medborgare, barnet föds utom äktenskap i Finland och faderskapet fastställs,
barnets far avled innan barnet föddes, men fadern var finsk medborgare och gift med barnets mor medan han levde eller
barnets far avled innan barnet föddes, barnet föds utom äktenskap i Finland och faderskapet fastställs.
Ett barn får finskt medborgarskap också om hen föds i Finland och inte får medborgarskap i något annan land av sina föräldrar.
I detta fall fastställer Migrationsverket barnets medborgarskap.
Ett barn kan samtidigt ha både finskt medborgarskap och medborgarskap i ett annat land, om det andra landet godkänner flerfaldigt medborgarskap.
Fråga mer om detta vid ditt eget lands beskickning.
Läs mer om finskt medborgarskap på InfoFinlands sida Finskt medborgarskap.
Finskt medborgarskap till barn med finsk farfinska _ svenska _ engelska
Att ansöka om finskt medborgarskapfinska _ svenska _ engelska
Om barnet inte får finskt medborgarskap
Om ditt barn inte får finskt medborgarskap vid födelsen ska du ansöka om ett pass för barnet vid ditt hemlands beskickning.
För detta behöver du barnets födelseattest från magistraten.
På InfoFinlands sida Ambassader i Finland hittar du information om andra länders beskickningar i Finland.
Därefter måste du ansöka om uppehållstillstånd eller registrering av EU-medborgares uppehållsrätt för barnet.
Om barnet får medborgarskap i ett EU-land, ska du ansöka om registrering av EU-medborgares uppehållsrätt för barnet i Migrationsverkets e-tjänst Enter Finland eller vid Migrationsverkets serviceställe.
Om barnet får medborgarskap i ett annat land, ska du ansöka om uppehållstillstånd för barnet i Migrationsverkets e-tjänst Enter Finland eller vid Migrationsverkets serviceställe.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Barnets sociala trygghet
Om barnet omfattas av Den sociala tryggheten i Finland får hen ett FPA-kort, det vill säga ett sjukförsäkringskort.
FPA skickar kortet hem efter att barnet har fått en personbeteckning och ett namn.
Du måste ansöka om familjeförmåner separat från FPA.
Läs mer om ämnet på InfoFinlands sidor Stöd till gravida och Stöd efter barnets födelse.
Erkännande av faderskap
Om barnets föräldrar är gifta behöver faderskapet inte erkännas separat.
Om barnets mor och far inte är gifta och faderskapet inte erkänns, är barnet officiellt faderlöst.
Faderskapet kan erkänns redan under graviditeten vid mödrarådgivningsbyrån eller efter barnets födelse hos barnatillsyningsmannen i den egna kommunen.
Om faderskapet erkänts före födelsen inleds behandlingen av faderskapsärendet först 30 dagar efter barnets födelse.
Magistraten bekräftar erkännandet av faderskapet.
Läs mer på InfoFinlands sida Samboförhållande.
linkkiSocial- och hälsovårdsministeriet:
Erkännande och fastställande av partnerskapfinska _ svenska
Barnet måste ha en vårdnadshavare
Enligt finländsk lag är en person som är under 18 år ett barn.
Personer under 18 år ska ha minst en vårdnadshavare.
Vanligtvis är barnets föräldrar dess vårdnadshavare.
Om ett barn föds inom äktenskap är båda föräldrarna tillsammans barnets vårdnadshavare.
Om föräldrarna inte är gifta och faderskapet inte har erkänts, är modern barnets vårdnadshavare och bestämmer ensam om alla barnets angelägenheter.
Detta innebär att modern ensam bestämmer om barnets angelägenheter även om föräldrarna bor tillsammans.
Fadern får vårdnad om barnet om föräldrarna ingår ett avtal om gemensam vårdnad och faderskapet har erkänts.
Vårdnadsavtalet ingås antingen på rådgivningsbyrån före barnets födelse eller hos barnatillsyningsmannen efter barnets födelse.
Barnets födelse registreras på sjukhuset
Vilket medborgarskap får barnet?
Om barnet inte får finskt medborgarskap
Barnets sociala trygghet
Erkännande av faderskap
Barnet måste ha en vårdnadshavare
Barnets födelse registreras på sjukhuset
När ett barn har fötts registrerar sjukhuset födelsen i Finlands befolkningsdatasystem, och barnet får en tillfällig personbeteckning.
Detta görs om
barnets mor har uppehållsrätt i Finland,
modern har en hemkommun i Finland och
modern har en finsk personbeteckning.
Om barnets mor inte är registrerad i Finland kan sjukhuset inte registrera födelsen och magistraten skickar ingen blankett till modern.
I detta fall ska du kontakta magistraten och be om anvisningar om hur barnet registreras.
Du kan läsa mer om registreringen av modern på InfoFinlands sida Registrering som invånare.
Kontaktuppgifter till magistratfinska _ svenska _ engelska
Inom två veckor efter att barnets födelse registrerats skickar magistraten en blankett hem till modern.
Med den här blanketten kan du meddela följande information till myndigheterna:
modersmål
religion.
Fyll i blanketten noggrant och underteckna den.
Om föräldrarna är gifta ska båda föräldrarna underteckna blanketten.
Returnera blanketten till magistraten inom två månader efter att barnet fötts.
Du kan skicka blanketten per post eller lämna den personligen till magistraten i ditt område.
Först efter detta registreras ditt barn i befolkningsdatasystemet.
I Finland finns en namnlag. Enligt den ska alla som har en hemort i Finland ha ett efternamn och 1–4 förnamn.
Förnamnen ska vara förenliga med Finlands namnlag.
Till exempel får syskon inte ha samma namn som första namn.
Barnet får efternamn av sina föräldrar.
Om föräldrarna har samma efternamn, blir detta även barnets efternamn.
Om föräldrarna har olika efternamn beror barnets efternamn på situationen.
Om föräldrarna är gifta kan de välja endera makens efternamn till barnet.
Om föräldrarna inte är gifta kan barnet få antingen moderns eller faderns efternamn, om faderskapet har fastställts.
Läs mer om fastställande av faderskap vid punkten Erkännande av faderskap på den här sidan.
Om föräldrarna har ett kombinerat efternamn, blir detta även barnets efternamn.
Om föräldrarna har gemensamma barn sedan tidigare, ska minderåriga syskon ha samma efternamn.
Om föräldrarna har separerat, bestämmer barnets vårdnadshavare vilket namn barnet får.
Om föräldrarna inte kommer överens om barnets efternamn, får barnet moderns efternamn.
Broschyren Makens efternamn och barnets efternamnfinska _ svenska _ engelska
Namnlagenfinska _ svenska
Barnets modersmål
När barnet föds måste man registrera dess modersmål.
Det är obligatoriskt att registrera språket.
Ditt barn kan endast ha ett språk som modersmål.
Du kan ändra språket senare om du vill.
Det är bra att fundera på vilket språk du vill registrera för ditt barn.
Språkvalet kan påverka barnets möjligheter att studera olika språk i skolan.
Barn, vars modersmål inte är finska eller svenska, studerar finska eller svenska som andraspråk i den så kallade S2-undervisningen.
Barnet kan även läsa sitt eget modersmål om man har registrerat något annat språk än finska eller svenska som modersmål för barnet.
Att delta i modersmålsundervisningen är frivilligt.
linkkiUtbildningsstyrelsen:
Eget språk, eget sinnefinska _ engelska _ ryska _ estniska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ burmesiska _ bosniska
Barnets religion
Barnets religion är familjens ensak.
Du får själv bestämma vilket trossamfund ditt barn ska höra till.
Det är inte obligatoriskt att ange barnets religion.
Om den ena föräldern har ensam vårdnad om barnet, kan den föräldern ensam bestämma vilket trossamfund barnet ska höra till.
linkkiUndervisnings- och kulturministeriet:
Religionsfrihetfinska _ svenska _ engelska
linkkiFritänkarförbundet r.f.:
Religionsfriheten för barn och ungafinska
Vilket medborgarskap får barnet?
Barnets medborgarskap beror på föräldrarnas medborgarskap.
När ett barn föds, får barnet finskt medborgarskap om
barnets mor är finsk medborgare,
barnets far är finsk medborgare och föräldrarna är gifta,
barnets far är finsk medborgare, barnet föds utom äktenskap i Finland och faderskapet fastställs,
barnets far avled innan barnet föddes, men fadern var finsk medborgare och gift med barnets mor medan han levde eller
barnets far avled innan barnet föddes, barnet föds utom äktenskap i Finland och faderskapet fastställs.
Ett barn får finskt medborgarskap också om hen föds i Finland och inte får medborgarskap i något annan land av sina föräldrar.
I detta fall fastställer Migrationsverket barnets medborgarskap.
Ett barn kan samtidigt ha både finskt medborgarskap och medborgarskap i ett annat land, om det andra landet godkänner flerfaldigt medborgarskap.
Fråga mer om detta vid ditt eget lands beskickning.
Läs mer om finskt medborgarskap på InfoFinlands sida Finskt medborgarskap.
Finskt medborgarskap till barn med finsk farfinska _ svenska _ engelska
Att ansöka om finskt medborgarskapfinska _ svenska _ engelska
Om barnet inte får finskt medborgarskap
Om ditt barn inte får finskt medborgarskap vid födelsen ska du ansöka om ett pass för barnet vid ditt hemlands beskickning.
För detta behöver du barnets födelseattest från magistraten.
På InfoFinlands sida Ambassader i Finland hittar du information om andra länders beskickningar i Finland.
Därefter måste du ansöka om uppehållstillstånd eller registrering av EU-medborgares uppehållsrätt för barnet.
Om barnet får medborgarskap i ett EU-land, ska du ansöka om registrering av EU-medborgares uppehållsrätt för barnet i Migrationsverkets e-tjänst Enter Finland eller vid Migrationsverkets serviceställe.
Om barnet får medborgarskap i ett annat land, ska du ansöka om uppehållstillstånd för barnet i Migrationsverkets e-tjänst Enter Finland eller vid Migrationsverkets serviceställe.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Barnets sociala trygghet
Om barnet omfattas av Den sociala tryggheten i Finland får hen ett FPA-kort, det vill säga ett sjukförsäkringskort.
FPA skickar kortet hem efter att barnet har fått en personbeteckning och ett namn.
Du måste ansöka om familjeförmåner separat från FPA.
Läs mer om ämnet på InfoFinlands sidor Stöd till gravida och Stöd efter barnets födelse.
Erkännande av faderskap
Om barnets föräldrar är gifta behöver faderskapet inte erkännas separat.
Om barnets mor och far inte är gifta och faderskapet inte erkänns, är barnet officiellt faderlöst.
Faderskapet kan erkänns redan under graviditeten vid mödrarådgivningsbyrån eller efter barnets födelse hos barnatillsyningsmannen i den egna kommunen.
Om faderskapet erkänts före födelsen inleds behandlingen av faderskapsärendet först 30 dagar efter barnets födelse.
Magistraten bekräftar erkännandet av faderskapet.
Läs mer på InfoFinlands sida Samboförhållande.
linkkiSocial- och hälsovårdsministeriet:
Erkännande och fastställande av partnerskapfinska _ svenska
Barnet måste ha en vårdnadshavare
Enligt finländsk lag är en person som är under 18 år ett barn.
Personer under 18 år ska ha minst en vårdnadshavare.
Vanligtvis är barnets föräldrar dess vårdnadshavare.
Om ett barn föds inom äktenskap är båda föräldrarna tillsammans barnets vårdnadshavare.
Om föräldrarna inte är gifta och faderskapet inte har erkänts, är modern barnets vårdnadshavare och bestämmer ensam om alla barnets angelägenheter.
Detta innebär att modern ensam bestämmer om barnets angelägenheter även om föräldrarna bor tillsammans.
Fadern får vårdnad om barnet om föräldrarna ingår ett avtal om gemensam vårdnad och faderskapet har erkänts.
Vårdnadsavtalet ingås antingen på rådgivningsbyrån före barnets födelse eller hos barnatillsyningsmannen efter barnets födelse.
Barnets födelse registreras på sjukhuset
Vilket medborgarskap får barnet?
Om barnet inte får finskt medborgarskap
Barnets sociala trygghet
Erkännande av faderskap
Barnet måste ha en vårdnadshavare
Barnets födelse registreras på sjukhuset
När ett barn har fötts registrerar sjukhuset födelsen i Finlands befolkningsdatasystem, och barnet får en tillfällig personbeteckning.
Detta görs om
barnets mor har uppehållsrätt i Finland,
modern har en hemkommun i Finland och
modern har en finsk personbeteckning.
Om barnets mor inte är registrerad i Finland kan sjukhuset inte registrera födelsen och magistraten skickar ingen blankett till modern.
I detta fall ska du kontakta magistraten och be om anvisningar om hur barnet registreras.
Du kan läsa mer om registreringen av modern på InfoFinlands sida Registrering som invånare.
Kontaktuppgifter till magistratfinska _ svenska _ engelska
Inom två veckor efter att barnets födelse registrerats skickar magistraten en blankett hem till modern.
Med den här blanketten kan du meddela följande information till myndigheterna:
modersmål
religion.
Fyll i blanketten noggrant och underteckna den.
Om föräldrarna är gifta ska båda föräldrarna underteckna blanketten.
Returnera blanketten till magistraten inom två månader efter att barnet fötts.
Du kan skicka blanketten per post eller lämna den personligen till magistraten i ditt område.
Först efter detta registreras ditt barn i befolkningsdatasystemet.
I Finland finns en namnlag. Enligt den ska alla som har en hemort i Finland ha ett efternamn och 1–4 förnamn.
Förnamnen ska vara förenliga med Finlands namnlag.
Till exempel får syskon inte ha samma namn som första namn.
Barnet får efternamn av sina föräldrar.
Om föräldrarna har samma efternamn, blir detta även barnets efternamn.
Om föräldrarna har olika efternamn beror barnets efternamn på situationen.
Om föräldrarna är gifta kan de välja endera makens efternamn till barnet.
Om föräldrarna inte är gifta kan barnet få antingen moderns eller faderns efternamn, om faderskapet har fastställts.
Läs mer om fastställande av faderskap vid punkten Erkännande av faderskap på den här sidan.
Om föräldrarna har ett kombinerat efternamn, blir detta även barnets efternamn.
Om föräldrarna har gemensamma barn sedan tidigare, ska minderåriga syskon ha samma efternamn.
Om föräldrarna har separerat, bestämmer barnets vårdnadshavare vilket namn barnet får.
Om föräldrarna inte kommer överens om barnets efternamn, får barnet moderns efternamn.
Broschyren Makens efternamn och barnets efternamnfinska _ svenska _ engelska
Namnlagenfinska _ svenska
Barnets modersmål
När barnet föds måste man registrera dess modersmål.
Det är obligatoriskt att registrera språket.
Ditt barn kan endast ha ett språk som modersmål.
Du kan ändra språket senare om du vill.
Det är bra att fundera på vilket språk du vill registrera för ditt barn.
Språkvalet kan påverka barnets möjligheter att studera olika språk i skolan.
Barn, vars modersmål inte är finska eller svenska, studerar finska eller svenska som andraspråk i den så kallade S2-undervisningen.
Barnet kan även läsa sitt eget modersmål om man har registrerat något annat språk än finska eller svenska som modersmål för barnet.
Att delta i modersmålsundervisningen är frivilligt.
linkkiUtbildningsstyrelsen:
Eget språk, eget sinne(pdf, 789.88 KB)finska
Barnets religion
Barnets religion är familjens ensak.
Du får själv bestämma vilket trossamfund ditt barn ska höra till.
Det är inte obligatoriskt att ange barnets religion.
Om den ena föräldern har ensam vårdnad om barnet, kan den föräldern ensam bestämma vilket trossamfund barnet ska höra till.
linkkiUndervisnings- och kulturministeriet:
Religionsfrihetfinska _ svenska _ engelska
linkkiFritänkarförbundet r.f.:
Religionsfriheten för barn och ungafinska
Vilket medborgarskap får barnet?
Barnets medborgarskap beror på föräldrarnas medborgarskap.
När ett barn föds, får barnet finskt medborgarskap om
barnets mor är finsk medborgare,
barnets far är finsk medborgare och föräldrarna är gifta,
barnets far är finsk medborgare, barnet föds utom äktenskap i Finland och faderskapet fastställs,
barnets far avled innan barnet föddes, men fadern var finsk medborgare och gift med barnets mor medan han levde eller
barnets far avled innan barnet föddes, barnet föds utom äktenskap i Finland och faderskapet fastställs.
Ett barn får finskt medborgarskap också om hen föds i Finland och inte får medborgarskap i något annan land av sina föräldrar.
I detta fall fastställer Migrationsverket barnets medborgarskap.
Ett barn kan samtidigt ha både finskt medborgarskap och medborgarskap i ett annat land, om det andra landet godkänner flerfaldigt medborgarskap.
Fråga mer om detta vid ditt eget lands beskickning.
Läs mer om finskt medborgarskap på InfoFinlands sida Finskt medborgarskap.
Finskt medborgarskap till barn med finsk farfinska _ svenska _ engelska
Att ansöka om finskt medborgarskapfinska _ svenska _ engelska
Om barnet inte får finskt medborgarskap
Om ditt barn inte får finskt medborgarskap vid födelsen ska du ansöka om ett pass för barnet vid ditt hemlands beskickning.
För detta behöver du barnets födelseattest från magistraten.
På InfoFinlands sida Ambassader i Finland hittar du information om andra länders beskickningar i Finland.
Därefter måste du ansöka om uppehållstillstånd eller registrering av EU-medborgares uppehållsrätt för barnet.
Om barnet får medborgarskap i ett EU-land, ska du ansöka om registrering av EU-medborgares uppehållsrätt för barnet i Migrationsverkets e-tjänst Enter Finland eller vid Migrationsverkets serviceställe.
Om barnet får medborgarskap i ett annat land, ska du ansöka om uppehållstillstånd för barnet i Migrationsverkets e-tjänst Enter Finland eller vid Migrationsverkets serviceställe.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Barnets sociala trygghet
Om barnet omfattas av Den sociala tryggheten i Finland får hen ett FPA-kort, det vill säga ett sjukförsäkringskort.
FPA skickar kortet hem efter att barnet har fått en personbeteckning och ett namn.
Du måste ansöka om familjeförmåner separat från FPA.
Läs mer om ämnet på InfoFinlands sidor Stöd till gravida och Stöd efter barnets födelse.
Erkännande av faderskap
Om barnets föräldrar är gifta behöver faderskapet inte erkännas separat.
Om barnets mor och far inte är gifta och faderskapet inte erkänns, är barnet officiellt faderlöst.
Faderskapet kan erkänns redan under graviditeten vid mödrarådgivningsbyrån eller efter barnets födelse hos barnatillsyningsmannen i den egna kommunen.
Om faderskapet erkänts före födelsen inleds behandlingen av faderskapsärendet först 30 dagar efter barnets födelse.
Magistraten bekräftar erkännandet av faderskapet.
Läs mer på InfoFinlands sida Samboförhållande.
linkkiSocial- och hälsovårdsministeriet:
Erkännande och fastställande av partnerskapfinska _ svenska
Barnet måste ha en vårdnadshavare
Enligt finländsk lag är en person som är under 18 år ett barn.
Personer under 18 år ska ha minst en vårdnadshavare.
Vanligtvis är barnets föräldrar dess vårdnadshavare.
Om ett barn föds inom äktenskap är båda föräldrarna tillsammans barnets vårdnadshavare.
Om föräldrarna inte är gifta och faderskapet inte har erkänts, är modern barnets vårdnadshavare och bestämmer ensam om alla barnets angelägenheter.
Detta innebär att modern ensam bestämmer om barnets angelägenheter även om föräldrarna bor tillsammans.
Fadern får vårdnad om barnet om föräldrarna ingår ett avtal om gemensam vårdnad och faderskapet har erkänts.
Vårdnadsavtalet ingås antingen på rådgivningsbyrån före barnets födelse eller hos barnatillsyningsmannen efter barnets födelse.
Förskoleundervisning
Mångkulturell barndagvård
Grundläggande utbildning
Förberedande utbildning inför yrkesutbildning
Yrkesutbildning
Högskolor
Medborgarinstitut
Hjälp i frågor om utbildning
Förskoleundervisning
Förskoleundervisningen är avsedd för sexåringar och den ges vid daghem.
I förskoleundervisningen skaffar sig barnet förberedande färdigheter inför grundskolan.
Förskoleundervisningen ges vanligen på förmiddagen och på eftermiddagen kan barnet vara i dagvården.
Förskoleundervisningen börjar i augusti och anmälan ska göras i februari.
Blivande förskolebarn får mer information om detta per post, på dagvårdens webbplats och i lokaltidningen.
Alla som ansöker om en förskoleplats ska lämna in en ansökan om förskoleundervisning.
Man kan anmäla sig till förskoleundervisningen antingen elektroniskt eller med en ansökningsblankett.
Läs mer:
Mångkulturell barndagvård
Mångkulturell barndagvård i Rovaniemi betyder att alla barn beaktas likvärdigt och rättvist oavsett ålder, kön eller hudfärg.
I tillgången till dagvårdstjänster är målet att uppfylla närserviceprincipen för varje barn.
I dagvården lär barnet känna den finländska kulturen, lär sig det finska språket och verkar i en social grupp.
Familjer med främmande modersmål har vid behov rätt till tolktjänster.
Dagvården samarbetar med invandrarbyrån i frågor som rör barnet och familjen.
När barnet börjar i dagvården fyller man tillsammans med familjen i blanketten Uppgifter om invandrarbarn.
Grundläggande utbildning
Anmälan till grundskolan
I Rovaniemi stad finns 23 skolor med årskurserna 1–6, Lapplands övningsskola som upprätthålls av
Lapplands universitet och Rovaniemi Steinerskola som är en privatskola.
Rovaniemi stads skoltjänster är indelade i fyra områden som även fungerar som elevantagningsområden.
Elevens närskola bestäms enligt gränserna för dessa områden.
Anmälan till grundskolan sker vid den skola som anges i ett brev som varje ny elev får hem eller per telefon till skolan.
Läs mer:
Anmälan till den grundläggande utbildningen
Undervisning för invandrare
Invandrarelever använder i huvudsak grundskolans och gymnasieskolans vanliga tjänster.
För barn som nyligen invandrat ordnas förberedande undervisning inför grundskolan som vanligtvis pågår i ett år.
För elever som nyligen invandrat finns en klass för förberedande undervisning inför grundskolan vid skolan
Särdrag i undervisningen
Modersmålsundervisning ges i ryska och i mån av möjlighet även i andra språk.
Finska undervisas som främmande språk och målet är en funktionell tvåspråkighet.
Om det finns minst tre elever som befriats från religionsundervisningen och deras föräldrar kräver detta, ordnas undervisning i elevernas egen religion.
Invandrareleverna bedöms som regel enligt grundskolans allmänna bedömningsgrunder med beaktande av elevens utgångsläge.
Under de tre första åren i landet får invandrareleverna en särskild stödundervisning avsedd för dem.
Också nya elever har rätt till denna stödundervisning.
Grundskolans övriga stödåtgärder omfattar den övriga stödundervisningen i grundskolan, specialundervisning, individuella studieplaner, flexibel bedömning,
Undervisning för invandrare
Förberedande utbildning inför yrkesutbildning
Lapplands yrkesinstitut
Lapplands yrkesinstitut erbjuder förberedande utbildning för invandrare som vill söka till yrkesutbildning.
Läs mer:
linkkiLapplands yrkeshögskola:
Lapplands yrkeshögskolafinska _ engelska
Rovala-institutets utbildning för invandrare
I Rovala-institutets utbildning för invandrare kan man studera det finska språket och den finska kulturen, arbetslivsfärdigheter och skaffa sig kunskaper om det finländska samhället.
Studerandena inom integrationsutbildningen kommer från tiotals olika länder och undervisningsspråket är finska. En kurs kan ha 8
–15 studeranden och vanligtvis finns det 8–10 undervisningsgrupper.
Integrationsutbildningen är arbetskraftsutbildning och man söker till kurserna via Rovaniemi TE-byrå.
De som är klienter vid FPA kan få utbildningsstöd under utbildningen.
Kursansökan kan lämnas in via Internet.
För den som flyttar till Finland är det viktigt att känna till de grundläggande reglerna som gäller i arbetslivet och det finländska samhället.
På kursen lär de studerande sig det grundläggande om arbetslivet, tränar på sin
jobbsökningsförmåga och planerar sin framtid.
Läs mer:
Utbildning för invandrare
Yrkesutbildning
Lapplands yrkesinstitut
Vid Lapplands yrkesinstitut kan du studera och skaffa dig yrkesinriktad grundutbildning och vuxenutbildning i alla studieområden förutom inom idrottsområdet och turism-, kosthålls- och ekonomibranschen.
Läs mer:
Lapplands yrkesinstitut
Läroavtalsutbildning
Lapplands läroavtalscenter
Lapplands läroavtalscenter ordnar läroavtalsutbildning enligt lagen om yrkesutbildning och lagen om yrkesinriktad vuxenutbildning samt stödtjänster för arbetslivet och regionutvecklingen.
Läs mer:
Lapplands läroavtalscenterfinska
Gymnasium
På Rovaniemi stads område finns det fyra gymnasiealternativ: gymnasieskolorna Lyseonpuiston lukio, Muurolan lukio och Ounasvaaran lukio samt yrkesgymnasiet Rovaniemen ammattilukio.
Läs mer:
Gymnasieskolorfinska
Högskolor
Rovaniemi yrkeshögskola
Rovaniemi yrkeshögskola eller RAMK är den nordligaste yrkeshögskolan inom EU. Skolan ingår i Lapplands högskolekoncern.
Vid RAMK finns det elva finskspråkiga och tre engelskspråkiga utbildningsprogram som leder till yrkeshögskoleexamen, fem utbildningsprogram som leder till högre
Läs mer:
Lapplands yrkeshögskola
Vid vårt vetenskaps- och konstuniversitet fås utbildning och idkas forskning inom pedagogik, turism och affärsverksamhet, juridik, konstindustri och samhällsvetenskaper.
Inom forskningen har universitetet två tvärvetenskapliga och internationella
profilområden: forskning i arktiska och nordliga frågor och forskning inom turism.
Läs mer
Lapplands universitetfinska _ engelska
Lapplands öppna universitet
Det öppna universitetet vid Lapplands universitet erbjuder studiemöjligheter enligt studiekraven vid de pedagogiska, juridiska, konst- och samhällsvetenskapliga fakulteterna.
Utbudet kompletteras av språk- och metodstudier.
Läs mer:
Lapplands öppna universitetfinska _ engelska
Medborgarinstitut
Vid medborgarinstitutet kan du studera och idka som hobby till exempel språk, konstämnen, motion med mera.
I Rovaniemi finns två medborgarinstitut. Mer information om dessa hittar du på följande adresser:
Läs mer:
Hjälp i frågor om utbildning
Arbetskraftsbyråns informationstjänst för utbildning och yrkesval
Informationstjänsten för utbildning och yrkesval vid arbetskraftsbyrån i Rovaniemi
Valtakatu 16
Arbetskraftsrådgivare 010 604 6590
MoniNet
MoniNet är ett mångkulturellt center i Rovaniemi, Lappland.
Det upprätthålls av föreningen Rovalan Setlementti ry.
Det erbjuder tjänster för invandrare som bor i Rovaniemi och andra områden i Lapplands län.
Vi betjänar på finska, engelska, ryska och svenska.
Kontaktuppgifter:
MoniNet
Etelärinne 32
tfn 040 559 6564
Läs mer:
MoniNet
Förskoleundervisning
Mångkulturell barndagvård
Grundläggande utbildning
Förberedande utbildning inför yrkesutbildning
Yrkesutbildning
Högskolor
Medborgarinstitut
Hjälp i frågor om utbildning
Förskoleundervisning
Förskoleundervisningen är avsedd för sexåringar och den ges vid daghem.
I förskoleundervisningen skaffar sig barnet förberedande färdigheter inför grundskolan.
Förskoleundervisningen ges vanligen på förmiddagen och på eftermiddagen kan barnet vara i dagvården.
Förskoleundervisningen börjar i augusti och anmälan ska göras i februari.
Blivande förskolebarn får mer information om detta per post, på dagvårdens webbplats och i lokaltidningen.
Alla som ansöker om en förskoleplats ska lämna in en ansökan om förskoleundervisning.
Man kan anmäla sig till förskoleundervisningen antingen elektroniskt eller med en ansökningsblankett.
Läs mer:
Mångkulturell barndagvård
Mångkulturell barndagvård i Rovaniemi betyder att alla barn beaktas likvärdigt och rättvist oavsett ålder, kön eller hudfärg.
I tillgången till dagvårdstjänster är målet att uppfylla närserviceprincipen för varje barn.
I dagvården lär barnet känna den finländska kulturen, lär sig det finska språket och verkar i en social grupp.
Familjer med främmande modersmål har vid behov rätt till tolktjänster.
Dagvården samarbetar med invandrarbyrån i frågor som rör barnet och familjen.
När barnet börjar i dagvården fyller man tillsammans med familjen i blanketten Uppgifter om invandrarbarn.
Grundläggande utbildning
Anmälan till grundskolan
I Rovaniemi stad finns 23 skolor med årskurserna 1–6, Lapplands övningsskola som upprätthålls av
Lapplands universitet och Rovaniemi Steinerskola som är en privatskola.
Rovaniemi stads skoltjänster är indelade i fyra områden som även fungerar som elevantagningsområden.
Elevens närskola bestäms enligt gränserna för dessa områden.
Anmälan till grundskolan sker vid den skola som anges i ett brev som varje ny elev får hem eller per telefon till skolan.
Läs mer:
Anmälan till den grundläggande utbildningen
Undervisning för invandrare
Invandrarelever använder i huvudsak grundskolans och gymnasieskolans vanliga tjänster.
För barn som nyligen invandrat ordnas förberedande undervisning inför grundskolan som vanligtvis pågår i ett år.
För elever som nyligen invandrat finns en klass för förberedande undervisning inför grundskolan vid skolan
Särdrag i undervisningen
Modersmålsundervisning ges i ryska och i mån av möjlighet även i andra språk.
Finska undervisas som främmande språk och målet är en funktionell tvåspråkighet.
Om det finns minst tre elever som befriats från religionsundervisningen och deras föräldrar kräver detta, ordnas undervisning i elevernas egen religion.
Invandrareleverna bedöms som regel enligt grundskolans allmänna bedömningsgrunder med beaktande av elevens utgångsläge.
Under de tre första åren i landet får invandrareleverna en särskild stödundervisning avsedd för dem.
Också nya elever har rätt till denna stödundervisning.
Grundskolans övriga stödåtgärder omfattar den övriga stödundervisningen i grundskolan, specialundervisning, individuella studieplaner, flexibel bedömning,
Undervisning för invandrare
Förberedande utbildning inför yrkesutbildning
Lapplands yrkesinstitut
Lapplands yrkesinstitut erbjuder förberedande utbildning för invandrare som vill söka till yrkesutbildning.
Läs mer:
linkkiLapplands yrkeshögskola:
Lapplands yrkeshögskolafinska _ engelska
Rovala-institutets utbildning för invandrare
I Rovala-institutets utbildning för invandrare kan man studera det finska språket och den finska kulturen, arbetslivsfärdigheter och skaffa sig kunskaper om det finländska samhället.
Studerandena inom integrationsutbildningen kommer från tiotals olika länder och undervisningsspråket är finska. En kurs kan ha 8
–15 studeranden och vanligtvis finns det 8–10 undervisningsgrupper.
Integrationsutbildningen är arbetskraftsutbildning och man söker till kurserna via Rovaniemi TE-byrå.
De som är klienter vid FPA kan få utbildningsstöd under utbildningen.
Kursansökan kan lämnas in via Internet.
För den som flyttar till Finland är det viktigt att känna till de grundläggande reglerna som gäller i arbetslivet och det finländska samhället.
På kursen lär de studerande sig det grundläggande om arbetslivet, tränar på sin
jobbsökningsförmåga och planerar sin framtid.
Läs mer:
Utbildning för invandrare
Yrkesutbildning
Lapplands yrkesinstitut
Vid Lapplands yrkesinstitut kan du studera och skaffa dig yrkesinriktad grundutbildning och vuxenutbildning i alla studieområden förutom inom idrottsområdet och turism-, kosthålls- och ekonomibranschen.
Läs mer:
Lapplands yrkesinstitut
Läroavtalsutbildning
Lapplands läroavtalscenter
Lapplands läroavtalscenter ordnar läroavtalsutbildning enligt lagen om yrkesutbildning och lagen om yrkesinriktad vuxenutbildning samt stödtjänster för arbetslivet och regionutvecklingen.
Läs mer:
Lapplands läroavtalscenterfinska
Gymnasium
På Rovaniemi stads område finns det fyra gymnasiealternativ: gymnasieskolorna Lyseonpuiston lukio, Muurolan lukio och Ounasvaaran lukio samt yrkesgymnasiet Rovaniemen ammattilukio.
Läs mer:
Gymnasieskolorfinska
Högskolor
Rovaniemi yrkeshögskola
Rovaniemi yrkeshögskola eller RAMK är den nordligaste yrkeshögskolan inom EU. Skolan ingår i Lapplands högskolekoncern.
Vid RAMK finns det elva finskspråkiga och tre engelskspråkiga utbildningsprogram som leder till yrkeshögskoleexamen, fem utbildningsprogram som leder till högre
Läs mer:
Lapplands yrkeshögskola
Vid vårt vetenskaps- och konstuniversitet fås utbildning och idkas forskning inom pedagogik, turism och affärsverksamhet, juridik, konstindustri och samhällsvetenskaper.
Inom forskningen har universitetet två tvärvetenskapliga och internationella
profilområden: forskning i arktiska och nordliga frågor och forskning inom turism.
Läs mer
Lapplands universitetfinska _ engelska
Lapplands öppna universitet
Det öppna universitetet vid Lapplands universitet erbjuder studiemöjligheter enligt studiekraven vid de pedagogiska, juridiska, konst- och samhällsvetenskapliga fakulteterna.
Utbudet kompletteras av språk- och metodstudier.
Läs mer:
Lapplands öppna universitetfinska _ engelska
Medborgarinstitut
Vid medborgarinstitutet kan du studera och idka som hobby till exempel språk, konstämnen, motion med mera.
I Rovaniemi finns två medborgarinstitut. Mer information om dessa hittar du på följande adresser:
Läs mer:
Hjälp i frågor om utbildning
Arbetskraftsbyråns informationstjänst för utbildning och yrkesval
Informationstjänsten för utbildning och yrkesval vid arbetskraftsbyrån i Rovaniemi
Valtakatu 16
Arbetskraftsrådgivare 010 604 6590
MoniNet
MoniNet är ett mångkulturellt center i Rovaniemi, Lappland.
Det upprätthålls av föreningen Rovalan Setlementti ry.
Det erbjuder tjänster för invandrare som bor i Rovaniemi och andra områden i Lapplands län.
Vi betjänar på finska, engelska, ryska och svenska.
Kontaktuppgifter:
MoniNet
Etelärinne 32
tfn 040 559 6564
Läs mer:
MoniNet
Förskoleundervisning Mångkulturell barndagvård
Grundläggande utbildning
Förberedande utbildning inför yrkesutbildning
Yrkesutbildning Högskolor
Medborgarinstitut
Hjälp i frågor om utbildning
Förskoleundervisning
Förskoleundervisningen är avsedd för sexåringar och den ges vid daghem.
I förskoleundervisningen skaffar sig barnet förberedande färdigheter inför grundskolan.
Förskoleundervisningen ges vanligen på förmiddagen och på eftermiddagen kan barnet vara i dagvården.
Förskoleundervisningen börjar i augusti och anmälan ska göras i februari.
Blivande förskolebarn får mer information om detta per post, på dagvårdens webbplats och i lokaltidningen.
Alla som ansöker om en förskoleplats ska lämna in en ansökan om förskoleundervisning.
Mångkulturell barndagvård i Rovaniemi betyder att alla barn beaktas likvärdigt och rättvist oavsett ålder, kön eller hudfärg.
I tillgången till dagvårdstjänster är målet att uppfylla närserviceprincipen för varje barn.
I dagvården lär barnet känna den finländska kulturen, lär sig det finska språket och verkar i en social grupp.
Familjer med främmande modersmål har vid behov rätt till tolktjänster.
Dagvården samarbetar med invandrarbyrån i frågor som rör barnet och familjen.
När barnet börjar i dagvården fyller man tillsammans med familjen i blanketten Uppgifter om invandrarbarn.
Anmälan till grundskolan
Lapplands universitet och Rovaniemi Steinerskola som är en privatskola.
Rovaniemi stads skoltjänster är indelade i fyra områden som även fungerar som elevantagningsområden.
Elevens närskola bestäms enligt gränserna för dessa områden. Närskolan är i regel den skola som ligger närmast elevens hem.
Anmälan till grundskolan sker vid den skola som anges i ett brev som varje ny elev får hem eller per telefon till skolan.
Grundläggande utbildning
Undervisning för invandrare
Invandrarelever använder i huvudsak grundskolans och gymnasieskolans vanliga tjänster.
För barn som nyligen invandrat ordnas förberedande undervisning inför grundskolan som vanligtvis pågår i ett år.
För elever som nyligen invandrat finns en klass för förberedande undervisning inför grundskolan vid skolan
Därefter placeras invandrareleverna i en finskspråkig klass i sin närskola.
Särdrag i undervisningen
Modersmålsundervisning ges i ryska och i mån av möjlighet även i andra språk.
Om det finns minst tre elever som befriats från religionsundervisningen och deras föräldrar kräver detta, ordnas undervisning i elevernas egen religion.
Invandrareleverna bedöms som regel enligt grundskolans allmänna bedömningsgrunder med beaktande av elevens utgångsläge.
Under de tre första åren i landet får invandrareleverna en särskild stödundervisning avsedd för dem.
Också nya elever har rätt till denna stödundervisning.
Undervisning för invandrare
Lapplands yrkesinstitut
Lapplands yrkesinstitut erbjuder förberedande utbildning för invandrare som vill söka till yrkesutbildning.
Lapplands yrkeshögskolafinska _ engelska
Rovala-institutets utbildning för invandrare
I Rovala-institutets utbildning för invandrare kan man studera det finska språket och den finska kulturen, arbetslivsfärdigheter och skaffa sig kunskaper om det finländska samhället.
I integrationsutbildningen studerar man finska, kommunikationsfärdigheter och mycket annat. För den som flyttar till
Finland är det viktigt att känna till de grundläggande reglerna som gäller i arbetslivet och det finländska samhället.
jobbsökningsförmåga och planerar sin framtid.
Utbildning för invandrare
Yrkesutbildning
Vid Lapplands yrkesinstitut kan du studera och skaffa dig yrkesinriktad grundutbildning och vuxenutbildning i alla studieområden förutom inom idrottsområdet och turism-, kosthålls- och ekonomibranschen.
Läs mer:
Lapplands yrkesinstitut
Lapplands läroavtalscenter
Lapplands läroavtalscenterfinska
Högskolor Rovaniemi yrkeshögskola
Rovaniemi yrkeshögskola eller RAMK är den nordligaste yrkeshögskolan inom EU. Skolan ingår i Lapplands högskolekoncern.
Vid RAMK finns det elva finskspråkiga och tre engelskspråkiga utbildningsprogram som leder till yrkeshögskoleexamen, fem utbildningsprogram som leder till högre
Vid vårt vetenskaps- och konstuniversitet fås utbildning och idkas forskning inom pedagogik, turism och affärsverksamhet, juridik, konstindustri och samhällsvetenskaper.
Inom forskningen har universitetet två tvärvetenskapliga och internationella
profilområden: forskning i arktiska och nordliga frågor och forskning inom turism.
Lapplands universitetfinska _ engelska
Lapplands öppna universitet
Utbudet kompletteras av språk- och metodstudier.
Lapplands öppna universitetfinska _ engelska
Medborgarinstitut
Hjälp i frågor om utbildning
MoniNet
MoniNet är ett mångkulturellt center i Rovaniemi, Lappland. Det upprätthålls av föreningen Rovalan Setlementti ry.
Det erbjuder tjänster för invandrare som bor i Rovaniemi och andra områden i Lapplands län.
Kontaktuppgifter:
I Finland är enligt lag personer under 18 år barn.
Barn under 18 år ska alltid ha en minst en vårdnadshavare.
Vanligtvis är barnets föräldrar dess vårdnadshavare.
När en person fyller 18 år blir han eller hon myndig.
Enligt Finlands lag är alla barn jämställda oavsett bakgrund eller ålder.
Rättigheterna och skyldigheterna enligt Finlands grundlag gäller alla barn som bor i Finland.
Enligt grundlagen ska barn bemötas som jämlika individer och de ska ha rätt till medinflytande i frågor som gäller dem själva.
Ta också del av InfoFinlands sidor Ekonomiskt stöd till familjer och Vård av barnet.
I Finland är enligt lag personer under 18 år barn.
Barn under 18 år ska alltid ha en minst en vårdnadshavare.
Vanligtvis är barnets föräldrar dess vårdnadshavare.
När en person fyller 18 år blir han eller hon myndig.
Enligt Finlands lag är alla barn jämställda oavsett bakgrund eller ålder.
Rättigheterna och skyldigheterna enligt Finlands grundlag gäller alla barn som bor i Finland.
Enligt grundlagen ska barn bemötas som jämlika individer och de ska ha rätt till medinflytande i frågor som gäller dem själva.
Ta också del av InfoFinlands sidor Ekonomiskt stöd till familjer och Vård av barnet.
I Finland är enligt lag personer under 18 år barn.
Barn under 18 år ska alltid ha en minst en vårdnadshavare.
Vanligtvis är barnets föräldrar dess vårdnadshavare.
När en person fyller 18 år blir han eller hon myndig.
Enligt Finlands lag är alla barn jämställda oavsett bakgrund eller ålder.
Rättigheterna och skyldigheterna enligt Finlands grundlag gäller alla barn som bor i Finland.
Enligt grundlagen ska barn bemötas som jämlika individer och de ska ha rätt till medinflytande i frågor som gäller dem själva.
Ta också del av InfoFinlands sidor Ekonomiskt stöd till familjer och Vård av barnet.
Ett samboförhållande upphör när parterna inte längre bor på samma adress.
Upphörandet av samboförhållandet kan påverka till exempel de stöd som FPA betalar och barnens dagvårdsavgifter.
Du ska själv meddela att samboförhållandet har upphört.
Om samborna har gemensamma minderåriga barn ska de tillsammans besluta om barnens situation på samma sätt som vid skilsmässa.
Också sambor kan få hjälp med att komma överens om saker och ting, till exempel genom medling i familjefrågor.
Läs mer på InfoFinlands sida Barn vid skilsmässa.
I ett samboförhållande kan makarna ha ett gemensamt efternamn.
Efternamnet påverkas inte av att samboförhållandet eventuellt upphör.
Om du vill byta efternamn ska du ansöka om namnändring hos magistraten.
I ett samboförhållande behåller vardera part sin egen egendom.
När samboförhållandet upphör delas egendomen vanligtvis så att båda parterna får sin egen egendom.
Om samborna förvärvar egendom tillsammans ska båda parterna antecknas som köpare och alla kvitton sparas.
Då delas denna egendom jämnt om samboförhållandet upphör.
Om bara en av parterna står som köpare är denne ägare till egendomen när samboförhållandet upphör.
Sambor kan ha sådan egendom om vars ägande de inte har en överenskommelse.
Då utgår man ifrån att båda äger en lika stor andel och denna egendom delas på hälft.
Om fördelningen av ägodelarna blir stridig, kan samborna i vissa fall ansöka om en bodelningsman hos tingsrätten som hjälper i bodelningen.
Man kan ansöka om bodelningsman om samboförhållandet har varat minst fem år och parterna har gemensamma barn.
I vissa fall kan den ena sambon få jämkning av den andra sambon när paret skiljer sig.
En sambo kan få jämkning om han eller hon till exempel genom arbete hjälpt den andra sambon att utöka sin egendom och för att det därför skulle vara orättvist att fördela egendomen enbart baserat på ägarskapet.
Om samboförhållandet upphör på grund av att den ena parten dör, ärver samborna inte varandra.
Sambor har till exempel inte rätt att bo kvar i familjens gemensamma hem om det tillhör den döda sambon.
Arvet går till den döda makens barn eller syskon.
Sambor kan dock upprätta ett testamente (testamentti) för det fall att någon avlider.
Genom testamente kan de säkerställa att en viss egendom, till exempel den gemensamma bostaden, ärvs av sambon.
Sambor kan även upprätta ett skriftligt avtal om hur egendomen ska fördelas om paret går isär.
Om du vill upprätta ett avtal eller ett testamente för fördelning av egendomen i ett samboförhållande, kan du be om råd till exempel vid rättshjälpsbyrån eller av en jurist.
linkkiRättsväsendet:
Rättshjälpsbyråerfinska _ svenska _ engelska
Ett samboförhållande upphör när parterna inte längre bor på samma adress.
Upphörandet av samboförhållandet kan påverka till exempel de stöd som FPA betalar och barnens dagvårdsavgifter.
Du ska själv meddela att samboförhållandet har upphört.
Om samborna har gemensamma minderåriga barn ska de tillsammans besluta om barnens situation på samma sätt som vid skilsmässa.
Också sambor kan få hjälp med att komma överens om saker och ting, till exempel genom medling i familjefrågor.
Läs mer på InfoFinlands sida Barn vid skilsmässa.
I ett samboförhållande kan makarna ha ett gemensamt efternamn.
Efternamnet påverkas inte av att samboförhållandet eventuellt upphör.
Om du vill byta efternamn ska du ansöka om namnändring hos magistraten.
I ett samboförhållande behåller vardera part sin egen egendom.
När samboförhållandet upphör delas egendomen vanligtvis så att båda parterna får sin egen egendom.
Om samborna förvärvar egendom tillsammans ska båda parterna antecknas som köpare och alla kvitton sparas.
Då delas denna egendom jämnt om samboförhållandet upphör.
Om bara en av parterna står som köpare är denne ägare till egendomen när samboförhållandet upphör.
Sambor kan ha sådan egendom om vars ägande de inte har en överenskommelse.
Då utgår man ifrån att båda äger en lika stor andel och denna egendom delas på hälft.
Om fördelningen av ägodelarna blir stridig, kan samborna i vissa fall ansöka om en bodelningsman hos tingsrätten som hjälper i bodelningen.
Man kan ansöka om bodelningsman om samboförhållandet har varat minst fem år och parterna har gemensamma barn.
I vissa fall kan den ena sambon få jämkning av den andra sambon när paret skiljer sig.
En sambo kan få jämkning om han eller hon till exempel genom arbete hjälpt den andra sambon att utöka sin egendom och för att det därför skulle vara orättvist att fördela egendomen enbart baserat på ägarskapet.
Om samboförhållandet upphör på grund av att den ena parten dör, ärver samborna inte varandra.
Sambor har till exempel inte rätt att bo kvar i familjens gemensamma hem om det tillhör den döda sambon.
Arvet går till den döda makens barn eller syskon.
Sambor kan dock upprätta ett testamente (testamentti) för det fall att någon avlider.
Genom testamente kan de säkerställa att en viss egendom, till exempel den gemensamma bostaden, ärvs av sambon.
Sambor kan även upprätta ett skriftligt avtal om hur egendomen ska fördelas om paret går isär.
Om du vill upprätta ett avtal eller ett testamente för fördelning av egendomen i ett samboförhållande, kan du be om råd till exempel vid rättshjälpsbyrån eller av en jurist.
linkkiRättsväsendet:
Rättshjälpsbyråerfinska _ svenska _ engelska
Ett samboförhållande upphör när parterna inte längre bor på samma adress.
Upphörandet av samboförhållandet kan påverka till exempel de stöd som FPA betalar och barnens dagvårdsavgifter.
Du ska själv meddela att samboförhållandet har upphört.
Om samborna har gemensamma minderåriga barn ska de tillsammans besluta om barnens situation på samma sätt som vid skilsmässa.
Också sambor kan få hjälp med att komma överens om saker och ting, till exempel genom medling i familjefrågor.
Läs mer på InfoFinlands sida Barn vid skilsmässa.
I ett samboförhållande kan makarna ha ett gemensamt efternamn.
Efternamnet påverkas inte av att samboförhållandet eventuellt upphör.
Om du vill byta efternamn ska du ansöka om namnändring hos magistraten.
I ett samboförhållande behåller vardera part sin egen egendom.
När samboförhållandet upphör delas egendomen vanligtvis så att båda parterna får sin egen egendom.
Om samborna förvärvar egendom tillsammans ska båda parterna antecknas som köpare och alla kvitton sparas.
Då delas denna egendom jämnt om samboförhållandet upphör.
Om bara en av parterna står som köpare är denne ägare till egendomen när samboförhållandet upphör.
Sambor kan ha sådan egendom om vars ägande de inte har en överenskommelse.
Då utgår man ifrån att båda äger en lika stor andel och denna egendom delas på hälft.
Om fördelningen av ägodelarna blir stridig, kan samborna i vissa fall ansöka om en bodelningsman hos tingsrätten som hjälper i bodelningen.
Man kan ansöka om bodelningsman om samboförhållandet har varat minst fem år och parterna har gemensamma barn.
I vissa fall kan den ena sambon få jämkning av den andra sambon när paret skiljer sig.
En sambo kan få jämkning om han eller hon till exempel genom arbete hjälpt den andra sambon att utöka sin egendom och för att det därför skulle vara orättvist att fördela egendomen enbart baserat på ägarskapet.
Om samboförhållandet upphör på grund av att den ena parten dör, ärver samborna inte varandra.
Sambor har till exempel inte rätt att bo kvar i familjens gemensamma hem om det tillhör den döda sambon.
Arvet går till den döda makens barn eller syskon.
Sambor kan dock upprätta ett testamente (testamentti) för det fall att någon avlider.
Genom testamente kan de säkerställa att en viss egendom, till exempel den gemensamma bostaden, ärvs av sambon.
Sambor kan även upprätta ett skriftligt avtal om hur egendomen ska fördelas om paret går isär.
Om du vill upprätta ett avtal eller ett testamente för fördelning av egendomen i ett samboförhållande, kan du be om råd till exempel vid rättshjälpsbyrån eller av en jurist.
linkkiRättsväsendet:
Rättshjälpsbyråerfinska _ svenska _ engelska
Ett samboförhållande är ett förhållande där ett par lever tillsammans utan att vara gifta.
I Finland får alla par själva bestämma om de inleder ett samboförhållande, om spelreglerna i sin relation och om de gör slut på samboförhållandet.
Ett samboförhållande registreras inte någonstans.
Till skillnad från äktenskap
har sambor inte underhållsskyldighet gentemot varandra
ärver sambor inte varandra
kan den ena sambon inte få änkepension om den andra sambon dör.
Ni kan ta ett gemensamt efternamn om
ni har gemensamma barn eller
om ni har bott tillsammans minst fem år.
Om ni vill ha ett gemensamt efternamn ska ni skicka in en anmälan om namnändring till magistraten.
Om ni bor stadigvarande tillsammans i samma bostad, hör ni till samma hushåll.
Detta har betydelse om ni till exempel ansöker om bostadsbidrag från FPA.
Läs mer om bostadsbidrag för sambor på InfoFinlands sida Bostadsbidrag.
Äktenskap som ingåtts utomlands
Ett samboförhållande kan utgöra ett hinder för att få uppehållstillstånd.
Myndigheterna överväger beviljandet av uppehållstillstånd alltid fall för fall.
Barn till föräldrar i samboförhållande
Fastställande av faderskap (Isyyden tunnustaminen)
Om ni lever i ett samboförhållande och får ett barn ska barnets far fastställas.
Om faderskapet inte fastställs är barnet officiellt faderlöst och då ansvarar modern ensam för underhåll och vård av barnet, även om ni bor tillsammans.
Faderskapet kan fastställas vid mödravården under graviditeten.
När barnet är fött kan faderskapet fastställas hos barntillsynsmannen i hemkommunen.
Faderskapet fastställs av magistratet.
När faderskapet har fastställts
kan barnet ges faderns efternamn
kan fadern vara barnets vårdnadshavare antingen tillsammans med barnets mor eller ensam.
Vårdnadshavaren (huoltaja) är den person som ansvarar för vården och uppfostran av barnet.
är fadern förpliktad att delta i underhåll av barnet
har barnet rätt att ärva sin far och släkten på sin fars sida och tvärtom
har barnet rätt till familjepension om fadern dör.
Om fadern inte erkänner sitt faderskap kan modern väcka talan för fastställande av faderskapet.
linkkiSocial- och hälsovårdsministeriet:
Erkännande och fastställande av partnerskapfinska _ svenska
Barnets efternamn vid samboende
När ett barn föds i ett samboförhållande, kan hen få
moderns efternamn eller
faderns efternamn, om faderskapet har fastställts, eller
föräldrarnas gemensamma efternamn eller
ett kombinerat efternamn som har bildats av föräldrarnas efternamn.
Om föräldrarna inte har ett gemensamt efternamn men de har gemensamma barn, får barnet samma efternamn som dess syskon har.
Du kan ansöka om ett gemensamt efternamn med din sambo
om ni har bott tillsammans minst fem år eller
Ett samboförhållande är ett förhållande där ett par lever tillsammans utan att vara gifta.
I Finland får alla par själva bestämma om de inleder ett samboförhållande, om spelreglerna i sin relation och om de gör slut på samboförhållandet.
Ett samboförhållande registreras inte någonstans.
Till skillnad från äktenskap
har sambor inte underhållsskyldighet gentemot varandra
ärver sambor inte varandra
kan den ena sambon inte få änkepension om den andra sambon dör.
Ni kan ta ett gemensamt efternamn om
ni har gemensamma barn eller
om ni har bott tillsammans minst fem år.
Om ni vill ha ett gemensamt efternamn ska ni skicka in en anmälan om namnändring till magistraten.
Om ni bor stadigvarande tillsammans i samma bostad, hör ni till samma hushåll.
Detta har betydelse om ni till exempel ansöker om bostadsbidrag från FPA.
Läs mer om bostadsbidrag för sambor på InfoFinlands sida Bostadsbidrag.
Äktenskap som ingåtts utomlands
Ett samboförhållande kan utgöra ett hinder för att få uppehållstillstånd.
Myndigheterna överväger beviljandet av uppehållstillstånd alltid fall för fall.
Barn till föräldrar i samboförhållande
Fastställande av faderskap (Isyyden tunnustaminen)
Om ni lever i ett samboförhållande och får ett barn ska barnets far fastställas.
Om faderskapet inte fastställs är barnet officiellt faderlöst och då ansvarar modern ensam för underhåll och vård av barnet, även om ni bor tillsammans.
Faderskapet kan fastställas vid mödravården under graviditeten.
När barnet är fött kan faderskapet fastställas hos barntillsynsmannen i hemkommunen.
Faderskapet fastställs av magistratet.
När faderskapet har fastställts
kan barnet ges faderns efternamn
kan fadern vara barnets vårdnadshavare antingen tillsammans med barnets mor eller ensam.
Vårdnadshavaren (huoltaja) är den person som ansvarar för vården och uppfostran av barnet.
är fadern förpliktad att delta i underhåll av barnet
har barnet rätt att ärva sin far och släkten på sin fars sida och tvärtom
har barnet rätt till familjepension om fadern dör.
Om fadern inte erkänner sitt faderskap kan modern väcka talan för fastställande av faderskapet.
linkkiSocial- och hälsovårdsministeriet:
Erkännande och fastställande av partnerskapfinska _ svenska
Barnets efternamn vid samboende
När ett barn föds i ett samboförhållande, kan hen få
moderns efternamn eller
faderns efternamn, om faderskapet har fastställts, eller
föräldrarnas gemensamma efternamn eller
ett kombinerat efternamn som har bildats av föräldrarnas efternamn.
Om föräldrarna inte har ett gemensamt efternamn men de har gemensamma barn, får barnet samma efternamn som dess syskon har.
Du kan ansöka om ett gemensamt efternamn med din sambo
om ni har bott tillsammans minst fem år eller
Ett samboförhållande är ett förhållande där ett par lever tillsammans utan att vara gifta.
I Finland får alla par själva bestämma om de inleder ett samboförhållande, om spelreglerna i sin relation och om de gör slut på samboförhållandet.
Ett samboförhållande registreras inte någonstans.
Till skillnad från äktenskap
har sambor inte underhållsskyldighet gentemot varandra
ärver sambor inte varandra
kan den ena sambon inte få änkepension om den andra sambon dör.
Ni kan ta ett gemensamt efternamn om
ni har gemensamma barn eller
om ni har bott tillsammans minst fem år.
Om ni vill ha ett gemensamt efternamn ska ni skicka in en anmälan om namnändring till magistraten.
Om ni bor stadigvarande tillsammans i samma bostad, hör ni till samma hushåll.
Detta har betydelse om ni till exempel ansöker om bostadsbidrag från FPA.
Läs mer om bostadsbidrag för sambor på InfoFinlands sida Bostadsbidrag.
Äktenskap som ingåtts utomlands
Ett samboförhållande kan utgöra ett hinder för att få uppehållstillstånd.
Myndigheterna överväger beviljandet av uppehållstillstånd alltid fall för fall.
Barn till föräldrar i samboförhållande
Fastställande av faderskap (Isyyden tunnustaminen)
Om ni lever i ett samboförhållande och får ett barn ska barnets far fastställas.
Om faderskapet inte fastställs är barnet officiellt faderlöst och då ansvarar modern ensam för underhåll och vård av barnet, även om ni bor tillsammans.
Faderskapet kan fastställas vid mödravården under graviditeten.
När barnet är fött kan faderskapet fastställas hos barntillsynsmannen i hemkommunen.
Faderskapet fastställs av magistratet.
När faderskapet har fastställts
kan barnet ges faderns efternamn
kan fadern vara barnets vårdnadshavare antingen tillsammans med barnets mor eller ensam.
Vårdnadshavaren (huoltaja) är den person som ansvarar för vården och uppfostran av barnet.
är fadern förpliktad att delta i underhåll av barnet
har barnet rätt att ärva sin far och släkten på sin fars sida och tvärtom
har barnet rätt till familjepension om fadern dör.
Om fadern inte erkänner sitt faderskap kan modern väcka talan för fastställande av faderskapet.
linkkiSocial- och hälsovårdsministeriet:
Erkännande och fastställande av partnerskapfinska _ svenska
Barnets efternamn vid samboende
När ett barn föds i ett samboförhållande, kan hen få
moderns efternamn eller
faderns efternamn, om faderskapet har fastställts, eller
föräldrarnas gemensamma efternamn eller
ett kombinerat efternamn som har bildats av föräldrarnas efternamn.
Om föräldrarna inte har ett gemensamt efternamn men de har gemensamma barn, får barnet samma efternamn som dess syskon har.
Du kan ansöka om ett gemensamt efternamn med din sambo
om ni har bott tillsammans minst fem år eller
Om familjen har barn under 18 år och äktenskapet slutar ska föräldrarna i samband med skilsmässan komma överens om följande:
Var ska barnet bo?
Vem är barnets vårdnadshavare?
Hur ordnas umgänget?
Underhållsbidrag.
När föräldrarna har kommit överens om barnets boende, vårdnad, umgängesrätt och underhållsbidrag kan socialväsendet på orten bekräfta avtalet.
När socialväsendet bekräftar avtalet är det lika officiellt som ett domstolsbeslut.
Mer information får du vid socialbyrån i din hemkommun.
Information för föräldrar som planerar att skiljasfinska
linkkiFöreningen för ensamstående föräldrar:
Skilsmässa i Finlandengelska _ ryska _ estniska
Om ni inte kommer överens
Om ni inte kan komma överens om boende, vårdnad, umgänge och underhåll kan ni ansöka om medling i familjefrågor (perheasioiden sovittelu).
Om ni inte får fram ett avtal där heller, måste ni låta tingsrätten lösa tvisten.
Domstolen tar hänsyn till barnets intressen och dess egna önskemål.
Domstolen kan även begära en utredning av kommunens socialväsen.
Fråga om medling i familjefrågor vid socialväsendet i din hemkommun.
Mer information om juristtjänster och rättshjälp hittar du på InfoFinlands sida Behöver du en jurist?.
Boende
Låt alltid barnets intressen gå först när ni beslutar om boendet.
Officiellt kan ett barn bara bo på ett ställe.
Vid skilsmässa kommer man överens om hos vilken förälder barnet har sin officiella adress.
I praktiken kan barnet dock bo en del av tiden hos sin andra förälder.
Barnbidraget betalas till den förälder hos vilken barnet bor officiellt.
Barnets officiella adress påverkar också till exempel FPA:s bostadsbidrag.
Vårdnad
Vårdnaden om ett barn innebär
att man uppfostrar barnet
att man tar hand om och beslutar om barnets angelägenheter.
Barnets vårdnadshavare har även rätt att få information om allt som berör barnet av myndigheter.
När ett äktenskap slutar beslutar barnets föräldrar hur vårdnaden ska ordnas.
Föräldrarna kan komma överens om gemensam vårdnad eller om att den ena föräldern har ensam vårdnad.
Vårdnaden är inte beroende av vem barnet bor med.
Läs mer om gemensam och ensam vårdnad på InfoFinlands sida Familjer med en förälder.
Gemensam vårdnad och ensam vårdnadfinska
Umgängesrätt
Barnet har rätt att ha kontakt med båda sina föräldrar efter skilsmässan.
Han eller hon har också rätt att träffa den förälder som han eller hon inte bor med.
Umgängesrätten kan till exempel innebära att barnet bor hos den ena föräldern och träffar den andra föräldern vartannat veckoslut och dessutom vissa tider under loven.
Om barnet är mycket litet kan umgänget ordnas bara över dagen.
Umgängesrätten kan också vara så omfattande att barnet bor lika mycket hos båda föräldrarna.
Officiellt kan barnet dock bara ha en adress.
Låt alltid barnets intressen gå först när ni fattar beslut.
När ni skiljer er kan ni på förhand komma överens om hur ofta barnet kan träffa den förälder som bor på ett annat ställe.
Om ni vill kan ni upprätta ett skriftligt avtal om umgängesarrangemanget.
Ni kan också besluta att ni kommer separat överens om alla träffar.
Hur ordnas umgängetfinska
Om umgänget blir problematiskt
Om ni har ingått ett avtal om umgänget, men den förälder som bor med barnet inte följer avtalet kan den förälder som bor annanstans kontakta barnatillsyningsmannen i kommunen.
Barnatillsyningsmannen ordnar ett möte med föräldrarna.
Om du misstänker att barnets hälsa eller säkerhet äventyras när barnet träffar den andra föräldern ska du meddela detta till socialmyndigheter.
Om misstanken är befogad, kan det beslutas att umgänget ska ske under socialmyndigheters uppsikt.
Underhållsbidrag för barn
Båda föräldrarna bär ansvaret för underhåll av ett barn under 18 år, även om de inte bor tillsammans.
Den förälder som inte bor med barnet betalar underhållsbidrag till den förälder hos vilken barnet bor.
Läs mer om underhållsbidrag på InfoFinlands sida Familjer med en förälder.
Information för underhållsskyldigafinska
Barnets efternamn vid skilsmässa
Barnet behåller sitt tidigare efternamn när föräldrarna skiljer sig.
Efternamnet kan även bytas.
Skicka in en ansökan om namnändring till magistraten.
Om barnet har fyllt tolv år måste man få barnets skriftliga tillstånd för att byta barnets efternamn.
Det är bra att diskutera bytet av efternamn även med barn som ännu inte har fyllt tolv år.
Barnkapningar (lapsikaappaus)
Det är fråga om barnkapning när
ett barn under 16 år som är bosatt i Finland förs utomlands utan vårdnadshavarens tillstånd
ett barn som förts utomlands inte har lämnats tillbaka till Finland vid avtalad tidpunkt.
I Finland är barnkapning ett brott.
Ta kontakt med polisen på din hemort.
Mer information och råd får du från föreningen Kaapatut Lapset ry.
Internationella bortföranden av barnfinska _ svenska _ engelska _ ryska _ franska
linkkiBortförda barn rf:
Stöd och information för offer för barnkidnappningfinska _ svenska _ engelska _ turkiska _ arabiska _ tyska _ italienska
_ danska
Kontaktuppgifter till polisstationernafinska _ svenska _ engelska
Om familjen har barn under 18 år och äktenskapet slutar ska föräldrarna i samband med skilsmässan komma överens om följande:
Var ska barnet bo?
Vem är barnets vårdnadshavare?
Hur ordnas umgänget?
Underhållsbidrag.
När föräldrarna har kommit överens om barnets boende, vårdnad, umgängesrätt och underhållsbidrag kan socialväsendet på orten bekräfta avtalet.
När socialväsendet bekräftar avtalet är det lika officiellt som ett domstolsbeslut.
Mer information får du vid socialbyrån i din hemkommun.
Information för föräldrar som planerar att skiljasfinska
linkkiFöreningen för ensamstående föräldrar:
Skilsmässa i Finlandengelska _ ryska _ estniska
Om ni inte kommer överens
Om ni inte kan komma överens om boende, vårdnad, umgänge och underhåll kan ni ansöka om medling i familjefrågor (perheasioiden sovittelu).
Om ni inte får fram ett avtal där heller, måste ni låta tingsrätten lösa tvisten.
Domstolen tar hänsyn till barnets intressen och dess egna önskemål.
Domstolen kan även begära en utredning av kommunens socialväsen.
Fråga om medling i familjefrågor vid socialväsendet i din hemkommun.
Mer information om juristtjänster och rättshjälp hittar du på InfoFinlands sida Behöver du en jurist?.
Boende
Låt alltid barnets intressen gå först när ni beslutar om boendet.
Officiellt kan ett barn bara bo på ett ställe.
Vid skilsmässa kommer man överens om hos vilken förälder barnet har sin officiella adress.
I praktiken kan barnet dock bo en del av tiden hos sin andra förälder.
Barnbidraget betalas till den förälder hos vilken barnet bor officiellt.
Barnets officiella adress påverkar också till exempel FPA:s bostadsbidrag.
Vårdnad
Vårdnaden om ett barn innebär
att man uppfostrar barnet
att man tar hand om och beslutar om barnets angelägenheter.
Barnets vårdnadshavare har även rätt att få information om allt som berör barnet av myndigheter.
När ett äktenskap slutar beslutar barnets föräldrar hur vårdnaden ska ordnas.
Föräldrarna kan komma överens om gemensam vårdnad eller om att den ena föräldern har ensam vårdnad.
Vårdnaden är inte beroende av vem barnet bor med.
Läs mer om gemensam och ensam vårdnad på InfoFinlands sida Familjer med en förälder.
Gemensam vårdnad och ensam vårdnadfinska
Umgängesrätt
Barnet har rätt att ha kontakt med båda sina föräldrar efter skilsmässan.
Han eller hon har också rätt att träffa den förälder som han eller hon inte bor med.
Umgängesrätten kan till exempel innebära att barnet bor hos den ena föräldern och träffar den andra föräldern vartannat veckoslut och dessutom vissa tider under loven.
Om barnet är mycket litet kan umgänget ordnas bara över dagen.
Umgängesrätten kan också vara så omfattande att barnet bor lika mycket hos båda föräldrarna.
Officiellt kan barnet dock bara ha en adress.
Låt alltid barnets intressen gå först när ni fattar beslut.
När ni skiljer er kan ni på förhand komma överens om hur ofta barnet kan träffa den förälder som bor på ett annat ställe.
Om ni vill kan ni upprätta ett skriftligt avtal om umgängesarrangemanget.
Ni kan också besluta att ni kommer separat överens om alla träffar.
Hur ordnas umgängetfinska
Om umgänget blir problematiskt
Om ni har ingått ett avtal om umgänget, men den förälder som bor med barnet inte följer avtalet kan den förälder som bor annanstans kontakta barnatillsyningsmannen i kommunen.
Barnatillsyningsmannen ordnar ett möte med föräldrarna.
Om du misstänker att barnets hälsa eller säkerhet äventyras när barnet träffar den andra föräldern ska du meddela detta till socialmyndigheter.
Om misstanken är befogad, kan det beslutas att umgänget ska ske under socialmyndigheters uppsikt.
Underhållsbidrag för barn
Båda föräldrarna bär ansvaret för underhåll av ett barn under 18 år, även om de inte bor tillsammans.
Den förälder som inte bor med barnet betalar underhållsbidrag till den förälder hos vilken barnet bor.
Läs mer om underhållsbidrag på InfoFinlands sida Familjer med en förälder.
Information för underhållsskyldigafinska
Barnets efternamn vid skilsmässa
Barnet behåller sitt tidigare efternamn när föräldrarna skiljer sig.
Efternamnet kan även bytas.
Skicka in en ansökan om namnändring till magistraten.
Om barnet har fyllt tolv år måste man få barnets skriftliga tillstånd för att byta barnets efternamn.
Det är bra att diskutera bytet av efternamn även med barn som ännu inte har fyllt tolv år.
Barnkapningar (lapsikaappaus)
Det är fråga om barnkapning när
ett barn under 16 år som är bosatt i Finland förs utomlands utan vårdnadshavarens tillstånd
ett barn som förts utomlands inte har lämnats tillbaka till Finland vid avtalad tidpunkt.
I Finland är barnkapning ett brott.
Ta kontakt med polisen på din hemort.
Mer information och råd får du från föreningen Kaapatut Lapset ry.
Internationella bortföranden av barnfinska _ svenska _ engelska _ ryska _ franska
linkkiBortförda barn rf:
Stöd och information för offer för barnkidnappningfinska _ svenska _ engelska _ turkiska _ arabiska _ tyska _ italienska
_ danska
Kontaktuppgifter till polisstationernafinska _ svenska _ engelska
Om familjen har barn under 18 år och äktenskapet slutar ska föräldrarna i samband med skilsmässan komma överens om följande:
Var ska barnet bo?
Vem är barnets vårdnadshavare?
Hur ordnas umgänget?
Underhållsbidrag.
När föräldrarna har kommit överens om barnets boende, vårdnad, umgängesrätt och underhållsbidrag kan socialväsendet på orten bekräfta avtalet.
När socialväsendet bekräftar avtalet är det lika officiellt som ett domstolsbeslut.
Mer information får du vid socialbyrån i din hemkommun.
Information för föräldrar som planerar att skiljasfinska
linkkiFöreningen för ensamstående föräldrar:
Skilsmässa i Finlandengelska _ ryska _ estniska
Om ni inte kommer överens
Om ni inte kan komma överens om boende, vårdnad, umgänge och underhåll kan ni ansöka om medling i familjefrågor (perheasioiden sovittelu).
Om ni inte får fram ett avtal där heller, måste ni låta tingsrätten lösa tvisten.
Domstolen tar hänsyn till barnets intressen och dess egna önskemål.
Domstolen kan även begära en utredning av kommunens socialväsen.
Fråga om medling i familjefrågor vid socialväsendet i din hemkommun.
Mer information om juristtjänster och rättshjälp hittar du på InfoFinlands sida Behöver du en jurist?.
Boende
Låt alltid barnets intressen gå först när ni beslutar om boendet.
Officiellt kan ett barn bara bo på ett ställe.
Vid skilsmässa kommer man överens om hos vilken förälder barnet har sin officiella adress.
I praktiken kan barnet dock bo en del av tiden hos sin andra förälder.
Barnbidraget betalas till den förälder hos vilken barnet bor officiellt.
Barnets officiella adress påverkar också till exempel FPA:s bostadsbidrag.
Vårdnad
Vårdnaden om ett barn innebär
att man uppfostrar barnet
att man tar hand om och beslutar om barnets angelägenheter.
Barnets vårdnadshavare har även rätt att få information om allt som berör barnet av myndigheter.
När ett äktenskap slutar beslutar barnets föräldrar hur vårdnaden ska ordnas.
Föräldrarna kan komma överens om gemensam vårdnad eller om att den ena föräldern har ensam vårdnad.
Vårdnaden är inte beroende av vem barnet bor med.
Läs mer om gemensam och ensam vårdnad på InfoFinlands sida Familjer med en förälder.
Gemensam vårdnad och ensam vårdnadfinska
Umgängesrätt
Barnet har rätt att ha kontakt med båda sina föräldrar efter skilsmässan.
Han eller hon har också rätt att träffa den förälder som han eller hon inte bor med.
Umgängesrätten kan till exempel innebära att barnet bor hos den ena föräldern och träffar den andra föräldern vartannat veckoslut och dessutom vissa tider under loven.
Om barnet är mycket litet kan umgänget ordnas bara över dagen.
Umgängesrätten kan också vara så omfattande att barnet bor lika mycket hos båda föräldrarna.
Officiellt kan barnet dock bara ha en adress.
Låt alltid barnets intressen gå först när ni fattar beslut.
När ni skiljer er kan ni på förhand komma överens om hur ofta barnet kan träffa den förälder som bor på ett annat ställe.
Om ni vill kan ni upprätta ett skriftligt avtal om umgängesarrangemanget.
Ni kan också besluta att ni kommer separat överens om alla träffar.
Hur ordnas umgängetfinska
Om umgänget blir problematiskt
Om ni har ingått ett avtal om umgänget, men den förälder som bor med barnet inte följer avtalet kan den förälder som bor annanstans kontakta barnatillsyningsmannen i kommunen.
Barnatillsyningsmannen ordnar ett möte med föräldrarna.
Om du misstänker att barnets hälsa eller säkerhet äventyras när barnet träffar den andra föräldern ska du meddela detta till socialmyndigheter.
Om misstanken är befogad, kan det beslutas att umgänget ska ske under socialmyndigheters uppsikt.
Underhållsbidrag för barn
Båda föräldrarna bär ansvaret för underhåll av ett barn under 18 år, även om de inte bor tillsammans.
Den förälder som inte bor med barnet betalar underhållsbidrag till den förälder hos vilken barnet bor.
Läs mer om underhållsbidrag på InfoFinlands sida Familjer med en förälder.
Information för underhållsskyldigafinska
Barnets efternamn vid skilsmässa
Barnet behåller sitt tidigare efternamn när föräldrarna skiljer sig.
Efternamnet kan även bytas.
Skicka in en ansökan om namnändring till magistraten.
Om barnet har fyllt tolv år måste man få barnets skriftliga tillstånd för att byta barnets efternamn.
Det är bra att diskutera bytet av efternamn även med barn som ännu inte har fyllt tolv år.
Barnkapningar (lapsikaappaus)
Det är fråga om barnkapning när
ett barn under 16 år som är bosatt i Finland förs utomlands utan vårdnadshavarens tillstånd
ett barn som förts utomlands inte har lämnats tillbaka till Finland vid avtalad tidpunkt.
I Finland är barnkapning ett brott.
Ta kontakt med polisen på din hemort.
Mer information och råd får du från föreningen Kaapatut Lapset ry.
Internationella bortföranden av barnfinska _ svenska _ engelska _ ryska _ franska
linkkiBortförda barn rf:
Stöd och information för offer för barnkidnappningfinska _ svenska _ engelska _ turkiska _ arabiska _ tyska _ italienska
_ danska
Kontaktuppgifter till polisstationernafinska _ svenska _ engelska
När äktenskapet slutar kan ni gemensamt komma överens om hur ni delar egendomen.
Ni kan även tillsammans besluta vem av er som tillsvidare ska bo kvar i det gemensamma hemmet.
Hjälp med att dela egendomen
Om ni inte kan komma överens om hur ni ska dela upp egendomen, kan vem som helst av makarna kräva egendomsfördelning, det vill säga bodelning (ositus).
Bodelningen kan göras direkt när man har lämnat in den första skilsmässoansökan.
Man behöver alltså inte vänta tills betänketiden på sex månader har gått ut.
När ni kräver bodelning förordnar tingsrätten en bodelningsman som delar egendomen.
Bodelningsmannen tar betalt för arbetet.
När bodelningen inleds ska man utreda hur mycket egendom och skulder vardera maka har.
På webbplatsen för Suomen lakiopas får du information om vilka handlingar du behöver för bodelningen.
Mer information om bodelningen får du på justitieministeriets webbplats.
Delas egendomen jämnt eller inte?
Vanligtvis delas egendomen vid skilsmässa jämnt mellan makarna.
I undantagsfall delas egendomen inte jämnt.
Då kan bodelningen jämkas.
Detta betyder att man i situationen beaktar vad som är rimligt.
Om äktenskapet till exempel har varat under fem år delas egendomen inte nödvändigtvis jämnt.
Bodelningen kan jämkas endast om någon av makarna separat kräver det.
Om ni har skrivit äktenskapsförord påverkar detta avtal egendomsfördelningen.
Mer information om äktenskapsförord får du på InfoFinlands sida Äktenskapsförord.
Bodelning mellan makarfinska _ svenska _ engelska
När äktenskapet slutar kan ni gemensamt komma överens om hur ni delar egendomen.
Ni kan även tillsammans besluta vem av er som tillsvidare ska bo kvar i det gemensamma hemmet.
Hjälp med att dela egendomen
Om ni inte kan komma överens om hur ni ska dela upp egendomen, kan vem som helst av makarna kräva egendomsfördelning, det vill säga bodelning (ositus).
Bodelningen kan göras direkt när man har lämnat in den första skilsmässoansökan.
Man behöver alltså inte vänta tills betänketiden på sex månader har gått ut.
När ni kräver bodelning förordnar tingsrätten en bodelningsman som delar egendomen.
Bodelningsmannen tar betalt för arbetet.
När bodelningen inleds ska man utreda hur mycket egendom och skulder vardera maka har.
På webbplatsen för Suomen lakiopas får du information om vilka handlingar du behöver för bodelningen.
Mer information om bodelningen får du på justitieministeriets webbplats.
Delas egendomen jämnt eller inte?
Vanligtvis delas egendomen vid skilsmässa jämnt mellan makarna.
I undantagsfall delas egendomen inte jämnt.
Då kan bodelningen jämkas.
Detta betyder att man i situationen beaktar vad som är rimligt.
Om äktenskapet till exempel har varat under fem år delas egendomen inte nödvändigtvis jämnt.
Bodelningen kan jämkas endast om någon av makarna separat kräver det.
Om ni har skrivit äktenskapsförord påverkar detta avtal egendomsfördelningen.
Mer information om äktenskapsförord får du på InfoFinlands sida Äktenskapsförord.
Bodelning mellan makarfinska _ svenska _ engelska
När äktenskapet slutar kan ni gemensamt komma överens om hur ni delar egendomen.
Ni kan även tillsammans besluta vem av er som tillsvidare ska bo kvar i det gemensamma hemmet.
Hjälp med att dela egendomen
Om ni inte kan komma överens om hur ni ska dela upp egendomen, kan vem som helst av makarna kräva egendomsfördelning, det vill säga bodelning (ositus).
Bodelningen kan göras direkt när man har lämnat in den första skilsmässoansökan.
Man behöver alltså inte vänta tills betänketiden på sex månader har gått ut.
När ni kräver bodelning förordnar tingsrätten en bodelningsman som delar egendomen.
Bodelningsmannen tar betalt för arbetet.
När bodelningen inleds ska man utreda hur mycket egendom och skulder vardera maka har.
På webbplatsen för Suomen lakiopas får du information om vilka handlingar du behöver för bodelningen.
Mer information om bodelningen får du på justitieministeriets webbplats.
Delas egendomen jämnt eller inte?
Vanligtvis delas egendomen vid skilsmässa jämnt mellan makarna.
I undantagsfall delas egendomen inte jämnt.
Då kan bodelningen jämkas.
Detta betyder att man i situationen beaktar vad som är rimligt.
Om äktenskapet till exempel har varat under fem år delas egendomen inte nödvändigtvis jämnt.
Bodelningen kan jämkas endast om någon av makarna separat kräver det.
Om ni har skrivit äktenskapsförord påverkar detta avtal egendomsfördelningen.
Mer information om äktenskapsförord får du på InfoFinlands sida Äktenskapsförord.
Bodelning mellan makarfinska _ svenska _ engelska
Om du eller din maka/make har hemort i Finland kan du ansöka om skilsmässa enligt Finlands lag.
Det finns även vissa andra fall där du kan ansöka om skilsmässa enligt Finlands lag.
Om skilsmässa stadgas i äktenskapslagen.
Att ansöka om skilsmässa
Skilsmässa kan sökas av den ena eller av båda makarna tillsammans.
Du kan ansöka om skilsmässa ensam även om din maka eller make inte vill skiljas.
Man ansöker om skilsmässa i tingsrätten.
Domstolen undersöker inte varför man ansöker om skilsmässa.
Inte heller relationen mellan makarna undersöks.
Man ansöker om skilsmässa med en skriftlig ansökan.
Du kan lämna in skilsmässoansökan i tingsrätten i din egen eller din maka/makes hemkommun.
Du kan även skicka in ansökan till tingsrättens kansli per post, som telegram eller via e-post.
Du hittar skilsmässoansökan på tjänsten suomi.fi.
Ansökan om skilsmässa görs i två steg.
Först lämnar man in skilsmässoansökan.
Efter betänketiden fullföljer man sin ansökan med en ny ansökan.
Domstolen dömer till skilsmässa först efter att den andra ansökan har lämnats in.
Parterna döms till skilsmässa även om den andra parten motsätter sig det.
Mer information om att ansöka om skilsmässa hittar du på justitieministeriets webbplats.
Äktenskapslagenfinska _ svenska _ engelska
Skilsmässoansökan(pdf, 100 kb)finska _ svenska
linkkiRättsväsendet:
Att ansöka om skilsmässafinska _ svenska _ engelska
linkkiFöreningen för ensamstående föräldrar:
Skilsmässa i Finlandengelska _ ryska _ estniska
Betänketid
När den första ansökan om skilsmässa har lämnats in börjar en sex månader lång betänketid.
Betänketiden är obligatorisk, förutom om du och din maka/make har bott på skilda adresser de senaste två åren.
Om du och din maka/make ansöker om skilsmässa tillsammans, börjar betänketiden direkt när er gemensamma ansökan har kommit in hos tingsrätten.
Om en av makarna ensam ansöker om skilsmässa, börjar betänketiden från den dag då ansökan delges den andra makan.
Tingsrätten ser till att ansökan delges den andra makan.
Efter betänketiden
Tingsrätten dömer makarna till skilsmässa när
betänketiden på sex månader har gått ut och
när den ena makan eller båda makarna tillsammans kräver att de ska dömas till skilsmässa.
Kravet om att äktenskapet ska dömas till skilsmässa efter betänketiden görs likadant som den första ansökan.
Det är viktigt att lämna in den andra ansökan om skilsmässa inom ett år efter att betänketiden började.
I annat fall förfaller ärendet.
Skilsmässa utan betänketid
Om du och din maka/make har bott på skilda adresser utan avbrott de senaste två åren innan ni ansöker om skilsmässa behövs ingen betänktetid.
Då kan domstolen döma till skilsmässa direkt.
Medling i familjefrågor
När ni överväger skilsmässa och behöver hjälp med att komma överens om saker och ting, kan ni ansöka om medling i familjefrågor (perheasioiden sovittelu).
Medling kan ofta vara nyttig och hjälpa er att komma överens i olika frågor utan rättegång.
Man kan till exempel prata om barnens situation i medlingen.
Medlaren är oftast en anställd vid socialbyrån, barnrådgivningen eller familjerådgivningen.
Du kan diskutera med dem konfidentiellt.
Fråga socialbyrån i din hemkommun hur medling i familjefrågor ordnas i din hemkommun.
Mer information om medling i familjefrågor får du på justitieministeriets webbplats.
Stöd under skilsmässan
Vid problem i parförhållandet kan du söka hjälp till exempel vid familjerådgivningen eller hälsovårdscentralen i din hemkommun.
Mer information får du på InfoFinlands sida Problem i äktenskap eller parförhållande.
I våldssituationer får du mer information på InfoFinlands sida Våld.
Många organisationer och församlingar ordnar stödgruppsverksamhet för personer som har skilt sig.
Mer information får du till exempel på Väestöliittos webbplats eller webbplatsen för kyrkans familjerådgivningscentral.
På webbplatsen för föreningen för familjer med en förälder, Yhden Vanhemman Perheiden Liitto ry, finns information och råd för föräldrar som överväger skilsmässa.
Miessakit rf strävar efter att sörja för mäns välbefinnande och erbjuder sociala aktiviteter och stöd.
Föreningen har verksamhet i Helsingfors, Tammerfors och Lahtis.
Du hittar mer information på föreningens webbplats på finska, svenska och engelska.
linkkiEvangelisk-lutherska kyrkan i Finland:
Information om kyrkans familjerådgivningfinska _ svenska
Stöd för mänfinska _ svenska _ engelska
linkkiDuo För bikulturella familjer:
Skilsmässa i ett bikulturellt äktenskapengelska
Efternamn vid skilsmässa
Om ditt äktenskap slutar med skilsmässa, ändras inte ditt efternamn.
Om du vill kan du ta ett annat efternamn.
Du kan till exempel ta vilket som helst namn som du har haft tidigare.
Skicka in en ansökan om namnändring till magistraten.
Skilsmässa och uppehållstillstånd
Om du har ett tidsbegränsat uppehållstillstånd som beviljats på grund av familjeband, kan skilsmässan inverka på uppehållstillståndet.
I sådana situationer avvägs alltid fall till fall om uppehållstillståndet förlängs efter skilsmässan eller om det återkallas.
Mer information får du på InfoFinlands sida Problem med uppehållstillståndet.
Egendom vid skilsmässa
Information om egendomsfördelning vid skilsmässa finns på InfoFinlands sida Egendom vid skilsmässa.
Barn vid skilsmässa
Mer information om barn vid skilsmässa finns på InfoFinlands sida Barn vid skilsmässa.
Om du eller din maka/make har hemort i Finland kan du ansöka om skilsmässa enligt Finlands lag.
Det finns även vissa andra fall där du kan ansöka om skilsmässa enligt Finlands lag.
Om skilsmässa stadgas i äktenskapslagen.
Att ansöka om skilsmässa
Skilsmässa kan sökas av den ena eller av båda makarna tillsammans.
Du kan ansöka om skilsmässa ensam även om din maka eller make inte vill skiljas.
Man ansöker om skilsmässa i tingsrätten.
Domstolen undersöker inte varför man ansöker om skilsmässa.
Inte heller relationen mellan makarna undersöks.
Man ansöker om skilsmässa med en skriftlig ansökan.
Du kan lämna in skilsmässoansökan i tingsrätten i din egen eller din maka/makes hemkommun.
Du kan även skicka in ansökan till tingsrättens kansli per post, som telegram eller via e-post.
Du hittar skilsmässoansökan på tjänsten suomi.fi.
Ansökan om skilsmässa görs i två steg.
Först lämnar man in skilsmässoansökan.
Efter betänketiden fullföljer man sin ansökan med en ny ansökan.
Domstolen dömer till skilsmässa först efter att den andra ansökan har lämnats in.
Parterna döms till skilsmässa även om den andra parten motsätter sig det.
Mer information om att ansöka om skilsmässa hittar du på justitieministeriets webbplats.
Äktenskapslagenfinska _ svenska _ engelska
Skilsmässoansökan(pdf, 100 kb)finska _ svenska
linkkiRättsväsendet:
Att ansöka om skilsmässafinska _ svenska _ engelska
linkkiFöreningen för ensamstående föräldrar:
Skilsmässa i Finlandengelska _ ryska _ estniska
Betänketid
När den första ansökan om skilsmässa har lämnats in börjar en sex månader lång betänketid.
Betänketiden är obligatorisk, förutom om du och din maka/make har bott på skilda adresser de senaste två åren.
Om du och din maka/make ansöker om skilsmässa tillsammans, börjar betänketiden direkt när er gemensamma ansökan har kommit in hos tingsrätten.
Om en av makarna ensam ansöker om skilsmässa, börjar betänketiden från den dag då ansökan delges den andra makan.
Tingsrätten ser till att ansökan delges den andra makan.
Efter betänketiden
Tingsrätten dömer makarna till skilsmässa när
betänketiden på sex månader har gått ut och
när den ena makan eller båda makarna tillsammans kräver att de ska dömas till skilsmässa.
Kravet om att äktenskapet ska dömas till skilsmässa efter betänketiden görs likadant som den första ansökan.
Det är viktigt att lämna in den andra ansökan om skilsmässa inom ett år efter att betänketiden började.
I annat fall förfaller ärendet.
Skilsmässa utan betänketid
Om du och din maka/make har bott på skilda adresser utan avbrott de senaste två åren innan ni ansöker om skilsmässa behövs ingen betänktetid.
Då kan domstolen döma till skilsmässa direkt.
Medling i familjefrågor
När ni överväger skilsmässa och behöver hjälp med att komma överens om saker och ting, kan ni ansöka om medling i familjefrågor (perheasioiden sovittelu).
Medling kan ofta vara nyttig och hjälpa er att komma överens i olika frågor utan rättegång.
Man kan till exempel prata om barnens situation i medlingen.
Medlaren är oftast en anställd vid socialbyrån, barnrådgivningen eller familjerådgivningen.
Du kan diskutera med dem konfidentiellt.
Fråga socialbyrån i din hemkommun hur medling i familjefrågor ordnas i din hemkommun.
Mer information om medling i familjefrågor får du på justitieministeriets webbplats.
Stöd under skilsmässan
Vid problem i parförhållandet kan du söka hjälp till exempel vid familjerådgivningen eller hälsovårdscentralen i din hemkommun.
Mer information får du på InfoFinlands sida Problem i äktenskap eller parförhållande.
I våldssituationer får du mer information på InfoFinlands sida Våld.
Många organisationer och församlingar ordnar stödgruppsverksamhet för personer som har skilt sig.
Mer information får du till exempel på Väestöliittos webbplats eller webbplatsen för kyrkans familjerådgivningscentral.
På webbplatsen för föreningen för familjer med en förälder, Yhden Vanhemman Perheiden Liitto ry, finns information och råd för föräldrar som överväger skilsmässa.
Miessakit rf strävar efter att sörja för mäns välbefinnande och erbjuder sociala aktiviteter och stöd.
Föreningen har verksamhet i Helsingfors, Tammerfors och Lahtis.
Du hittar mer information på föreningens webbplats på finska, svenska och engelska.
linkkiEvangelisk-lutherska kyrkan i Finland:
Information om kyrkans familjerådgivningfinska _ svenska
Stöd för mänfinska _ svenska _ engelska
linkkiDuo För bikulturella familjer:
Skilsmässa i ett bikulturellt äktenskapengelska
Efternamn vid skilsmässa
Om ditt äktenskap slutar med skilsmässa, ändras inte ditt efternamn.
Om du vill kan du ta ett annat efternamn.
Du kan till exempel ta vilket som helst namn som du har haft tidigare.
Skicka in en ansökan om namnändring till magistraten.
Skilsmässa och uppehållstillstånd
Om du har ett tidsbegränsat uppehållstillstånd som beviljats på grund av familjeband, kan skilsmässan inverka på uppehållstillståndet.
I sådana situationer avvägs alltid fall till fall om uppehållstillståndet förlängs efter skilsmässan eller om det återkallas.
Mer information får du på InfoFinlands sida Problem med uppehållstillståndet.
Egendom vid skilsmässa
Information om egendomsfördelning vid skilsmässa finns på InfoFinlands sida Egendom vid skilsmässa.
Barn vid skilsmässa
Mer information om barn vid skilsmässa finns på InfoFinlands sida Barn vid skilsmässa.
Om du eller din maka/make har hemort i Finland kan du ansöka om skilsmässa enligt Finlands lag.
Det finns även vissa andra fall där du kan ansöka om skilsmässa enligt Finlands lag.
Om skilsmässa stadgas i äktenskapslagen.
Att ansöka om skilsmässa
Skilsmässa kan sökas av den ena eller av båda makarna tillsammans.
Du kan ansöka om skilsmässa ensam även om din maka eller make inte vill skiljas.
Man ansöker om skilsmässa i tingsrätten.
Domstolen undersöker inte varför man ansöker om skilsmässa.
Inte heller relationen mellan makarna undersöks.
Man ansöker om skilsmässa med en skriftlig ansökan.
Du kan lämna in skilsmässoansökan i tingsrätten i din egen eller din maka/makes hemkommun.
Du kan även skicka in ansökan till tingsrättens kansli per post, som telegram eller via e-post.
Du hittar skilsmässoansökan på tjänsten suomi.fi.
Ansökan om skilsmässa görs i två steg.
Först lämnar man in skilsmässoansökan.
Efter betänketiden fullföljer man sin ansökan med en ny ansökan.
Domstolen dömer till skilsmässa först efter att den andra ansökan har lämnats in.
Parterna döms till skilsmässa även om den andra parten motsätter sig det.
Mer information om att ansöka om skilsmässa hittar du på justitieministeriets webbplats.
Äktenskapslagenfinska _ svenska _ engelska
Skilsmässoansökan(pdf, 100 kb)finska _ svenska
linkkiRättsväsendet:
Att ansöka om skilsmässafinska _ svenska _ engelska
linkkiFöreningen för ensamstående föräldrar:
Skilsmässa i Finlandengelska _ ryska _ estniska
Betänketid
När den första ansökan om skilsmässa har lämnats in börjar en sex månader lång betänketid.
Betänketiden är obligatorisk, förutom om du och din maka/make har bott på skilda adresser de senaste två åren.
Om du och din maka/make ansöker om skilsmässa tillsammans, börjar betänketiden direkt när er gemensamma ansökan har kommit in hos tingsrätten.
Om en av makarna ensam ansöker om skilsmässa, börjar betänketiden från den dag då ansökan delges den andra makan.
Tingsrätten ser till att ansökan delges den andra makan.
Efter betänketiden
Tingsrätten dömer makarna till skilsmässa när
betänketiden på sex månader har gått ut och
när den ena makan eller båda makarna tillsammans kräver att de ska dömas till skilsmässa.
Kravet om att äktenskapet ska dömas till skilsmässa efter betänketiden görs likadant som den första ansökan.
Det är viktigt att lämna in den andra ansökan om skilsmässa inom ett år efter att betänketiden började.
I annat fall förfaller ärendet.
Skilsmässa utan betänketid
Om du och din maka/make har bott på skilda adresser utan avbrott de senaste två åren innan ni ansöker om skilsmässa behövs ingen betänktetid.
Då kan domstolen döma till skilsmässa direkt.
Medling i familjefrågor
När ni överväger skilsmässa och behöver hjälp med att komma överens om saker och ting, kan ni ansöka om medling i familjefrågor (perheasioiden sovittelu).
Medling kan ofta vara nyttig och hjälpa er att komma överens i olika frågor utan rättegång.
Man kan till exempel prata om barnens situation i medlingen.
Medlaren är oftast en anställd vid socialbyrån, barnrådgivningen eller familjerådgivningen.
Du kan diskutera med dem konfidentiellt.
Fråga socialbyrån i din hemkommun hur medling i familjefrågor ordnas i din hemkommun.
Mer information om medling i familjefrågor får du på justitieministeriets webbplats.
Stöd under skilsmässan
Vid problem i parförhållandet kan du söka hjälp till exempel vid familjerådgivningen eller hälsovårdscentralen i din hemkommun.
Mer information får du på InfoFinlands sida Problem i äktenskap eller parförhållande.
I våldssituationer får du mer information på InfoFinlands sida Våld.
Många organisationer och församlingar ordnar stödgruppsverksamhet för personer som har skilt sig.
Mer information får du till exempel på Väestöliittos webbplats eller webbplatsen för kyrkans familjerådgivningscentral.
På webbplatsen för föreningen för familjer med en förälder, Yhden Vanhemman Perheiden Liitto ry, finns information och råd för föräldrar som överväger skilsmässa.
Miessakit rf strävar efter att sörja för mäns välbefinnande och erbjuder sociala aktiviteter och stöd.
Föreningen har verksamhet i Helsingfors, Tammerfors och Lahtis.
Du hittar mer information på föreningens webbplats på finska, svenska och engelska.
linkkiEvangelisk-lutherska kyrkan i Finland:
Information om kyrkans familjerådgivningfinska _ svenska
Stöd för mänfinska _ svenska _ engelska
linkkiDuo För bikulturella familjer:
Skilsmässa i ett bikulturellt äktenskapengelska
Efternamn vid skilsmässa
Om ditt äktenskap slutar med skilsmässa, ändras inte ditt efternamn.
Om du vill kan du ta ett annat efternamn.
Du kan till exempel ta vilket som helst namn som du har haft tidigare.
Skicka in en ansökan om namnändring till magistraten.
Skilsmässa och uppehållstillstånd
Om du har ett tidsbegränsat uppehållstillstånd som beviljats på grund av familjeband, kan skilsmässan inverka på uppehållstillståndet.
I sådana situationer avvägs alltid fall till fall om uppehållstillståndet förlängs efter skilsmässan eller om det återkallas.
Mer information får du på InfoFinlands sida Problem med uppehållstillståndet.
Egendom vid skilsmässa
Information om egendomsfördelning vid skilsmässa finns på InfoFinlands sida Egendom vid skilsmässa.
Barn vid skilsmässa
Mer information om barn vid skilsmässa finns på InfoFinlands sida Barn vid skilsmässa.
Äkta makar är sinsemellan likvärdiga.
De bör i äktenskapet visa varandra förtroende och i samråd verka för familjens bästa.
Vardera maken har rätt att själv besluta om sitt deltagande i förvärvsarbete samt i samhällelig och annan verksamhet utanför familjen.
Läs mer om föräldrarnas skyldigheter gentemot sina barn på InfoFinlands sida Fostran av barn i Finland.
Makarnas underhållsskyldighet
Vardera maken ska efter förmåga bidra till familjens gemensamma hushåll och makarnas underhåll.
Om den ena maken inte förvärvsarbetar ska den förmögnare maken stå för kostnader för till exempel mat och kläder.
Barn i äktenskapet
När en gift kvinna får ett barn registreras kvinnans make automatiskt som barnets far i befolkningsregistret.
Båda föräldrarna registreras som barnets vårdnadshavare.
Gifta par kan adoptera barn tillsammans.
Om du är intresserad av adoption, fråga om råd vid socialbyrån i din hemkommun.
Egendom
Den egendom som maken har vid ingående av äktenskap eller förvärvar under äktenskapet förblir hans tillhörighet.
Makarna kan också förvärva egendom som de äger tillsammans.
Makar har giftorätt till varandras egendom.
Om äktenskapet slutar i skilsmässa delas makarnas sammanlagda egendom jämnt mellan makarna.
Om äktenskapet slutar med att en av makarna dör, delas makarnas sammanlagda egendom mellan arvingarna till den avlidna makan och den maka som fortfarande lever.
Giftorätten kan inte upphävas med testamente.
Om makarna har upprättat ett äktenskapsförord delas egendomen vid skilsmässa eller när den ena makan avlider i enlighet med det. Om makarna har upprättat ett äktenskapsförord delas egendomen i enlighet med det.
Läs mer på InfoFinlands sida Ingående av äktenskap i Finland, komihåglista och Äktenskapsförord.
Skulder
Vardera maken ansvarar ensam för den skuld som de har tagit före äktenskapet eller under det.
Om den ena maken har tagit lån för att försörja familjen, till exempel för att köpa mat, ansvarar båda makarna för denna skuld.
Om makarna vill, kan de åta sig gemensamma skulder. Då måste de också återbetala skulderna tillsammans.
Gemensam bostad
Den ena maken kan inte utan den andra makens tillstånd sälja familjens gemensamma bostad eller tillhörande lös egendom, såsom möbler.
Problem i äktenskapet?
Om du har problem i parförhållandet kan du söka hjälp vid till exempel familjerådgivningen eller hälsovårdscentralen i din hemkommun.
Mer information får du på InfoFinlands sida Problem i äktenskap eller parförhållande.
På InfoFinlands sida Våld hittar du information om vad du kan göra om din partner utövar våld eller hotar med våld.
Många organisationer och församlingar ordnar stödgruppsverksamhet för personer som har skilt sig.
Mer information får du till exempel på Väestöliittos webbplats eller webbplatsen för kyrkans familjerådgivningscentral.
Ibland kan ett äktenskap sluta med skilsmässa.
Läs mer på InfoFinlands sida Skilsmässa.
linkkiEvangelisk-lutherska kyrkan i Finland:
Information om kyrkans familjerådgivningfinska _ svenska
Stöd vid skilsmässafinska
En familjemedlems död
Vad ska man göra och var får man hjälp när en familjemedlem dör?
Läs mer på InfoFinlands sida Dödsfall.
Äkta makar är sinsemellan likvärdiga.
De bör i äktenskapet visa varandra förtroende och i samråd verka för familjens bästa.
Vardera maken har rätt att själv besluta om sitt deltagande i förvärvsarbete samt i samhällelig och annan verksamhet utanför familjen.
Läs mer om föräldrarnas skyldigheter gentemot sina barn på InfoFinlands sida Fostran av barn i Finland.
Makarnas underhållsskyldighet
Vardera maken ska efter förmåga bidra till familjens gemensamma hushåll och makarnas underhåll.
Om den ena maken inte förvärvsarbetar ska den förmögnare maken stå för kostnader för till exempel mat och kläder.
Barn i äktenskapet
När en gift kvinna får ett barn registreras kvinnans make automatiskt som barnets far i befolkningsregistret.
Båda föräldrarna registreras som barnets vårdnadshavare.
Gifta par kan adoptera barn tillsammans.
Om du är intresserad av adoption, fråga om råd vid socialbyrån i din hemkommun.
Egendom
Den egendom som maken har vid ingående av äktenskap eller förvärvar under äktenskapet förblir hans tillhörighet.
Makarna kan också förvärva egendom som de äger tillsammans.
Makar har giftorätt till varandras egendom.
Om äktenskapet slutar i skilsmässa delas makarnas sammanlagda egendom jämnt mellan makarna.
Om äktenskapet slutar med att en av makarna dör, delas makarnas sammanlagda egendom mellan arvingarna till den avlidna makan och den maka som fortfarande lever.
Giftorätten kan inte upphävas med testamente.
Om makarna har upprättat ett äktenskapsförord delas egendomen vid skilsmässa eller när den ena makan avlider i enlighet med det. Om makarna har upprättat ett äktenskapsförord delas egendomen i enlighet med det.
Läs mer på InfoFinlands sida Ingående av äktenskap i Finland, komihåglista och Äktenskapsförord.
Skulder
Vardera maken ansvarar ensam för den skuld som de har tagit före äktenskapet eller under det.
Om den ena maken har tagit lån för att försörja familjen, till exempel för att köpa mat, ansvarar båda makarna för denna skuld.
Om makarna vill, kan de åta sig gemensamma skulder. Då måste de också återbetala skulderna tillsammans.
Gemensam bostad
Den ena maken kan inte utan den andra makens tillstånd sälja familjens gemensamma bostad eller tillhörande lös egendom, såsom möbler.
Problem i äktenskapet?
Om du har problem i parförhållandet kan du söka hjälp vid till exempel familjerådgivningen eller hälsovårdscentralen i din hemkommun.
Mer information får du på InfoFinlands sida Problem i äktenskap eller parförhållande.
På InfoFinlands sida Våld hittar du information om vad du kan göra om din partner utövar våld eller hotar med våld.
Många organisationer och församlingar ordnar stödgruppsverksamhet för personer som har skilt sig.
Mer information får du till exempel på Väestöliittos webbplats eller webbplatsen för kyrkans familjerådgivningscentral.
Ibland kan ett äktenskap sluta med skilsmässa.
Läs mer på InfoFinlands sida Skilsmässa.
linkkiEvangelisk-lutherska kyrkan i Finland:
Information om kyrkans familjerådgivningfinska _ svenska
Stöd vid skilsmässafinska
En familjemedlems död
Vad ska man göra och var får man hjälp när en familjemedlem dör?
Läs mer på InfoFinlands sida Dödsfall.
Äkta makar är sinsemellan likvärdiga.
De bör i äktenskapet visa varandra förtroende och i samråd verka för familjens bästa.
Vardera maken har rätt att själv besluta om sitt deltagande i förvärvsarbete samt i samhällelig och annan verksamhet utanför familjen.
Läs mer om föräldrarnas skyldigheter gentemot sina barn på InfoFinlands sida Fostran av barn i Finland.
Makarnas underhållsskyldighet
Vardera maken ska efter förmåga bidra till familjens gemensamma hushåll och makarnas underhåll.
Om den ena maken inte förvärvsarbetar ska den förmögnare maken stå för kostnader för till exempel mat och kläder.
Barn i äktenskapet
När en gift kvinna får ett barn registreras kvinnans make automatiskt som barnets far i befolkningsregistret.
Båda föräldrarna registreras som barnets vårdnadshavare.
Gifta par kan adoptera barn tillsammans.
Om du är intresserad av adoption, fråga om råd vid socialbyrån i din hemkommun.
Egendom
Den egendom som maken har vid ingående av äktenskap eller förvärvar under äktenskapet förblir hans tillhörighet.
Makarna kan också förvärva egendom som de äger tillsammans.
Makar har giftorätt till varandras egendom.
Om äktenskapet slutar i skilsmässa delas makarnas sammanlagda egendom jämnt mellan makarna.
Om äktenskapet slutar med att en av makarna dör, delas makarnas sammanlagda egendom mellan arvingarna till den avlidna makan och den maka som fortfarande lever.
Giftorätten kan inte upphävas med testamente.
Om makarna har upprättat ett äktenskapsförord delas egendomen vid skilsmässa eller när den ena makan avlider i enlighet med det. Om makarna har upprättat ett äktenskapsförord delas egendomen i enlighet med det.
Läs mer på InfoFinlands sida Ingående av äktenskap i Finland, komihåglista och Äktenskapsförord.
Skulder
Vardera maken ansvarar ensam för den skuld som de har tagit före äktenskapet eller under det.
Om den ena maken har tagit lån för att försörja familjen, till exempel för att köpa mat, ansvarar båda makarna för denna skuld.
Om makarna vill, kan de åta sig gemensamma skulder. Då måste de också återbetala skulderna tillsammans.
Gemensam bostad
Den ena maken kan inte utan den andra makens tillstånd sälja familjens gemensamma bostad eller tillhörande lös egendom, såsom möbler.
Problem i äktenskapet?
Om du har problem i parförhållandet kan du söka hjälp vid till exempel familjerådgivningen eller hälsovårdscentralen i din hemkommun.
Mer information får du på InfoFinlands sida Problem i äktenskap eller parförhållande.
På InfoFinlands sida Våld hittar du information om vad du kan göra om din partner utövar våld eller hotar med våld.
Många organisationer och församlingar ordnar stödgruppsverksamhet för personer som har skilt sig.
Mer information får du till exempel på Väestöliittos webbplats eller webbplatsen för kyrkans familjerådgivningscentral.
Ibland kan ett äktenskap sluta med skilsmässa.
Läs mer på InfoFinlands sida Skilsmässa.
linkkiEvangelisk-lutherska kyrkan i Finland:
Information om kyrkans familjerådgivningfinska _ svenska
Stöd vid skilsmässafinska
En familjemedlems död
Vad ska man göra och var får man hjälp när en familjemedlem dör?
Läs mer på InfoFinlands sida Dödsfall.
Vigseln kan förrättas
som en kyrklig vigsel.
Personerna som ska gifta sig ska båda vara närvarande vid vigseln.
Dessutom måste minst två vittnen vara närvarande.
Civilvigsel
Civilvigsel kan enligt lag förrättas av en häradsskrivare som arbetar vid magistraten (maistraatti) eller en lagman eller tingsdomare som arbetar i tingsrätten (käräjäoikeus).
Boka vigseltiden i magistraten eller tingsrätten i god tid för bröllopsdagen.
Civilvigseln är avgiftsfri om den förrättas i magistraten eller tingsrätten under tjänstetid.
På separat överenskommelse kan vigseln också förrättas någon annanstans, till exempel hemma eller i en festlokal.
Var och en har rätt till civilvigsel, också de som tillhör något religionssamfund.
Grundläggande information om vigseln finns på magistratens webbplats.
Vigselfinska _ svenska _ engelska
Kontaktuppgifter till magistratfinska _ svenska _ engelska
linkkiRättsväsendet:
Kontaktuppgifter till tingsrättfinska _ svenska _ engelska
Kyrklig vigsel
Kyrklig vigsel kan förrättas i
evangelisk-lutherska kyrkan (evankelis-luterilainen kirkko)
ortodoxa kyrkan (ortodoksinen kirkko) eller
i något annat religiöst samfund som är registrerat i Finland.
Varje religiöst samfund bestämmer själv vilka villkor som gäller för vigseln och hurudan vigselceremonin är.
Om makarna inte bekänner sig till samma religion förrättas vigseln i magistraten och äktenskapet kan välsignas i kyrkan.
I den lutherska kyrkan kan medlemmar i kristna religionssamfund, till exempel en lutheran och en ortodox, vigas.
linkkiEvangelisk-lutherska kyrkan:
Information om äktenskapfinska _ svenska _ engelska
linkkiFinska ortodoxa kyrkan:
Finska ortodoxa kyrkanfinska _ svenska _ ryska
linkkiFritänkarförbundet r.f.:
Registrerade religiösa samfund med vigselrättfinska
Utländska medborgare
I magistraten vigs även utländska medborgare.
I Finland görs alltid en hindersprövning innan äktenskapet ingås.
Läs mer på InfoFinlands sida Prövning av hinder mot äktenskap.
Inverkan på uppehållstillstånd och medborgarskap
Maken, makan, sambon eller den registrerade partnern till en finsk eller en utländsk medborgare som är bosatt i Finland kan få ett uppehållstillstånd i Finland.
De kan få ett permanent uppehållstillstånd när äktenskapet har varat fem år.
Läs mer på InfoFinlands sida Uppehållstillstånd för make eller maka.
Finskt medborgarskap kan inte fås via äktenskap.
Äktenskap som ingåtts utomlands ska registreras i magistraten
Ett äktenskap som ingåtts utomlands är officiellt i Finland först när det registrerats i Finland.
Om äktenskapet har ingåtts utomlands måste man uppvisa ett legaliserat och översatt vigselintyg i magistraten för registrering.
Finska medborgare som är bosatta utomlands kan också skicka vigselhandlingarna till den lokala finska beskickningen som skickar handlingarna till magistraten i Finland.
Om personer som är bosatta i Finland antecknas grundläggande uppgifter i befolkningsdatasystemet.
Uppgifter som registreras är bland annat namn, födelsedatum, medborgarskap, familjeförhållanden och adress.
Utlänningar ska enligt lag anmäla till registret samma uppgifter som finska medborgare om deras vistelse i Finland varar över ett år.
Blanketten för registrering av ett äktenskap som ingåtts utomlandsfinska _ engelska
Vigseln kan förrättas
som en kyrklig vigsel.
Personerna som ska gifta sig ska båda vara närvarande vid vigseln.
Dessutom måste minst två vittnen vara närvarande.
Civilvigsel
Civilvigsel kan enligt lag förrättas av en häradsskrivare som arbetar vid magistraten (maistraatti) eller en lagman eller tingsdomare som arbetar i tingsrätten (käräjäoikeus).
Boka vigseltiden i magistraten eller tingsrätten i god tid för bröllopsdagen.
Civilvigseln är avgiftsfri om den förrättas i magistraten eller tingsrätten under tjänstetid.
På separat överenskommelse kan vigseln också förrättas någon annanstans, till exempel hemma eller i en festlokal.
Var och en har rätt till civilvigsel, också de som tillhör något religionssamfund.
Grundläggande information om vigseln finns på magistratens webbplats.
Vigselfinska _ svenska _ engelska
Kontaktuppgifter till magistratfinska _ svenska _ engelska
linkkiRättsväsendet:
Kontaktuppgifter till tingsrättfinska _ svenska _ engelska
Kyrklig vigsel
Kyrklig vigsel kan förrättas i
evangelisk-lutherska kyrkan (evankelis-luterilainen kirkko)
ortodoxa kyrkan (ortodoksinen kirkko) eller
i något annat religiöst samfund som är registrerat i Finland.
Varje religiöst samfund bestämmer själv vilka villkor som gäller för vigseln och hurudan vigselceremonin är.
Om makarna inte bekänner sig till samma religion förrättas vigseln i magistraten och äktenskapet kan välsignas i kyrkan.
I den lutherska kyrkan kan medlemmar i kristna religionssamfund, till exempel en lutheran och en ortodox, vigas.
linkkiEvangelisk-lutherska kyrkan:
Information om äktenskapfinska _ svenska _ engelska
linkkiFinska ortodoxa kyrkan:
Finska ortodoxa kyrkanfinska _ svenska _ ryska
linkkiFritänkarförbundet r.f.:
Registrerade religiösa samfund med vigselrättfinska
Utländska medborgare
I magistraten vigs även utländska medborgare.
I Finland görs alltid en hindersprövning innan äktenskapet ingås.
Läs mer på InfoFinlands sida Prövning av hinder mot äktenskap.
Inverkan på uppehållstillstånd och medborgarskap
Maken, makan, sambon eller den registrerade partnern till en finsk eller en utländsk medborgare som är bosatt i Finland kan få ett uppehållstillstånd i Finland.
De kan få ett permanent uppehållstillstånd när äktenskapet har varat fem år.
Läs mer på InfoFinlands sida Uppehållstillstånd för make eller maka.
Finskt medborgarskap kan inte fås via äktenskap.
Äktenskap som ingåtts utomlands ska registreras i magistraten
Ett äktenskap som ingåtts utomlands är officiellt i Finland först när det registrerats i Finland.
Om äktenskapet har ingåtts utomlands måste man uppvisa ett legaliserat och översatt vigselintyg i magistraten för registrering.
Finska medborgare som är bosatta utomlands kan också skicka vigselhandlingarna till den lokala finska beskickningen som skickar handlingarna till magistraten i Finland.
Om personer som är bosatta i Finland antecknas grundläggande uppgifter i befolkningsdatasystemet.
Uppgifter som registreras är bland annat namn, födelsedatum, medborgarskap, familjeförhållanden och adress.
Utlänningar ska enligt lag anmäla till registret samma uppgifter som finska medborgare om deras vistelse i Finland varar över ett år.
Blanketten för registrering av ett äktenskap som ingåtts utomlandsfinska _ engelska
På den här sidan hittar du information om sådana ärenden som du måste sköta om du vill gifta dig i Finland.
Prövning av hinder mot äktenskap
Före äktenskapet måste en prövning av hinder mot äktenskap (avioliiton esteiden tutkinta) göras.
Vid hindersprövningen utreder myndigheterna om det finns hinder för äktenskapet enligt Finlands lag.
Du kan begära hindersprövning vid vilken magistrat (maistraatti) som helst.
Du måste själv skriftligt begära hindersprövning.
Prövningen tar ungefär en vecka.
När hindersprövningen är klar får du ett intyg om det.
Intyget är giltigt i fyra månader.
Du måste ta med dig intyget om hindersprövning till vigseltillfället.
Magistraten undersöker om det finns hinder mot äktenskapet utifrån de uppgifter som finns registrerade i Finlands befolkningsdatasystem.
Om det inte finns någon uppgift om ditt civilstånd i Finlands befolkningsdatasystem, ska du lämna in ett ämbetsbevis (siviilisäätytodistus) från myndigheten i ditt hemland till magistraten.
Du kan även skaffa intyget från ditt lands ambassad eller konsulat i Finland.
Om varken maken eller makan är finska medborgare och inte bor i Finland, ska de lämna in förutom ett ämbetsbevis till magistraten även en utredning över att lagen i deras hemland tillåter giftermål i Finland.
Observera att hindersprövningen kan ta flera veckor om den kräver intyg från andra länder.
Legalisering och översättning av intyg
Utländska intyg ska vanligtvis legaliseras och översättas till antingen svenska, finska eller engelska.
Även översättningen ska legaliseras.
Om översättningen görs av en auktoriserad översättare i Finland eller ett annat EU-land, behöver översättningen inte legaliseras.
Intyg som utfärdats av en myndighet i ett nordiskt land eller EU-land behöver inte legaliseras.
Inte heller intyg som utfärdats av en ambassad eller ett konsulat i Finland behöver legaliseras.
Om intyget har utfärdats av en myndighet i ett EU-land och åtföljs av blankett EU 2016/1191, behöver intyget inte översättas.
Anhållan om prövning av hinder mot äktenskapfinska _ svenska _ engelska
Beslut om efternamn
I Finland kan makarna byta efternamn när de gifter sig.
När du gifter dig kan du
behålla ditt nuvarande efternamn
ta din makes eller makas efternamn
bilda ett kombinerat efternamn av era efternamn.
I ett kombinerat efternamn syns båda efternamnen, till exempel Virtanen-Smith.
Namnen kan även skrivas isär, utan bindestreck.
Makarna kan även ansöka om ett helt nytt efternamn som deras gemensamma namn.
Ett nytt efternamn ansöks hos magistraten.
Ansökan är avgiftsbelagd.
Ett efternamn som maken eller makan har fått från sitt tidigare äktenskap kan inte väljas som efternamn.
Välj efternamnet tillsammans med din make eller maka redan när ni ansöker om prövning av hinder mot äktenskap.
Om du vill byta efternamn ska du meddela detta till magistraten.
Du får blanketten från magistraten eller på magistratens webbplats.
Om du inte meddelar att du vill byta efternamn, behåller du ditt efternamn.
Broschyren Makens efternamn och barnets efternamnfinska _ svenska _ engelska
Äktenskapsförord
Äktenskapsförord är frivilligt.
Med äktenskapsförord kan makarna utesluta giftorätten i den andras egendom antingen helt eller delvis om de skiljer sig eller om den ena av makarna dör.
Äktenskapsförord kan upprättas före äktenskapet eller under det.
Båda makarna ska underteckna äktenskapsförordet och två vittnen ska vidimera underskrifterna.
Äktenskapsförordet ska registreras hos magistraten, så att det kan träda i kraft.
Mer information om makarnas egendom hittar du på InfoFinlands sida Äkta makars rättigheter och skyldigheter.
Äktenskapsförordfinska _ svenska
Val av vigselform
Borgerlig vigsel sker hos magistraten (maistraatti) eller tingsrätten (käräjäoikeus).
Religiös vigsel sker i kyrkan eller ett annat religiöst samfund som har rätt att viga till äktenskap.
Båda makarna måste vara på plats vid vigseltillfället.
Dessutom ska minst två vittnen som har fyllt 15 år vara på plats.
Borgerlig vigsel
Boka tid för vigseln hos magistraten eller tingsrätten i god tid före bröllopsdagen.
En borgerlig vigsel är avgiftsfri om den sker i magistratens eller tingsrättens lokaler under tjänstetid.
Vigseln kan även ske på andra ställen, till exempel i hemmet eller en festlokal.
Alla har rätt till borgerlig vigsel, även de som tillhör ett trossamfund.
Religiös vigsel
Varje religiöst samfund bestämmer själv vilka villkor vigseln omfattas av och hurdan tillställning vigseln är.
Om du vill ha en religiös vigsel kommer du överens om detta med ett religiöst samfund.
Vigselfinska _ svenska _ engelska
Äktenskapsförord (avioehtosopimus) påverkar delningen av makarnas egendom vid skilsmässa eller dödsfall.
Om makarna inte har upprättat ett äktenskapsförord, räknas båda parternas egendom med i bodelningen och egendomen delas jämnt mellan makarna.
Vanligast är att äktenskapsförordet fastställer att ingendera maken har rätt till den andras egendom.
Äktenskapsförordet kan upprättas före eller under äktenskapet.
För det behövs båda makarnas medgivande.
Äktenskapsförordet görs skriftligt. Det dateras och undertecknas.
Därtill måste två ojäviga personer bevittna det.
Äktenskapsförordet skickas till magistraten för registrering.
Det är bra att anlita en kunnig jurist för upprättandet av avtalet.
Äktenskapsförordet är frivilligt.
Äktenskapsförordfinska _ svenska
Äktenskapsförord (avioehtosopimus) påverkar delningen av makarnas egendom vid skilsmässa eller dödsfall.
Om makarna inte har upprättat ett äktenskapsförord, räknas båda parternas egendom med i bodelningen och egendomen delas jämnt mellan makarna.
Vanligast är att äktenskapsförordet fastställer att ingendera maken har rätt till den andras egendom.
Äktenskapsförordet kan upprättas före eller under äktenskapet.
För det behövs båda makarnas medgivande.
Äktenskapsförordet görs skriftligt. Det dateras och undertecknas.
Därtill måste två ojäviga personer bevittna det.
Äktenskapsförordet skickas till magistraten för registrering.
Det är bra att anlita en kunnig jurist för upprättandet av avtalet.
Äktenskapsförordet är frivilligt.
Äktenskapsförordfinska _ svenska
Medborgare i alla länder kan gifta sig i Finland.
är minst 18 år gammal
inte är gift eller i registrerat parförhållande sedan tidigare.
Även samkönade par kan gifta sig i Finland.
Nära släktingar får inte gifta sig enligt Finlands lag.
Äktenskapet är alltid ett frivilligt val som ingen kan tvingas till.
Till exempel föräldrarna får inte tvinga sitt barn att gifta sig.
Att tvinga någon till äktenskap är ett brott i Finland.
I Finland kan kvinnor och män själva besluta vem de ska gifta sig med.
Man behöver inte be om tillstånd från till exempel släktingar.
Mer information om giftermål i Finland hittar du på InfoFinlands sida Ingående av äktenskap i Finland, komihåglista.
Äktenskap och uppehållstillstånd
Om din make eller maka bor stadigvarande i Finland, kan du få uppehållstillstånd i Finland på grund av äktenskapet.
Äktenskapet är dock ingen garanti för uppehållstillstånd.
Läs mer på InfoFinlands sida Uppehållstillstånd för make eller maka.
Du kan inte få finskt medborgarskap via ett äktenskap.
Äktenskap som ingåtts utomlands
Ett äktenskap som ingåtts utomlands är officiellt i Finland först när det har registrerats i befolkningsdatasystemet i Finland.
För registreringen ska du lämna in ett legaliserat äktenskapsintyg i original till magistraten (maistraatti) i din hemkommun.
Intyg som utfärdats av en myndighet i ett nordiskt land eller EU-land behöver inte legaliseras.
Om intyget är på ett annat språk än svenska, engelska eller finska, måste det översättas till ett av dessa språk. Även översättningen måste legaliseras.
Om översättningen görs av en auktoriserad översättare i Finland behöver den inte legaliseras.
Om intyget har utfärdats av en myndighet i ett EU-land och åtföljs av blankett EU 2016/1191, behöver intyget inte översättas.
Broschyr Information om äktenskapslagenfinska _ svenska _ engelska _ ryska _ arabiska
Om du har din hemvist i Finland bestäms ditt efternamn enligt finsk lag.
Detta görs även om du inte är finsk medborgare.
När ni ska gifta er måste ni fatta beslut om ert efternamn.
Ni
kan ta ett gemensamt efternamn eller
ha kvar era egna efternamn eller
bilda ett kombinerat efternamn av era efternamn.
I ett kombinerat efternamn syns bådas efternamn, till exempel Virtanen-Smith.
Namnen kan även skrivas isär, utan bindestreck.
Ni kan även välja att ta ett helt nytt efternamn som ert gemensamma namn.
Ansök om det nya efternamnet hos magistraten med ansökan om namnändring.
Ett efternamn som maken eller makan har fått från sitt tidigare äktenskap kan inte väljas som efternamn.
Välj efternamnet redan när ni ansöker om prövning av hinder mot äktenskap.
Meddela namnet till magistraten.
Ni får blanketten från magistraten eller på magistratens webbplats.
Broschyren Makens efternamn och barnets efternamnfinska _ svenska _ engelska
Ändring av efternamnet under äktenskap
Om du har ett kombinerat efternamn, till exempel Virtanen-Smith, kan du under äktenskapet lämna bort ettdera namnet.
Du kan också börja använda ett kombinerat efternamn under äktenskapet.
Du ansöker om detta skriftligt hos magistraten.
Uppgift till myndigheterna i det egna landet (utländska medborgare)
Om ditt efternamn ändras ska du meddela detta även till beskickningen för ditt eget land så att du får ett nytt pass med det nya namnet och så att myndigheterna i båda länderna har samma uppgifter.
Du får mer information om detta vid ditt eget lands beskickning.
Du hittar kontaktuppgifterna till beskickningarna på utrikesministeriets webbplats.
Läs mer om barnets efternamn på sidan När ett barn föds i Finland.
Läs mer om efternamn vid skilsmässa på sidan Skilsmässa.
Andra länders beskickningar i Finlandfinska _ svenska _ engelska
Om du har din hemvist i Finland bestäms ditt efternamn enligt finsk lag.
Detta görs även om du inte är finsk medborgare.
När ni ska gifta er måste ni fatta beslut om ert efternamn.
Ni
kan ta ett gemensamt efternamn eller
ha kvar era egna efternamn eller
bilda ett kombinerat efternamn av era efternamn.
I ett kombinerat efternamn syns bådas efternamn, till exempel Virtanen-Smith.
Namnen kan även skrivas isär, utan bindestreck.
Ni kan även välja att ta ett helt nytt efternamn som ert gemensamma namn.
Ansök om det nya efternamnet hos magistraten med ansökan om namnändring.
Ett efternamn som maken eller makan har fått från sitt tidigare äktenskap kan inte väljas som efternamn.
Välj efternamnet redan när ni ansöker om prövning av hinder mot äktenskap.
Meddela namnet till magistraten.
Ni får blanketten från magistraten eller på magistratens webbplats.
Broschyren Makens efternamn och barnets efternamnfinska _ svenska _ engelska
Ändring av efternamnet under äktenskap
Om du har ett kombinerat efternamn, till exempel Virtanen-Smith, kan du under äktenskapet lämna bort ettdera namnet.
Du kan också börja använda ett kombinerat efternamn under äktenskapet.
Du ansöker om detta skriftligt hos magistraten.
Uppgift till myndigheterna i det egna landet (utländska medborgare)
Om ditt efternamn ändras ska du meddela detta även till beskickningen för ditt eget land så att du får ett nytt pass med det nya namnet och så att myndigheterna i båda länderna har samma uppgifter.
Du får mer information om detta vid ditt eget lands beskickning.
Du hittar kontaktuppgifterna till beskickningarna på utrikesministeriets webbplats.
Läs mer om barnets efternamn på sidan När ett barn föds i Finland.
Läs mer om efternamn vid skilsmässa på sidan Skilsmässa.
Andra länders beskickningar i Finlandfinska _ svenska _ engelska
I Finland är det vanligt med familjer med en förälder.
Ett barn kan födas utom äktenskapet eller också är dess föräldrar skilda.
I familjer med en förälder bor en av föräldrarna med sina barn utan make eller maka.
Föräldern kan då ha antingen ensam eller gemensam vårdnad om barnet.
Som ensamstående förälder har man själv ansvaret för fostran av barnet.
Om föräldrarna däremot har gemensam vårdnad (yhteishuoltaja) kommer föräldrarna tillsammans överens om barnets angelägenheter.
Föräldrar som har gemensam vårdnad beslutar tillsammans om många saker. Dessa är barnets
bostadsort
fostran
språk
religion
utbildning
hälsovård
disponering av barnets egendom
Gemensam vårdnad förutsätter att barnets föräldrar klarar av att tillsammans agera för barnets bästa.
Till exempel för en passansökan behövs båda föräldrarnas tillstånd.
En ensamstående förälder fattar på egen hand alla beslut som rör barnet.
Myndigheter såsom daghem eller skola ger information om barnet endast till vårdnadshavaren.
Den andra föräldern får dock bestämma om vården och fostran av barnet när barnet är hos honom eller henne.
Vid skilsmässa eller när sambor flyttar isär måste föräldrarna besluta om barnets vårdnad, underhåll, boende och umgängesrätt.
Läs mer på InfoFinlands sida Barn vid skilsmässa.
Man kan också adoptera ett barn ensam.
Om du vill adoptera ett barn på egen hand, fråga om råd vid socialbyrån i din hemkommun.
Föreningen för familjer med en förälder (Yhden Vanhemman Perheiden Liitto) ger information och ordnar aktiviteter för familjer med en förälder.
På Finlex webbplats kan du läsa lagen angående vårdnad om barn och umgängesrätt.
Föreningen för små familjer är en medborgarorganisation som grundats av ensamstående föräldrar och som erbjuder aktiviteter för medlemsfamiljerna.
Lagen angående vårdnad om barn och umgängesrättfinska _ svenska _ engelska
linkkiFöreningen för familjer med en förälder r.f.:
Information för familjer med en förälderfinska
linkkiFöreningen för små familjer r.f.:
Verksamhet för små familjerfinska _ engelska
Underhållsbidrag
Båda föräldrarna bär ansvaret för underhållet av ett barn under 18 år, även om de inte bor tillsammans.
När föräldrarna skiljer sig ska de komma överens om underhållet av barnet samt om eventuellt underhållsbidrag (elatusapu).
Underhållsbidragets belopp beräknas utifrån barnets underhållsbehov och föräldrarnas underhållsförmåga.
Med barnets underhållsbehov avses det penningbelopp som försörjningen av barnet kostar varje månad.
I beloppet ingår till exempel utgifter för mat och kläder samt eventuella dagvårdsavgifter.
Barnets underhållsbehov delas mellan föräldrarna enligt deras underhållsförmåga.
Underhållsförmågan beräknas genom att dra av skatter och övriga obligatoriska utgifter av inkomsterna.
Du kan be om hjälp med att beräkna underhållsbehovet hos barnatillsyningsmannen (lastenvalvoja) i din hemkommun.
Det är bra att upprätta ett skriftligt avtal om underhållsbidraget som socialnämnden bekräftar.
Ett avtal som bekräftats på detta sätt är lika officiellt som ett domstolsbeslut.
Begär bekräftande av avtalet hos barnatillsyningsmannen i din hemkommun.
Om föräldrarna inte kan enas om underhållsbidraget kan de få hjälp i form av medling i familjefrågor.
I sista hand avgörs ärendet i tingsrätten.
Mer information om medling i familjefrågor hittar du på InfoFinlands sida Skilsmässa.
Underhållsstöd
I vissa situationer kan den förälder som bor med barnet ansöka om underhållsstöd (elatustuki) vid FPA.
Du kan ansöka om underhållsstöd från Fpa i följande situationer:
Den underhållsskyldiga föräldern har inte betalat det bekräftade underhållsbidraget (Fpa indriver det hos denne senare).
Underhållsbidraget har på grund av förälderns ekonomiska situation fastställts till ett belopp som underskrider underhållsstödet.
Det har på grund av förälderns ekonomiska situation fastställts att inget underhållsbidrag betalas.
Faderskapet har inte fastställts för ett barn fött utom äktenskapet.
Du kan få underhållsstöd om du bor stadigvarande i Finland.
Du kan få underhållsstöd också om du har flyttat till Finland från ett annat EU- eller EES-land eller Schweiz för att arbeta.
Också barnet för vilket man söker underhållsstöd ska bo i Finland.
Du får mer information om underhållsstödet på Fpa.
Underhållsbidrag och underhållsstödfinska _ svenska _ engelska
Skilsmässa i Finlandengelska _ ryska _ estniska
På den här sidan finns information om tjänsterna i Rovaniemi.
Annan viktig information om boendet i Finland finns på InfoFinlands sida Boende.
Hyresboende
Kunta-asunnot Oy:s bostäder
Övriga hyresbostäder
Bostäder för ungdomar och studerande
Boende i ägarbostad
Boende i bostadsrättsbostad
Napapiirin Residuum
Oy
Hyresboende
Förfrågningar om hyresbostäder på Rovaniemi stads område kan ställas direkt till fastighetsägare eller till bostadsförmedlingar.
Kunta-asunnot Oy:s bostäder
Via Rovanapa Oy kan du ansöka om en bostad vid Kunta-asunnot Oy.
Lediga bostäder och ansökningsblanketter hittar du även på Kunta-asunnot Oy:s webbplats..
Adress:
Kontaktuppgifter till enheten som väljer hyresgästerna, telefontid kl. 12–15:
tfn 016 3223 412
tfn 016 3223 414
Övriga hyresbostäder
hittar du en lista över webbsidor där du kan ansöka om bostad.
På sidan finns även information om att bo i hyresbostad och om sådant som rör flytten.
Information om boendefinska _ engelska
Bostäder för ungdomar och studerande
Också ungdomar och studerande kan söka Kunta-asunnot Oy:s bostäder och andra hyresbostäder.
Ungdomar kan även söka bostad via ungdomsbostadsföreningen Rovaniemen nuorisoasunnot ry.
Om du studerar vid gymnasium, yrkesläroanstalt, yrkeshögskola eller universitet kan du söka bostad hos Domus Arctica-stiftelsen.
Ungdomsbostadsföreningen Rovaniemen nuorisoasunnot ry:s webbplatsfinska
Domus Arctica-stiftelsens webbplatsfinska _ engelska
Studentkåren vid Lapplands universitet informerar också om bostäder som hyrs ut till studerande.
Dessa bostäder hittar du på studentkårens webbplats.
Mer information om boende hittar du under följande länkar.
linkkiRovaniemi stads ungdomstjänster:
Hyresbostäder i Rovaniemifinska
linkkiFörbundet för ungdomsbostäder rf:
Boendeguide för ungafinska
Privatpersoner lägger även ut tidningsannonser om bostäder som de hyr ut.
Boende i ägarbostad
De flesta invånarna i Rovaniemi äger sin bostad. De har tagit lån eller finansierat sin bostad på andra sätt.
Staten stöder boende i ägarbostad genom att gå i borgen för privatpersoners bostadslån.
Dessutom är en del av räntan på bostadslånet avdragsgill i beskattningen.
Mer information om att köpa en egen bostad får du på banken eller hos fastighetsförmedlare.
Fastighetsförmedlare och privatpersoner annonserar bostäder som de säljer i lokaltidningar (såsom Lapin Kansa) och på Internet.
Allmän information om boende:
Miljöministeriet linkkiMiljöministeriet:
Webbplatsen asuminen.fifinska _ svenska _ engelska
Boende i bostadsrättsbostad
Att bo i en bostadsrättsbostad är ett alternativ till att köpa eller hyra sin bostad.
Genom att betala en bostadsrättsavgift, som är 15 procent av bostadens anskaffningspris, och därefter varje månad ett rimligt bruksvederlag får man rätt att förvalta över bostaden precis som om den vore en ägarbostad.
Man kan inte lösa in bostaden, men man kan sälja bostadsrätten eller byta till en annan bostad.
I Rovaniemi finns 400 bostadsrättsbostäder.
Om du är intresserad av en bostad ska du kontakta något av de företag som tillhandahåller bostadsrättsbostäder:
Webbplats för Asokoditfinska
Oyfinska
Oy finska
Mer information om hur man ansöker om en bostadsrättsbostad (Rovaniemi stad, miljötillsyn):
tfn 016 322 8091 eller tfn 016 322 8014
Byggande och tomter
Mer information om bygglov och tomter samt om vatten, el och hushållsavfall hittar du under länkarna nedan.
Napapiirin Residuum
Oy
Sopsortering och avfallsåtervinningfinska
På den här sidan finns information om tjänsterna i Rovaniemi.
Annan viktig information om boendet i Finland finns på InfoFinlands sida Boende.
Hyresboende
Kunta-asunnot Oy:s bostäder
Övriga hyresbostäder
Bostäder för ungdomar och studerande
Boende i ägarbostad
Boende i bostadsrättsbostad
Napapiirin Residuum
Oy
Hyresboende
Förfrågningar om hyresbostäder på Rovaniemi stads område kan ställas direkt till fastighetsägare eller till bostadsförmedlingar.
Kunta-asunnot Oy:s bostäder
Via Rovanapa Oy kan du ansöka om en bostad vid Kunta-asunnot Oy.
Lediga bostäder och ansökningsblanketter hittar du även på Kunta-asunnot Oy:s webbplats..
Adress:
Kontaktuppgifter till enheten som väljer hyresgästerna, telefontid kl. 12–15:
tfn 016 3223 412
tfn 016 3223 414
Övriga hyresbostäder
hittar du en lista över webbsidor där du kan ansöka om bostad.
På sidan finns även information om att bo i hyresbostad och om sådant som rör flytten.
Information om boendefinska _ engelska
Bostäder för ungdomar och studerande
Också ungdomar och studerande kan söka Kunta-asunnot Oy:s bostäder och andra hyresbostäder.
Ungdomar kan även söka bostad via ungdomsbostadsföreningen Rovaniemen nuorisoasunnot ry.
Om du studerar vid gymnasium, yrkesläroanstalt, yrkeshögskola eller universitet kan du söka bostad hos Domus Arctica-stiftelsen.
Ungdomsbostadsföreningen Rovaniemen nuorisoasunnot ry:s webbplatsfinska
Domus Arctica-stiftelsens webbplatsfinska _ engelska
Studentkåren vid Lapplands universitet informerar också om bostäder som hyrs ut till studerande.
Dessa bostäder hittar du på studentkårens webbplats.
Mer information om boende hittar du under följande länkar.
linkkiRovaniemi stads ungdomstjänster:
Hyresbostäder i Rovaniemifinska
linkkiFörbundet för ungdomsbostäder rf:
Boendeguide för ungafinska
Privatpersoner lägger även ut tidningsannonser om bostäder som de hyr ut.
Boende i ägarbostad
De flesta invånarna i Rovaniemi äger sin bostad. De har tagit lån eller finansierat sin bostad på andra sätt.
Staten stöder boende i ägarbostad genom att gå i borgen för privatpersoners bostadslån.
Dessutom är en del av räntan på bostadslånet avdragsgill i beskattningen.
Mer information om att köpa en egen bostad får du på banken eller hos fastighetsförmedlare.
Fastighetsförmedlare och privatpersoner annonserar bostäder som de säljer i lokaltidningar (såsom Lapin Kansa) och på Internet.
Allmän information om boende:
Miljöministeriet linkkiMiljöministeriet:
Webbplatsen asuminen.fifinska _ svenska _ engelska
Boende i bostadsrättsbostad
Att bo i en bostadsrättsbostad är ett alternativ till att köpa eller hyra sin bostad.
Genom att betala en bostadsrättsavgift, som är 15 procent av bostadens anskaffningspris, och därefter varje månad ett rimligt bruksvederlag får man rätt att förvalta över bostaden precis som om den vore en ägarbostad.
Man kan inte lösa in bostaden, men man kan sälja bostadsrätten eller byta till en annan bostad.
I Rovaniemi finns 400 bostadsrättsbostäder.
Om du är intresserad av en bostad ska du kontakta något av de företag som tillhandahåller bostadsrättsbostäder:
Webbplats för Asokoditfinska
Oyfinska
Oy finska
Mer information om hur man ansöker om en bostadsrättsbostad (Rovaniemi stad, miljötillsyn):
tfn 016 322 8091 eller tfn 016 322 8014
Byggande och tomter
Mer information om bygglov och tomter samt om vatten, el och hushållsavfall hittar du under länkarna nedan.
Napapiirin Residuum
Oy
På den här sidan finns information om tjänsterna i Rovaniemi.
Hyresboende
Kunta-asunnot Oy:s bostäder
Boende i ägarbostad
Boende i bostadsrättsbostad
Napapiirin Residuum
Oy Hyresboende
Förfrågningar om hyresbostäder på Rovaniemi stads område kan ställas direkt till fastighetsägare eller till bostadsförmedlingar.
Kunta-asunnot Oy:s bostäder
Via Rovanapa Oy kan du ansöka om en bostad vid Kunta-asunnot Oy. Lediga bostäder och ansökningsblanketter hittar du även på Kunta-asunnot Oy:s webbplats..
tfn 016 3223 412 tfn 016 3223 414
Övriga hyresbostäder
hittar du en lista över webbsidor där du kan ansöka om bostad.
På sidan finns även information om att bo i hyresbostad och om sådant som rör flytten.
Information om boendefinska _ engelska
Bostäder för ungdomar och studerande
Också ungdomar och studerande kan söka Kunta-asunnot Oy:s bostäder och andra hyresbostäder.
Domus Arctica-stiftelsens webbplatsfinska _ engelska
Studentkåren vid Lapplands universitet informerar också om bostäder som hyrs ut till studerande.
Dessa bostäder hittar du på studentkårens webbplats.
Mer information om boende hittar du under följande länkar.
linkkiRovaniemi stads ungdomstjänster: Hyresbostäder i Rovaniemifinska
linkkiFörbundet för ungdomsbostäder rf: Boendehandbok för ungdomarfinska
Privatpersoner lägger även ut tidningsannonser om bostäder som de hyr ut.
Boende i ägarbostad
De har tagit lån eller finansierat sin bostad på andra sätt.
Dessutom är en del av räntan på bostadslånet avdragsgill i beskattningen.
Mer information om att köpa en egen bostad får du på banken eller hos fastighetsförmedlare.
Fastighetsförmedlare och privatpersoner annonserar bostäder som de säljer i lokaltidningar (såsom Lapin Kansa) och på Internet.
Allmän information om boende:
Miljöministeriet linkkiMiljöministeriet:
Webbplatsen asuminen.fifinska _ svenska _ engelska
Boende i bostadsrättsbostad
Att bo i en bostadsrättsbostad är ett alternativ till att köpa eller hyra sin bostad.
Genom att betala en bostadsrättsavgift, som är 15 procent av bostadens anskaffningspris, och därefter varje månad ett rimligt bruksvederlag får man rätt att förvalta över bostaden precis som om den vore en ägarbostad.
Man kan inte lösa in bostaden, men man kan sälja bostadsrätten eller byta till en annan bostad.
Om du är intresserad av en bostad ska du kontakta något av de företag som tillhandahåller bostadsrättsbostäder:
Webbplats för Asokoditfinska
Avainboendefinska
Oy finska
Förfrågningar om bostadsrättsavgifter och bruksvederlag samt om lediga bostäder eller bostäder som kommer att bli lediga ställs direkt till ägaren.
Mer information om hur man ansöker om en bostadsrättsbostad (Rovaniemi stad, miljötillsyn):
tfn 016 322 8091 eller tfn 016 322 8014
Byggande och tomter
Mer information om bygglov och tomter samt om vatten, el och hushållsavfall hittar du under länkarna nedan.
Napapiirin Residuum
Oy
Före äktenskapet ska ni tillsammans skriftligt begära hindersprövning (esteiden tutkiminen).
Hindersprövningen görs i magistraten (maistraatti).
Skriftlig begäran kan lämnas in till vilken magistrat som helst.
Hindersprövningen kostar ingenting.
Om endera parten hör till den evangelisk-lutherska kyrkan eller ortodoxa kyrkan kan ni också begära hindersprövning i den egna församlingen.
Hindersprövningen är obligatorisk och utan den kan vigseln inte förrättas.
Av hindersprövningen framgår till exempel om den ena parten redan är gift med någon annan.
I Finland tar hindersprövningen ungefär en vecka.
Intyget över hindersprövningen är i kraft fyra månader.
Om äktenskapet inte ingås inom denna tid måste hindersprövningen göras på nytt.
Intyget över hindersprövningen ska finnas med vid vigselförrättningen.
Till Finland genom giftermål
Enligt Finlands lag ska hinder mot äktenskap prövas om du är finsk medborgare eller permanent bosatt i Finland och uppgifterna om dig finns i befolkningsregistret.
Om uppgifterna om en utländsk maka eller make inte kan kontrolleras i befolkningsdatasystemet måste personen lämna ett intyg från myndigheterna i sitt eget land för prövning av äktenskapshinder till magistraten.
Det är bra att reservera tid för detta eftersom förfaringssätten varierar i olika länder.
Du kan fråga mer om vilka intyg som behövs vid magistraten.
Den utländska partnern behöver dessutom ett identitetsbevis, ett civilståndsintyg (ogift, skild, änka/änkling) och ett Apostilleintyg för dessa.
Apostilleintyget bevisar att myndighetshandlingen är utfärdad av en behörig person.
Myndigheter som utfärdar Apostilleintyg finns i alla länder som är anslutna till Haagkonventionen.
En engelskspråkig förteckning över konventionsstaterna finns på webbplatsen för internationella domstolen i Haag.
Dokument som införs från andra länder ska dessutom ha en stämpel som bestyrker dokumentet.
Stämpeln ska begäras vid utrikesministeriet i det ifrågavarande landet och dessutom vid Finlands beskickning i landet.
Fråga mer om detta vid beskickningen för ditt eget land.
Kontaktuppgifter till magistratfinska _ svenska _ engelska
Anhållan om prövning av hinder mot äktenskapfinska _ svenska
Länder som är anslutna till Apostilleavtaletengelska _ franska _ spanska _ tyska _ portugisiska
Före äktenskapet ska ni tillsammans skriftligt begära hindersprövning (esteiden tutkiminen).
Hindersprövningen görs i magistraten (maistraatti).
Skriftlig begäran kan lämnas in till vilken magistrat som helst.
Hindersprövningen kostar ingenting.
Om endera parten hör till den evangelisk-lutherska kyrkan eller ortodoxa kyrkan kan ni också begära hindersprövning i den egna församlingen.
Hindersprövningen är obligatorisk och utan den kan vigseln inte förrättas.
Av hindersprövningen framgår till exempel om den ena parten redan är gift med någon annan.
I Finland tar hindersprövningen ungefär en vecka.
Intyget över hindersprövningen är i kraft fyra månader.
Om äktenskapet inte ingås inom denna tid måste hindersprövningen göras på nytt.
Intyget över hindersprövningen ska finnas med vid vigselförrättningen.
Till Finland genom giftermål
Enligt Finlands lag ska hinder mot äktenskap prövas om du är finsk medborgare eller permanent bosatt i Finland och uppgifterna om dig finns i befolkningsregistret.
Om uppgifterna om en utländsk maka eller make inte kan kontrolleras i befolkningsdatasystemet måste personen lämna ett intyg från myndigheterna i sitt eget land för prövning av äktenskapshinder till magistraten.
Det är bra att reservera tid för detta eftersom förfaringssätten varierar i olika länder.
Du kan fråga mer om vilka intyg som behövs vid magistraten.
Den utländska partnern behöver dessutom ett identitetsbevis, ett civilståndsintyg (ogift, skild, änka/änkling) och ett Apostilleintyg för dessa.
Apostilleintyget bevisar att myndighetshandlingen är utfärdad av en behörig person.
Myndigheter som utfärdar Apostilleintyg finns i alla länder som är anslutna till Haagkonventionen.
En engelskspråkig förteckning över konventionsstaterna finns på webbplatsen för internationella domstolen i Haag.
Dokument som införs från andra länder ska dessutom ha en stämpel som bestyrker dokumentet.
Stämpeln ska begäras vid utrikesministeriet i det ifrågavarande landet och dessutom vid Finlands beskickning i landet.
Fråga mer om detta vid beskickningen för ditt eget land.
Kontaktuppgifter till magistratfinska _ svenska _ engelska
Anhållan om prövning av hinder mot äktenskapfinska _ svenska
Länder som är anslutna till Apostilleavtaletengelska _ franska _ spanska _ tyska _ portugisiska
Definition av en familj
I Finland utgörs en familj av
makar
sambor
ogifta barn under 18 och deras vårdnadshavare som bor i Finland
I Finland uppfattas en familj i snävare bemärkelse än i många andra länder.
I Finland anses oftast kärnfamiljen, d.v.s. föräldrarna och barnen utgöra en familj.
Till exempel om mor- eller farföräldrarna, föräldrarna och barnen bor i samma lägenhet räknas officiellt bara föräldrarna och barnen till samma familj.
Mor- eller farföräldrarna bildar en egen familj.
En familj kan ha barn eller bestå av ett barnlöst par.
De vuxna i familjen kan vara av samma eller olika kön.
En familj bildas också av en ensamstående mor eller far och hens barn.
Med ombildade familjer avses ett par som bor tillsammans med ett eller flera barn från parets tidigare förhållanden.
Också parets gemensamma barn kan bo med familjen.
Om du är frånskild kan du gifta om dig utan tillstånd från din före detta maka eller make.
Du behöver inte tillstånd från din före detta maka eller make för att ingå ett nytt äktenskap även om du och din före detta maka eller make har barn tillsammans.
Regnbågsfamiljer
Regnbågsfamiljer är familjer som bildas av homosexuella, lesbiska, bi- och transsexuella föräldrar och deras barn.
De är till exempel familjer som bildas av två kvinnor eller två män samt familjer med fler än två föräldrar
Gifta makar av samma kön har rätt att adoptera ett barn och rätt till adoption inom familjen.
Adoption inom familjen betyder att makan/maken adopterar sin makas/makes barn och blir officiellt barnets andra förälder.
I Finland kan ett barn ha högst två juridiska föräldrar.
Om du planerar adoption inom familjen ska du kontakta socialbyrån i din hemkommun.
Regnbågsfamiljer rf är en organisation som stöder regnbågsfamiljer samt ger råd och ordnar verksamhet för dem.
Kontaktuppgifterna hittar du på organisationens webbplats.
linkkiRegnbågsfamiljer:
Stöd och verksamhet för regnbågsfamiljerfinska
Underhållsskyldighet
Enligt Finlands lag är föräldrarna förpliktade att ta hand om sina minderåriga barn ekonomiskt och gifta par om varandra.
Familjemedlemmarnas underhållsskyldighet sträcker sig inte till släktingar, till exempel vuxna syskon eller mor- eller farföräldrar.
I Finland utgår man alltså inte från att enskilda människor tar hand om sådana släktingar som har det dåligt ställt ekonomiskt.
Stödet kommer från samhället i form av den sociala tryggheten.
Hushåll
Till samma hushåll hör alla som stadigvarande bor i samma bostad.
Mer information om ämnet hushåll finns på InfoFinlands sida boende.
Parförhållande
Ett par kan välja om de vill leva tillsammans i ett samboförhållande eller i ett äktenskap.
Det är bra att beakta att parförhållandets form påverkar makarnas rättigheter och skyldigheter, frågor som rör egendom och arv, vårdnad om och underhåll av barn samt adoption.
Råd i frågor som rör familjen
Väestöliitto tillhandahåller rådgivning telefonledes och via e-post när du behöver samtalsstöd i frågor som rör barnuppfostran eller relationerna i familjen.
Samtal tas emot på följande språk:
ryska och engelska tfn 050 325 7173
Läs mer på InfoFinlands sida Fostran av barn i Finland.
Läs mer på InfoFinlands sida Problem i familjen.
Till Finland på grund av familjebandfinska _ svenska _ engelska
linkkiBefolkningsförbundet:
Rådgivning till invandrare telefonledes och via e-postfinska _ svenska _ engelska
Handbok för familjer med två kulturer (pdf, 4,74 Mt)finska _ engelska _ ryska _ franska _ spanska _ thai
På den här sidan hittar du information om ärenden som du måste sköta då du vill ingå äktenskap i Finland.
Prövning av äktenskapshinder
Före äktenskapet måste hinder mot äktenskapet prövas.
Detta görs antingen av den magistrat eller den församling som förrättar vigseln.
Läs mer om prövning av äktenskapshinder på InfoFinlands sida Prövning av hinder mot äktenskap.
Välja efternamn
När du gifter dig kan du och din make eller maka ta ett gemensamt efternamn.
Du kan också behålla ditt eget efternamn eller ta ett dubbelnamn.
Mer information hittar du på InfoFinlands sida Välja efternamn.
Civilvigsel eller religiös vigsel
I Finland kan äktenskap ingås
i ett religiöst samfund som har rätt att förrätta vigsel
Civilvigsel förrättas i magistraten, religiös vigsel förrättas i en kyrka eller i något annat religiöst samfund.
Mer information hittar du på InfoFinlands sida Vigsel.
På den här sidan hittar du information om ärenden som du måste sköta då du vill ingå äktenskap i Finland.
Prövning av äktenskapshinder
Före äktenskapet måste hinder mot äktenskapet prövas.
Detta görs antingen av den magistrat eller den församling som förrättar vigseln.
Läs mer om prövning av äktenskapshinder på InfoFinlands sida Prövning av hinder mot äktenskap.
Välja efternamn
När du gifter dig kan du och din make eller maka ta ett gemensamt efternamn.
Du kan också behålla ditt eget efternamn eller ta ett dubbelnamn.
Mer information hittar du på InfoFinlands sida Välja efternamn.
Civilvigsel eller religiös vigsel
I Finland kan äktenskap ingås
i ett religiöst samfund som har rätt att förrätta vigsel
Civilvigsel förrättas i magistraten, religiös vigsel förrättas i en kyrka eller i något annat religiöst samfund.
Mer information hittar du på InfoFinlands sida Vigsel.
Handikappbidrag för barn under 16 år
Ett barn under 16 år kan få handikappbidrag (vammaistuki) om hen på grund av sitt handikapp eller sin sjukdom behöver regelbunden vård, omsorg och rehabilitering under minst sex månaders tid.
Du ansöker om handikappbidrag för barn under 16 år vid FPA.
Handikappbidraget beviljas vanligtvis för en bestämd period.
När perioden har gått kan man ansöka om förlängning för bidraget.
Handikappbidrag för barnfinska _ svenska _ engelska
Specialvårdspenning
Du kan få specialvårdspenning från FPA om
ditt barn är under 16 år och vårdas på sjukhus eller
om du tar hand om barnet i hemmet och hemvården ansluter sig till barnets sjukhusvård eller
om utbetalningen av ditt arbetsmarknadsstöd avbryts tillfälligt eftersom du på grund av vården av ditt barn inte kan delta i integrationsåtgärderna eller
ditt barn provar på att återvända till skolan eller barnomsorgen.
Specialvårdspenning för barn under 16 årfinska _ svenska _ engelska
Rehabilitering för barn
FPA ordnar rehabiliteringen och ersätter kostnaderna för den.
Rehabiliteringen kan omfatta många olika slags aktiviteter.
Den kan till exempel bestå av fysioterapi eller olika kurser där man lär sig att leva med sitt handikapp.
FPA kan även ordna rehabilitering som behovsprövad rehabilitering (harkinnanvarainen kuntoutus).
Behovsprövad rehabilitering har som mål att förbättra arbets- eller funktionsförmågan.
Om barnet inte kan få krävande medicinska rehabilitering från FPA, ska rehabiliteringen ordnas av hemkommunen.
Krävande medicinsk rehabiliteringfinska _ svenska _ engelska
Handikappade barns skolgång
Ett handikappat barn har rätt till skolgång i närliggande skola.
Ett handikappat barn kan få specialundervisning om barnets handikapp försvårar inlärningen.
Barnet kan vid behov även få ett skolgångsbiträde (koulunkäyntiavustaja).
FPA kan betala dyra och krävande hjälpmedel (apuväline) som det handikappade barnet behöver för sin skolgång.
Sådana hjälpmedel är till exempel datorer och tilläggsutrustning till datorer.
Barnet kan också få hjälpmedel om han eller hon inte kan studera utan dem eller om det är mycket svårt utan dem.
Hjälpmedel kan fås tidigast när barnet går i grundskolans årskurs sju.
Hjälpmedel för arbete och studierfinska _ svenska _ engelska
Handikappade barns fritid
Information om hobbymöjligheterna på din hemort får du till exempel vid idrotts- och kulturförvaltningen i din hemkommun.
Också handikapporganisationer tillhandahåller många slags hobbyverksamheter.
Till exempel föreningen för handikappidrott och -motion i Finland, VAU ry, ordnar olika idrotts- och motionsevenemang.
linkkiDe Utvecklingsstördas Stödförbund (VAU):
Motion för handikappade barn och ungafinska _ svenska _ engelska
Enligt Finlands lag är äktenskapet (avioliitto) ett lagstadgat förhållande mellan två människor.
Äktenskap ingås genom vigsel.
Det är vanligt att par lever i ett samboförhållande före äktenskapet.
Läs mer på InfoFinlands sida Samboförhållande.
Förlovning
Före äktenskapet kan ett par förlova sig.
Förlovningen är ett löfte om äktenskap.
Förlovningen är frivillig och krävs inte i lag.
Paret kan hålla förlovningen privat eller offentliggöra den till andra människor.
Vem kan ingå äktenskap?
I Finland kan alla gifta sig som
har fyllt 18 år och
inte är gifta eller under förmynderskap.
En person som står under förmynderskap klarar inte av att sköta sina angelägenheter utan de sköts av en intressebevakare.
Äktenskap mellan två personer av samma kön har varit tillåtet i Finland sedan 1.3.2017.
Innan dess kunde två personer av samma kön endast ingå ett registrerat partnerskap.
Nya registrerade partnerskap kan inte längre ingås i Finland, men tidigare registrerad partnerskap förblir i kraft.
Ett registrerat partnerskap kan ändras till äktenskap vid magistraten.
Äktenskap mellan följande nära släktingar är förbjudet:
barn och föräldrar
syskon eller halvsyskon
adoptivföräldrar och adoptivbarn samt
barn till syskon (till exempel morbror och systerdotter).
Justitieministeriet kan på synnerligen vägande skäl ge tillstånd till äktenskap i de två sistnämnda fallen.
Äktenskapet är alltid ett frivilligt val som ingen kan tvingas till.
När äktenskapets lagliga villkor uppfylls kan ett par gifta sig.
De behöver till exempel inte be om tillstånd av släktingar.
På justitieministeriets webbplats beskrivs kortfattat bestämmelserna om giftermål och skilsmässa samt äktenskapets rättsverkningar.
Äktenskapslagen finns i sin helhet på Finlex webbplats.
Broschyr Information om äktenskapslagenfinska _ svenska _ engelska _ ryska _ arabiska
Äktenskapslagenfinska _ svenska _ engelska
Enligt Finlands lag är äktenskapet (avioliitto) ett lagstadgat förhållande mellan två människor.
Äktenskap ingås genom vigsel.
Det är vanligt att par lever i ett samboförhållande före äktenskapet.
Läs mer på InfoFinlands sida Samboförhållande.
Förlovning
Före äktenskapet kan ett par förlova sig.
Förlovningen är ett löfte om äktenskap.
Förlovningen är frivillig och krävs inte i lag.
Paret kan hålla förlovningen privat eller offentliggöra den till andra människor.
Vem kan ingå äktenskap?
I Finland kan alla gifta sig som
har fyllt 18 år och
inte är gifta eller under förmynderskap.
En person som står under förmynderskap klarar inte av att sköta sina angelägenheter utan de sköts av en intressebevakare.
Äktenskap mellan två personer av samma kön har varit tillåtet i Finland sedan 1.3.2017.
Innan dess kunde två personer av samma kön endast ingå ett registrerat partnerskap.
Nya registrerade partnerskap kan inte längre ingås i Finland, men tidigare registrerad partnerskap förblir i kraft.
Ett registrerat partnerskap kan ändras till äktenskap vid magistraten.
Äktenskap mellan följande nära släktingar är förbjudet:
barn och föräldrar
syskon eller halvsyskon
adoptivföräldrar och adoptivbarn samt
barn till syskon (till exempel morbror och systerdotter).
Justitieministeriet kan på synnerligen vägande skäl ge tillstånd till äktenskap i de två sistnämnda fallen.
Äktenskapet är alltid ett frivilligt val som ingen kan tvingas till.
När äktenskapets lagliga villkor uppfylls kan ett par gifta sig.
De behöver till exempel inte be om tillstånd av släktingar.
På justitieministeriets webbplats beskrivs kortfattat bestämmelserna om giftermål och skilsmässa samt äktenskapets rättsverkningar.
Äktenskapslagen finns i sin helhet på Finlex webbplats.
Broschyr Information om äktenskapslagenfinska _ svenska _ engelska _ ryska _ arabiska
Äktenskapslagenfinska _ svenska _ engelska
Om du på grund av skada eller sjukdom inte kan arbeta kan du få invalidpension (työkyvyttömyyseläke).
Om du är blind eller rörelsehindrad kan du få invalidpension även om du skulle kunna arbeta.
Invalidpension betalas till 16–64-åringar.
Huruvida du får pensionen beror på hur länge du har bott i Finland.
Vanligtvis kan du få invalidpension när du har bott tre år i Finland.
Du kan söka invalidpension hos FPA.
Sjukpensionfinska _ svenska _ engelska
Handikappbidrag för vuxna
Om du har ett handikapp eller en sjukdom som försämrar din funktionsförmåga sammanhängande under minst ett år kan du få handikappbidrag (vammaistuki).
Du måste ha ett läkarintyg för att få handikappbidrag.
Handikappbidrag för vuxna betalas till 16–64-åringar.
Huruvida du får bidraget beror på hur länge du har bott i Finland.
Vanligtvis kan du få handikappbidrag när du har bott tre år i Finland.
Handikappbidragets storlek beror på hur svårt ditt handikapp är.
Du kan söka handikappbidrag hos FPA.
Handikappbidrag för vuxnafinska _ svenska _ engelska
Hälsa och rehabiliteringfinska _ svenska _ ryska _ estniska
Stöd för vård av en handikappad anhörig
Om du vårdar en handikappad närstående i hemmet kan du få stöd för närståendevård (omaishoidontuki) från din hemkommun.
För att få stöd måste du göra ett avtal om närståendevård med din kommun.
Du kan ansöka om stödet vid socialbyrån i din egen kommun.
linkkiNärståendevårdare och Vänner -Förbundet rf:
Handikappbidrag för barn och specialvårdpenning
Läs mer om handikappbidrag för barn och specialvårdpenning på InfoFinlands sida Ett handikappat barn.
Vårdbidrag för pensionstagare
En pensionär vars funktionsförmåga försämrats under sammanlagt minst ett år på grund av sjukdom eller skada kan få vårdbidrag för pensionstagare (eläkettä saavan hoitotuki).
Du kan få stöd om du på grund av ditt handikapp eller din sjukdom behöver kontinuerligt hjälp.
Hur stort stöd du får beror på hur mycket hjälp du behöver.
Vårdbidrag för pensionstagare kan sökas hos FPA.
Vårdbidrag för pensionstagarefinska _ svenska _ engelska
Bidrag för kläder och mat
Om ditt handikapp eller din sjukdom orsakar dig extra kostnader för mat eller kläder kan du ansöka om bidrag för kläder och mat (vaatetus- ja ravitsemustuki).
Du kan ansöka om bidraget vid socialbyrån i din hemkommun.
linkkiInstitutet för hälsa och välfärd:
Extra kostnader för kläder och matfinska _ svenska
I Finland är det vanligt med familjer med en förälder.
Ett barn kan födas utom äktenskapet eller också är dess föräldrar skilda.
I familjer med en förälder bor en av föräldrarna med sina barn utan make eller maka.
Föräldern kan då ha antingen ensam eller gemensam vårdnad om barnet.
Som ensamstående förälder har man själv ansvaret för fostran av barnet.
Om föräldrarna däremot har gemensam vårdnad (yhteishuoltaja) kommer föräldrarna tillsammans överens om barnets angelägenheter.
Föräldrar som har gemensam vårdnad beslutar tillsammans om många saker. Dessa är barnets
bostadsort
fostran
språk
religion
utbildning
hälsovård
disponering av barnets egendom
Gemensam vårdnad förutsätter att barnets föräldrar klarar av att tillsammans agera för barnets bästa.
Till exempel för en passansökan behövs båda föräldrarnas tillstånd.
En ensamstående förälder fattar på egen hand alla beslut som rör barnet.
Myndigheter såsom daghem eller skola ger information om barnet endast till vårdnadshavaren.
Den andra föräldern får dock bestämma om vården och fostran av barnet när barnet är hos honom eller henne.
Vid skilsmässa eller när sambor flyttar isär måste föräldrarna besluta om barnets vårdnad, underhåll, boende och umgängesrätt.
Läs mer på InfoFinlands sida Barn vid skilsmässa.
Man kan också adoptera ett barn ensam.
Om du vill adoptera ett barn på egen hand, fråga om råd vid socialbyrån i din hemkommun.
Föreningen för familjer med en förälder (Yhden Vanhemman Perheiden Liitto) ger information och ordnar aktiviteter för familjer med en förälder.
På Finlex webbplats kan du läsa lagen angående vårdnad om barn och umgängesrätt.
Föreningen för små familjer är en medborgarorganisation som grundats av ensamstående föräldrar och som erbjuder aktiviteter för medlemsfamiljerna.
Lagen angående vårdnad om barn och umgängesrättfinska _ svenska _ engelska
linkkiFöreningen för familjer med en förälder r.f.:
Information för familjer med en förälderfinska
linkkiFöreningen för små familjer r.f.:
Verksamhet för små familjerfinska _ engelska
Underhållsbidrag
Båda föräldrarna bär ansvaret för underhållet av ett barn under 18 år, även om de inte bor tillsammans.
När föräldrarna skiljer sig ska de komma överens om underhållet av barnet samt om eventuellt underhållsbidrag (elatusapu).
Underhållsbidragets belopp beräknas utifrån barnets underhållsbehov och föräldrarnas underhållsförmåga.
Med barnets underhållsbehov avses det penningbelopp som försörjningen av barnet kostar varje månad.
I beloppet ingår till exempel utgifter för mat och kläder samt eventuella dagvårdsavgifter.
Barnets underhållsbehov delas mellan föräldrarna enligt deras underhållsförmåga.
Underhållsförmågan beräknas genom att dra av skatter och övriga obligatoriska utgifter av inkomsterna.
Du kan be om hjälp med att beräkna underhållsbehovet hos barnatillsyningsmannen (lastenvalvoja) i din hemkommun.
Det är bra att upprätta ett skriftligt avtal om underhållsbidraget som socialnämnden bekräftar.
Ett avtal som bekräftats på detta sätt är lika officiellt som ett domstolsbeslut.
Begär bekräftande av avtalet hos barnatillsyningsmannen i din hemkommun.
Om föräldrarna inte kan enas om underhållsbidraget kan de få hjälp i form av medling i familjefrågor.
I sista hand avgörs ärendet i tingsrätten.
Mer information om medling i familjefrågor hittar du på InfoFinlands sida Skilsmässa.
Underhållsstöd
I vissa situationer kan den förälder som bor med barnet ansöka om underhållsstöd (elatustuki) vid FPA.
Du kan ansöka om underhållsstöd från Fpa i följande situationer:
Den underhållsskyldiga föräldern har inte betalat det bekräftade underhållsbidraget (Fpa indriver det hos denne senare).
Underhållsbidraget har på grund av förälderns ekonomiska situation fastställts till ett belopp som underskrider underhållsstödet.
Det har på grund av förälderns ekonomiska situation fastställts att inget underhållsbidrag betalas.
Faderskapet har inte fastställts för ett barn fött utom äktenskapet.
Du kan få underhållsstöd om du bor stadigvarande i Finland.
Du kan få underhållsstöd också om du har flyttat till Finland från ett annat EU- eller EES-land eller Schweiz för att arbeta.
Också barnet för vilket man söker underhållsstöd ska bo i Finland.
Du får mer information om underhållsstödet på Fpa.
Underhållsbidrag och underhållsstödfinska _ svenska _ engelska
Skilsmässa i Finlandengelska _ ryska _ estniska
I Finland är det vanligt med familjer med en förälder.
Ett barn kan födas utom äktenskapet eller också är dess föräldrar skilda.
I familjer med en förälder bor en av föräldrarna med sina barn utan make eller maka.
Föräldern kan då ha antingen ensam eller gemensam vårdnad om barnet.
Som ensamstående förälder har man själv ansvaret för fostran av barnet.
Om föräldrarna däremot har gemensam vårdnad (yhteishuoltaja) kommer föräldrarna tillsammans överens om barnets angelägenheter.
Föräldrar som har gemensam vårdnad beslutar tillsammans om många saker. Dessa är barnets
bostadsort
fostran
språk
religion
utbildning
hälsovård
disponering av barnets egendom
Gemensam vårdnad förutsätter att barnets föräldrar klarar av att tillsammans agera för barnets bästa.
Till exempel för en passansökan behövs båda föräldrarnas tillstånd.
En ensamstående förälder fattar på egen hand alla beslut som rör barnet.
Myndigheter såsom daghem eller skola ger information om barnet endast till vårdnadshavaren.
Den andra föräldern får dock bestämma om vården och fostran av barnet när barnet är hos honom eller henne.
Vid skilsmässa eller när sambor flyttar isär måste föräldrarna besluta om barnets vårdnad, underhåll, boende och umgängesrätt.
Läs mer på InfoFinlands sida Barn vid skilsmässa.
Man kan också adoptera ett barn ensam.
Om du vill adoptera ett barn på egen hand, fråga om råd vid socialbyrån i din hemkommun.
Föreningen för familjer med en förälder (Yhden Vanhemman Perheiden Liitto) ger information och ordnar aktiviteter för familjer med en förälder.
På Finlex webbplats kan du läsa lagen angående vårdnad om barn och umgängesrätt.
Föreningen för små familjer är en medborgarorganisation som grundats av ensamstående föräldrar och som erbjuder aktiviteter för medlemsfamiljerna.
Lagen angående vårdnad om barn och umgängesrättfinska _ svenska _ engelska
linkkiFöreningen för familjer med en förälder r.f.:
Information för familjer med en förälderfinska
linkkiFöreningen för små familjer r.f.:
Verksamhet för små familjerfinska _ engelska
Underhållsbidrag
Båda föräldrarna bär ansvaret för underhållet av ett barn under 18 år, även om de inte bor tillsammans.
När föräldrarna skiljer sig ska de komma överens om underhållet av barnet samt om eventuellt underhållsbidrag (elatusapu).
Underhållsbidragets belopp beräknas utifrån barnets underhållsbehov och föräldrarnas underhållsförmåga.
Med barnets underhållsbehov avses det penningbelopp som försörjningen av barnet kostar varje månad.
I beloppet ingår till exempel utgifter för mat och kläder samt eventuella dagvårdsavgifter.
Barnets underhållsbehov delas mellan föräldrarna enligt deras underhållsförmåga.
Underhållsförmågan beräknas genom att dra av skatter och övriga obligatoriska utgifter av inkomsterna.
Du kan be om hjälp med att beräkna underhållsbehovet hos barnatillsyningsmannen (lastenvalvoja) i din hemkommun.
Det är bra att upprätta ett skriftligt avtal om underhållsbidraget som socialnämnden bekräftar.
Ett avtal som bekräftats på detta sätt är lika officiellt som ett domstolsbeslut.
Begär bekräftande av avtalet hos barnatillsyningsmannen i din hemkommun.
Om föräldrarna inte kan enas om underhållsbidraget kan de få hjälp i form av medling i familjefrågor.
I sista hand avgörs ärendet i tingsrätten.
Mer information om medling i familjefrågor hittar du på InfoFinlands sida Skilsmässa.
Underhållsstöd
I vissa situationer kan den förälder som bor med barnet ansöka om underhållsstöd (elatustuki) vid FPA.
Du kan ansöka om underhållsstöd från Fpa i följande situationer:
Den underhållsskyldiga föräldern har inte betalat det bekräftade underhållsbidraget (Fpa indriver det hos denne senare).
Underhållsbidraget har på grund av förälderns ekonomiska situation fastställts till ett belopp som underskrider underhållsstödet.
Det har på grund av förälderns ekonomiska situation fastställts att inget underhållsbidrag betalas.
Faderskapet har inte fastställts för ett barn fött utom äktenskapet.
Du kan få underhållsstöd om du bor stadigvarande i Finland.
Du kan få underhållsstöd också om du har flyttat till Finland från ett annat EU- eller EES-land eller Schweiz för att arbeta.
Också barnet för vilket man söker underhållsstöd ska bo i Finland.
Du får mer information om underhållsstödet på Fpa.
Underhållsbidrag och underhållsstödfinska _ svenska _ engelska
Skilsmässa i Finlandengelska _ ryska _ estniska
Kommunerna måste ordna de särskilda tjänster som handikappade behöver.
Dessa särskilda tjänster är till exempel färdtjänst, hjälpmedel eller en personlig assistent.
Syftet med tjänsterna är att hjälpa den handikappade att vara delaktig i samhället och underlätta livet med handikappet.
Om du har uppehållstillstånd och hemkommun i Finland har du rätt att använda de tjänster som kommunen tillhandahåller.
Du får mer information om rätten till hemkommun på InfoFinlands sida Hemkommun i Finland.
linkkiStödcentralen Hilma för handikappade invandrare:
Serviceguide för handikappade invandrare(pdf, 797,26)finska _ engelska _ ryska _ arabiska
linkkiInstitutet för hälsa och välfärd:
Handbok för handikappservicefinska _ svenska
linkkiSocial- och hälsovårdsministeriet:
Handikappservice och stödåtgärderfinska _ svenska _ engelska
Söka tjänster
Tjänsterna för handikappade fås oftast endast med ett läkarintyg (lääkärintodistus).
Besök till exempel din egen hälsostation för en hälsoundersökning.
När du har ett läkarintyg ska du kontakta socialbyrån i din hemkommun.
I kommunen finns en socialarbetare som ansvarar för tjänsterna för handikappade.
Han eller hon ger dig råd och hjälp när du ansöker om tjänster.
Syftet med serviceplanen är att reda ut vilken handikappservice du behöver.
Därefter tas beslut om tjänsterna, och du kan överklaga beslutet om du inte är nöjd med de tjänster som du har beviljats.
Boende
Kommunerna ordnar stödboende och serviceboende för handikappade personer som behöver stöd och hjälp i sitt boende.
Läs mer på InfoFinlands sida Stöd- och serviceboende.
Hjälpmedel
Hälsostationen och centralsjukhuset bekostar de hjälpmedel som ges som medicinsk rehabilitering (lääkinnällinen kuntoutus).
Det innebär att du inte behöver betala för de hjälpmedel som du behöver för att klara dig i vardagen.
Sådana kostnadsfria hjälpmedel är till exempel rullstolar, hörselskadades hörselapparater samt synskadades vita käppar och ledahundar.
Om du måste låta utföra ändringsarbeten i din bostad eller montera fasta hjälpmedel i bostaden kan du få ersättning för dessa av kommunen.
Ändringsarbetena kan vara till exempel ombyggnad av bostaden så att den blir tillgänglig för rullstol.
Fasta hjälpmedel kan till exempel vara olika typer av lyftanordningar samt brandvarnare och dörrklocka för hörselskadade, där ljudet har ersatts med lampor.
Socialarbetaren som ansvarar för handikapptjänster i din hemkommun bedömer tillsammans med dig om du behöver göra ändringsarbeten i din bostad.
FPA kan betala sådana hjälpmedel som du behöver för arbete eller studier.
Hjälpmedel ges till personer som inte klarar av arbete eller studier utan dem eller om det är mycket svårt att studera utan hjälpmedel.
Du kan fråga vid närmaste FPA-byrå hur du kan få hjälpmedel.
linkkiInstitutet för hälsa och välfärd:
Hjälpmedel för att röra sigfinska _ svenska
Hjälpmedel för arbete och studierfinska _ svenska _ engelska
Att röra sig
Om du på grund av ditt handikapp inte kan använda kollektivtrafiken kan du ha rätt till färdtjänst (kuljetuspalvelu).
Vid behov kan du även få en följeslagare (saattaja), d.v.s. en person som assisterar dig på resor.
Du kan få färdtjänst och följeslagare på resor som anknyter till arbete, studier eller fritid.
Du kan söka färdtjänst hos en socialarbetare inom handikappservicen i din hemkommun.
Du betalar för färdtjänsten enligt kollektivtrafikens taxa.
På grund av ditt handikapp kan du även få rabatt på kollektivtrafikens biljettpriser.
Du kan fråga om detta på socialbyrån i din hemkommun.
linkkiInstitutet för hälsa och välfärd:
Färdtjänst och följeslagartjänstfinska _ svenska
Assistentservice
Om du på grund av ditt handikapp behöver mycket hjälp med det vanliga livet kan du få en personlig assistent (henkilökohtainen avustaja).
Assistenten kan hjälpa dig till exempel med att laga mat, handla, på din arbetsplats, i dina studier eller dina hobbyer.
Din hemkommun betalar assistentens lön.
Du kan ansöka om en assistent vid socialbyrån i din hemkommun.
linkkiInstitutet för hälsa och välfärd:
Personlig assistansfinska _ svenska
Tolktjänster
Tolkning för en handikappad är inte det samma som språktolkning.
Du har rätt att använda tolktjänst (tulkkauspalvelu) för handikappade om du har
en hörselskada eller
en syn- och hörselskada eller
en talskada
och om du på grund av din skada behöver hjälp av en tolk
för att arbeta,
studera efter grundläggande studier,
uträtta ärenden,
vid social delaktighet,
Du kan ansöka om tolktjänst vid FPA.
Om du inte förstår finska eller det finska teckenspråket kan du också behöva en annan tolk.
Finländska handikapptolkar kan inte nödvändigtvis de teckenspråk som används i andra länder.
FPA ordnar inte en annan tolk.
När du sköter ärenden med myndigheter, kom alltid ihåg att bekräfta tolksbehovet.
Det åligger myndigheten med vilken du sköter ärenden att ordna tolktjänsten.
Om du blir kallad till hälsovården, kom ihåg att på förhand ange att du behöver en tolk.
Om du söker dig till jourmottagnignen eller läkaren, kan du beställa en tolk vid FPA.
Tolktjänster för handikappadefinska _ svenska
Rehabilitering
Om du har ett gravt handikapp och är under 65 år kan FPA ordna krävande medicinsk rehabilitering (vaativa lääkinnällinen kuntoutus) och ersätta en del av kostnaderna för rehabiliteringen.
Du kan få rehabilitering om ditt handikapp orsakar stora svårigheter att klara av vardagen i hemmet, skolan eller arbetet.
Medicinsk rehabilitering kan ordnas i ett rehabiliteringscenter eller som öppen terapi. Under den öppna terapin kan du bo hemma.
Målet med rehabiliteringen är att hjälpa dig att klara dig bättre i vardagen.
Om du inte kan få krävande medicinsk rehabilitering via FPA ska din hemkommun ordna rehabilitering för dig.
Läs mer på InfoFinlands sida Rehabilitering.
Krävande medicinsk rehabiliteringfinska _ svenska _ engelska
Att ansöka om medicinsk rehabiliteringfinska _ svenska _ engelska
Särskilda tjänster för utvecklingsstörda
Särskilda tjänster för utvecklingsstörda är bland annat
boendetjänster
familjevård
anstaltsvård
arbetsverksamhet och dagverksamhet.
Boendetjänster (asumispalvelu) innebär att en utvecklingsstörd person kan bo i sin egen bostad och där få olika typer av hjälp och stöd.
Läs mer på InfoFinlands sida Stöd- och serviceboende.
Familjevård (perhehoito) innebär att en person vårdas, fostras eller omhändertas i ett privat hem utanför det egna hemmet.
En utvecklingsstörd person som behöver vård kan bo i ett familjehem.
Man kan också bo tillfälligt i ett familjehem.
Familjevård kan även ordnas i den vårdbehövandes eget hem.
Om en utvecklingsstörd person behöver kontinuerlig vård och inte kan få det hemma eller i en servicebostad kan han eller hon även bo på en anstalt (laitos).
Man kan också bo korta tider i en anstalt.
Kommunerna ordnar arbetsverksamhet och dagverksamhet för handikappade personer.
I arbetsverksamheten (työtoiminta) ingår lätt arbete.
Dagverksamheten (päivätoiminta) är avsedd för svårt handikappade personer som inte kan delta i arbetsverksamheten.
Dagverksamheten kan omfatta till exempel matlagning, motion, samtal och friluftsliv.
På internet finns en databank för utvecklingsstörda (Kehitysvammahuollon tietopankki) med mycket nyttig information om utvecklingsstörningar och tjänster för handikappade.
Tjänsten är finskspråkig.
Boendeservice för utvecklingsstördafinska
Utvecklingsstörda och arbetefinska
Dagverksamhetfinska
Definition av en familj
I Finland utgörs en familj av
makar
sambor
ogifta barn under 18 och deras vårdnadshavare som bor i Finland
I Finland uppfattas en familj i snävare bemärkelse än i många andra länder.
I Finland anses oftast kärnfamiljen, d.v.s. föräldrarna och barnen utgöra en familj.
Till exempel om mor- eller farföräldrarna, föräldrarna och barnen bor i samma lägenhet räknas officiellt bara föräldrarna och barnen till samma familj.
Mor- eller farföräldrarna bildar en egen familj.
En familj kan ha barn eller bestå av ett barnlöst par.
De vuxna i familjen kan vara av samma eller olika kön.
En familj bildas också av en ensamstående mor eller far och hens barn.
Med ombildade familjer avses ett par som bor tillsammans med ett eller flera barn från parets tidigare förhållanden.
Också parets gemensamma barn kan bo med familjen.
Om du är frånskild kan du gifta om dig utan tillstånd från din före detta maka eller make.
Du behöver inte tillstånd från din före detta maka eller make för att ingå ett nytt äktenskap även om du och din före detta maka eller make har barn tillsammans.
Regnbågsfamiljer
Regnbågsfamiljer är familjer som bildas av homosexuella, lesbiska, bi- och transsexuella föräldrar och deras barn.
De är till exempel familjer som bildas av två kvinnor eller två män samt familjer med fler än två föräldrar
Gifta makar av samma kön har rätt att adoptera ett barn och rätt till adoption inom familjen.
Adoption inom familjen betyder att makan/maken adopterar sin makas/makes barn och blir officiellt barnets andra förälder.
I Finland kan ett barn ha högst två juridiska föräldrar.
Om du planerar adoption inom familjen ska du kontakta socialbyrån i din hemkommun.
Regnbågsfamiljer rf är en organisation som stöder regnbågsfamiljer samt ger råd och ordnar verksamhet för dem.
Kontaktuppgifterna hittar du på organisationens webbplats.
linkkiRegnbågsfamiljer:
Stöd och verksamhet för regnbågsfamiljerfinska
Underhållsskyldighet
Enligt Finlands lag är föräldrarna förpliktade att ta hand om sina minderåriga barn ekonomiskt och gifta par om varandra.
Familjemedlemmarnas underhållsskyldighet sträcker sig inte till släktingar, till exempel vuxna syskon eller mor- eller farföräldrar.
I Finland utgår man alltså inte från att enskilda människor tar hand om sådana släktingar som har det dåligt ställt ekonomiskt.
Stödet kommer från samhället i form av den sociala tryggheten.
Hushåll
Till samma hushåll hör alla som stadigvarande bor i samma bostad.
Mer information om ämnet hushåll finns på InfoFinlands sida boende.
Parförhållande
Ett par kan välja om de vill leva tillsammans i ett samboförhållande eller i ett äktenskap.
Det är bra att beakta att parförhållandets form påverkar makarnas rättigheter och skyldigheter, frågor som rör egendom och arv, vårdnad om och underhåll av barn samt adoption.
Råd i frågor som rör familjen
Väestöliitto tillhandahåller rådgivning telefonledes och via e-post när du behöver samtalsstöd i frågor som rör barnuppfostran eller relationerna i familjen.
Samtal tas emot på följande språk:
ryska och engelska tfn 050 325 7173
Läs mer på InfoFinlands sida Fostran av barn i Finland.
Läs mer på InfoFinlands sida Problem i familjen.
Till Finland på grund av familjebandfinska _ svenska _ engelska
linkkiBefolkningsförbundet:
Rådgivning till invandrare telefonledes och via e-postfinska _ svenska _ engelska
Handbok för familjer med två kulturer (pdf, 4,74 Mt)finska _ engelska _ ryska _ franska _ spanska _ thai
Definition av en familj
I Finland utgörs en familj av
makar
sambor
ogifta barn under 18 och deras vårdnadshavare som bor i Finland
I Finland uppfattas en familj i snävare bemärkelse än i många andra länder.
I Finland anses oftast kärnfamiljen, d.v.s. föräldrarna och barnen utgöra en familj.
Till exempel om mor- eller farföräldrarna, föräldrarna och barnen bor i samma lägenhet räknas officiellt bara föräldrarna och barnen till samma familj.
Mor- eller farföräldrarna bildar en egen familj.
En familj kan ha barn eller bestå av ett barnlöst par.
De vuxna i familjen kan vara av samma eller olika kön.
En familj bildas också av en ensamstående mor eller far och hens barn.
Med ombildade familjer avses ett par som bor tillsammans med ett eller flera barn från parets tidigare förhållanden.
Också parets gemensamma barn kan bo med familjen.
Om du är frånskild kan du gifta om dig utan tillstånd från din före detta maka eller make.
Du behöver inte tillstånd från din före detta maka eller make för att ingå ett nytt äktenskap även om du och din före detta maka eller make har barn tillsammans.
Regnbågsfamiljer
Regnbågsfamiljer är familjer som bildas av homosexuella, lesbiska, bi- och transsexuella föräldrar och deras barn.
De är till exempel familjer som bildas av två kvinnor eller två män samt familjer med fler än två föräldrar
Gifta makar av samma kön har rätt att adoptera ett barn och rätt till adoption inom familjen.
Adoption inom familjen betyder att makan/maken adopterar sin makas/makes barn och blir officiellt barnets andra förälder.
I Finland kan ett barn ha högst två juridiska föräldrar.
Om du planerar adoption inom familjen ska du kontakta socialbyrån i din hemkommun.
Regnbågsfamiljer rf är en organisation som stöder regnbågsfamiljer samt ger råd och ordnar verksamhet för dem.
Kontaktuppgifterna hittar du på organisationens webbplats.
linkkiRegnbågsfamiljer:
Stöd och verksamhet för regnbågsfamiljerfinska
Underhållsskyldighet
Enligt Finlands lag är föräldrarna förpliktade att ta hand om sina minderåriga barn ekonomiskt och gifta par om varandra.
Familjemedlemmarnas underhållsskyldighet sträcker sig inte till släktingar, till exempel vuxna syskon eller mor- eller farföräldrar.
I Finland utgår man alltså inte från att enskilda människor tar hand om sådana släktingar som har det dåligt ställt ekonomiskt.
Stödet kommer från samhället i form av den sociala tryggheten.
Hushåll
Till samma hushåll hör alla som stadigvarande bor i samma bostad.
Mer information om ämnet hushåll finns på InfoFinlands sida boende.
Parförhållande
Ett par kan välja om de vill leva tillsammans i ett samboförhållande eller i ett äktenskap.
Det är bra att beakta att parförhållandets form påverkar makarnas rättigheter och skyldigheter, frågor som rör egendom och arv, vårdnad om och underhåll av barn samt adoption.
Råd i frågor som rör familjen
Väestöliitto tillhandahåller rådgivning telefonledes och via e-post när du behöver samtalsstöd i frågor som rör barnuppfostran eller relationerna i familjen.
Samtal tas emot på följande språk:
ryska och engelska tfn 050 325 7173
Läs mer på InfoFinlands sida Fostran av barn i Finland.
Läs mer på InfoFinlands sida Problem i familjen.
Till Finland på grund av familjebandfinska _ svenska _ engelska
linkkiBefolkningsförbundet:
Rådgivning till invandrare telefonledes och via e-postfinska _ svenska _ engelska
Handbok för familjer med två kulturer (pdf, 4,74 Mt)finska _ engelska _ ryska _ franska _ spanska _ thai
Enligt finsk lag får ingen diskrimineras på grund av ett handikapp.
Handikappade personer har rätt att leva ett normalt liv, till exempel studera, arbeta och bilda familj.
Finland har ratificerat FN:s konvention om rättigheter för personer med funktionshinder.
Handikappade personer kan ha svårt att klara av det dagliga livet på grund av sitt handikapp eller sin sjukdom.
Kommunerna måste tillhandahålla handikappade de tjänster som de behöver.
Sådana tjänster är till exempel färd- och assistenttjänsterna.
Om du har uppehållstillstånd och hemkommun i Finland, har du rätt till kommunens tjänster för handikappade.
Läs mer om tjänsterna för handikappade och om att ansöka dem på InfoFinlands sida Tjänster för handikappade.
Handikapporganisationer
I Finland finns flera organisationer som arbetar för att förbättra handikappade personers ställning i samhället.
Hos dessa organisationer kan du få råd och hjälp till exempel vid ansökan om tjänster.
Många organisationer erbjuder fritidsverksamhet och kamratstöd till personer i alla åldrar.
Du hittar kontaktuppgifterna till organisationerna på Handikappforums webbplats.
I Finland finns även stödcentret
Hilma för handikappade invandrare som erbjuder servicevägledning och rådgivning för handikappade invandrare och långtidssjuka.
linkkiStödcentralen Hilma för handikappade invandrare:
Stöd och hjälp för handikappade invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ persiska _ arabiska _ kurdiska
Handikapporganisationer i Finlandfinska _ svenska
Synskadade
Om du är blind eller har nedsatt syn kan du få tjänster för synskadade.
Om du behöver hjälpmedel ska du först besöka din egen hälsostation för en läkarundersökning.
Läkaren bedömer din synskada och därefter kan du få hjälpmedel i form av medicinsk rehabilitering.
Läs mer på InfoFinlands sida Tjänster för handikappade.
Om du på grund av ditt handikapp behöver till exempel en speciell dator eller särskilda hushållsapparater kan du få understöd för detta vid socialbyrån i din hemkommun.
Detta är dock prövningsbaserat, med andra ord är det inte säkert att du får stödet.
På biblioteket för synskadade Celia kan du låna ljudböcker, punktskriftsböcker, e-böcker och reliefbilder.
Biblioteket producerar även läroböcker för synskadade skolelevers och studerandes behov.
Synskadades förbund är en organisation som arbetar för att förbättra synskadades ställning i samhället.
Förbundet erbjuder även mycket nyttig information och tjänster till synskadade.
De vanligaste hjälpmedlen för synskadadefinska
linkkiCelia:
De synskadades bibliotekfinska _ svenska _ engelska
Hörselskadade
Personer med en hörselskada är döva eller har nedsatt hörsel.
Många kommunicerar med teckenspråk.
I Finland används det finska och det finlandssvenska teckenspråket.
Personer med en hörselskada använder ofta även hörapparater.
Om du behöver hjälpmedel ska du först besöka din egen hälsostation för en läkarundersökning.
Läkaren bedömer din hörselskada och därefter kan du få hjälpmedel i form av medicinsk rehabilitering.
Du kan till exempel få ett brandlarm avsett för hörselskadade och en texttelefon för att kunna bo tryggt i ditt hem.
Ansök om dessa hjälpmedel vid socialbyrån i din hemkommun.
Om du behöver det på grund av din hörselskada kan du få tolktjänster till exempel i arbetet, studierna eller när du ska sköta ärenden.
Tolkning kan ges på teckenspråk eller vara skrivtolkning.
Ansök om rätten att använda tolktjänster hos FPA.
Läs mer om hjälpmedel och tolktjänster på InfoFinlands sida Tjänster för handikappade.
På internet finns ordboken för det finska teckenspråket, Suvi.
Hörselförbundet och Finlands Dövas Förbund är organisationer som arbetar för att förbättra hörselskadade personers ställning i samhället.
De erbjuder även mycket nyttig information och tjänster till hörselskadade.
linkkiFinska Hörselförbundet rf:
Hjälpmedel för hörselnfinska
linkkiFinska Hörselförbundet rf:
Hörselapparatfinska
Tolktjänster för handikappadefinska _ svenska
Ordbok i det finska teckenspråketfinska
linkkiFinska Hörselförbundet rf:
Information om Hörselförbundetfinska
linkkiFinlands Dövas Förbund rf:
Information om Finlands Dövas Förbundfinska _ svenska _ engelska
linkkiDövas folkhögskola:
Utbildning för döva invandrarefinska _ svenska _ engelska
Rörelsehandikappade
En rörelsehandikappad person kan inte röra sig självständigt eller utan hjälpmedel.
En rörelsenedsättning kan bero på en sjukdom, ett olycksfall eller genetiska orsaker.
Om du behöver hjälpmedel ska du först besöka din egen hälsostation för en läkarundersökning.
Läkaren bedömer din rörelsenedsättning och därefter kan du få hjälpmedel i form av medicinsk rehabilitering.
Om det måste göras förändringsarbeten eller installeras fasta hjälpmedel i din bostad kan du få ersättning för detta av din hemkommun.
Bostaden kan till exempel byggas om så att du kan röra dig med en rullstol i den.
Fasta hjälpmedel är till exempel stödhandtag, ramper och elektriska dörrar.
Läs mer om hjälpmedel och förändringsarbeten på InfoFinlands sida Tjänster för handikappade.
linkkiInvalidförbundet:
Stöd och verksamhet för rörelsehindradefinska
Utvecklingsstörda
En utvecklingsstörning gör det svårare att lära sig och förstå nya saker.
För en utvecklingsstörd person är det svårare att lära sig och minnas saker än för andra.
Utvecklingsstörningen upptäcks ofta i barndomen eller ungdomen.
För en utvecklingsstörd person finns olika slags specialtjänster.
Sådana är till exempel boendetjänster, arbetsverksamhet och dagverksamhet.
Läs mer om tjänsterna för utvecklingsstörda på InfoFinlands sida Tjänster för handikappade.
Det finns även många organisationer där du kan få information och stöd.
Du hittar mer information till exempel på Kehitysvammaliittos och Kehitysvammaisten Tukiliittos webbplatser.
Information för utvecklingsstörda och anhörigafinska
linkkiFörbundet Utvecklingsstörning:
Utvecklingsstördas intressebevakningsorganisationfinska _ engelska
linkkiUtvecklingsstördas intressebevakningsorganisation:
Utvecklingsstördas intressebevakningsorganisationfinska _ svenska _ engelska
Handikappbidrag för barn under 16 år
Ett barn under 16 år kan få handikappbidrag (vammaistuki) om hen på grund av sitt handikapp eller sin sjukdom behöver regelbunden vård, omsorg och rehabilitering under minst sex månaders tid.
Du ansöker om handikappbidrag för barn under 16 år vid FPA.
Handikappbidraget beviljas vanligtvis för en bestämd period.
När perioden har gått kan man ansöka om förlängning för bidraget.
Handikappbidrag för barnfinska _ svenska _ engelska
Specialvårdspenning
Du kan få specialvårdspenning från FPA om
ditt barn är under 16 år och vårdas på sjukhus eller
om du tar hand om barnet i hemmet och hemvården ansluter sig till barnets sjukhusvård eller
om utbetalningen av ditt arbetsmarknadsstöd avbryts tillfälligt eftersom du på grund av vården av ditt barn inte kan delta i integrationsåtgärderna eller
ditt barn provar på att återvända till skolan eller barnomsorgen.
Specialvårdspenning för barn under 16 årfinska _ svenska _ engelska
Rehabilitering för barn
FPA ordnar rehabiliteringen och ersätter kostnaderna för den.
Rehabiliteringen kan omfatta många olika slags aktiviteter.
Den kan till exempel bestå av fysioterapi eller olika kurser där man lär sig att leva med sitt handikapp.
FPA kan även ordna rehabilitering som behovsprövad rehabilitering (harkinnanvarainen kuntoutus).
Behovsprövad rehabilitering har som mål att förbättra arbets- eller funktionsförmågan.
Om barnet inte kan få krävande medicinska rehabilitering från FPA, ska rehabiliteringen ordnas av hemkommunen.
Krävande medicinsk rehabiliteringfinska _ svenska _ engelska
Handikappade barns skolgång
Ett handikappat barn har rätt till skolgång i närliggande skola.
Ett handikappat barn kan få specialundervisning om barnets handikapp försvårar inlärningen.
Barnet kan vid behov även få ett skolgångsbiträde (koulunkäyntiavustaja).
FPA kan betala dyra och krävande hjälpmedel (apuväline) som det handikappade barnet behöver för sin skolgång.
Sådana hjälpmedel är till exempel datorer och tilläggsutrustning till datorer.
Barnet kan också få hjälpmedel om han eller hon inte kan studera utan dem eller om det är mycket svårt utan dem.
Hjälpmedel kan fås tidigast när barnet går i grundskolans årskurs sju.
Hjälpmedel för arbete och studierfinska _ svenska _ engelska
Handikappade barns fritid
Information om hobbymöjligheterna på din hemort får du till exempel vid idrotts- och kulturförvaltningen i din hemkommun.
Också handikapporganisationer tillhandahåller många slags hobbyverksamheter.
Till exempel föreningen för handikappidrott och -motion i Finland, VAU ry, ordnar olika idrotts- och motionsevenemang.
linkkiDe Utvecklingsstördas Stödförbund (VAU):
Motion för handikappade barn och ungafinska _ svenska _ engelska
Handikappbidrag för barn under 16 år
Ett barn under 16 år kan få handikappbidrag (vammaistuki) om hen på grund av sitt handikapp eller sin sjukdom behöver regelbunden vård, omsorg och rehabilitering under minst sex månaders tid.
Du ansöker om handikappbidrag för barn under 16 år vid FPA.
Handikappbidraget beviljas vanligtvis för en bestämd period.
När perioden har gått kan man ansöka om förlängning för bidraget.
Handikappbidrag för barnfinska _ svenska _ engelska
Specialvårdspenning
Du kan få specialvårdspenning från FPA om
ditt barn är under 16 år och vårdas på sjukhus eller
om du tar hand om barnet i hemmet och hemvården ansluter sig till barnets sjukhusvård eller
om utbetalningen av ditt arbetsmarknadsstöd avbryts tillfälligt eftersom du på grund av vården av ditt barn inte kan delta i integrationsåtgärderna eller
ditt barn provar på att återvända till skolan eller barnomsorgen.
Specialvårdspenning för barn under 16 årfinska _ svenska _ engelska
Rehabilitering för barn
FPA ordnar rehabiliteringen och ersätter kostnaderna för den.
Rehabiliteringen kan omfatta många olika slags aktiviteter.
Den kan till exempel bestå av fysioterapi eller olika kurser där man lär sig att leva med sitt handikapp.
FPA kan även ordna rehabilitering som behovsprövad rehabilitering (harkinnanvarainen kuntoutus).
Behovsprövad rehabilitering har som mål att förbättra arbets- eller funktionsförmågan.
Om barnet inte kan få krävande medicinska rehabilitering från FPA, ska rehabiliteringen ordnas av hemkommunen.
Krävande medicinsk rehabiliteringfinska _ svenska _ engelska
Handikappade barns skolgång
Ett handikappat barn har rätt till skolgång i närliggande skola.
Ett handikappat barn kan få specialundervisning om barnets handikapp försvårar inlärningen.
Barnet kan vid behov även få ett skolgångsbiträde (koulunkäyntiavustaja).
FPA kan betala dyra och krävande hjälpmedel (apuväline) som det handikappade barnet behöver för sin skolgång.
Sådana hjälpmedel är till exempel datorer och tilläggsutrustning till datorer.
Barnet kan också få hjälpmedel om han eller hon inte kan studera utan dem eller om det är mycket svårt utan dem.
Hjälpmedel kan fås tidigast när barnet går i grundskolans årskurs sju.
Hjälpmedel för arbete och studierfinska _ svenska _ engelska
Handikappade barns fritid
Information om hobbymöjligheterna på din hemort får du till exempel vid idrotts- och kulturförvaltningen i din hemkommun.
Också handikapporganisationer tillhandahåller många slags hobbyverksamheter.
Till exempel föreningen för handikappidrott och -motion i Finland, VAU ry, ordnar olika idrotts- och motionsevenemang.
linkkiDe Utvecklingsstördas Stödförbund (VAU):
Motion för handikappade barn och ungafinska _ svenska _ engelska
Rehabilitering som ordnas av kommunerna
Kommunerna ordnar medicinsk rehabilitering till exempel vid hälsovårdscentraler och i sjukhus.
Du kan få kommunal rehabilitering om du har hemkommun i Finland.
Kommunernas rehabilitering omfattar:
rådgivning om rehabilitering
undersökningar för att fastställa rehabiliteringsbehovet
vård för att förbättra arbets- och funktionsförmågan
rehabiliteringsperioder
hjälpmedelstjänster
anpassningsträning
rehabiliteringshandledning
Mer information om kommunens rehabiliteringstjänster får du vid din egen hälsostation.
Rehabilitering som ordnas av FPA
FPA:s rehabilitering kan vara:
rehabilitering för gravt handikappade
behovsprövad rehabilitering
rehabiliteringspsykoterapi
Yrkesinriktad rehabilitering ordnas av arbetspensionsanstalter (työeläkelaitokset) och FPA (Kela).
Medicinsk rehabilitering ordnas av kommunerna och FPA.
Om du lider av en yrkessjukdom eller har blivit skadad i ett olycksfall, kan du få rehabilitering från försäkringsbolaget (vakuutusyhtiö).
FPA kan betala ut understöd för psykoterapin, men du måste själv hitta en lämplig terapeut.
FPA:s rehabilitering är avsedd för personer som omfattas av den finländska sjukförsäkringen (sairausvakuutus).
Mer information om sjukförsäkringen får du på InfoFinlands sida Den sociala tryggheten i Finland.
Rehabilitering för arbete
Du kan få yrkesinriktad rehabilitering om du har sådana hälsoproblem som hindrar dig från att arbeta.
Du kan också få rehabilitering om du riskerar att tvingas sluta arbeta på grund av dina hälsoproblem.
Du har rätt till rehabilitering efter ett arbetsolycksfall.
Arbetspensionsanstalter ordnar yrkesinriktad rehabilitering för arbetstagare.
Du kan ansöka om rehabilitering vid arbetspensionsanstalten om du har arbetat fem år eller längre.
Fråga mer av de sakkunniga inom rehabiliteringsfrågor vid din arbetspensionsanstalt.
FPA ordnar yrkesinriktad rehabilitering för unga personer och vuxna som inte arbetar.
Yrkesinriktad rehabiliteringfinska _ svenska _ engelska
Att ansöka om yrkesinriktad rehabiliteringfinska _ svenska _ engelska
Rehabilitering för gravt handikappade
Om du är under 65 år och har på grund av sjukdom eller funktionsnedsättning stora svårigheter att klara av vardagen, till exempel om du har svårt att röra dig eller ta hand om dig själv, kan FPA ordna krävande medicinsk rehabilitering (vaativa lääkinnällinen kuntoutus) för dig.
Rehabiliteringen genomförs på ett sätt som passar just dig.
Du kan få rehabilitering till exempel vid en rehabiliteringsinrättning (kuntoutuslaitos).
Du kan också bo hemma och gå på rehabilitering därifrån.
Målet med rehabiliteringen är att stöda dig och dina närstående så att du kan föra ett aktivt liv.
Mer information om krävande medicinsk rehabilitering fås av FPA.
Krävande medicinsk rehabiliteringfinska _ svenska _ engelska
Att ansöka om medicinsk rehabiliteringfinska _ svenska _ engelska
Behovsprövad rehabilitering
Du kan få behovsprövad rehabilitering om ditt mål är att fortsätta arbeta, återgå till arbetet eller börja arbeta.
Du kan få behovsprövad rehabilitering om hälso- och sjukvården konstaterar att du har en skada eller sjukdom som kräver rehabilitering.
Behovsprövad rehabilitering kan till exempel omfatta
rehabiliteringskurser för personer med en viss sjukdom
kurser för anpassningsträning
Läs mer om de olika alternativen för behovsprövad rehabilitering på FPA:s webbplats.
Behovsprövad rehabiliteringfinska _ svenska
Psykoterapi som rehabilitering
Om du behöver psykoterapi som stöd för din arbets- eller studieförmåga, kan du eventuellt ansöka om rehabiliterande psykoterapi (kuntoutuspsykoterapia).
Villkor för att du ska få rehabiliterande psykoterapi är att
du har fått psykiatrisk vård i minst tre månader och
den vårdande psykiatern skriver ett utlåtande med rekommendation om rehabiliterande psykoterapi.
Lär mer om mentala tjänster på InfoFinlands sida Mental hälsa.
För personer i åldern 16–25 år kan den också omfatta musikterapi.
Terapi för unga kan också omfatta besök av föräldrar.
Du kan få understöd för terapin ett år i taget under högst tre år.
FPA ersätter högst 80 terapibesök om året och högst 200 besök under tre år.
För att få FPA:s bidrag för psykoterapi ska terapeuten ha rätt att använda psykoterapeutens yrkesbenämning och vara godkänd av FPA.
Rehabiliterande psykoterapifinska _ svenska _ engelska
linkkiFinlands Psykologiförbund:
Hur söker du dig till rehabilitering
När du behöver rehabilitering behöver du först ett läkarutlåtande.
Ta kontakt med din läkare, företagsläkare eller FPA.
Om du ansöker om krävande medicinsk rehabilitering behöver du dessutom en rehabiliteringsplan (kuntoutussuunnitelma).
När du har fått ett läkarutlåtande eller en rehabiliteringsplan kan du ansöka om rehabilitering vid din arbetspensionsanstalt eller FPA.
Du kan fråga vid kommunens hälsovårdstjänster arbetspensionsanstalten eller FPA om olika rehabiliteringsmöjligheter.
Mer information om FPA:s rehabiliteringar hittar du också på FPA:s webbplats.
Om du söker till rehabilitering som ordnas av FPA ska du lämna in din ansökan om rehabilitering till FPA innan rehabiliteringen börjar.
FPA ger ett skriftligt beslut om rehabilitering.
Sköta ärenden på Internetfinska _ svenska _ engelska
Kontaktuppgifter till FPAfinska _ svenska _ engelska
Elektronisk tidsbeställningfinska _ svenska _ engelska
Under rehabiliteringen kan du få rehabiliteringspenning (kuntoutusraha), om du är 16–67 år och om rehabiliteringen har som syfte att bevara din arbetsförmåga eller göra det möjligt för dig att återvända till arbetslivet eller komma in i arbetslivet.
För att få rehabiliteringspenning måste du också få ett rehabiliteringsbeslut (kuntoutuspäätös) till exempel från FPA eller företagshälsovården.
Du kan få rehabiliteringspenning på samma villkor också när din hemkommun ordnar din rehabilitering.
FPA kan delvis ersätta resorna till rehabiliteringen.
Rehabiliteringspenningfinska _ svenska _ engelska
Om du på grund av skada eller sjukdom inte kan arbeta kan du få invalidpension (työkyvyttömyyseläke).
Om du är blind eller rörelsehindrad kan du få invalidpension även om du skulle kunna arbeta.
Invalidpension betalas till 16–64-åringar.
Huruvida du får pensionen beror på hur länge du har bott i Finland.
Vanligtvis kan du få invalidpension när du har bott tre år i Finland.
Du kan söka invalidpension hos FPA.
Sjukpensionfinska _ svenska _ engelska
Handikappbidrag för vuxna
Om du har ett handikapp eller en sjukdom som försämrar din funktionsförmåga sammanhängande under minst ett år kan du få handikappbidrag (vammaistuki).
Du måste ha ett läkarintyg för att få handikappbidrag.
Handikappbidrag för vuxna betalas till 16–64-åringar.
Huruvida du får bidraget beror på hur länge du har bott i Finland.
Vanligtvis kan du få handikappbidrag när du har bott tre år i Finland.
Handikappbidragets storlek beror på hur svårt ditt handikapp är.
Du kan söka handikappbidrag hos FPA.
Handikappbidrag för vuxnafinska _ svenska _ engelska
Hälsa och rehabiliteringfinska _ svenska _ ryska _ estniska
Stöd för vård av en handikappad anhörig
Om du vårdar en handikappad närstående i hemmet kan du få stöd för närståendevård (omaishoidontuki) från din hemkommun.
För att få stöd måste du göra ett avtal om närståendevård med din kommun.
Du kan ansöka om stödet vid socialbyrån i din egen kommun.
linkkiNärståendevårdare och Vänner -Förbundet rf:
Handikappbidrag för barn och specialvårdpenning
Läs mer om handikappbidrag för barn och specialvårdpenning på InfoFinlands sida Ett handikappat barn.
Vårdbidrag för pensionstagare
En pensionär vars funktionsförmåga försämrats under sammanlagt minst ett år på grund av sjukdom eller skada kan få vårdbidrag för pensionstagare (eläkettä saavan hoitotuki).
Du kan få stöd om du på grund av ditt handikapp eller din sjukdom behöver kontinuerligt hjälp.
Hur stort stöd du får beror på hur mycket hjälp du behöver.
Vårdbidrag för pensionstagare kan sökas hos FPA.
Vårdbidrag för pensionstagarefinska _ svenska _ engelska
Bidrag för kläder och mat
Om ditt handikapp eller din sjukdom orsakar dig extra kostnader för mat eller kläder kan du ansöka om bidrag för kläder och mat (vaatetus- ja ravitsemustuki).
Du kan ansöka om bidraget vid socialbyrån i din hemkommun.
linkkiInstitutet för hälsa och välfärd:
Extra kostnader för kläder och matfinska _ svenska
Om du på grund av skada eller sjukdom inte kan arbeta kan du få invalidpension (työkyvyttömyyseläke).
Om du är blind eller rörelsehindrad kan du få invalidpension även om du skulle kunna arbeta.
Invalidpension betalas till 16–64-åringar.
Huruvida du får pensionen beror på hur länge du har bott i Finland.
Vanligtvis kan du få invalidpension när du har bott tre år i Finland.
Du kan söka invalidpension hos FPA.
Sjukpensionfinska _ svenska _ engelska
Handikappbidrag för vuxna
Om du har ett handikapp eller en sjukdom som försämrar din funktionsförmåga sammanhängande under minst ett år kan du få handikappbidrag (vammaistuki).
Du måste ha ett läkarintyg för att få handikappbidrag.
Handikappbidrag för vuxna betalas till 16–64-åringar.
Huruvida du får bidraget beror på hur länge du har bott i Finland.
Vanligtvis kan du få handikappbidrag när du har bott tre år i Finland.
Handikappbidragets storlek beror på hur svårt ditt handikapp är.
Du kan söka handikappbidrag hos FPA.
Handikappbidrag för vuxnafinska _ svenska _ engelska
Hälsa och rehabiliteringfinska _ svenska _ ryska _ estniska
Stöd för vård av en handikappad anhörig
Om du vårdar en handikappad närstående i hemmet kan du få stöd för närståendevård (omaishoidontuki) från din hemkommun.
För att få stöd måste du göra ett avtal om närståendevård med din kommun.
Du kan ansöka om stödet vid socialbyrån i din egen kommun.
linkkiNärståendevårdare och Vänner -Förbundet rf:
Handikappbidrag för barn och specialvårdpenning
Läs mer om handikappbidrag för barn och specialvårdpenning på InfoFinlands sida Ett handikappat barn.
Vårdbidrag för pensionstagare
En pensionär vars funktionsförmåga försämrats under sammanlagt minst ett år på grund av sjukdom eller skada kan få vårdbidrag för pensionstagare (eläkettä saavan hoitotuki).
Du kan få stöd om du på grund av ditt handikapp eller din sjukdom behöver kontinuerligt hjälp.
Hur stort stöd du får beror på hur mycket hjälp du behöver.
Vårdbidrag för pensionstagare kan sökas hos FPA.
Vårdbidrag för pensionstagarefinska _ svenska _ engelska
Bidrag för kläder och mat
Om ditt handikapp eller din sjukdom orsakar dig extra kostnader för mat eller kläder kan du ansöka om bidrag för kläder och mat (vaatetus- ja ravitsemustuki).
Du kan ansöka om bidraget vid socialbyrån i din hemkommun.
linkkiInstitutet för hälsa och välfärd:
Extra kostnader för kläder och matfinska _ svenska
Om du blir sjuk eller råkar ut för en olycka har du rätt att stanna hemma från arbetet.
Om du omfattas av den finländska sjukförsäkringen (sairausvakuutus) har du efter en självrisktid (omavastuuaika) rätt att söka sjukdagpenning (sairauspäiväraha) hos FPA (Kela).
Självrisktiden är vanligen den dag då du insjuknade och därpå följande nio vardagar.
Om din anställning har varat över en månad före insjuknandet betalar din arbetsgivare full lön för självrisktiden.
Sjukdagpenning betalas för högst 300 vardagar.
Den ska sökas inom två månader efter insjuknandet.
Du kan söka sjukdagpenning om du:
omfattas av den finländska sjukförsäkringen (sairausvakuutus): läs mer på InfoFinlands sida Den sociala tryggheten i Finland
är 16–67 år
är arbetsoförmögen på grund av din sjukdom
har arbetat tre månader som anställd, företagare eller yrkesutövare tre månader innan du insjuknade eller har tre månader innan du insjuknade varit heltidsstuderande, arbetslös arbetssökande, d.v.s. kund vid arbets- och näringsbyrån (työ- ja elinkeinotoimisto), sabbatsledig (sapattivapaa) eller alterneringsledig (vuorotteluvapaa).
Om du får lön under sjukledigheten, ansöker din arbetsgivare om sjukdagpenningen och då betalas sjukdagpenningen till din arbetsgivare.
Om du är sjuk en lång tid och din arbetsgivare inte längre betalar dig lön under sjukledigheten kan du söka FPA:s sjukdagpenning när lönen inte längre utbetalas.
Sjukdagpenningens belopp beror på inkomsterna.
Den beräknas oftast på basis av de arbetsinkomster som bekräftats i beskattningen.
Till exempel beaktas inte royaltyn och anställningsoptioner vid beräkning av dagpenningens belopp.
Om din inkomst har ökat kan du söka sjukdagpenning på basis av arbetsinkomsten under de senaste sex månaderna.
Du ska då bifoga till ansökan ett löneintyg för löner som du har fått.
Be om intyget av din arbetsgivare.
När du söker sjukdagpenning ska du bifoga till ansökan:
ett läkarintyg om arbetsoförmögenhet
ett löneintyg för de senaste sex månaderna om dina inkomster har ökat.
Mer information om sjukdagpenningen får du på FPA:s webbplats.
Om du är sjuk en lång tid ska du ta reda på om rehabilitering kan vara till nytta för dig.
Sjukdagpenningfinska _ svenska _ engelska
Att ansöka om sjukdagpenningfinska _ svenska _ engelska
Hälsa och rehabiliteringfinska _ svenska _ ryska _ estniska
Partiell sjukdagpenning
Den partiella sjukdagpenningen (osasairauspäiväraha) är avsedd för 16–67-åriga heltidsarbetande anställda eller företagare som omfattas av den sociala tryggheten i Finland.
Syftet med den partiella sjukdagpenningen är att du kan fortsätta att arbeta eller att återgå till arbetet trots att du har blivit sjuk.
Diskutera först med din läkare inom företagshälsovården och din arbetsgivare om möjligheten att söka partiell sjukdagpenning.
Företagshälsovårdsläkaren avgör om du kan deltidsarbeta medan du är sjuk.
När du söker partiell sjukdagpenning ska du bifoga till ansökan:
ett läkarintyg om arbetsoförmögenhet
ansökan om sjukdagpenning
en kopia av överenskommelsen mellan dig och din arbetsgivare om att du under en viss tid ska arbeta på deltid.
Arbetstidsarrangemanget och lönen ska framgå ur avtalet.
ett löneintyg för de senaste sex månaderna före insjuknandet om dina inkomster har ökat.
Partiell sjukdagpenning ska sökas inom två månader efter att du börjar arbeta på deltid.
Mer information om den partiella sjukdagpenningen får du på FPA:s webbplats.
Partiell sjukdagpenningfinska _ svenska _ engelska
Att ansöka om partiell sjukdagpenningfinska _ svenska _ engelska
Kommunerna måste ordna de särskilda tjänster som handikappade behöver.
Dessa särskilda tjänster är till exempel färdtjänst, hjälpmedel eller en personlig assistent.
Syftet med tjänsterna är att hjälpa den handikappade att vara delaktig i samhället och underlätta livet med handikappet.
Om du har uppehållstillstånd och hemkommun i Finland har du rätt att använda de tjänster som kommunen tillhandahåller.
Du får mer information om rätten till hemkommun på InfoFinlands sida Hemkommun i Finland.
linkkiStödcentralen Hilma för handikappade invandrare:
Serviceguide för handikappade invandrare(pdf, 797,26)finska _ svenska _ engelska _ ryska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ thai _ burmesiska
linkkiInstitutet för hälsa och välfärd:
Handbok för handikappservicefinska _ svenska
linkkiSocial- och hälsovårdsministeriet:
Handikappservice och stödåtgärderfinska _ svenska _ engelska
Söka tjänster
Tjänsterna för handikappade fås oftast endast med ett läkarintyg (lääkärintodistus).
Besök till exempel din egen hälsostation för en hälsoundersökning.
När du har ett läkarintyg ska du kontakta socialbyrån i din hemkommun.
I kommunen finns en socialarbetare som ansvarar för tjänsterna för handikappade.
Han eller hon ger dig råd och hjälp när du ansöker om tjänster.
Syftet med serviceplanen är att reda ut vilken handikappservice du behöver.
Därefter tas beslut om tjänsterna, och du kan överklaga beslutet om du inte är nöjd med de tjänster som du har beviljats.
Boende
Kommunerna ordnar stödboende och serviceboende för handikappade personer som behöver stöd och hjälp i sitt boende.
Läs mer på InfoFinlands sida Stöd- och serviceboende.
Hjälpmedel
Hälsostationen och centralsjukhuset bekostar de hjälpmedel som ges som medicinsk rehabilitering (lääkinnällinen kuntoutus).
Det innebär att du inte behöver betala för de hjälpmedel som du behöver för att klara dig i vardagen.
Sådana kostnadsfria hjälpmedel är till exempel rullstolar, hörselskadades hörselapparater samt synskadades vita käppar och ledahundar.
Om du måste låta utföra ändringsarbeten i din bostad eller montera fasta hjälpmedel i bostaden kan du få ersättning för dessa av kommunen.
Ändringsarbetena kan vara till exempel ombyggnad av bostaden så att den blir tillgänglig för rullstol.
Fasta hjälpmedel kan till exempel vara olika typer av lyftanordningar samt brandvarnare och dörrklocka för hörselskadade, där ljudet har ersatts med lampor.
Socialarbetaren som ansvarar för handikapptjänster i din hemkommun bedömer tillsammans med dig om du behöver göra ändringsarbeten i din bostad.
FPA kan betala sådana hjälpmedel som du behöver för arbete eller studier.
Hjälpmedel ges till personer som inte klarar av arbete eller studier utan dem eller om det är mycket svårt att studera utan hjälpmedel.
Du kan fråga vid närmaste FPA-byrå hur du kan få hjälpmedel.
linkkiInstitutet för hälsa och välfärd:
Hjälpmedel för att röra sigfinska _ svenska
Hjälpmedel för arbete och studierfinska _ svenska _ engelska
Att röra sig
Om du på grund av ditt handikapp inte kan använda kollektivtrafiken kan du ha rätt till färdtjänst (kuljetuspalvelu).
Vid behov kan du även få en följeslagare (saattaja), d.v.s. en person som assisterar dig på resor.
Du kan få färdtjänst och följeslagare på resor som anknyter till arbete, studier eller fritid.
Du kan söka färdtjänst hos en socialarbetare inom handikappservicen i din hemkommun.
Du betalar för färdtjänsten enligt kollektivtrafikens taxa.
På grund av ditt handikapp kan du även få rabatt på kollektivtrafikens biljettpriser.
Du kan fråga om detta på socialbyrån i din hemkommun.
Färdtjänst och följeslagartjänstfinska _ svenska
Assistentservice
Om du på grund av ditt handikapp behöver mycket hjälp med det vanliga livet kan du få en personlig assistent (henkilökohtainen avustaja).
Assistenten kan hjälpa dig till exempel med att laga mat, handla, på din arbetsplats, i dina studier eller dina hobbyer.
Din hemkommun betalar assistentens lön.
Du kan ansöka om en assistent vid socialbyrån i din hemkommun.
linkkiInstitutet för hälsa och välfärd:
Personlig assistansfinska _ svenska
Tolktjänster
Tolkning för en handikappad är inte det samma som språktolkning.
Du har rätt att använda tolktjänst (tulkkauspalvelu) för handikappade om du har
en hörselskada eller
en syn- och hörselskada eller
en talskada
och om du på grund av din skada behöver hjälp av en tolk
för att arbeta,
studera efter grundläggande studier,
uträtta ärenden,
vid social delaktighet,
Du kan ansöka om tolktjänst vid FPA.
Om du inte förstår finska eller det finska teckenspråket kan du också behöva en annan tolk.
Finländska handikapptolkar kan inte nödvändigtvis de teckenspråk som används i andra länder.
FPA ordnar inte en annan tolk.
När du sköter ärenden med myndigheter, kom alltid ihåg att bekräfta tolksbehovet.
Det åligger myndigheten med vilken du sköter ärenden att ordna tolktjänsten.
Om du blir kallad till hälsovården, kom ihåg att på förhand ange att du behöver en tolk.
Om du söker dig till jourmottagnignen eller läkaren, kan du beställa en tolk vid FPA.
Tolktjänster för handikappadefinska _ svenska
Rehabilitering
Om du har ett gravt handikapp och är under 65 år kan FPA ordna krävande medicinsk rehabilitering (vaativa lääkinnällinen kuntoutus) och ersätta en del av kostnaderna för rehabiliteringen.
Du kan få rehabilitering om ditt handikapp orsakar stora svårigheter att klara av vardagen i hemmet, skolan eller arbetet.
Medicinsk rehabilitering kan ordnas i ett rehabiliteringscenter eller som öppen terapi. Under den öppna terapin kan du bo hemma.
Målet med rehabiliteringen är att hjälpa dig att klara dig bättre i vardagen.
Om du inte kan få krävande medicinsk rehabilitering via FPA ska din hemkommun ordna rehabilitering för dig.
Läs mer på InfoFinlands sida Rehabilitering.
Krävande medicinsk rehabiliteringfinska _ svenska _ engelska
Att ansöka om medicinsk rehabiliteringfinska _ svenska _ engelska
Särskilda tjänster för utvecklingsstörda
Särskilda tjänster för utvecklingsstörda är bland annat
boendetjänster
familjevård
anstaltsvård
arbetsverksamhet och dagverksamhet.
Boendetjänster (asumispalvelu) innebär att en utvecklingsstörd person kan bo i sin egen bostad och där få olika typer av hjälp och stöd.
Läs mer på InfoFinlands sida Stöd- och serviceboende.
Familjevård (perhehoito) innebär att en person vårdas, fostras eller omhändertas i ett privat hem utanför det egna hemmet.
En utvecklingsstörd person som behöver vård kan bo i ett familjehem.
Man kan också bo tillfälligt i ett familjehem.
Familjevård kan även ordnas i den vårdbehövandes eget hem.
Om en utvecklingsstörd person behöver kontinuerlig vård och inte kan få det hemma eller i en servicebostad kan han eller hon även bo på en anstalt (laitos).
Man kan också bo korta tider i en anstalt.
Kommunerna ordnar arbetsverksamhet och dagverksamhet för handikappade personer.
I arbetsverksamheten (työtoiminta) ingår lätt arbete.
Dagverksamheten (päivätoiminta) är avsedd för svårt handikappade personer som inte kan delta i arbetsverksamheten.
Dagverksamheten kan omfatta till exempel matlagning, motion, samtal och friluftsliv.
På internet finns en databank för utvecklingsstörda (Kehitysvammahuollon tietopankki) med mycket nyttig information om utvecklingsstörningar och tjänster för handikappade.
Tjänsten är finskspråkig.
Boendeservice för utvecklingsstördafinska
Utvecklingsstörda och arbetefinska
Dagverksamhetfinska
Kommunerna måste ordna de särskilda tjänster som handikappade behöver.
Dessa särskilda tjänster är till exempel färdtjänst, hjälpmedel eller en personlig assistent.
Syftet med tjänsterna är att hjälpa den handikappade att vara delaktig i samhället och underlätta livet med handikappet.
Om du har uppehållstillstånd och hemkommun i Finland har du rätt att använda de tjänster som kommunen tillhandahåller.
Du får mer information om rätten till hemkommun på InfoFinlands sida Hemkommun i Finland.
linkkiStödcentralen Hilma för handikappade invandrare:
Serviceguide för handikappade invandrare(pdf, 797,26)finska _ svenska _ engelska _ ryska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ thai _ burmesiska
linkkiInstitutet för hälsa och välfärd:
Handbok för handikappservicefinska _ svenska
linkkiSocial- och hälsovårdsministeriet:
Handikappservice och stödåtgärderfinska _ svenska _ engelska
Söka tjänster
Tjänsterna för handikappade fås oftast endast med ett läkarintyg (lääkärintodistus).
Besök till exempel din egen hälsostation för en hälsoundersökning.
När du har ett läkarintyg ska du kontakta socialbyrån i din hemkommun.
I kommunen finns en socialarbetare som ansvarar för tjänsterna för handikappade.
Han eller hon ger dig råd och hjälp när du ansöker om tjänster.
Syftet med serviceplanen är att reda ut vilken handikappservice du behöver.
Därefter tas beslut om tjänsterna, och du kan överklaga beslutet om du inte är nöjd med de tjänster som du har beviljats.
Boende
Kommunerna ordnar stödboende och serviceboende för handikappade personer som behöver stöd och hjälp i sitt boende.
Läs mer på InfoFinlands sida Stöd- och serviceboende.
Hjälpmedel
Hälsostationen och centralsjukhuset bekostar de hjälpmedel som ges som medicinsk rehabilitering (lääkinnällinen kuntoutus).
Det innebär att du inte behöver betala för de hjälpmedel som du behöver för att klara dig i vardagen.
Sådana kostnadsfria hjälpmedel är till exempel rullstolar, hörselskadades hörselapparater samt synskadades vita käppar och ledahundar.
Om du måste låta utföra ändringsarbeten i din bostad eller montera fasta hjälpmedel i bostaden kan du få ersättning för dessa av kommunen.
Ändringsarbetena kan vara till exempel ombyggnad av bostaden så att den blir tillgänglig för rullstol.
Fasta hjälpmedel kan till exempel vara olika typer av lyftanordningar samt brandvarnare och dörrklocka för hörselskadade, där ljudet har ersatts med lampor.
Socialarbetaren som ansvarar för handikapptjänster i din hemkommun bedömer tillsammans med dig om du behöver göra ändringsarbeten i din bostad.
FPA kan betala sådana hjälpmedel som du behöver för arbete eller studier.
Hjälpmedel ges till personer som inte klarar av arbete eller studier utan dem eller om det är mycket svårt att studera utan hjälpmedel.
Du kan fråga vid närmaste FPA-byrå hur du kan få hjälpmedel.
linkkiInstitutet för hälsa och välfärd:
Hjälpmedel för att röra sigfinska _ svenska
Hjälpmedel för arbete och studierfinska _ svenska _ engelska
Att röra sig
Om du på grund av ditt handikapp inte kan använda kollektivtrafiken kan du ha rätt till färdtjänst (kuljetuspalvelu).
Vid behov kan du även få en följeslagare (saattaja), d.v.s. en person som assisterar dig på resor.
Du kan få färdtjänst och följeslagare på resor som anknyter till arbete, studier eller fritid.
Du kan söka färdtjänst hos en socialarbetare inom handikappservicen i din hemkommun.
Du betalar för färdtjänsten enligt kollektivtrafikens taxa.
På grund av ditt handikapp kan du även få rabatt på kollektivtrafikens biljettpriser.
Du kan fråga om detta på socialbyrån i din hemkommun.
Färdtjänst och följeslagartjänstfinska _ svenska
Assistentservice
Om du på grund av ditt handikapp behöver mycket hjälp med det vanliga livet kan du få en personlig assistent (henkilökohtainen avustaja).
Assistenten kan hjälpa dig till exempel med att laga mat, handla, på din arbetsplats, i dina studier eller dina hobbyer.
Din hemkommun betalar assistentens lön.
Du kan ansöka om en assistent vid socialbyrån i din hemkommun.
linkkiInstitutet för hälsa och välfärd:
Personlig assistansfinska _ svenska
Tolktjänster
Tolkning för en handikappad är inte det samma som språktolkning.
Du har rätt att använda tolktjänst (tulkkauspalvelu) för handikappade om du har
en hörselskada eller
en syn- och hörselskada eller
en talskada
och om du på grund av din skada behöver hjälp av en tolk
för att arbeta,
studera efter grundläggande studier,
uträtta ärenden,
vid social delaktighet,
Du kan ansöka om tolktjänst vid FPA.
Om du inte förstår finska eller det finska teckenspråket kan du också behöva en annan tolk.
Finländska handikapptolkar kan inte nödvändigtvis de teckenspråk som används i andra länder.
FPA ordnar inte en annan tolk.
När du sköter ärenden med myndigheter, kom alltid ihåg att bekräfta tolksbehovet.
Det åligger myndigheten med vilken du sköter ärenden att ordna tolktjänsten.
Om du blir kallad till hälsovården, kom ihåg att på förhand ange att du behöver en tolk.
Om du söker dig till jourmottagnignen eller läkaren, kan du beställa en tolk vid FPA.
Tolktjänster för handikappadefinska _ svenska
Rehabilitering
Om du har ett gravt handikapp och är under 65 år kan FPA ordna krävande medicinsk rehabilitering (vaativa lääkinnällinen kuntoutus) och ersätta en del av kostnaderna för rehabiliteringen.
Du kan få rehabilitering om ditt handikapp orsakar stora svårigheter att klara av vardagen i hemmet, skolan eller arbetet.
Medicinsk rehabilitering kan ordnas i ett rehabiliteringscenter eller som öppen terapi. Under den öppna terapin kan du bo hemma.
Målet med rehabiliteringen är att hjälpa dig att klara dig bättre i vardagen.
Om du inte kan få krävande medicinsk rehabilitering via FPA ska din hemkommun ordna rehabilitering för dig.
Läs mer på InfoFinlands sida Rehabilitering.
Krävande medicinsk rehabiliteringfinska _ svenska _ engelska
Att ansöka om medicinsk rehabiliteringfinska _ svenska _ engelska
Särskilda tjänster för utvecklingsstörda
Särskilda tjänster för utvecklingsstörda är bland annat
boendetjänster
familjevård
anstaltsvård
arbetsverksamhet och dagverksamhet.
Boendetjänster (asumispalvelu) innebär att en utvecklingsstörd person kan bo i sin egen bostad och där få olika typer av hjälp och stöd.
Läs mer på InfoFinlands sida Stöd- och serviceboende.
Familjevård (perhehoito) innebär att en person vårdas, fostras eller omhändertas i ett privat hem utanför det egna hemmet.
En utvecklingsstörd person som behöver vård kan bo i ett familjehem.
Man kan också bo tillfälligt i ett familjehem.
Familjevård kan även ordnas i den vårdbehövandes eget hem.
Om en utvecklingsstörd person behöver kontinuerlig vård och inte kan få det hemma eller i en servicebostad kan han eller hon även bo på en anstalt (laitos).
Man kan också bo korta tider i en anstalt.
Kommunerna ordnar arbetsverksamhet och dagverksamhet för handikappade personer.
I arbetsverksamheten (työtoiminta) ingår lätt arbete.
Dagverksamheten (päivätoiminta) är avsedd för svårt handikappade personer som inte kan delta i arbetsverksamheten.
Dagverksamheten kan omfatta till exempel matlagning, motion, samtal och friluftsliv.
På internet finns en databank för utvecklingsstörda (Kehitysvammahuollon tietopankki) med mycket nyttig information om utvecklingsstörningar och tjänster för handikappade.
Tjänsten är finskspråkig.
Boendeservice för utvecklingsstördafinska
Utvecklingsstörda och arbetefinska
Dagverksamhetfinska
Egenvårdsläkemedel (itsehoitolääke) kan köpas utan läkarrecept.
Exempel på egenvårdsläkemedel är de flesta värkmediciner.
För många läkemedel behöver du dock ett recept, d.v.s. en läkemedelsförskrivning (lääkemääräys) för att köpa dem.
Receptet skrivs ut av en läkare.
Också många sjukskötare har rätt att skriva ut vissa läkemedel.
Till exempel antibiotika är receptbelagda läkemedel.
Om du har en långvarig sjukdom ska du ta med dina gamla recept till läkarmottagningen så kan läkaren beakta dessa när han eller hon skriver ut ett recept.
Om läkaren har skrivit ut ett elektroniskt recept (sähköinen resepti), kan du ta ut medicinerna på apoteket utan pappersrecept.
Receptet är giltigt två år från den dag det skrivits ut.
Ett recept som du skaffat utomlands är inte giltigt i Finland.
Undantag är recept som är utskrivna i de övriga nordiska länderna och europeiska recept. De är giltiga i Finland.
Du måste begära ett europeiskt recept särskilt av din läkare.
Europeiska recept kan skrivas ut av yrkesutbildade personer inom hälso- och sjukvården som arbetar i ett EU- eller EES-land eller Schweiz och har förskrivningsrätt.
På läkemedelsförpackningen står det sista användningsdatumet.
Om läkemedlet har föråldrats kan det inte längre användas.
Släng inte föråldrade läkemedel utan lämna dem alltid till apoteket (apteekki), eftersom de är problemavfall.
Information om läkemedelspreparatfinska
linkkiKanta:
Elektroniskt receptfinska _ svenska _ engelska
Var får jag läkemedel?
Du kan köpa läkemedel på apoteket.
Till apotekets tjänster hör också sidoapotek och apotekens tjänsteställen samt apotekets egen webbtjänst.
I Finland får läkemedel inte säljas annanstans.
Vitaminer och naturprodukter säljs också i vanliga butiker.
Apoteken har vanligen öppet från morgon till kväll.
I större städer kan det finnas apotek som har öppet till sent på kvällen.
På Apotekareförbundets (Apteekkariliitto) webbplats kan du söka information om apoteken på din hemort och deras öppettider.
På apoteket kan du byta ut det läkemedel som föreskrivs på receptet mot ett annat, förmånligare läkemedel om det verksamma ämnet är detsamma i båda preparaten.
Den anställda på apoteket berättar för kunden om det finns ett billigare alternativ.
linkkiSocial- och hälsovårdsministeriet:
Apotekfinska _ svenska _ engelska _ ryska
linkkiApotekareförbundet:
Apotekens kontaktuppgifterfinska
FPA-ersättning för läkemedel
Om du omfattas av den finländska sjukförsäkringen (sairausvakuutus) ersätter FPA (Kela) en del av kostnaderna för många läkemedel.
Du får ingen ersättning för läkemedel som du köper utan recept.
Man kan få ersättning först efter att den initiala självrisken (alkuomavastuu) har överskridits, det vill säga efter att du har köpt ersättningsgilla mediciner för över 50 euro under ett år.
Den initiala självrisken gäller inte mediciner för personer under 18 år.
Du kan få ersättningen redan på apoteket.
Ersättningen dras av läkemedlets pris i kassan.
Du kan också söka ersättning i efterhand med en blankett.
Bifoga apotekets utredning över de köpta läkemedlen och kassakvittot.
Mer information om vem som omfattas den finländska sjukförsäkringen får du på InfoFinlands sida Den sociala tryggheten i Finland.
Läkemedelsersättningarfinska _ svenska _ engelska
Hälsa och rehabiliteringfinska _ svenska _ ryska _ estniska
Läkemedel från utlandet
Vissa läkemedel kan du ta med dig från utlandet till Finland för eget bruk.
Importen är dock begränsad.
Begränsningarna beror på vilken sorts läkemedel det är fråga om och från vilket land du tar med dig läkemedlet till Finland.
Du måste också till exempel med ett recept eller ett läkarintyg kunna bevisa att läkemedlet är avsett för eget bruk.
Ta reda på begränsningarna innan du för in läkemedel i Finland.
Ta reda på begränsningarna också om du vill beställa läkemedel till Finland per post.
Från EES-länderna får du ta med dig den mängd läkemedel för eget bruk som motsvarar ett års förbrukning.
Per post får du från EES-länderna beställa den mängd läkemedel som motsvarar högst tre månaders förbrukning.
Från länder utanför EES-området får du ta med dig till Finland den mängd läkemedel för eget bruk som motsvarar högst tre månaders förbrukning.
Enligt lag får man inte beställa läkemedel per post från länder utanför EES-området.
Om läkemedlet har klassificerats som narkotika är begränsningarna strängare.
Om du är osäker på om ett visst läkemedel får föras in i Finland ska du fråga råd vid Tullen (Tulli).
Om du beställer läkemedel från utlandet får du ingen ersättning från FPA (Kela) för dem.
I EU-länderna finns några webbapotek där man kan lagligt köpa egenvårdsläkemedel.
Största delen av läkemedelsbutikerna på internet är dock illegala.
Det kan också vara en hälsorisk att köpa läkemedel i en olaglig webbutik.
linkkiTullen:
Personliga läkemedelfinska _ svenska _ engelska
linkkiFimea:
Införsel av läkemedel till Finlandfinska _ svenska _ engelska
linkkiFimea:
Läkemedelshandel på internetfinska _ svenska _ engelska
Enligt finsk lag får ingen diskrimineras på grund av ett handikapp.
Handikappade personer har rätt att leva ett normalt liv, till exempel studera, arbeta och bilda familj.
Finland har ratificerat FN:s konvention om rättigheter för personer med funktionshinder.
Handikappade personer kan ha svårt att klara av det dagliga livet på grund av sitt handikapp eller sin sjukdom.
Kommunerna måste tillhandahålla handikappade de tjänster som de behöver.
Sådana tjänster är till exempel färd- och assistenttjänsterna.
Om du har uppehållstillstånd och hemkommun i Finland, har du rätt till kommunens tjänster för handikappade.
Läs mer om tjänsterna för handikappade och om att ansöka dem på InfoFinlands sida Tjänster för handikappade.
Handikapporganisationer
I Finland finns flera organisationer som arbetar för att förbättra handikappade personers ställning i samhället.
Hos dessa organisationer kan du få råd och hjälp till exempel vid ansökan om tjänster.
Många organisationer erbjuder fritidsverksamhet och kamratstöd till personer i alla åldrar.
Du hittar kontaktuppgifterna till organisationerna på Handikappforums webbplats.
I Finland finns även stödcentret
Hilma för handikappade invandrare som erbjuder servicevägledning och rådgivning för handikappade invandrare och långtidssjuka.
linkkiStödcentralen Hilma för handikappade invandrare:
Stöd och hjälp för handikappade invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ persiska _ arabiska _ kurdiska
Handikapporganisationer i Finlandfinska _ svenska
Synskadade
Om du är blind eller har nedsatt syn kan du få tjänster för synskadade.
Om du behöver hjälpmedel ska du först besöka din egen hälsostation för en läkarundersökning.
Läkaren bedömer din synskada och därefter kan du få hjälpmedel i form av medicinsk rehabilitering.
Läs mer på InfoFinlands sida Tjänster för handikappade.
Om du på grund av ditt handikapp behöver till exempel en speciell dator eller särskilda hushållsapparater kan du få understöd för detta vid socialbyrån i din hemkommun.
Detta är dock prövningsbaserat, med andra ord är det inte säkert att du får stödet.
På biblioteket för synskadade Celia kan du låna ljudböcker, punktskriftsböcker, e-böcker och reliefbilder.
Biblioteket producerar även läroböcker för synskadade skolelevers och studerandes behov.
Synskadades förbund är en organisation som arbetar för att förbättra synskadades ställning i samhället.
Förbundet erbjuder även mycket nyttig information och tjänster till synskadade.
De vanligaste hjälpmedlen för synskadadefinska
linkkiCelia:
De synskadades bibliotekfinska _ svenska _ engelska
Hörselskadade
Personer med en hörselskada är döva eller har nedsatt hörsel.
Många kommunicerar med teckenspråk.
I Finland används det finska och det finlandssvenska teckenspråket.
Personer med en hörselskada använder ofta även hörapparater.
Om du behöver hjälpmedel ska du först besöka din egen hälsostation för en läkarundersökning.
Läkaren bedömer din hörselskada och därefter kan du få hjälpmedel i form av medicinsk rehabilitering.
Du kan till exempel få ett brandlarm avsett för hörselskadade och en texttelefon för att kunna bo tryggt i ditt hem.
Ansök om dessa hjälpmedel vid socialbyrån i din hemkommun.
Om du behöver det på grund av din hörselskada kan du få tolktjänster till exempel i arbetet, studierna eller när du ska sköta ärenden.
Tolkning kan ges på teckenspråk eller vara skrivtolkning.
Ansök om rätten att använda tolktjänster hos FPA.
Läs mer om hjälpmedel och tolktjänster på InfoFinlands sida Tjänster för handikappade.
På internet finns ordboken för det finska teckenspråket, Suvi.
Hörselförbundet och Finlands Dövas Förbund är organisationer som arbetar för att förbättra hörselskadade personers ställning i samhället.
De erbjuder även mycket nyttig information och tjänster till hörselskadade.
linkkiFinska Hörselförbundet rf:
Hjälpmedel för hörselnfinska
linkkiFinska Hörselförbundet rf:
Hörselapparatfinska
Tolktjänster för handikappadefinska _ svenska
Ordbok i det finska teckenspråketfinska
linkkiFinska Hörselförbundet rf:
Information om Hörselförbundetfinska
linkkiFinlands Dövas Förbund rf:
Information om Finlands Dövas Förbundfinska _ svenska _ engelska
linkkiDövas folkhögskola:
Utbildning för döva invandrarefinska _ svenska _ engelska
Rörelsehandikappade
En rörelsehandikappad person kan inte röra sig självständigt eller utan hjälpmedel.
En rörelsenedsättning kan bero på en sjukdom, ett olycksfall eller genetiska orsaker.
Om du behöver hjälpmedel ska du först besöka din egen hälsostation för en läkarundersökning.
Läkaren bedömer din rörelsenedsättning och därefter kan du få hjälpmedel i form av medicinsk rehabilitering.
Om det måste göras förändringsarbeten eller installeras fasta hjälpmedel i din bostad kan du få ersättning för detta av din hemkommun.
Bostaden kan till exempel byggas om så att du kan röra dig med en rullstol i den.
Fasta hjälpmedel är till exempel stödhandtag, ramper och elektriska dörrar.
Läs mer om hjälpmedel och förändringsarbeten på InfoFinlands sida Tjänster för handikappade.
linkkiInvalidförbundet:
Stöd och verksamhet för rörelsehindradefinska
Utvecklingsstörda
En utvecklingsstörning gör det svårare att lära sig och förstå nya saker.
För en utvecklingsstörd person är det svårare att lära sig och minnas saker än för andra.
Utvecklingsstörningen upptäcks ofta i barndomen eller ungdomen.
För en utvecklingsstörd person finns olika slags specialtjänster.
Sådana är till exempel boendetjänster, arbetsverksamhet och dagverksamhet.
Läs mer om tjänsterna för utvecklingsstörda på InfoFinlands sida Tjänster för handikappade.
Det finns även många organisationer där du kan få information och stöd.
Du hittar mer information till exempel på Kehitysvammaliittos och Kehitysvammaisten Tukiliittos webbplatser.
Information för utvecklingsstörda och anhörigafinska
linkkiFörbundet Utvecklingsstörning:
Utvecklingsstördas intressebevakningsorganisationfinska _ engelska
linkkiUtvecklingsstördas intressebevakningsorganisation:
Utvecklingsstördas intressebevakningsorganisationfinska _ svenska _ engelska
Enligt finsk lag får ingen diskrimineras på grund av ett handikapp.
Handikappade personer har rätt att leva ett normalt liv, till exempel studera, arbeta och bilda familj.
Finland har ratificerat FN:s konvention om rättigheter för personer med funktionshinder.
Handikappade personer kan ha svårt att klara av det dagliga livet på grund av sitt handikapp eller sin sjukdom.
Kommunerna måste tillhandahålla handikappade de tjänster som de behöver.
Sådana tjänster är till exempel färd- och assistenttjänsterna.
Om du har uppehållstillstånd och hemkommun i Finland, har du rätt till kommunens tjänster för handikappade.
Läs mer om tjänsterna för handikappade och om att ansöka dem på InfoFinlands sida Tjänster för handikappade.
Handikapporganisationer
I Finland finns flera organisationer som arbetar för att förbättra handikappade personers ställning i samhället.
Hos dessa organisationer kan du få råd och hjälp till exempel vid ansökan om tjänster.
Många organisationer erbjuder fritidsverksamhet och kamratstöd till personer i alla åldrar.
Du hittar kontaktuppgifterna till organisationerna på Handikappforums webbplats.
I Finland finns även stödcentret
Hilma för handikappade invandrare som erbjuder servicevägledning och rådgivning för handikappade invandrare och långtidssjuka.
linkkiStödcentralen Hilma för handikappade invandrare:
Stöd och hjälp för handikappade invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ persiska _ arabiska _ kurdiska
Handikapporganisationer i Finlandfinska _ svenska
Synskadade
Om du är blind eller har nedsatt syn kan du få tjänster för synskadade.
Om du behöver hjälpmedel ska du först besöka din egen hälsostation för en läkarundersökning.
Läkaren bedömer din synskada och därefter kan du få hjälpmedel i form av medicinsk rehabilitering.
Läs mer på InfoFinlands sida Tjänster för handikappade.
Om du på grund av ditt handikapp behöver till exempel en speciell dator eller särskilda hushållsapparater kan du få understöd för detta vid socialbyrån i din hemkommun.
Detta är dock prövningsbaserat, med andra ord är det inte säkert att du får stödet.
På biblioteket för synskadade Celia kan du låna ljudböcker, punktskriftsböcker, e-böcker och reliefbilder.
Biblioteket producerar även läroböcker för synskadade skolelevers och studerandes behov.
Synskadades förbund är en organisation som arbetar för att förbättra synskadades ställning i samhället.
Förbundet erbjuder även mycket nyttig information och tjänster till synskadade.
De vanligaste hjälpmedlen för synskadadefinska
linkkiCelia:
De synskadades bibliotekfinska _ svenska _ engelska
Hörselskadade
Personer med en hörselskada är döva eller har nedsatt hörsel.
Många kommunicerar med teckenspråk.
I Finland används det finska och det finlandssvenska teckenspråket.
Personer med en hörselskada använder ofta även hörapparater.
Om du behöver hjälpmedel ska du först besöka din egen hälsostation för en läkarundersökning.
Läkaren bedömer din hörselskada och därefter kan du få hjälpmedel i form av medicinsk rehabilitering.
Du kan till exempel få ett brandlarm avsett för hörselskadade och en texttelefon för att kunna bo tryggt i ditt hem.
Ansök om dessa hjälpmedel vid socialbyrån i din hemkommun.
Om du behöver det på grund av din hörselskada kan du få tolktjänster till exempel i arbetet, studierna eller när du ska sköta ärenden.
Tolkning kan ges på teckenspråk eller vara skrivtolkning.
Ansök om rätten att använda tolktjänster hos FPA.
Läs mer om hjälpmedel och tolktjänster på InfoFinlands sida Tjänster för handikappade.
På internet finns ordboken för det finska teckenspråket, Suvi.
Hörselförbundet och Finlands Dövas Förbund är organisationer som arbetar för att förbättra hörselskadade personers ställning i samhället.
De erbjuder även mycket nyttig information och tjänster till hörselskadade.
linkkiFinska Hörselförbundet rf:
Hjälpmedel för hörselnfinska
linkkiFinska Hörselförbundet rf:
Hörselapparatfinska
Tolktjänster för handikappadefinska _ svenska
Ordbok i det finska teckenspråketfinska
linkkiFinska Hörselförbundet rf:
Information om Hörselförbundetfinska
linkkiFinlands Dövas Förbund rf:
Information om Finlands Dövas Förbundfinska _ svenska _ engelska
linkkiDövas folkhögskola:
Utbildning för döva invandrarefinska _ svenska _ engelska
Rörelsehandikappade
En rörelsehandikappad person kan inte röra sig självständigt eller utan hjälpmedel.
En rörelsenedsättning kan bero på en sjukdom, ett olycksfall eller genetiska orsaker.
Om du behöver hjälpmedel ska du först besöka din egen hälsostation för en läkarundersökning.
Läkaren bedömer din rörelsenedsättning och därefter kan du få hjälpmedel i form av medicinsk rehabilitering.
Om det måste göras förändringsarbeten eller installeras fasta hjälpmedel i din bostad kan du få ersättning för detta av din hemkommun.
Bostaden kan till exempel byggas om så att du kan röra dig med en rullstol i den.
Fasta hjälpmedel är till exempel stödhandtag, ramper och elektriska dörrar.
Läs mer om hjälpmedel och förändringsarbeten på InfoFinlands sida Tjänster för handikappade.
linkkiInvalidförbundet:
Stöd och verksamhet för rörelsehindradefinska
Utvecklingsstörda
En utvecklingsstörning gör det svårare att lära sig och förstå nya saker.
För en utvecklingsstörd person är det svårare att lära sig och minnas saker än för andra.
Utvecklingsstörningen upptäcks ofta i barndomen eller ungdomen.
För en utvecklingsstörd person finns olika slags specialtjänster.
Sådana är till exempel boendetjänster, arbetsverksamhet och dagverksamhet.
Läs mer om tjänsterna för utvecklingsstörda på InfoFinlands sida Tjänster för handikappade.
Det finns även många organisationer där du kan få information och stöd.
Du hittar mer information till exempel på Kehitysvammaliittos och Kehitysvammaisten Tukiliittos webbplatser.
Information för utvecklingsstörda och anhörigafinska
linkkiFörbundet Utvecklingsstörning:
Utvecklingsstördas intressebevakningsorganisationfinska _ engelska
linkkiUtvecklingsstördas intressebevakningsorganisation:
Utvecklingsstördas intressebevakningsorganisationfinska _ svenska _ engelska
Du kan köpa ett graviditetstest på apoteket.
Även stora mataffärer säljer graviditetstest.
När du är gravid:
Boka en tid på mödrarådgivningen.
Besök läkaren före slutet av den fjärde graviditetsmånaden.
Om du arbetar, meddela arbetsgivaren skriftligt senast två månader innan du går på moderskapsledighet.
Boka en tid på mödrarådgivningen
När du upptäcker att du är gravid, kontakta mödrarådgivningen eller familjecentret i din hemkommun.
Du kan använda tjänsterna vid rådgivningsbyrån eller familjecentret om du har en hemkommun i Finland.
Läs mer på InfoFinlands sida Hemkommun i Finland.
Också asylsökande kan använda tjänsterna vid mödrarådgivningen.
I vissa städer får du använda tjänsterna vid mödrarådgivningen även om du vistas i Finland utan uppehållstillstånd.
På rådgivningsbyrån följer en hälsovårdare ditt hälsotillstånd och babyns hälsa.
På rådgivningsbyrån får du anvisningar för en trygg graviditet och förlossning.
Du får även viktig information om tjänsterna för barnfamiljer i Finland.
Du behöver inte betala för tjänsterna vid rådgivningsbyrån.
Barnets båda föräldrar är välkomna till rådgivningsbyrån.
Om du vill kan du även be en stödperson att följa med.
Om du behöver tolk kan sköterskan på rådgivningsbyrån be en tolk att närvara vid besöken.
Tolken ska vara vuxen.
linkkiInstitutet för hälsa och välfärd:
Broschyren Vi väntar barn(pdf, 1,46 Mt)finska _ svenska _ engelska _ ryska _ somaliska
linkkiSocial- och hälsovårdsministeriet:
Information om rådgivningsbyråernas tjänsterfinska _ svenska _ engelska _ ryska
Besök läkaren
Besök läkaren vid rådgivningsbyrån före slutet av den fjärde graviditetsmånaden.
Du kan ofta boka läkartiden via mödrarådgivningen.
När du har gjort en läkarkontroll får du ett graviditetsintyg.
Du behöver intyget om du ansöker om moderskapsledighet av din arbetsgivare.
Du behöver intyget även om du ansöker om moderskapsunderstödet och moderskapspenning hos FPA.
Läs mer om dessa förmåner på InfoFinlands sida Stöd till gravida.
På sidan Den sociala tryggheten i Finland finns information om vem som har rätt till FPA:s förmåner.
Privata mödrarådgivningar
I Finland finns även privata mödrarådgivningar.
Tänk på att privata hälso- och sjukvårdstjänster är avgiftsbelagda.
Läs mer på sidan Hälsovårdstjänster Finland.
Könsstympning och graviditet
Om du har blivit utsatt för könsstympning kan du få en öppningsoperation.
Den underlättar undersökningarna under graviditeten.
Också förlossningen blir lättare.
Öppningsoperationen kan göras före graviditeten, när graviditeten är halvvägs eller i samband med förlossningen.
Hälsovårdaren på rådgivningsbyrån frågar om du har blivit utsatt för könsstympning.
Det är viktigt att du berättar detta så att hälsovårdaren kan hänvisa dig till öppningsoperation.
Förlossningen
I Finland föder kvinnorna oftast på sjukhus.
Fråga på mödrarådgivningen på vilket sjukhus du ska föda.
Om du har en hemkommun i Finland kostar förlossningen inte särskilt mycket.
Barnets andra förälder kan vara med på förlossningen.
Om du vill kan du även be någon annan släkting eller en vän att följa med.
I Finland föder de flesta kvinnorna vaginalt.
Det är vanligtvis det tryggaste sättet.
Om det inte är möjligt fattar läkaren beslut om kejsarsnitt.
Om du är rädd inför förlossningen, prata om det på rådgivningsbyrån.
Du kan få hjälp med rädslan till exempel på polikliniken för förlossningsrädsla.
Efter förlossningen stannar du oftast några dagar på sjukhuset med barnet.
Den andra föräldern eller din stödperson kan vara på sjukhuset hela dagen för att hjälpa dig.
Om du har fått ditt första barn kan stödpersonen ofta även tillbringa nätterna på sjukhuset.
När du åker till sjukhuset ska du ta med dig tillräckligt varma kläder för barnet för hemresan.
Om du åker hem med barnet i bil, behöver du ett babyskydd i bilen.
Tolkning vid förlossningen
Man vet inte i förväg när förlossningen börjar.
Därför kan det vara svårt att få en tolk till förlossningen.
En del tolkcentraler har jour på veckoslut samt kvällar och nätter.
Du får mer information om tolktjänsterna i din kommun på rådgivningsbyrån.
Läs mer om tolktjänsterna på InfoFinlands sida Behöver du en tolk?
När barnet har fötts
På sidan När ett barn föds i Finland finns viktig information om de praktiska ärenden som du måste ta hand om när barnet har fötts.
På sidan finns till exempel information om registrering av barnet i befolkningsdatasystemet, om namnlagen i Finland och om barnets sociala trygghet.
Hjälp med babyn
Om du känner att du inte klarar dig med babyn utan hjälp kan du bo på ett mödrahem och lära dig hur du tar hand om barnet där.
Fråga om verksamheten vid din mödrarådgivning.
För mödrahemmet behöver du en remiss som utfärdas av kommunen.
Rehabilitering som ordnas av kommunerna
Kommunerna ordnar medicinsk rehabilitering till exempel vid hälsovårdscentraler och i sjukhus.
Du kan få kommunal rehabilitering om du har hemkommun i Finland.
Kommunernas rehabilitering omfattar:
rådgivning om rehabilitering
undersökningar för att fastställa rehabiliteringsbehovet
vård för att förbättra arbets- och funktionsförmågan
rehabiliteringsperioder
hjälpmedelstjänster
anpassningsträning
rehabiliteringshandledning
Mer information om kommunens rehabiliteringstjänster får du vid din egen hälsostation.
Rehabilitering som ordnas av FPA
FPA:s rehabilitering kan vara:
rehabilitering för gravt handikappade
behovsprövad rehabilitering
rehabiliteringspsykoterapi
Yrkesinriktad rehabilitering ordnas av arbetspensionsanstalter (työeläkelaitokset) och FPA (Kela).
Medicinsk rehabilitering ordnas av kommunerna och FPA.
Om du lider av en yrkessjukdom eller har blivit skadad i ett olycksfall, kan du få rehabilitering från försäkringsbolaget (vakuutusyhtiö).
FPA kan betala ut understöd för psykoterapin, men du måste själv hitta en lämplig terapeut.
FPA:s rehabilitering är avsedd för personer som omfattas av den finländska sjukförsäkringen (sairausvakuutus).
Mer information om sjukförsäkringen får du på InfoFinlands sida Den sociala tryggheten i Finland.
Rehabilitering för arbete
Du kan få yrkesinriktad rehabilitering om du har sådana hälsoproblem som hindrar dig från att arbeta.
Du kan också få rehabilitering om du riskerar att tvingas sluta arbeta på grund av dina hälsoproblem.
Du har rätt till rehabilitering efter ett arbetsolycksfall.
Arbetspensionsanstalter ordnar yrkesinriktad rehabilitering för arbetstagare.
Du kan ansöka om rehabilitering vid arbetspensionsanstalten om du har arbetat fem år eller längre.
Fråga mer av de sakkunniga inom rehabiliteringsfrågor vid din arbetspensionsanstalt.
FPA ordnar yrkesinriktad rehabilitering för unga personer och vuxna som inte arbetar.
Yrkesinriktad rehabiliteringfinska _ svenska _ engelska
Att ansöka om yrkesinriktad rehabiliteringfinska _ svenska _ engelska
Rehabilitering för gravt handikappade
Om du är under 65 år och har på grund av sjukdom eller funktionsnedsättning stora svårigheter att klara av vardagen, till exempel om du har svårt att röra dig eller ta hand om dig själv, kan FPA ordna krävande medicinsk rehabilitering (vaativa lääkinnällinen kuntoutus) för dig.
Rehabiliteringen genomförs på ett sätt som passar just dig.
Du kan få rehabilitering till exempel vid en rehabiliteringsinrättning (kuntoutuslaitos).
Du kan också bo hemma och gå på rehabilitering därifrån.
Målet med rehabiliteringen är att stöda dig och dina närstående så att du kan föra ett aktivt liv.
Mer information om krävande medicinsk rehabilitering fås av FPA.
Krävande medicinsk rehabiliteringfinska _ svenska _ engelska
Att ansöka om medicinsk rehabiliteringfinska _ svenska _ engelska
Behovsprövad rehabilitering
Du kan få behovsprövad rehabilitering om ditt mål är att fortsätta arbeta, återgå till arbetet eller börja arbeta.
Du kan få behovsprövad rehabilitering om hälso- och sjukvården konstaterar att du har en skada eller sjukdom som kräver rehabilitering.
Behovsprövad rehabilitering kan till exempel omfatta
rehabiliteringskurser för personer med en viss sjukdom
kurser för anpassningsträning
Läs mer om de olika alternativen för behovsprövad rehabilitering på FPA:s webbplats.
Behovsprövad rehabiliteringfinska _ svenska
Psykoterapi som rehabilitering
Om du behöver psykoterapi som stöd för din arbets- eller studieförmåga, kan du eventuellt ansöka om rehabiliterande psykoterapi (kuntoutuspsykoterapia).
Villkor för att du ska få rehabiliterande psykoterapi är att
du har fått psykiatrisk vård i minst tre månader och
den vårdande psykiatern skriver ett utlåtande med rekommendation om rehabiliterande psykoterapi.
Lär mer om mentala tjänster på InfoFinlands sida Mental hälsa.
För personer i åldern 16–25 år kan den också omfatta musikterapi.
Terapi för unga kan också omfatta besök av föräldrar.
Du kan få understöd för terapin ett år i taget under högst tre år.
FPA ersätter högst 80 terapibesök om året och högst 200 besök under tre år.
För att få FPA:s bidrag för psykoterapi ska terapeuten ha rätt att använda psykoterapeutens yrkesbenämning och vara godkänd av FPA.
Rehabiliterande psykoterapifinska _ svenska _ engelska
linkkiFinlands Psykologiförbund:
Hur söker du dig till rehabilitering
När du behöver rehabilitering behöver du först ett läkarutlåtande.
Ta kontakt med din läkare, företagsläkare eller FPA.
Om du ansöker om krävande medicinsk rehabilitering behöver du dessutom en rehabiliteringsplan (kuntoutussuunnitelma).
När du har fått ett läkarutlåtande eller en rehabiliteringsplan kan du ansöka om rehabilitering vid din arbetspensionsanstalt eller FPA.
Du kan fråga vid kommunens hälsovårdstjänster arbetspensionsanstalten eller FPA om olika rehabiliteringsmöjligheter.
Mer information om FPA:s rehabiliteringar hittar du också på FPA:s webbplats.
Om du söker till rehabilitering som ordnas av FPA ska du lämna in din ansökan om rehabilitering till FPA innan rehabiliteringen börjar.
FPA ger ett skriftligt beslut om rehabilitering.
Sköta ärenden på Internetfinska _ svenska _ engelska
Kontaktuppgifter till FPAfinska _ svenska _ engelska
Elektronisk tidsbeställningfinska _ svenska _ engelska
Under rehabiliteringen kan du få rehabiliteringspenning (kuntoutusraha), om du är 16–67 år och om rehabiliteringen har som syfte att bevara din arbetsförmåga eller göra det möjligt för dig att återvända till arbetslivet eller komma in i arbetslivet.
För att få rehabiliteringspenning måste du också få ett rehabiliteringsbeslut (kuntoutuspäätös) till exempel från FPA eller företagshälsovården.
Du kan få rehabiliteringspenning på samma villkor också när din hemkommun ordnar din rehabilitering.
FPA kan delvis ersätta resorna till rehabiliteringen.
Rehabiliteringspenningfinska _ svenska _ engelska
Rehabilitering som ordnas av kommunerna
Kommunerna ordnar medicinsk rehabilitering till exempel vid hälsovårdscentraler och i sjukhus.
Du kan få kommunal rehabilitering om du har hemkommun i Finland.
Kommunernas rehabilitering omfattar:
rådgivning om rehabilitering
undersökningar för att fastställa rehabiliteringsbehovet
vård för att förbättra arbets- och funktionsförmågan
rehabiliteringsperioder
hjälpmedelstjänster
anpassningsträning
rehabiliteringshandledning
Mer information om kommunens rehabiliteringstjänster får du vid din egen hälsostation.
Rehabilitering som ordnas av FPA
FPA:s rehabilitering kan vara:
rehabilitering för gravt handikappade
behovsprövad rehabilitering
rehabiliteringspsykoterapi
Yrkesinriktad rehabilitering ordnas av arbetspensionsanstalter (työeläkelaitokset) och FPA (Kela).
Medicinsk rehabilitering ordnas av kommunerna och FPA.
Om du lider av en yrkessjukdom eller har blivit skadad i ett olycksfall, kan du få rehabilitering från försäkringsbolaget (vakuutusyhtiö).
FPA kan betala ut understöd för psykoterapin, men du måste själv hitta en lämplig terapeut.
FPA:s rehabilitering är avsedd för personer som omfattas av den finländska sjukförsäkringen (sairausvakuutus).
Mer information om sjukförsäkringen får du på InfoFinlands sida Den sociala tryggheten i Finland.
Rehabilitering för arbete
Du kan få yrkesinriktad rehabilitering om du har sådana hälsoproblem som hindrar dig från att arbeta.
Du kan också få rehabilitering om du riskerar att tvingas sluta arbeta på grund av dina hälsoproblem.
Du har rätt till rehabilitering efter ett arbetsolycksfall.
Arbetspensionsanstalter ordnar yrkesinriktad rehabilitering för arbetstagare.
Du kan ansöka om rehabilitering vid arbetspensionsanstalten om du har arbetat fem år eller längre.
Fråga mer av de sakkunniga inom rehabiliteringsfrågor vid din arbetspensionsanstalt.
FPA ordnar yrkesinriktad rehabilitering för unga personer och vuxna som inte arbetar.
Yrkesinriktad rehabiliteringfinska _ svenska _ engelska
Att ansöka om yrkesinriktad rehabiliteringfinska _ svenska _ engelska
Rehabilitering för gravt handikappade
Om du är under 65 år och har på grund av sjukdom eller funktionsnedsättning stora svårigheter att klara av vardagen, till exempel om du har svårt att röra dig eller ta hand om dig själv, kan FPA ordna krävande medicinsk rehabilitering (vaativa lääkinnällinen kuntoutus) för dig.
Rehabiliteringen genomförs på ett sätt som passar just dig.
Du kan få rehabilitering till exempel vid en rehabiliteringsinrättning (kuntoutuslaitos).
Du kan också bo hemma och gå på rehabilitering därifrån.
Målet med rehabiliteringen är att stöda dig och dina närstående så att du kan föra ett aktivt liv.
Mer information om krävande medicinsk rehabilitering fås av FPA.
Krävande medicinsk rehabiliteringfinska _ svenska _ engelska
Att ansöka om medicinsk rehabiliteringfinska _ svenska _ engelska
Behovsprövad rehabilitering
Du kan få behovsprövad rehabilitering om ditt mål är att fortsätta arbeta, återgå till arbetet eller börja arbeta.
Du kan få behovsprövad rehabilitering om hälso- och sjukvården konstaterar att du har en skada eller sjukdom som kräver rehabilitering.
Behovsprövad rehabilitering kan till exempel omfatta
rehabiliteringskurser för personer med en viss sjukdom
kurser för anpassningsträning
Läs mer om de olika alternativen för behovsprövad rehabilitering på FPA:s webbplats.
Behovsprövad rehabiliteringfinska _ svenska
Psykoterapi som rehabilitering
Om du behöver psykoterapi som stöd för din arbets- eller studieförmåga, kan du eventuellt ansöka om rehabiliterande psykoterapi (kuntoutuspsykoterapia).
Villkor för att du ska få rehabiliterande psykoterapi är att
du har fått psykiatrisk vård i minst tre månader och
den vårdande psykiatern skriver ett utlåtande med rekommendation om rehabiliterande psykoterapi.
Lär mer om mentala tjänster på InfoFinlands sida Mental hälsa.
För personer i åldern 16–25 år kan den också omfatta musikterapi.
Terapi för unga kan också omfatta besök av föräldrar.
Du kan få understöd för terapin ett år i taget under högst tre år.
FPA ersätter högst 80 terapibesök om året och högst 200 besök under tre år.
För att få FPA:s bidrag för psykoterapi ska terapeuten ha rätt att använda psykoterapeutens yrkesbenämning och vara godkänd av FPA.
Rehabiliterande psykoterapifinska _ svenska _ engelska
linkkiFinlands Psykologiförbund:
Hur söker du dig till rehabilitering
När du behöver rehabilitering behöver du först ett läkarutlåtande.
Ta kontakt med din läkare, företagsläkare eller FPA.
Om du ansöker om krävande medicinsk rehabilitering behöver du dessutom en rehabiliteringsplan (kuntoutussuunnitelma).
När du har fått ett läkarutlåtande eller en rehabiliteringsplan kan du ansöka om rehabilitering vid din arbetspensionsanstalt eller FPA.
Du kan fråga vid kommunens hälsovårdstjänster arbetspensionsanstalten eller FPA om olika rehabiliteringsmöjligheter.
Mer information om FPA:s rehabiliteringar hittar du också på FPA:s webbplats.
Om du söker till rehabilitering som ordnas av FPA ska du lämna in din ansökan om rehabilitering till FPA innan rehabiliteringen börjar.
FPA ger ett skriftligt beslut om rehabilitering.
Sköta ärenden på Internetfinska _ svenska _ engelska
Kontaktuppgifter till FPAfinska _ svenska _ engelska
Elektronisk tidsbeställningfinska _ svenska _ engelska
Under rehabiliteringen kan du få rehabiliteringspenning (kuntoutusraha), om du är 16–67 år och om rehabiliteringen har som syfte att bevara din arbetsförmåga eller göra det möjligt för dig att återvända till arbetslivet eller komma in i arbetslivet.
För att få rehabiliteringspenning måste du också få ett rehabiliteringsbeslut (kuntoutuspäätös) till exempel från FPA eller företagshälsovården.
Du kan få rehabiliteringspenning på samma villkor också när din hemkommun ordnar din rehabilitering.
FPA kan delvis ersätta resorna till rehabiliteringen.
Rehabiliteringspenningfinska _ svenska _ engelska
I Finland kan du avbryta en graviditet i tidigt skede i följande fall:
om förlossningen kan utgöra en risk för din hälsa
om du är under 17 eller över 40 år gammal
om du redan har fött fyra barn
om du inte kan ta hand om barnet på grund av en sjukdom.
Som orsak för abort (abortti) räcker även att det med tanke på din livssituation skulle vara en alltför stor belastning att föda barnet eller att ta hand om det.
I praktiken kan orsaken vara någon av följande:
familjeförhållanden
arbetssituation
boende
Kvinnan har rätt att själv besluta om hon vill göra abort.
Partnern kan delta i beslutsfattandet om kvinnan vill ta hänsyn till hans åsikt.
Om du är minderårig och vill göra abort behöver du inte tillstånd av dina föräldrar.
Det är dock ofta bra att diskutera saken med föräldrarna.
Om du ändå inte vill göra det har de yrkesutbildade personerna inom hälsovården tystnadsplikt.
Aborten ska göras före den tolfte graviditetsveckan.
Av speciellt vägande skäl kan abort göras även senare men då behöver du ett specialtillstånd från Valvira (Valvira).
Du behöver tillstånd från Valvira även om aborten görs på grund av att fostret har en svår sjukdom eller ett handikapp.
Fråga mer av läkaren vid din egen hälsostation (terveysasema).
Om du vill avbryta graviditeten ska du kontakta hälsostationen i ditt eget område så fort som möjligt och boka tid hos en läkare.
Du kan också boka tid hos en privatläkare, men kontrollera när du bokar tiden att läkaren har Valviras tillstånd att ge ett utlåtande för abort.
Om du vill kan du ta med dig din partner till läkarmottagningen.
Läkaren skriver en remiss till det sjukhus där aborten görs.
På sjukhuset samtalar en skötare och en läkare med dig.
Ni fattar gemensamt beslutet om på vilket sätt graviditeten avbryts.
På detta inverkar hur långt graviditeten har gått och din egen åsikt.
Graviditeten avbryts med läkemedel eller med skrapning (kaavinta).
Skrapning görs vanligtvis i narkos och därefter ska du stanna några timmar på sjukhuset.
Om aborten görs medicinskt doseras läkemedlet med 1–3 dagars mellanrum via slidan så att livmoderns börjar dras samman och töms.
Var förberedd på att du behöver smärtlindring när livmodern dras samman.
Ibland behövs det skrapning efter medicinsk abort.
2–4 veckor efter aborten görs en efterkontroll på hälsostationen.
När du ska fatta beslut om abort får du stöd till exempel av en hälsovårdare eller en läkare vid hälsostationen.
Mer information om olika ställen där du får hjälp i en krävande livssituation finns på InfoFinlands sida Mental hälsa.
Abortfinska
Tillstånd till att avbryta graviditetenfinska _ svenska
På den här sidan finns information om tjänsterna i Rovaniemi.
Allmän information om studier i finska och svenska i Finland hittar du på InfoFinlands sida Finska och svenska språket.
Kurser i finska språket
Kurser i finska språket vid öppna universitetet
Moninets webbplats
Kurser i finska språket
Medborgarinstitutet i Rovaniemi erbjuder kurser i finska språket.
Du hittar en lista över kurserna i finska på medborgarinstitutets webbplats.
Studier i finska språket på Internetfinska _ engelska
Du ska anmäla dig till kursen i förväg: fyll i anmälningsblanketten, lämna den till Rovalas kontor och betala kursavgiften.
Du kan också betala kursavgiften på Internet om du har webbankkoder till Handelsbanken, Sparbanken Optia, Nordea, Andelsbanken eller Danske Bank.
Du kan inte anmäla dig per telefon.M
kursanmälanfinska
Kontaktuppgifter:
Rovala 5
tfn 040 4873 010
Kontorets öppettider
linkkiRovala:
Medborgarinstitutetfinska
Kurser i finska språket vid öppna universitetet
Språkcentret vid Lapplands universitet ordnar kurser i finska språket på engelska.
Du kan söka till Finnish for Foreigners-kurserna via öppna universitetet.
Kurserna är avgiftsbelagda.
Information om nya kurser och ansökan till kurserna finns på öppna universitetets webbplats.
Öppna universitetet
Moninets webbplats
På MoniNets webbplats finns en studiemiljö för finska språket där du kan studera finska på egen hand.
I studiemiljön finns sju avsnitt som handlar om invandrarens liv i Finland.
Varje avsnitt innehåller vokabulär- och grammatikövningar.
Settlementföreningen Rovalan Setlementti ry/MoniNet
Studier i finska språket på Internetfinska _ engelska
På MoniNets webbplats finns länkar till olika webbsidor där du kan studera finska på egen hand.
Settlementföreningen Rovalan Setlementti ry/MoniNet
Studier i finska språket på Internetfinska _ engelska
På den här sidan finns information om tjänsterna i Rovaniemi.
Allmän information om studier i finska och svenska i Finland hittar du på InfoFinlands sida Finska och svenska språket.
Kurser i finska språket
Kurser i finska språket vid öppna universitetet
Moninets webbplats
Kurser i finska språket
Medborgarinstitutet i Rovaniemi erbjuder kurser i finska språket.
Du hittar en lista över kurserna i finska på medborgarinstitutets webbplats.
Studier i finska språket på Internetfinska _ engelska
Du ska anmäla dig till kursen i förväg: fyll i anmälningsblanketten, lämna den till Rovalas kontor och betala kursavgiften.
Du kan också betala kursavgiften på Internet om du har webbankkoder till Handelsbanken, Sparbanken Optia, Nordea, Andelsbanken eller Danske Bank.
Du kan inte anmäla dig per telefon.M
kursanmälanfinska
Kontaktuppgifter:
Rovala 5
tfn 040 4873 010
Kontorets öppettider
linkkiRovala:
Medborgarinstitutetfinska
Kurser i finska språket vid öppna universitetet
Språkcentret vid Lapplands universitet ordnar kurser i finska språket på engelska.
Du kan söka till Finnish for Foreigners-kurserna via öppna universitetet.
Kurserna är avgiftsbelagda.
Information om nya kurser och ansökan till kurserna finns på öppna universitetets webbplats.
Öppna universitetet
Moninets webbplats
På MoniNets webbplats finns en studiemiljö för finska språket där du kan studera finska på egen hand.
I studiemiljön finns sju avsnitt som handlar om invandrarens liv i Finland.
Varje avsnitt innehåller vokabulär- och grammatikövningar.
Settlementföreningen Rovalan Setlementti ry/MoniNet
Studier i finska språket på Internetfinska _ engelska
På MoniNets webbplats finns länkar till olika webbsidor där du kan studera finska på egen hand.
På den här sidan finns information om tjänsterna i Rovaniemi.
Allmän information om studier i finska och svenska i Finland hittar du på InfoFinlands sida Finska och svenska språket.
Kurser i finska språket
Kurser i finska språket vid öppna universitetet
Medborgarinstitutet i Rovaniemi erbjuder kurser i finska språket.
Du hittar en lista över kurserna i finska på medborgarinstitutets webbplats.
Studier i finska språket på Internetfinska _ engelska
Du kan också betala kursavgiften på Internet om du har webbankkoder till Handelsbanken, Sparbanken Optia, Nordea, Andelsbanken eller Danske Bank.
kursanmälanfinska
Kontaktuppgifter:
Kurser i finska språket vid öppna universitetet
Språkcentret vid Lapplands universitet ordnar kurser i finska språket på engelska.
Du kan söka till Finnish for Foreigners-kurserna via öppna universitetet.
Kurserna är avgiftsbelagda.
Information om nya kurser och ansökan till kurserna finns på öppna universitetets webbplats.
Moninets webbplats
På MoniNets webbplats finns en studiemiljö för finska språket där du kan studera finska på egen hand.
I studiemiljön finns sju avsnitt som handlar om invandrarens liv i Finland.
Varje avsnitt innehåller vokabulär- och grammatikövningar.
Settlementföreningen Rovalan Setlementti ry/MoniNet
Studier i finska språket på Internetfinska _ engelska
På MoniNets webbplats finns länkar till olika webbsidor där du kan studera finska på egen hand.
Settlementföreningen Rovalan Setlementti ry/MoniNet
Studier i finska språket på Internetfinska _ engelska
Rättigheterna för klienter inom hälsovården tryggas i lag.
Patienternas rättigheter gäller offentliga och privata hälsovårdstjänster samt hälsovårdstjänster till exempel för åldringar och handikappade.
Om du har hemkommun (kotikunta) i Finland har du rätt att utnyttja de offentliga hälsovårdstjänsterna.
Mer information finns på InfoFinlands sida Hemkommun i Finland.
Vårdgaranti (hoitotakuu)
Om du behöver brådskande vård, till exempel om du råkar ut för en olycka, har du rätt att genast få vård på jourmottagningen vid den närmaste hälsovårdscentralen eller det närmaste sjukhuset.
Om du inte har hemkommun i Finland och inte heller någon annan grund ger dig rätt att utnyttja de offentliga hälsovårdstjänsterna i Finland måste du betala ett pris som motsvarar de faktiska kostnaderna för dessa hälsovårdstjänster.
Om du har hemkommun i Finland kan du utnyttja de offentliga hälsovårdstjänsterna i din kommun.
Hälsovårdscentralen måste besvara patienternas samtal eller ha öppet så att patienterna kan besöka hälsovårdscentralen alla vardagar under tjänstetid.
Om situationen kräver det har du rätt att besöka hälsostationen inom tre vardagar efter att du kontaktade hälsostationen.
Hälsostationen måste inleda även icke-brådskande vård senast inom tre månader.
Du kan bli intagen på sjukhus med en läkarremiss.
Sjukhuset måste bedöma vårdbehovet inom tre veckor efter att läkarremissen har kommit till sjukhuset.
Om det konstateras att en patient behöver vård på sjukhus måste vården inledas senast inom sex månader efter att vårdbehovet har bedömts.
Om den egna hälsostationen eller det egna sjukhuset inte kan ge patienten vård inom utsatt tid måste de ordna möjlighet för patienten att få vård på ett annat ställe.
Detta får inte orsaka extra kostnader för patienten.
linkkiSocial- och hälsovårdsministeriet:
Vårdgarantifinska _ svenska
Övriga rättigheter
Patienten har rätt:
till vård av hög kvalitet
till ett gott bemötande: patientens människovärde, övertygelse och integritet ska respekteras
till att patientens modersmål och kultur beaktas i den mån det är möjligt
att alltid när det är möjligt bli tillfrågad om sitt medgivande innan behandlingen påbörjas
att få upplysningar om sitt hälsotillstånd, vårdens omfattning, riskfaktorer och alternativa behandlingsmetoder
att kontrollera sina egna uppgifter i patientjournalen och rätta till dem
att få veta tidpunkten för intagning för vård om patienten måsta köa till vården
att vägra vård
att göra en anmärkning till den vårdande enheten om patienten är missnöjd
att vid behov få hjälp av patientombudsmannen (potilasasiamies).
En minderårig patients åsikt beaktas när barnet är tillräckligt utvecklat för att uttrycka sin åsikt.
En läkare eller någon annan yrkesutbildad person avgör detta.
Barnets föräldrar eller vårdnadshavare kan inte vägra vård om barnet behöver den.
Jämlikhet inom hälsovården
Enligt Finlands grundlag är alla människor lika inför lagen.
Ingen får utan godtagbar orsak behandlas olika på grund av kön, ålder, ursprung, språk, religion, övertygelse, åsikt, hälsotillstånd, funktionshinder, sexuell läggning eller annat som rör ens person.
I Finland gäller även en lag om likabehandling.
Denna lag tillämpas bland annat på diskriminering på grund av etniskt ursprung inom offentliga och privata social- och hälsovårdstjänster.
Diskrimineringsombudsmannen och diskriminerings- och jämställdhetsnämnden övervakar att människor inte diskrimineras på grund av sitt etniska ursprung.
Alla klienter inom hälsovården har rätt till likabehandling utan diskriminering.
Om du inte har rätt att använda de offentliga hälsovårdstjänsterna, har du rätt att behandlas jämlikt inom den privata hälsovården.
Diskriminering och dåligt bemötande inom hälsovården
Om du upplever att du blivit fel bemött inom hälsovården kan du ta kontakt med patientombudsmannen (potilasasiamies).
Patientombudsmannens tjänster är tillgängliga på alla ställen där hälsovårdstjänster tillhandahålls, till exempel på hälsostationer, sjukhus, privata läkarstationer, åldringshem och vårdanstalter för handikappade.
Patientombudsmannens tjänster är kostnadsfria.
Be om kontaktuppgifterna till patientombudsmannen vid den vårdenhet där du har varit klient.
Patientombudsmannen bistår i att reda ut missförstånd samt ger råd och hjälper dig om du vill göra en anmärkning eller söka patientskadeersättning.
Patientombudsmannen ger också information om patientens rättigheter och främjar förverkligandet av dessa.
linkkiSocial- och hälsovårdsministeriet:
Patientombudsmannenfinska _ svenska _ engelska _ ryska
Hjälp till diskrimineringsofferfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ thai _ vietnamesiska _ portugisiska _ tagalog _ polska
Tolktjänster
Inom hälsovården har du rätt att bli betjänad på finska och svenska.
Om inte talar dessa språk kan du i Finland få tolktjänster på många olika språk.
I en del situationer kan myndigheten beställa en tolk och betala för tolkningen. Detta är inte alltid möjligt.
Fråga myndigheten på förhand.
Tolkningen kan också ordnas per telefon.
Tolken ska vara myndig, så egna minderåriga barn kan inte användas som tolk.
Du får mer information på InfoFinlands sida Behöver du en tolk?.
Patientföreningar
I Finland finns många patientföreningar som tillhandahåller information och rådgivning för människor med en viss sjukdom.
Via en patientförening kan man också hitta kamratstöd.
Kontaktuppgifter till patientorganisationerfinska
Om du blir sjuk eller råkar ut för en olycka har du rätt att stanna hemma från arbetet.
Om du omfattas av den finländska sjukförsäkringen (sairausvakuutus) har du efter en självrisktid (omavastuuaika) rätt att söka sjukdagpenning (sairauspäiväraha) hos FPA (Kela).
Självrisktiden är vanligen den dag då du insjuknade och därpå följande nio vardagar.
Om din anställning har varat över en månad före insjuknandet betalar din arbetsgivare full lön för självrisktiden.
Sjukdagpenning betalas för högst 300 vardagar.
Den ska sökas inom två månader efter insjuknandet.
Du kan söka sjukdagpenning om du:
omfattas av den finländska sjukförsäkringen (sairausvakuutus): läs mer på InfoFinlands sida Den sociala tryggheten i Finland
är 16–67 år
är arbetsoförmögen på grund av din sjukdom
har arbetat tre månader som anställd, företagare eller yrkesutövare tre månader innan du insjuknade eller har tre månader innan du insjuknade varit heltidsstuderande, arbetslös arbetssökande, d.v.s. kund vid arbets- och näringsbyrån (työ- ja elinkeinotoimisto), sabbatsledig (sapattivapaa) eller alterneringsledig (vuorotteluvapaa).
Om du får lön under sjukledigheten, ansöker din arbetsgivare om sjukdagpenningen och då betalas sjukdagpenningen till din arbetsgivare.
Om du är sjuk en lång tid och din arbetsgivare inte längre betalar dig lön under sjukledigheten kan du söka FPA:s sjukdagpenning när lönen inte längre utbetalas.
Sjukdagpenningens belopp beror på inkomsterna.
Den beräknas oftast på basis av de arbetsinkomster som bekräftats i beskattningen.
Till exempel beaktas inte royaltyn och anställningsoptioner vid beräkning av dagpenningens belopp.
Om din inkomst har ökat kan du söka sjukdagpenning på basis av arbetsinkomsten under de senaste sex månaderna.
Du ska då bifoga till ansökan ett löneintyg för löner som du har fått.
Be om intyget av din arbetsgivare.
När du söker sjukdagpenning ska du bifoga till ansökan:
ett läkarintyg om arbetsoförmögenhet
ett löneintyg för de senaste sex månaderna om dina inkomster har ökat.
Mer information om sjukdagpenningen får du på FPA:s webbplats.
Om du är sjuk en lång tid ska du ta reda på om rehabilitering kan vara till nytta för dig.
Sjukdagpenningfinska _ svenska _ engelska
Att ansöka om sjukdagpenningfinska _ svenska _ engelska
Hälsa och rehabiliteringfinska _ svenska _ ryska _ estniska
Partiell sjukdagpenning
Den partiella sjukdagpenningen (osasairauspäiväraha) är avsedd för 16–67-åriga heltidsarbetande anställda eller företagare som omfattas av den sociala tryggheten i Finland.
Syftet med den partiella sjukdagpenningen är att du kan fortsätta att arbeta eller att återgå till arbetet trots att du har blivit sjuk.
Diskutera först med din läkare inom företagshälsovården och din arbetsgivare om möjligheten att söka partiell sjukdagpenning.
Företagshälsovårdsläkaren avgör om du kan deltidsarbeta medan du är sjuk.
När du söker partiell sjukdagpenning ska du bifoga till ansökan:
ett läkarintyg om arbetsoförmögenhet
ansökan om sjukdagpenning
en kopia av överenskommelsen mellan dig och din arbetsgivare om att du under en viss tid ska arbeta på deltid.
Arbetstidsarrangemanget och lönen ska framgå ur avtalet.
ett löneintyg för de senaste sex månaderna före insjuknandet om dina inkomster har ökat.
Partiell sjukdagpenning ska sökas inom två månader efter att du börjar arbeta på deltid.
Mer information om den partiella sjukdagpenningen får du på FPA:s webbplats.
Partiell sjukdagpenningfinska _ svenska _ engelska
Att ansöka om partiell sjukdagpenningfinska _ svenska _ engelska
I Finland tillhandahåller både den offentliga och den privata hälso- och sjukvården tjänster inom graviditetsprevention, gynekologi, tidig upptäckt av cancer, sexuell hälsa hos män, barnlöshet och könssjukdomar.
Har du rätt till de offentliga hälsovårdstjänsterna?
Läs mer på sidan Hälsovårdstjänster Finland.
Ungas sexualitetfinska _ engelska
Vuxnas sexualitetfinska _ svenska _ engelska
Du kan köpa kondomer i affärer, på bensinstationer, kiosker och apotek.
Du behöver inget recept.
För hormonella preventivmedel behöver du ett recept av en läkare.
Sådana preventivmedel är till exempel p-piller och minipiller.
De säljs på apoteket.
Du kan boka en tid på hälsostationen eller vid en privat läkarstation.
Även minderåriga barn kan boka tid hos läkaren och få ett recept för preventivmedel.
Du behöver inte tillstånd av dina föräldrar för receptet.
Vissa kommuner erbjuder unga kostnadsfria preventivmedel.
Du kan fråga om detta på hälsostationen eller av skolhälsovårdaren.
Om preventionen misslyckades eller om du glömde att använda preventivmedel kan du köpa ett akut p-piller på apoteket utan recept.
Du ska ta pillret så snart som möjligt efter samlaget, i regel senast inom 72 timmar.
Vissa preparat kan tas inom 120 timmar efter samlaget.
linkkiSHVS:
Graviditetspreventionfinska _ svenska _ engelska
Sexuell hälsa hos kvinnor
Alla läkare på hälsostationen gör gynekologiska undersökningar.
Fråga mer på din hälsostation.
Om du vill träffa en kvinnlig läkare, ange detta när du bokar tiden.
Läkaren kan vid behov skriva remiss till en specialist på gynekologiska polikliniken.
Du kan även boka tid hos en privat gynekolog.
Då kan du välja läkaren själv.
Tjänsterna hos privatläkare är mycket dyrare för klienten.
I Finland ordnas regelbundna screeningundersökningar för kvinnor i vissa åldrar.
På så sätt försöker man i ett tidigt skede hitta bröstcancer och livmoderhalscancer.
Undersökning av bröstcancer görs på kvinnor i åldern 50–69 år ungefär vartannat år.
Undersökning av livmoderhalscancer görs på kvinnor i åldern 30–60 år vart femte år.
linkkiSocial- och hälsovårdsministeriet:
Screeningsundersökningarfinska _ svenska _ engelska _ ryska
linkkiInstitutet för hälsa och välfärd:
Information om bröstcancerscreeningfinska _ svenska
Anvisning för identifiering av bröstcancer(pdf, 440kt)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ kinesiska _ thai _ rumänska _ samiska
Information om cancerscreeningfinska _ svenska _ engelska
Sexuell hälsa hos män
Du kan boka en läkartid på din egen hälsostation.
Om du vill kan du be om att få träffa en manlig läkare.
Läkaren kan vid behov skriva remiss till en specialist på urologiska polikliniken.
Du kan även boka tid på en privat läkarstation.
Tjänsterna hos privatläkare är mycket dyrare för klienten.
Barnlöshet
Barnlöshet kan oftast behandlas.
Orsaken till barnlöshet kan finnas hos kvinnan eller hos mannen.
Ibland hittar man ingen medicinsk orsak till den.
Om du har slutat använda preventivmedel, men en graviditet inte har börjat inom ett år, boka tid på hälsostationen eller hos en privat gynekolog.
Det är bra om paret besöker mottagningen tillsammans.
Läkaren skriver en remiss till undersökningar på barnlöshetspolikliniken.
Med undersökningarna utreds varför en graviditet inte har börjat.
Fertilitetsbehandlingar tillhandahålls av både offentliga och privata kliniker. till exempel kvinnans ålder påverkar rätten till fertilitetsbehandling inom de offentliga hälsovårdstjänsterna.
Könssjukdomar
Om du misstänker att du har en könssjukdom kan du boka en läkartid på hälsostationen eller en privat läkarstation.
I vissa städer finns en poliklinik för könssjukdomar där könssjukdomar behandlas.
Fråga mer på din hälsostation.
Du kan skydda dig mot de flesta könssjukdomarna med kondom eller slicklapp.
Också papperslösa och asylsökande har rätt att få behandling för könssjukdomar.
Om du vistas i Finland utan uppehållstillstånd kan du emellertid bli tvungen att betala för vården.
linkkiHivpoint:
Broschyren Information om sexuellt överförda sjukdomar(pdf, 1500kt)finska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
linkkiHivpoint:
Info om HIVfinska _ engelska _ ryska
linkkiHivpoint:
Broschyren Ett gott liv med HIVfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ thai
linkkiHivpoint:
Broschyren HIV i familjen(pdf, 881 kb)finska _ engelska _ ryska
Manlig omskärelse
Fundera noga på om omskärelse behövs.
Om pojken är gammal nog för att säga sin åsikt ska han tillfrågas om han samtycker till operationen.
Operationen får inte göras om pojken motsätter sig.
Om pojken har två vårdnadshavare måste båda ge sitt skriftliga samtycke till operationen.
Om det inte finns några medicinska skäl till omskärelsen kan den inte utföras inom den offentliga hälsovården.
Då måste du betala för operationen själv.
Endast en läkare får utföra operationen.
Den ska göras i steril miljö.
Läkaren ska se till att patienten får smärtlindring.
Fråga mer om omskärelse på rådgivningsbyrån, en hälsostationsläkare, skolhälsovårdaren eller skolläkaren.
Kvinnlig könsstympning
Könsstympning av flickor är ett brott i Finland.
Man kan få ett flerårigt fängelsestraff för det.
Det är likaså brottsligt att ta flickan utomlands för könsstympning.
Om du har blivit utsatt för detta kan du få en öppningsoperation.
Även en korrigerande operation är möjlig.
Fråga mer på din hälsostation.
Omskärelse av kvinnor och flickorfinska _ engelska _ somaliska _ arabiska
Om du blir sjuk eller råkar ut för en olycka har du rätt att stanna hemma från arbetet.
Om du omfattas av den finländska sjukförsäkringen (sairausvakuutus) har du efter en självrisktid (omavastuuaika) rätt att söka sjukdagpenning (sairauspäiväraha) hos FPA (Kela).
Självrisktiden är vanligen den dag då du insjuknade och därpå följande nio vardagar.
Om din anställning har varat över en månad före insjuknandet betalar din arbetsgivare full lön för självrisktiden.
Sjukdagpenning betalas för högst 300 vardagar.
Den ska sökas inom två månader efter insjuknandet.
Du kan söka sjukdagpenning om du:
omfattas av den finländska sjukförsäkringen (sairausvakuutus): läs mer på InfoFinlands sida Den sociala tryggheten i Finland
är 16–67 år
är arbetsoförmögen på grund av din sjukdom
har arbetat tre månader som anställd, företagare eller yrkesutövare tre månader innan du insjuknade eller har tre månader innan du insjuknade varit heltidsstuderande, arbetslös arbetssökande, d.v.s. kund vid arbets- och näringsbyrån (työ- ja elinkeinotoimisto), sabbatsledig (sapattivapaa) eller alterneringsledig (vuorotteluvapaa).
Om du får lön under sjukledigheten, ansöker din arbetsgivare om sjukdagpenningen och då betalas sjukdagpenningen till din arbetsgivare.
Om du är sjuk en lång tid och din arbetsgivare inte längre betalar dig lön under sjukledigheten kan du söka FPA:s sjukdagpenning när lönen inte längre utbetalas.
Sjukdagpenningens belopp beror på inkomsterna.
Den beräknas oftast på basis av de arbetsinkomster som bekräftats i beskattningen.
Till exempel beaktas inte royaltyn och anställningsoptioner vid beräkning av dagpenningens belopp.
Om din inkomst har ökat kan du söka sjukdagpenning på basis av arbetsinkomsten under de senaste sex månaderna.
Du ska då bifoga till ansökan ett löneintyg för löner som du har fått.
Be om intyget av din arbetsgivare.
När du söker sjukdagpenning ska du bifoga till ansökan:
ett läkarintyg om arbetsoförmögenhet
ett löneintyg för de senaste sex månaderna om dina inkomster har ökat.
Mer information om sjukdagpenningen får du på FPA:s webbplats.
Om du är sjuk en lång tid ska du ta reda på om rehabilitering kan vara till nytta för dig.
Sjukdagpenningfinska _ svenska _ engelska
Att ansöka om sjukdagpenningfinska _ svenska _ engelska
Hälsa och rehabiliteringfinska _ svenska _ ryska _ estniska
Partiell sjukdagpenning
Den partiella sjukdagpenningen (osasairauspäiväraha) är avsedd för 16–67-åriga heltidsarbetande anställda eller företagare som omfattas av den sociala tryggheten i Finland.
Syftet med den partiella sjukdagpenningen är att du kan fortsätta att arbeta eller att återgå till arbetet trots att du har blivit sjuk.
Diskutera först med din läkare inom företagshälsovården och din arbetsgivare om möjligheten att söka partiell sjukdagpenning.
Företagshälsovårdsläkaren avgör om du kan deltidsarbeta medan du är sjuk.
När du söker partiell sjukdagpenning ska du bifoga till ansökan:
ett läkarintyg om arbetsoförmögenhet
ansökan om sjukdagpenning
en kopia av överenskommelsen mellan dig och din arbetsgivare om att du under en viss tid ska arbeta på deltid.
Arbetstidsarrangemanget och lönen ska framgå ur avtalet.
ett löneintyg för de senaste sex månaderna före insjuknandet om dina inkomster har ökat.
Partiell sjukdagpenning ska sökas inom två månader efter att du börjar arbeta på deltid.
Mer information om den partiella sjukdagpenningen får du på FPA:s webbplats.
Partiell sjukdagpenningfinska _ svenska _ engelska
Att ansöka om partiell sjukdagpenningfinska _ svenska _ engelska
Egenvårdsläkemedel (itsehoitolääke) kan köpas utan läkarrecept.
Exempel på egenvårdsläkemedel är de flesta värkmediciner.
För många läkemedel behöver du dock ett recept, d.v.s. en läkemedelsförskrivning (lääkemääräys) för att köpa dem.
Receptet skrivs ut av en läkare.
Också många sjukskötare har rätt att skriva ut vissa läkemedel.
Till exempel antibiotika är receptbelagda läkemedel.
Om du har en långvarig sjukdom ska du ta med dina gamla recept till läkarmottagningen så kan läkaren beakta dessa när han eller hon skriver ut ett recept.
Om läkaren har skrivit ut ett elektroniskt recept (sähköinen resepti), kan du ta ut medicinerna på apoteket utan pappersrecept.
Receptet är giltigt två år från den dag det skrivits ut.
Ett recept som du skaffat utomlands är inte giltigt i Finland.
Undantag är recept som är utskrivna i de övriga nordiska länderna och europeiska recept. De är giltiga i Finland.
Du måste begära ett europeiskt recept särskilt av din läkare.
Europeiska recept kan skrivas ut av yrkesutbildade personer inom hälso- och sjukvården som arbetar i ett EU- eller EES-land eller Schweiz och har förskrivningsrätt.
På läkemedelsförpackningen står det sista användningsdatumet.
Om läkemedlet har föråldrats kan det inte längre användas.
Släng inte föråldrade läkemedel utan lämna dem alltid till apoteket (apteekki), eftersom de är problemavfall.
Information om läkemedelspreparatfinska
linkkiKanta:
Elektroniskt receptfinska _ svenska _ engelska
Var får jag läkemedel?
Du kan köpa läkemedel på apoteket.
Till apotekets tjänster hör också sidoapotek och apotekens tjänsteställen samt apotekets egen webbtjänst.
I Finland får läkemedel inte säljas annanstans.
Vitaminer och naturprodukter säljs också i vanliga butiker.
Apoteken har vanligen öppet från morgon till kväll.
I större städer kan det finnas apotek som har öppet till sent på kvällen.
På Apotekareförbundets (Apteekkariliitto) webbplats kan du söka information om apoteken på din hemort och deras öppettider.
På apoteket kan du byta ut det läkemedel som föreskrivs på receptet mot ett annat, förmånligare läkemedel om det verksamma ämnet är detsamma i båda preparaten.
Den anställda på apoteket berättar för kunden om det finns ett billigare alternativ.
linkkiSocial- och hälsovårdsministeriet:
Apotekfinska _ svenska _ engelska _ ryska
linkkiApotekareförbundet:
Apotekens kontaktuppgifterfinska
FPA-ersättning för läkemedel
Om du omfattas av den finländska sjukförsäkringen (sairausvakuutus) ersätter FPA (Kela) en del av kostnaderna för många läkemedel.
Du får ingen ersättning för läkemedel som du köper utan recept.
Man kan få ersättning först efter att den initiala självrisken (alkuomavastuu) har överskridits, det vill säga efter att du har köpt ersättningsgilla mediciner för över 50 euro under ett år.
Den initiala självrisken gäller inte mediciner för personer under 18 år.
Du kan få ersättningen redan på apoteket.
Ersättningen dras av läkemedlets pris i kassan.
Du kan också söka ersättning i efterhand med en blankett.
Bifoga apotekets utredning över de köpta läkemedlen och kassakvittot.
Mer information om vem som omfattas den finländska sjukförsäkringen får du på InfoFinlands sida Den sociala tryggheten i Finland.
Läkemedelsersättningarfinska _ svenska _ engelska
Hälsa och rehabiliteringfinska _ svenska _ ryska _ estniska
Läkemedel från utlandet
Vissa läkemedel kan du ta med dig från utlandet till Finland för eget bruk.
Importen är dock begränsad.
Begränsningarna beror på vilken sorts läkemedel det är fråga om och från vilket land du tar med dig läkemedlet till Finland.
Du måste också till exempel med ett recept eller ett läkarintyg kunna bevisa att läkemedlet är avsett för eget bruk.
Ta reda på begränsningarna innan du för in läkemedel i Finland.
Ta reda på begränsningarna också om du vill beställa läkemedel till Finland per post.
Från EES-länderna får du ta med dig den mängd läkemedel för eget bruk som motsvarar ett års förbrukning.
Per post får du från EES-länderna beställa den mängd läkemedel som motsvarar högst tre månaders förbrukning.
Från länder utanför EES-området får du ta med dig till Finland den mängd läkemedel för eget bruk som motsvarar högst tre månaders förbrukning.
Enligt lag får man inte beställa läkemedel per post från länder utanför EES-området.
Om läkemedlet har klassificerats som narkotika är begränsningarna strängare.
Om du är osäker på om ett visst läkemedel får föras in i Finland ska du fråga råd vid Tullen (Tulli).
Om du beställer läkemedel från utlandet får du ingen ersättning från FPA (Kela) för dem.
I EU-länderna finns några webbapotek där man kan lagligt köpa egenvårdsläkemedel.
Största delen av läkemedelsbutikerna på internet är dock illegala.
Det kan också vara en hälsorisk att köpa läkemedel i en olaglig webbutik.
linkkiTullen:
Personliga läkemedelfinska _ svenska _ engelska
linkkiFimea:
Införsel av läkemedel till Finlandfinska _ svenska _ engelska
linkkiFimea:
Läkemedelshandel på internetfinska _ svenska _ engelska
När ska jag söka hjälp?
Vem som helst kan behöva hjälp om livssituationen är påfrestande.
Livet kan vara svårt till exempel när man flyttar från ett land till ett annat, har problem på arbetsplatsen, förlorar sin arbetsplats, har problem i familjen, går igenom skilsmässa, förlorar en anhörig, blir sjuk eller när livet förändras på andra sätt.
Också positiva saker, t.ex. att man får barn, kan ändra livet så mycket att man behöver stöd i den nya situationen.
Ibland kan man må dåligt först i efterhand när man redan har lagt den svåra erfarenheten bakom sig och situationen har lugnat ner sig.
Det lönar sig att söka hjälp, om du har något av följande symptom:
sömnlöshet
ingen aptit
vardagen känns tung
du orkar inte arbeta eller träffa människor
fysiska symptom, utan att medicinska orsaker hittas för dessa
ökad alkohol- eller droganvändning
Det är inte ovanligt att söka hjälp för att få stöd med den mentala hälsan.
I Finland lider 20 % av befolkningen av depression i något skede av livet.
Depression(pdf, 110,37 kt)finska _ engelska _ ryska _ franska _ somaliska _ turkiska _ persiska _ arabiska _ kurdiska _ albanska _ vietnamesiska _ burmesiska _ bosniska _ serbiska _ swahili
Var får jag hjälp?
Ofta hjälper det redan att tala om dessa saker med familjen eller vänner. Ibland behövs det även annan hjälp.
Det kan hjälpa att tala med en hälsovårdare (terveydenhoitaja), läkare (lääkäri) eller en psykoterapeut (psykoterapeutti).
Tillsammans kan ni fundera på vilken sorts stöd som skulle passa just dig.
Ofta hjälper terapi, medicinering eller en kombination av båda.
Ibland behövs sjukhusvård.
Sjukhusvården räcker vanligen några veckor.
Målsättningen är att patienten kan återvända hem så fort som möjligt.
Därefter fortsätter vården som öppenvård.r.
Om du har hemkommun i Finland ska du först kontakta din egen hälsostation (terveysasema).
Hälsostationerna har vanligen öppet från måndag till fredag, ungefär kl. 8–16.
Ring hälsostationen genast på morgonen för att boka tid.
Om du behöver hjälp genast ska du tala om det när du ringer.
Läkaren skriver vid behov en remiss till psykiatriska polikliniken (psykiatrian poliklinikka) eller en annan vårdenhet för psykisk hälsa.
Du kan inte gå till polikliniken utan en läkarremiss.
Med läkaren eller psykologen kan du samtala konfidentiellt. De har tystnadsplikt.
De berättar inte om dina saker för andra myndigheter.
Om någon annan hälsovårdsenhet behöver dina uppgifter, ombeds du ge ditt medgivande för överlåtelse av dessa.
På din egen hälsostation får du mer information om hur mentalvårdstjänsterna är ordnade i din hemkommun.
Om du är orolig för en närstående person och tror att han eller hon kan vara i behov av hjälp, kan du rådfråga till exempel hälsovårdaren eller läkaren vid hälsocentralen.
linkkiSocial- och hälsovårdsministeriet:
Mentalvårdstjänsterfinska _ svenska _ engelska _ ryska
Privata mentalvårdstjänster
Du kan också boka tid hos en psykiater eller en psykolog vid en privat läkarstation.
Där får man ibland fortare en tid, men besöket kostar avsevärt mer för kunden.
FPA (Kela) ersätter en del av kostnaderna för besök hos privatläkare om du omfattas av den finländska sjukförsäkringen.
Fråga mer hos FPA.
FPA:s ersättning kan ibland dras av direkt på det belopp som du betalar vid kassan.
Ta med ett intyg över att du omfattas av den finländska sjukförsäkringen.
Du kan också söka ersättning från FPA även i efterhand.
Läs mer om vem som omfattas av den finländska sjukförsäkringen på InfoFinlands sida Den sociala tryggheten i Finland.
Sjukvårdsersättningarfinska _ svenska _ engelska
Privat psykoterapitjänst på Internetfinska _ svenska _ engelska _ ryska _ franska _ spanska _ turkiska _ kinesiska _ tyska _ portugisiska _ norska
_ holländska _ japanska _ italienska
_ danska
Privat läkarstationfinska _ svenska _ engelska
Privat läkarstationfinska _ svenska _ engelska
När hjälpbehovet är brådskande
Om du känner att du behöver hjälp omedelbart kan du kontakta den närmaste jourhavande hälsovårdscentralen eller sjukhusjouren.
Brådskande psykiatrisk sjukvård ges på jourenheter vid psykiatriska sjukhus.
Om din närstående utgör en fara för sig själv eller för andra och inte går med på att träffa en läkare kan du ringa hälstocentralen eller sjukhuset.
Om det behövs hjälp snabbt ska du berätta det vid samtalet.
Nämn också om du är rädd för att din närstående kommer att skada sig själv.
Om din närstående är i mycket dåligt skick och behöver akut psykiatrisk sjukhusvård kan han eller hon intas för vård mot sin vilja.
För detta behövs läkarens remiss för tvångsvård (pakkohoitolähete).
Om någon är i omedelbar livsfara kan du ringa nödnumret 112.
Ring inte nödnumret om situationen inte är akut.
Hjälp telefonledes
Kristelefon på finska: 09 2525 0111
Kristelefon för arabisktalande: 09 2525 0113.
Du kan även ringa och prata på engelska.
MIELI rf:s kristelefon erbjuder omedelbar samtalshjälp för människor i kris och deras närstående.
Samtalen besvaras av krisarbetare och utbildade frivilliga stödpersoner.
Du behöver inte uppge ditt namn när du ringer.
På kristelefonen kan du prata om en oväntad händelse eller en svår livssituation i en tillåtande och stödande atmosfär.
linkkiMIELI Psykisk Hälsa Finland rf:
Riksomfattande kristelefonfinska _ svenska _ engelska
Barn och unga
Om ditt barn är i en psykiskt påfrestande situation kan du kontakta familjerådgivningen (perheneuvola) i din hemkommun.
På familjerådgivningen kartläggs barnets situation så att barnet får den hjälp som det behöver.
Du kan också boka tid hos barnrådgivningens (lastenneuvola) psykolog eller en läkare på din egen hälsostation.
Om barnet är i skolåldern kan du kontakta skolpsykologen eller skolläkaren.
Mer information om hjälp för barn i problematiska situationer får du på InfoFinlands sida Var hittar jag hjälp när barn eller unga har problem?
Om du är ung kan du berätta om det som bekymrar dig till exempel för skolhälsovårdaren, skolpsykologen eller skolkuratorn.
Du kan också kontakta din egen hälsostation.
Läkaren kan vid behov skriva en remiss till ungdomspsykiatriska polikliniken (nuorisopsykiatrian poliklinikka).
Mer information om hjälp för unga i problematiska situationer får du på InfoFinlands sida Var hittar jag hjälp när barn eller unga har problem?
linkkiMannerheims barnskyddsförbund:
Nätstöd för ungdomar, Nuortennettifinska
linkkiMannerheims Barnskyddsförbund rf:
Stöd för föräldrarfinska
Studerande
I hälsovårdstjänsterna vid läroanstalter ordnas också mentalvårdstjänster för studerande.
Företagshälsovårdens tjänster
Om du har en anställning kan du tala med företagshälsovårdens läkare om sådant som rör den mentala hälsan.
Du kan även ha möjlighet att träffa en psykolog vid företagshälsovården.
Traumatiska upplevelser
Människor som blivit utsatta för traumatiska situationer löper risk att insjukna i posttraumatiskt stressyndrom (traumaperäinen stressihäiriö).
Upplevelser som kan orsaka ett trauma är exempelvis:
förföljelse och diskriminering
fängelse och tortyr
misshandel och våldtäkt
att bevittna våldsamma situationer
krigserfarenheter.
Vid posttraumatiskt stressyndrom väcker olika situationer minnesbilderna från den traumatiska situationen, vilket orsakar kraftig ångest.
I en sådan situation är det viktigt att man skaffar sig hjälp.
Posttraumatiskt stressyndrom påverkar inte bara den som insjuknat utan även dennes närstående.
De flesta som har insjuknat i posttraumatiskt stressyndrom återhämtar sig med rätt behandling.
Rehabiliteringscentret för tortyroffer (Kidutettujen kuntoutuskeskus) hjälper de flyktingar och asylsökande som har blivit utsatta för tortyr i sitt hemland.
Du kan kontakta centret vardagar kl. 8.30–13.30 Telefonnumret är (09) 7750 4584.
Rehabiliteringscentret för tortyrofferfinska _ engelska
Information om posttraumatiskt stressyndromfinska _ engelska _ ryska _ franska _ somaliska _ turkiska _ persiska _ arabiska _ kurdiska _ albanska _ vietnamesiska _ burmesiska _ bosniska _ serbiska _ swahili
Information på olika språk om mental hälsa på webben
På webbplatsen för MIELI Psykisk Hälsa Finland rf (MIELI Suomen Mielenterveys ry) hittar du information om
svåra livssituationer
problem med den mentala hälsan
kriser
om hur du kan söka hjälp
om hur du kan återhämta dig.
linkkiMIELI Psykisk Hälsa Finland rf:
Information om mental hälsafinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Egenvårdsläkemedel (itsehoitolääke) kan köpas utan läkarrecept.
Exempel på egenvårdsläkemedel är de flesta värkmediciner.
För många läkemedel behöver du dock ett recept, d.v.s. en läkemedelsförskrivning (lääkemääräys) för att köpa dem.
Receptet skrivs ut av en läkare.
Också många sjukskötare har rätt att skriva ut vissa läkemedel.
Till exempel antibiotika är receptbelagda läkemedel.
Om du har en långvarig sjukdom ska du ta med dina gamla recept till läkarmottagningen så kan läkaren beakta dessa när han eller hon skriver ut ett recept.
Om läkaren har skrivit ut ett elektroniskt recept (sähköinen resepti), kan du ta ut medicinerna på apoteket utan pappersrecept.
Receptet är giltigt två år från den dag det skrivits ut.
Ett recept som du skaffat utomlands är inte giltigt i Finland.
Undantag är recept som är utskrivna i de övriga nordiska länderna och europeiska recept. De är giltiga i Finland.
Du måste begära ett europeiskt recept särskilt av din läkare.
Europeiska recept kan skrivas ut av yrkesutbildade personer inom hälso- och sjukvården som arbetar i ett EU- eller EES-land eller Schweiz och har förskrivningsrätt.
På läkemedelsförpackningen står det sista användningsdatumet.
Om läkemedlet har föråldrats kan det inte längre användas.
Släng inte föråldrade läkemedel utan lämna dem alltid till apoteket (apteekki), eftersom de är problemavfall.
Information om läkemedelspreparatfinska
linkkiKanta:
Elektroniskt receptfinska _ svenska _ engelska
Var får jag läkemedel?
Du kan köpa läkemedel på apoteket.
Till apotekets tjänster hör också sidoapotek och apotekens tjänsteställen samt apotekets egen webbtjänst.
I Finland får läkemedel inte säljas annanstans.
Vitaminer och naturprodukter säljs också i vanliga butiker.
Apoteken har vanligen öppet från morgon till kväll.
I större städer kan det finnas apotek som har öppet till sent på kvällen.
På Apotekareförbundets (Apteekkariliitto) webbplats kan du söka information om apoteken på din hemort och deras öppettider.
På apoteket kan du byta ut det läkemedel som föreskrivs på receptet mot ett annat, förmånligare läkemedel om det verksamma ämnet är detsamma i båda preparaten.
Den anställda på apoteket berättar för kunden om det finns ett billigare alternativ.
linkkiSocial- och hälsovårdsministeriet:
Apotekfinska _ svenska _ engelska _ ryska
linkkiApotekareförbundet:
Apotekens kontaktuppgifterfinska
FPA-ersättning för läkemedel
Om du omfattas av den finländska sjukförsäkringen (sairausvakuutus) ersätter FPA (Kela) en del av kostnaderna för många läkemedel.
Du får ingen ersättning för läkemedel som du köper utan recept.
Man kan få ersättning först efter att den initiala självrisken (alkuomavastuu) har överskridits, det vill säga efter att du har köpt ersättningsgilla mediciner för över 50 euro under ett år.
Den initiala självrisken gäller inte mediciner för personer under 18 år.
Du kan få ersättningen redan på apoteket.
Ersättningen dras av läkemedlets pris i kassan.
Du kan också söka ersättning i efterhand med en blankett.
Bifoga apotekets utredning över de köpta läkemedlen och kassakvittot.
Mer information om vem som omfattas den finländska sjukförsäkringen får du på InfoFinlands sida Den sociala tryggheten i Finland.
Läkemedelsersättningarfinska _ svenska _ engelska
Hälsa och rehabiliteringfinska _ svenska _ ryska _ estniska
Läkemedel från utlandet
Vissa läkemedel kan du ta med dig från utlandet till Finland för eget bruk.
Importen är dock begränsad.
Begränsningarna beror på vilken sorts läkemedel det är fråga om och från vilket land du tar med dig läkemedlet till Finland.
Du måste också till exempel med ett recept eller ett läkarintyg kunna bevisa att läkemedlet är avsett för eget bruk.
Ta reda på begränsningarna innan du för in läkemedel i Finland.
Ta reda på begränsningarna också om du vill beställa läkemedel till Finland per post.
Från EES-länderna får du ta med dig den mängd läkemedel för eget bruk som motsvarar ett års förbrukning.
Per post får du från EES-länderna beställa den mängd läkemedel som motsvarar högst tre månaders förbrukning.
Från länder utanför EES-området får du ta med dig till Finland den mängd läkemedel för eget bruk som motsvarar högst tre månaders förbrukning.
Enligt lag får man inte beställa läkemedel per post från länder utanför EES-området.
Om läkemedlet har klassificerats som narkotika är begränsningarna strängare.
Om du är osäker på om ett visst läkemedel får föras in i Finland ska du fråga råd vid Tullen (Tulli).
Om du beställer läkemedel från utlandet får du ingen ersättning från FPA (Kela) för dem.
I EU-länderna finns några webbapotek där man kan lagligt köpa egenvårdsläkemedel.
Största delen av läkemedelsbutikerna på internet är dock illegala.
Det kan också vara en hälsorisk att köpa läkemedel i en olaglig webbutik.
linkkiTullen:
Personliga läkemedelfinska _ svenska _ engelska
linkkiFimea:
Införsel av läkemedel till Finlandfinska _ svenska _ engelska
linkkiFimea:
Läkemedelshandel på internetfinska _ svenska _ engelska
Du kan köpa ett graviditetstest på apoteket.
Även stora mataffärer säljer graviditetstest.
När du är gravid:
Boka en tid på mödrarådgivningen.
Besök läkaren före slutet av den fjärde graviditetsmånaden.
Om du arbetar, meddela arbetsgivaren skriftligt senast två månader innan du går på moderskapsledighet.
Boka en tid på mödrarådgivningen
När du upptäcker att du är gravid, kontakta mödrarådgivningen eller familjecentret i din hemkommun.
Du kan använda tjänsterna vid rådgivningsbyrån eller familjecentret om du har en hemkommun i Finland.
Läs mer på InfoFinlands sida Hemkommun i Finland.
Också asylsökande kan använda tjänsterna vid mödrarådgivningen.
I vissa städer får du använda tjänsterna vid mödrarådgivningen även om du vistas i Finland utan uppehållstillstånd.
På rådgivningsbyrån följer en hälsovårdare ditt hälsotillstånd och babyns hälsa.
På rådgivningsbyrån får du anvisningar för en trygg graviditet och förlossning.
Du får även viktig information om tjänsterna för barnfamiljer i Finland.
Du behöver inte betala för tjänsterna vid rådgivningsbyrån.
Barnets båda föräldrar är välkomna till rådgivningsbyrån.
Om du vill kan du även be en stödperson att följa med.
Om du behöver tolk kan sköterskan på rådgivningsbyrån be en tolk att närvara vid besöken.
Tolken ska vara vuxen.
linkkiInstitutet för hälsa och välfärd:
Broschyren Vi väntar barn(pdf, 1,46 Mt)finska _ svenska _ engelska _ ryska _ somaliska
linkkiSocial- och hälsovårdsministeriet:
Information om rådgivningsbyråernas tjänsterfinska _ svenska _ engelska _ ryska
Besök läkaren
Besök läkaren vid rådgivningsbyrån före slutet av den fjärde graviditetsmånaden.
Du kan ofta boka läkartiden via mödrarådgivningen.
När du har gjort en läkarkontroll får du ett graviditetsintyg.
Du behöver intyget om du ansöker om moderskapsledighet av din arbetsgivare.
Du behöver intyget även om du ansöker om moderskapsunderstödet och moderskapspenning hos FPA.
Läs mer om dessa förmåner på InfoFinlands sida Stöd till gravida.
På sidan Den sociala tryggheten i Finland finns information om vem som har rätt till FPA:s förmåner.
Privata mödrarådgivningar
I Finland finns även privata mödrarådgivningar.
Tänk på att privata hälso- och sjukvårdstjänster är avgiftsbelagda.
Läs mer på sidan Hälsovårdstjänster Finland.
Könsstympning och graviditet
Om du har blivit utsatt för könsstympning kan du få en öppningsoperation.
Den underlättar undersökningarna under graviditeten.
Också förlossningen blir lättare.
Öppningsoperationen kan göras före graviditeten, när graviditeten är halvvägs eller i samband med förlossningen.
Hälsovårdaren på rådgivningsbyrån frågar om du har blivit utsatt för könsstympning.
Det är viktigt att du berättar detta så att hälsovårdaren kan hänvisa dig till öppningsoperation.
Förlossningen
I Finland föder kvinnorna oftast på sjukhus.
Fråga på mödrarådgivningen på vilket sjukhus du ska föda.
Om du har en hemkommun i Finland kostar förlossningen inte särskilt mycket.
Barnets andra förälder kan vara med på förlossningen.
Om du vill kan du även be någon annan släkting eller en vän att följa med.
I Finland föder de flesta kvinnorna vaginalt.
Det är vanligtvis det tryggaste sättet.
Om det inte är möjligt fattar läkaren beslut om kejsarsnitt.
Om du är rädd inför förlossningen, prata om det på rådgivningsbyrån.
Du kan få hjälp med rädslan till exempel på polikliniken för förlossningsrädsla.
Efter förlossningen stannar du oftast några dagar på sjukhuset med barnet.
Den andra föräldern eller din stödperson kan vara på sjukhuset hela dagen för att hjälpa dig.
Om du har fått ditt första barn kan stödpersonen ofta även tillbringa nätterna på sjukhuset.
När du åker till sjukhuset ska du ta med dig tillräckligt varma kläder för barnet för hemresan.
Om du åker hem med barnet i bil, behöver du ett babyskydd i bilen.
Tolkning vid förlossningen
Man vet inte i förväg när förlossningen börjar.
Därför kan det vara svårt att få en tolk till förlossningen.
En del tolkcentraler har jour på veckoslut samt kvällar och nätter.
Du får mer information om tolktjänsterna i din kommun på rådgivningsbyrån.
Läs mer om tolktjänsterna på InfoFinlands sida Behöver du en tolk?
När barnet har fötts
På sidan När ett barn föds i Finland finns viktig information om de praktiska ärenden som du måste ta hand om när barnet har fötts.
På sidan finns till exempel information om registrering av barnet i befolkningsdatasystemet, om namnlagen i Finland och om barnets sociala trygghet.
Hjälp med babyn
Om du känner att du inte klarar dig med babyn utan hjälp kan du bo på ett mödrahem och lära dig hur du tar hand om barnet där.
Fråga om verksamheten vid din mödrarådgivning.
För mödrahemmet behöver du en remiss som utfärdas av kommunen.
Även om du inte har värk eller andra symptom, lönar det sig att regelbundet låta undersöka dina tänder.
Tandsjukdomar behandlas på bästa sätt då de upptäcks innan symptom uppkommer.
Mun- och tandhälsan påverkar hälsan i hela din kropps hälsa.
Om du har hemkommun (kotikunta) i Finland kan du utnyttja de offentliga tandvårdstjänsterna.
Mer information finns på InfoFinlands sida Hemkommun i Finland .
I nödfall får du behandling även om du inte har en hemkommun i eller uppehållstillstånd till Finland.
Det är möjligt att vårdutgifterna tas ut av dig i efterskott.
Hälso- och sjukvårdstjänster lämnas på finska och svenska i Finland.
Ofta klarar du dig också på engelska.
Om du inte kan något av dessa språk, ska du fråga om det är möjligt att anlita tolk när du bokar tid till tandvården.
Läs mer på InfoFinlands sida Behöver du en tolk?
När du har bokat tid till tandvård, är det viktigt att komma i tid.
Om du har bokat tid, men inte kan komma, är det väldigt viktigt att du avbokar besöket i tid, vanligen senast dagen innan.
Om du inte kommer och inte har avbokat tiden, måste du betala en ersättning.
linkkiSocial- och hälsovårdsministeriet:
Munhälsafinska _ svenska
Den offentliga tandvården
Kommunerna tillhandahåller tandvård vid hälsostationer (terveysasema) och tandkliniker (hammashoitola).
När du vill boka tid i tandvården ska du ringa tandvårdens tidsbeställning i din hemkommun.
Vårdbehovet bedöms ofta på telefon.
Om du inte behöver brådskande vård kan du tvingas vänta flera månader på en tid.
Intagning för vård måste ske inom sex månader.
När du vill boka tid för akut tandvård ska du ringa tandvårdens jourtidsbeställning (päivystysajanvaraus) i din hemkommun.
Kraftig värk, svullnad eller en olycka är orsaker för att få akut vård.
Brådskande fall sköts så fort som möjligt.
Kvällar och veckoslut är jourmottagningen centraliserad till större vårdenheter.
Om du bor på en liten ort kan du bli tvungen att åka till jourmottagningen i en närliggande stad.
Om du behöver mer krävande vårdåtgärder, som till exempel tandkirurgi, ska du först boka tid hos en tandläkare.
Vid behov skriver tandläkaren en remiss till specialtandvården.
Privata tandvårdstjänster
Du kan också boka tid hos en privat tandläkare.
Privat tandvård är dyrare än offentlig tandvård.
Om du omfattas av den sociala tryggheten i Finland ersätter FPA en del av kostnaderna.
FPA ersätter dock inte till exempel sådan vård som enbart har en kosmetisk effekt.
Mer information hittar du på FPA:s webbplats.
På InfoFinlands sida den sociala tryggheten i Finland får du mer information om vem som omfattas den finländska sjukförsäkringen.
Privat tandvård och ersättningarfinska _ svenska _ engelska
Jämför läkarpriserfinska _ engelska
Barn
Kommunen ordnar regelbundna tandläkarkontroller för barn.
För barn under skolåldern görs en tandläkarkontroll med ett par års mellanrum.
I en del städer kallas barnet till tandläkarkontrollen med ett brev som skickas hem.
Om tiden inte passar ska du ringa tidsbokningen och boka om tiden.
I en del städer måste man själv boka tid för kontrollen.
Barn i skolåldern går på tandläkarkontroll under skoldagen vid tandkliniken i området.
Kontroller görs i åk 1, 5 och 8.
Det är bra om föräldrarna är med på kontrollen åtminstone i åk 1.
Tandvården vid hälsovårdscentralen är kostnadsfri för barn under 18 år.
Munhälsa hos små barnfinska _ engelska
Munhälsa hos barn i skolåldernfinska _ svenska _ engelska
I Finland föder kvinnorna vanligen på sjukhus.
På rådgivningen får du information om sjukhuset eller sjukhusen i ditt område.
Om du har hemkommun i Finland får du sjukvården förmånligare.
Också en hemförlossning är möjlig, men den omfattas inte av den allmänna hälsovården och rekommenderas inte.
Detta innebär att föräldrarna själva måste sköta arrangemangen kring förlossningen.
Föräldrarna bär också ansvaret för att förlossningen förlöper bra.
Fadern är vanligtvis med på förlossningen. Stödpersonen kan också vara en släkting eller en vän.
Om du vill kan du även be att en frivillig stödperson som utbildats i att vara stödperson är med på förlossningen.
En sådan stödperson kallas doula.
Du kan fråga om doulaverksamheten på din hemort vid rådgivningen.
I Finland föder de flesta mammor vaginalt.
Det är ofta det tryggaste sättet.
Om det inte är möjligt till exempel på grund av barnets läge, fattar läkaren beslut om kejsarsnitt.
Om allt är väl i övrigt kan operationen planeras i förväg.
Ibland inleds förlossningen normalt men akut kejsarsnitt blir nödvändigt på grund av barnets tillstånd.
Om du är ängslig inför förlossningen ska du tala om det vid mödrarådgivningen.
Du kan få hjälp med din rädsla till exempel vid polikliniken för förlossningsrädsla (synnytyspelkopoliklinikka).
På mödrarådgivningen och på vissa förlossningssjukhus ordnas familjeträning som ska hjälpa modern och familjen att förbereda sig för den kommande förlossningen och att ta hand om babyn.
På familjeträningen får du också information om hur förlossningen sätter i gång och när det är dags att åka till sjukhuset.
Om ditt fostervatten går eller du har tätt återkommande smärtsamma värkar ska du ringa sjukhuset och fråga om det är dags att åka.
När du åker till sjukhuset ska du ta med dig tillräckligt varma kläder för barnet för hemresan.
Om du planerar att köra bil hem med barnet behöver du ett babyskydd (turvakaukalo) i bilen.
Tolkning vid förlossningen
Det kan vara svårt att få en tolk till förlossningen eftersom den exakta tidpunkten är svår att veta på förhand.
Vissa tolkcentraler håller vid behov jour på veckoslut och kvälls- och nattetid och även med kort varsel.
Du får mer information om tolktjänsterna i din kommun på rådgivningen.
Du kan också komma överens med personalen om att din språkkunniga make eller vän tolkar under förlossningen.
Beslutet om att använda tolk fattas av föräldrarna.
Läs mer på InfoFinlands sida Behöver du en tolk?
Omskärelse och förlossning
Om du har omskurits (ympärileikkaus) innan du kom till Finland öppnas din slidmynning med operation (avausleikkaus) i samband med förlossningen.
Öppningsoperationen kan även göras i mitten av graviditeten.
Det är bra att informera förlossningssjukhuset på förhand om omskärelsen så att det kan beaktas vid förlossningen.
linkkiInstitutet för hälsa och välfärd:
Broschyren Vi väntar barn(pdf, 1,46 Mt)finska _ svenska _ engelska _ ryska _ somaliska
I Finland kan du avbryta en graviditet i tidigt skede i följande fall:
om förlossningen kan utgöra en risk för din hälsa
om du är under 17 eller över 40 år gammal
om du redan har fött fyra barn
om du inte kan ta hand om barnet på grund av en sjukdom.
Som orsak för abort (abortti) räcker även att det med tanke på din livssituation skulle vara en alltför stor belastning att föda barnet eller att ta hand om det.
I praktiken kan orsaken vara någon av följande:
familjeförhållanden
arbetssituation
boende
Kvinnan har rätt att själv besluta om hon vill göra abort.
Partnern kan delta i beslutsfattandet om kvinnan vill ta hänsyn till hans åsikt.
Om du är minderårig och vill göra abort behöver du inte tillstånd av dina föräldrar.
Det är dock ofta bra att diskutera saken med föräldrarna.
Om du ändå inte vill göra det har de yrkesutbildade personerna inom hälsovården tystnadsplikt.
Aborten ska göras före den tolfte graviditetsveckan.
Av speciellt vägande skäl kan abort göras även senare men då behöver du ett specialtillstånd från Valvira (Valvira).
Du behöver tillstånd från Valvira även om aborten görs på grund av att fostret har en svår sjukdom eller ett handikapp.
Fråga mer av läkaren vid din egen hälsostation (terveysasema).
Om du vill avbryta graviditeten ska du kontakta hälsostationen i ditt eget område så fort som möjligt och boka tid hos en läkare.
Du kan också boka tid hos en privatläkare, men kontrollera när du bokar tiden att läkaren har Valviras tillstånd att ge ett utlåtande för abort.
Om du vill kan du ta med dig din partner till läkarmottagningen.
Läkaren skriver en remiss till det sjukhus där aborten görs.
På sjukhuset samtalar en skötare och en läkare med dig.
Ni fattar gemensamt beslutet om på vilket sätt graviditeten avbryts.
På detta inverkar hur långt graviditeten har gått och din egen åsikt.
Graviditeten avbryts med läkemedel eller med skrapning (kaavinta).
Skrapning görs vanligtvis i narkos och därefter ska du stanna några timmar på sjukhuset.
Om aborten görs medicinskt doseras läkemedlet med 1–3 dagars mellanrum via slidan så att livmoderns börjar dras samman och töms.
Var förberedd på att du behöver smärtlindring när livmodern dras samman.
Ibland behövs det skrapning efter medicinsk abort.
2–4 veckor efter aborten görs en efterkontroll på hälsostationen.
När du ska fatta beslut om abort får du stöd till exempel av en hälsovårdare eller en läkare vid hälsostationen.
Mer information om olika ställen där du får hjälp i en krävande livssituation finns på InfoFinlands sida Mental hälsa.
Abortfinska
Tillstånd till att avbryta graviditetenfinska _ svenska
Om ditt barn har hemkommun (kotikunta) i Finland har han eller hon rätt att utnyttja de offentliga hälsovårdstjänsterna.
Läs mer på InfoFinlands sida Hemkommun i Finland.
Om du omfattas av den finländska sjukförsäkringen (sairausvakuutus) kan du teckna en försäkring för ditt barn som täcker en del av kostnaderna för privata hälsovårdstjänster.
När ett barn insjuknar
Om barnet har feber eller annars är sjukt ska det inte tas till dagvården.
Om barnet har hosta eller snuva, men annars mår bra, kan barnet vara i dagvården.
Om ett barn under 10 år insjuknar akut kan barnets mamma eller pappa stanna hemma för att ta hand om barnet.
Vårdledigheten kan vara högst fyra dagar.
I kollektivavtalet bestäms om man får lön för denna tid eller inte.
Om ett barn blir sjukt under skoldagen vårdas han eller hon i skolan.
Vid behov förs barnet till stadens hälsostation.
Om ett sjukt barn behöver läkarhjälp eller uppsöka hälsovårdare ska du kontakta hälsostationen (terveysasema) eller en privat läkarstation i din hemkommun.
Hälsostationerna har öppet från måndag till fredag, vanligen kl. 8–16.
Det är bäst att ringa hälsostationen genast på morgonen när tidsbeställningen öppnar.
Vid tidsbeställningen bedöms vilken slags vård barnet behöver.
Kvällstid och under veckoslut har hälsostationerna stängt.
Då vårdas akuta sjukfall och olycksfall på jourmottagningen (päivystys).
Om barnets sjukdom inte kräver omedelbar vård ska du vänta tills din hälsostation har öppet igen.
Jourmottagningen för barn och unga finns ofta i en separat enhet.
Du kan också boka tid till läkare på en privat hälsostation.
De har ofta öppet också på kvällarna och ibland får man fortare en tid där.
Privata hälsovårdstjänster är dock avsevärt dyrare för kunden än offentliga.
Om du misstänker att ett barn har förgiftats kan du fråga råd vid Giftinformationscentralen (Myrkytystietokeskus).
Giftinformationscentralens telefontjänst är öppen 24 timmar om dygnet. Telefonnumret är (09) 471 977.
Om ett barn är i livsfara eller har hamnat i en olycka ska du ringa nödnumret (hätänumero) 112.
Ambulanser är endast avsedda för allvarliga och brådskande situationer.
Ring inte nödnumret vid vanliga sjukdomsfall.
Om barnet insjuknarfinska _ svenska _ engelska
Sjukvårdsersättningarfinska _ svenska _ engelska
Småbarns hälsa
Hälsotillståndet hos barn under skolåldern följs i barnrådgivningen (lastenneuvola).
Barnrådgivningen följer och stöder den fysiska, psykiska och sociala tillväxten och utvecklingen av barn under skolåldern.
På barnrådgivningen besöker barnen en läkare eller en hälsovårdare.
Familjen till ett barn som är under ett år gammalt kallas till barnrådgivningen minst nio gånger.
Efter det första året kallas man till barnrådgivningen ännu minst sex gånger.
Hälsovårdaren följer barnets utveckling, vaccinerar barnet och ger information om rätt kost.
Hälsovården besöket barnet också hemma direkt efter födseln.
Rådgivningsbyråns tjänster i den egna kommunen är kostnadsfria.
Du kan utnyttja barnrådgivningsbyråns tjänster i din egen kommun om du har hemkommun i Finland.
Mer information finns på InfoFinlands sida Hemkommun i Finland.
Du ska ha med dig kortet på varje besök till rådgivningen.
Hälsovårdaren antecknar uppgifter om barnets hälsa och vaccinationer på kortet.
linkkiSocial- och hälsovårdsministeriet:
Information om rådgivningsbyråernas tjänsterfinska _ svenska _ engelska _ ryska
Skolbarns hälsa
Varje skola har en läkare och en hälsovårdare.
Hälsovårdaren undersöker barnen i skolan.
Hälsovårdaren är på plats i skolan vissa dagar i veckan.
Eleverna kan själva besöka hälsovårdarens mottagning om de har problem.
Vid ett olycksfall i skolan får barnet första hjälpen.
Mer information om skolhälsovården finns på social- och hälsovårdsministeriets (Sosiaali- ja terveysministeriö) webbplats.
linkkiSocial- och hälsovårdsministeriet:
Skolhälsovårdfinska _ svenska
Vaccinationer
I Finland kan barnen vaccineras (rokotus) mot många smittsamma sjukdomar.
Vaccinationerna ges på barnrådgivningen (lastenneuvola) och inom skolhälsovården.
De vaccinationer som ingår i vaccinationsprogrammet är avgiftsfria för familjen.
Vaccinationerna är frivilliga.
De flesta barn i Finland får de vaccinationer som ingår i vaccinationsprogrammet.
Berätta för hälsovårdaren vilka vaccinationer ditt barn har fått innan ni kom till Finland.
Om du vill att ditt barn ska få en vaccination som inte ingår i vaccinationsprogrammet ska du beställa tid till en läkare.
Läkaren kan skriva ett recept på vaccinationen och hälsovårdaren kan vaccinera ditt barn.
Du köper själv vaccinationen på apoteket.
linkkiInstitutet för hälsa och välfärd:
Vaccinationsprogrammet i Finlandfinska _ svenska
Långvarig sjukdom och vård av ett handikappat barn
Om du under en lång tid tar hand om ett sjukt eller handikappat barn under 16 år kan du söka specialvårdpenning (erityishoitoraha) från FPA.
Från FPA kan du även få bidrag för rehabilitering (kuntoutus) av barnet.
Ett barn med en svår sjukdom eller ett handikapp kan även få FPA:s handikappbidrag för barn under 16 år (alle 16-vuotiaan vammaistuki).
FPA:s bidrag är avsedda för personer som omfattas av Den sociala tryggheten i Finland.
Du får mer information om att leva i Finland med ett handikappat barn på InfoFinlands sida Ett handikappat barn.
Specialvårdspenning för barn under 16 årfinska _ svenska _ engelska
Handikappbidrag för barnfinska _ svenska _ engelska
Omskärelse av pojkar
Omskärelse (ympärileikkaus) är alltid ett oåterkalleligt ingrepp.
Om det görs av icke-medicinska orsaker, inkräktar man på en pojkes fysiska integritet.
Omskärelse får endast göras av en legitimerad läkare.
För omskärelse behövs ett skriftligt samtycke av pojkens vårdnadshavare.
Om barnet har två vårdnadshavare, behövs varderas samtycke, i annat fall kan ingreppet inte göras.
Pojken har rätt att vägra att gå med på operationen.
Omskärelse får inte göras utan smärtlindring som ges av läkare, och det ska göras i en steril miljö.
Icke-medicinsk omskärelse omfattas inte av den offentligt finansierade hälsovården, och kan därför inte göras på en offentlig hälsostation, och man måste själv betala det.
Fråga mer om omskärelse på rådgivningen, av läkaren på hälsostationen, skolhälsovårdaren eller skolläkaren.
Omskärelse av flickor
Omskärelse (ympärileikkaus) av flickor är ett brott i Finland. Man kan få ett flera års fängelsestraff för det.
Det är också ett brott att föra en flicka till ett annat land, för att låta henne genomgå omskärelse där.
Omskärelse av kvinnor och flickorfinska _ engelska _ somaliska _ arabiska
Om du misstänker att du är gravid kan du göra ett graviditetstest (raskaustesti).
Graviditetstest kan köpas till exempel på apoteket.
När du är gravid:
Ta kontakt med mödrarådgivningen (äitiysneuvola) i din hemkommun.
Låt göra en läkarundersökning före utgången av den fjärde graviditetsmånaden.
Gör en skriftlig anmälan till din arbetsgivare senast två månader innan du blir moderskapsledig.
Mödrarådgivningen
På mödrarådgivningen får du handledning i allt som rör din graviditet och information om olika tjänster som samhället tillhandahåller.
På mödrarådgivningen följs också moderns och fostrets hälsotillstånd.
Rådgivningstjänsterna i den egna hemkommunen är gratis.
Du kan använda mödrarådgivningstjänsterna i din hemkommun om du har hemkommun (kotikunta) i Finland.
Mer information finns på InfoFinlands sida Hemkommun i Finland.
Också pappor är välkomna till rådgivningen.
På rådgivningen diskuteras parförhållandet och föräldraskapet samt papparollen och föräldrarnas ansvar.
Rådgivningen ordnar också förlossningsförberedelse och familjeträning för blivande mammor och pappor.
De flesta finländska pappor och mammor deltar i denna utbildning.
Rådgivningens skötare kan vid behov beställa en tolk som deltar i rådgivningsmötena.
Tolken ska vara vuxen, egna minderåriga barn kan alltså inte användas som tolk.
Mödrarådgivningen ger alla blivande föräldrar broschyren Vi väntar barn som ges ut av Institutet för hälsa och välfärd (Terveyden ja hyvinvoinnin laitos).
Det är bra att gå på läkarundersökning första gången före utgången av den fjärde graviditetsmånaden.
Då får du ett graviditetsintyg av läkaren eller från rådgivningen.
Det behöver du när du ansöker om moderskapsunderstöd (äitiysavustus) och moderskapspenning (äitiysraha) hos FPA (Kela).
Mer information finns på InfoFinlands sida Stöd till gravida.
På social- och hälsovårdsministeriets (Sosiaali- ja terveysministeriö) sidor finns allmän information om rådgivningsverksamheten i Finland.
linkkiInstitutet för hälsa och välfärd:
Broschyren Vi väntar barn(pdf, 1,46 Mt)finska _ svenska _ engelska _ ryska _ somaliska
linkkiSocial- och hälsovårdsministeriet:
Information om rådgivningsbyråernas tjänsterfinska _ svenska _ engelska _ ryska
Smärtor och blödningar under graviditeten
Små smärtor hör till en normal graviditet när livmodern växer.
Om du är osäker på om smärtan är normal ska du fråga råd vid din egen rådgivningsbyrå.
Om du har kraftiga smärtor eller blödningar ska du kontakta sjukhuset.
Vid behov kallas du till undersökning.
I brådskande fall behöver du ingen remiss.
Omskärelse och graviditet
Om du har omskurits innan du kom till Finland öppnas din slidmynning med operation (avausleikkaus) i samband med förlossningen.
Öppningsoperationen kan även göras i mitten av eller före graviditeten.
Öppningsoperationen gör förlossningen och undersökningarna under graviditeten lättare.
Operationen görs på sjukhus och återhämtningen tar vanligtvis 1–2 dagar.
Fråga mer av mödrarådgivningens hälsovårdare.
Stöd till gravida
Om du omfattas av den sociala tryggheten i Finland har du rätt till olika understöd från FPA under och efter graviditeten.
Läs mer på InfoFinlands sida Stöd till gravida och Stöd efter barnets födelse.
Sköta ärenden på Internetfinska _ svenska _ engelska
Kontaktuppgifter till kontorenfinska _ svenska _ engelska
Elektronisk tidsbeställningfinska _ svenska _ engelska
Vad ska jag göra om jag inte har hemkommun i Finland?
Ta kontakt med en privat läkarstation.
På de största orterna finns flera privatläkare och på somliga orter också privata rådgivningsbyråer.
Beakta att den privata hälsovården är dyr.
Du kan inte få en finsk personförsäkring om du inte omfattas av den sociala tryggheten i Finland.
Väntar du barn ensam eller i en svår livssituation?
Om du väntar barn och känner att du inte klarar dig på egen hand kan du kontakta ett mödrahem (ensikoti).
På mödrahemmet får du hjälp med föräldraskapet och livskompetensen.
Fråga om mödrahemsverksamheten på din egen rådgivningsbyrå.
Mödrahemmets tjänster är avsedda för personer som har hemkommun i Finland.
Du behöver också ett följebrev från kommunens socialväsen.
Mer information om rätten till hemkommun finns på InfoFinlands sida Hemkommun i Finland.
Överväger du att avbryta graviditeten?
Läs mer på InfoFinlands sida Abort.
linkkiFörbundet för mödra- och skyddshem:
Kontaktuppgifter till mödrahemfinska
I Finland tillhandahåller både den offentliga och den privata hälso- och sjukvården tjänster inom graviditetsprevention, gynekologi, tidig upptäckt av cancer, sexuell hälsa hos män, barnlöshet och könssjukdomar.
Har du rätt till de offentliga hälsovårdstjänsterna?
Läs mer på sidan Hälsovårdstjänster Finland.
Ungas sexualitetfinska _ engelska
Vuxnas sexualitetfinska _ svenska _ engelska
Du kan köpa kondomer i affärer, på bensinstationer, kiosker och apotek.
Du behöver inget recept.
För hormonella preventivmedel behöver du ett recept av en läkare.
Sådana preventivmedel är till exempel p-piller och minipiller.
De säljs på apoteket.
Du kan boka en tid på hälsostationen eller vid en privat läkarstation.
Även minderåriga barn kan boka tid hos läkaren och få ett recept för preventivmedel.
Du behöver inte tillstånd av dina föräldrar för receptet.
Vissa kommuner erbjuder unga kostnadsfria preventivmedel.
Du kan fråga om detta på hälsostationen eller av skolhälsovårdaren.
Om preventionen misslyckades eller om du glömde att använda preventivmedel kan du köpa ett akut p-piller på apoteket utan recept.
Du ska ta pillret så snart som möjligt efter samlaget, i regel senast inom 72 timmar.
Vissa preparat kan tas inom 120 timmar efter samlaget.
linkkiSHVS:
Graviditetspreventionfinska _ svenska _ engelska
Sexuell hälsa hos kvinnor
Alla läkare på hälsostationen gör gynekologiska undersökningar.
Fråga mer på din hälsostation.
Om du vill träffa en kvinnlig läkare, ange detta när du bokar tiden.
Läkaren kan vid behov skriva remiss till en specialist på gynekologiska polikliniken.
Du kan även boka tid hos en privat gynekolog.
Då kan du välja läkaren själv.
Tjänsterna hos privatläkare är mycket dyrare för klienten.
I Finland ordnas regelbundna screeningundersökningar för kvinnor i vissa åldrar.
På så sätt försöker man i ett tidigt skede hitta bröstcancer och livmoderhalscancer.
Undersökning av bröstcancer görs på kvinnor i åldern 50–69 år ungefär vartannat år.
Undersökning av livmoderhalscancer görs på kvinnor i åldern 30–60 år vart femte år.
linkkiSocial- och hälsovårdsministeriet:
Screeningsundersökningarfinska _ svenska _ engelska _ ryska
linkkiInstitutet för hälsa och välfärd:
Information om bröstcancerscreeningfinska _ svenska
Anvisning för identifiering av bröstcancer(pdf, 440kt)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ kinesiska _ thai _ rumänska _ samiska
Information om cancerscreeningfinska _ svenska _ engelska
Sexuell hälsa hos män
Du kan boka en läkartid på din egen hälsostation.
Om du vill kan du be om att få träffa en manlig läkare.
Läkaren kan vid behov skriva remiss till en specialist på urologiska polikliniken.
Du kan även boka tid på en privat läkarstation.
Tjänsterna hos privatläkare är mycket dyrare för klienten.
Barnlöshet
Barnlöshet kan oftast behandlas.
Orsaken till barnlöshet kan finnas hos kvinnan eller hos mannen.
Ibland hittar man ingen medicinsk orsak till den.
Om du har slutat använda preventivmedel, men en graviditet inte har börjat inom ett år, boka tid på hälsostationen eller hos en privat gynekolog.
Det är bra om paret besöker mottagningen tillsammans.
Läkaren skriver en remiss till undersökningar på barnlöshetspolikliniken.
Med undersökningarna utreds varför en graviditet inte har börjat.
Fertilitetsbehandlingar tillhandahålls av både offentliga och privata kliniker. till exempel kvinnans ålder påverkar rätten till fertilitetsbehandling inom de offentliga hälsovårdstjänsterna.
Könssjukdomar
Om du misstänker att du har en könssjukdom kan du boka en läkartid på hälsostationen eller en privat läkarstation.
I vissa städer finns en poliklinik för könssjukdomar där könssjukdomar behandlas.
Fråga mer på din hälsostation.
Du kan skydda dig mot de flesta könssjukdomarna med kondom eller slicklapp.
Också papperslösa och asylsökande har rätt att få behandling för könssjukdomar.
Om du vistas i Finland utan uppehållstillstånd kan du emellertid bli tvungen att betala för vården.
linkkiHivpoint:
Broschyren Information om sexuellt överförda sjukdomar(pdf, 1500kt)finska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
linkkiHivpoint:
Info om HIVfinska _ engelska _ ryska
linkkiHivpoint:
Broschyren Ett gott liv med HIVfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ thai
linkkiHivpoint:
Broschyren HIV i familjen(pdf, 881 kb)finska _ engelska _ ryska
Manlig omskärelse
Fundera noga på om omskärelse behövs.
Om pojken är gammal nog för att säga sin åsikt ska han tillfrågas om han samtycker till operationen.
Operationen får inte göras om pojken motsätter sig.
Om pojken har två vårdnadshavare måste båda ge sitt skriftliga samtycke till operationen.
Om det inte finns några medicinska skäl till omskärelsen kan den inte utföras inom den offentliga hälsovården.
Då måste du betala för operationen själv.
Endast en läkare får utföra operationen.
Den ska göras i steril miljö.
Läkaren ska se till att patienten får smärtlindring.
Fråga mer om omskärelse på rådgivningsbyrån, en hälsostationsläkare, skolhälsovårdaren eller skolläkaren.
Kvinnlig könsstympning
Könsstympning av flickor är ett brott i Finland.
Man kan få ett flerårigt fängelsestraff för det.
Det är likaså brottsligt att ta flickan utomlands för könsstympning.
Om du har blivit utsatt för detta kan du få en öppningsoperation.
Även en korrigerande operation är möjlig.
Fråga mer på din hälsostation.
Omskärelse av kvinnor och flickorfinska _ engelska _ somaliska _ arabiska
Vilka hälsotjänster kan du använda?
Offentliga hälsovårdstjänster
Privata hälsovårdstjänster
Hälsovård för medborgare i de nordiska länderna
Hälsovård för EU-medborgare
Hälsovård för anställda och företagare
Hälsovård för studerande
Hälsovård för invandrare och asylsökande
Hälsovård för papperslösa
Information på webben
Vilka hälsotjänster kan du använda?
Du kan utnyttja de offentliga hälsovårdstjänsterna i Finland om du har hemkommun (kotikunta) i Finland.
Rätten till hemkommun beror på följande:
från vilket land du kommer till Finland
varför du kommer till Finland (t.ex. arbete, studier)
om du ska bo stadigvarande i Finland eller vistas här tillfälligt
om din vistelse i Finland är tillfällig, beroende på hur länge vistelsen varar.
Om du inte är säker på om du har hemkommun i Finland kan du ta reda på din situation vid magistraten (maistraatti).
Mer information finns på InfoFinlands sida Hemkommun i Finland.
Om du inte har en hemkommun i Finland eller om du inte omfattas av sjukförsäkringen i Finland, kan du ändå ha rätt till vård eller ersättningar från FPA på någon annan grund.
Du måste ansöka separat om denna rätt.
Fråga mer hos FPA:s center för internationella ärenden.
Tfn 020 634 0200 (finska och engelska), 020 634 0300 (svenska)
Så här ansöker du om rätt till sjukvård hos FPAfinska _ svenska _ engelska
I nödfall får du vård inom den offentliga hälso- och sjukvården fastän du inte har en hemkommun i Finland eller rätt till vård på grund av arbete.
Du kan krävas på vårdkostnaderna i efterhand.
Om du inte har rätt till de offentliga hälsovårdstjänsterna, kan du boka tid på en privat läkarstation.
Privata hälsovårdstjänster är avsevärt dyrare för kunden än de offentliga.
Hälsovårdstjänster ges i Finland på finska och svenska.
Ofta klarar man sig även på engelska.
När du bokar tid till hälsovårdstjänster kan du fråga om möjligheten att använda en tolk (tulkki) om du inte behärskar dessa språk.
Läs mer på InfoFinlands sida Behöver du en tolk?
När du har bokat tid för ett läkarbesök ska du vara punktligt på plats.
Om du har bokat tid för ett läkarbesök men får förhinder är det mycket viktigt att du avbokar besöket i god tid, helst dagen innan.
Om du inte kommer och inte heller har avbokat din tidsbeställning måste du betala en avgift.
Hälsa och rehabiliteringfinska _ svenska _ ryska _ estniska
Sjukvård för utlänningar i Finlandfinska _ svenska _ engelska
Kontaktpunkt för gränsöverskridande hälso- och sjukvårdfinska _ svenska _ engelska
linkkiStödcentralen Hilma för funktionshindrade invandrare :
Handbok med ordlista i hälso- och sjukvård på finska(pdf, 341,02 kt)finska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska
Offentliga hälsovårdstjänster
När du blir sjuk ska du först kontakta din egen hälsostation (terveysasema). Där kan du boka tid hos en allmänläkare eller en hälsovårdare.
Mer information om hälsovårdstjänsterna i olika kommuner hittar du på InfoFinlands sida på de lokala informationssidorna eller på din egen kommuns sida.
Hälsostationens tjänster är relativt förmånliga för klienten eftersom de finansieras med skattemedel.
Hälsostationerna har vanligen öppet från måndag till fredag kl. 310 1671.
Det är klokt att ringa tidsbeställningen genast på morgonen när hälsostationen öppnar.
Om ditt besvär kräver brådskande vård får du en tid snabbt.
Om du inte behöver brådskande vård måste du vänta längre på att få en läkartid.
Vid tidsbeställningen får du veta hur snabbt du kommer att få vård.
Vid tidsbeställningen bedöms även om du behöver vård av läkare eller hälsovårdare.
I Finland kan hälsovårdare ge vård vid flera sjukdomar.
Vid behov kan hälsovårdaren ge remiss till läkare.
Om du har ett FPA-kort (Kela-kortti) ska du ta det med när du besöker hälsovårdsstationen.
Om du behöver en specialist, ska du först boka tid hos en allmänläkare.
Vid behov skriver hälsostationsläkaren en remiss till en specialist.
Specialister finns på vissa hälsostationer, på polikliniker och sjukhus.
Specialsjukvård ges på centralsjukhus och universitetssjukhus.
I Finland gör läkare inom de offentliga hälsovårdstjänsterna inga hembesök.
En del privata läkarstationer erbjuder denna tjänst. Ett hembesök av en privatläkare är dock dyrt.
Om din sjukdom är långvarig och du inte kan arbeta finns det mer information om FPA:s sjukpenning på InfoFinlands sida Stöd när du är sjuk.
Jour inom offentliga hälsovårdstjänster
Hälsostationerna har stängt kvällstid och under veckoslut.
Då vårdas akuta sjukfall på jourmottagningen (päivystys).
Jourmottagningen är avsedd för situationer där man behöver omedelbar vård.
Om din sjukdom inte kräver omedelbar vård ska du beställa tid på din egen hälsostation nästa gång den har öppet.
Jourmottagningen finns ofta i anslutning till sjukhus, i små städer också i en närliggande stad.
Jourmottagningen för barn och unga finns ofta separat.
Fråga mer vid din egen hälsostation under dess öppettider eller leta upp informationen på din hemkommuns webbplats.
Privata hälsovårdstjänster
Kontaktuppgifter till privata läkarstationer hittar du till exempel på internet.
Förmodligen får du en tid snabbare på en privat hälsostation än inom den offentliga hälsovården.
Privata hälsotjänster är avsevärt dyrare för klienten än de offentliga.
Olika läkarstationer erbjuder olika tjänster.
Privata hälsotjänster kan användas av alla, även personer som inte har en hemkommun i Finland.
Om du omfattas av den finländska sjukförsäkringen (sairausvakuutus) ersätter FPA en liten del av kostnaderna för privat sjukvård och tandvård.
Ibland kan också personer som inte omfattas av den finländska sjukförsäkringen ha rätt till ersättning från FPA.
Fråga mer hos FPA.
FPA:s ersättning kan ibland dras av direkt på det belopp som du betalar vid kassan.
Du kan också söka ersättning från FPA i efterhand.
Läs mer om sjukförsäkringen i Finland på InfoFinlands sida Den sociala tryggheten i Finland.
Sjukvårdsersättningarfinska _ svenska _ engelska
Jämför läkarpriserfinska _ engelska
Privat läkarstationfinska _ svenska _ engelska
Privat läkarstationfinska _ svenska _ engelska
linkkiAava:
Privat läkarstationfinska _ svenska _ engelska
Hälsovård för medborgare i de nordiska länderna
Om du har en sjukförsäkring i ett annat nordiskt land har du rätt till nödvändig sjukvård i Finland.
Du får vård på samma villkor och till samma kostnad som finländarna.
Ta med dig ett officiellt identitetsbevis när du använder hälsovårdstjänsterna.
Hälsovård för EU-medborgare
Om du har en sjukförsäkring i ett annat EU-land, EES-land eller i Schweiz har du rätt till nödvändig sjukvård i Finland.
För att få vård måste du ha ett europeiskt sjukvårdskort.
Du ska skaffa dig det europeiska sjukvårdskortet i det land där du har din sjukförsäkring.
Det europeiska sjukvårdskortet ger dig rätt till vård om du blir sjuk eller råkar ut för en olycka.
Du får vård även vid en långvarig sjukdom.
Med kortet får du även vård i samband med graviditet och förlossning.
Du får vård till samma kostnad som personer som är stadigvarande bosatta i Finland.
Information om det europeiska sjukvårdskortetfinska _ svenska _ engelska
Hälsovård för anställda och företagare
Om du har kommit till Finland för att arbeta kan du ha rätt att använda de offentliga hälsovårdstjänsterna i Finland.
Detta beror på hurdant och hur långt arbetsavtal du har samt från vilket land du har kommit till Finland.
I Finland är arbetsgivare skyldiga att ordna förebyggande företagshälsovård för sina anställda.
Företagare kan ordna sin egen företagshälsovård om de vill.
Företagare måste alltså inte ordna företagshälsovård för sig.
Företagare måste ändå ordna företagshälsovård för sina anställda.
Företagshälsovården kan ordnas vid den lokala hälsovårdscentralen eller till exempel på en privat läkarcentral.
Mer information får du på InfoFinlands sida Företagshälsovården och på social- och hälsovårdsministeriets webbplats.
linkkiSocial- och hälsovårdsministeriet:
Företagshälsovårdfinska _ svenska _ engelska
Hälsovård för studerande
Om du kommer från ett land som inte är ett EU-land, ett EES-land eller Schweiz till Finland för att studera behöver du vanligtvis ha en täckande sjukförsäkring i ditt hemland för att få uppehållstillstånd i Finland.
Om dina studier beräknas pågå i minst två år får du vanligen en hemkommun i Finland och rätt till de kommunala hälsovårdstjänsterna.
I detta fall räcker det om din sjukförsäkring i första hand täcker läkemedelskostnaderna.
Om du inte är säker på om du har rätt till hemkommun i Finland kan du kontrollera detta vid magistraten.
Du får mer information om hemkommun på InfoFinlands sida Hemkommun i Finland.
Mer information om uppehållstillstånd för studerande och om den sjukförsäkring som krävs för att få uppehållstillstånd får du på Migrationsverkets (Maahanmuuttovirasto) webbplats.
I Finland omfattas högskolestuderande av studerandehälsovården.
Fråga mer vid din egen läroanstalt.
Mer information om studerandehälsovården får du på Studenternas hälsovårdsstiftelses (SHVS) (YTHS) och social- och hälsovårdsministeriets (Sosiaali- ja terveysministeriö) webbplatser.
Information om uppehållstillstånd för studierfinska _ svenska _ engelska
linkkiSHVS:
Hälsovård för högskolestuderandefinska _ svenska _ engelska
linkkiSocial- och hälsovårdsministeriet:
Studerandehälsovårdfinska _ svenska
Hälsovård för invandrare och asylsökande
Om du har kommit till Finland som kvotflykting har du hemkommun i Finland och rätt att utnyttja de offentliga hälsovårdstjänsterna.
Om du är asylsökande och din ansökan inte ännu har behandlats kan du inte registrera dig i magistraten som kommuninvånare och inte heller utnyttja kommunens hälsovårdstjänster.
Fråga mer vid din förläggning.
Om du har fått uppehållstillstånd på grund av behovet av skydd och får rätt till hemkommun i Finland, kan du utnyttja hälsovårdstjänsterna i din egen kommun.
Läs mer om rätten till hemkommun på InfoFinlands sida Hemkommun i Finland.
Hälsovård för papperslösa
Global Clinic är en klinik där du kan få hjälp eller råd av en läkare eller sjukskötare om du vistas i Finland utan uppehållstillstånd.
Global Clinic bedriver verksamhet i följande städer:
Åbo
Uleåborg
Joensuu
Tammerfors
Du kan ringa eller skicka e-post.
En sjukskötare eller läkare besvarar ditt samtal.
Du hittar kontaktinformation på Global Clinic:s hemsidor.
Global Clinic:s tjänster är avgiftsfria för kunderna.
Global Clinic anmäler inte sina kunder till polisen eller andra myndigheter.
Klinikens adress eller öppettider meddelas inte offentligt.
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Information på webben
linkkiTuberkuloosi.fi:
Information om tuberkulosfinska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska _ portugisiska _ tagalog _ polska _ bosniska _ rumänska _ swahili
_ lettiska
_ litauiska
I Finland kan du avbryta en graviditet i tidigt skede i följande fall:
om förlossningen kan utgöra en risk för din hälsa
om du är under 17 eller över 40 år gammal
om du redan har fött fyra barn
om du inte kan ta hand om barnet på grund av en sjukdom.
Som orsak för abort (abortti) räcker även att det med tanke på din livssituation skulle vara en alltför stor belastning att föda barnet eller att ta hand om det.
I praktiken kan orsaken vara någon av följande:
familjeförhållanden
arbetssituation
boende
Kvinnan har rätt att själv besluta om hon vill göra abort.
Partnern kan delta i beslutsfattandet om kvinnan vill ta hänsyn till hans åsikt.
Om du är minderårig och vill göra abort behöver du inte tillstånd av dina föräldrar.
Det är dock ofta bra att diskutera saken med föräldrarna.
Om du ändå inte vill göra det har de yrkesutbildade personerna inom hälsovården tystnadsplikt.
Aborten ska göras före den tolfte graviditetsveckan.
Av speciellt vägande skäl kan abort göras även senare men då behöver du ett specialtillstånd från Valvira (Valvira).
Du behöver tillstånd från Valvira även om aborten görs på grund av att fostret har en svår sjukdom eller ett handikapp.
Fråga mer av läkaren vid din egen hälsostation (terveysasema).
Om du vill avbryta graviditeten ska du kontakta hälsostationen i ditt eget område så fort som möjligt och boka tid hos en läkare.
Du kan också boka tid hos en privatläkare, men kontrollera när du bokar tiden att läkaren har Valviras tillstånd att ge ett utlåtande för abort.
Om du vill kan du ta med dig din partner till läkarmottagningen.
Läkaren skriver en remiss till det sjukhus där aborten görs.
På sjukhuset samtalar en skötare och en läkare med dig.
Ni fattar gemensamt beslutet om på vilket sätt graviditeten avbryts.
På detta inverkar hur långt graviditeten har gått och din egen åsikt.
Graviditeten avbryts med läkemedel eller med skrapning (kaavinta).
Skrapning görs vanligtvis i narkos och därefter ska du stanna några timmar på sjukhuset.
Om aborten görs medicinskt doseras läkemedlet med 1–3 dagars mellanrum via slidan så att livmoderns börjar dras samman och töms.
Var förberedd på att du behöver smärtlindring när livmodern dras samman.
Ibland behövs det skrapning efter medicinsk abort.
2–4 veckor efter aborten görs en efterkontroll på hälsostationen.
När du ska fatta beslut om abort får du stöd till exempel av en hälsovårdare eller en läkare vid hälsostationen.
Mer information om olika ställen där du får hjälp i en krävande livssituation finns på InfoFinlands sida Mental hälsa.
Abortfinska
Tillstånd till att avbryta graviditetenfinska _ svenska
När ska jag söka hjälp?
Vem som helst kan behöva hjälp om livssituationen är påfrestande.
Livet kan vara svårt till exempel när man flyttar från ett land till ett annat, har problem på arbetsplatsen, förlorar sin arbetsplats, har problem i familjen, går igenom skilsmässa, förlorar en anhörig, blir sjuk eller när livet förändras på andra sätt.
Också positiva saker, t.ex. att man får barn, kan ändra livet så mycket att man behöver stöd i den nya situationen.
Ibland kan man må dåligt först i efterhand när man redan har lagt den svåra erfarenheten bakom sig och situationen har lugnat ner sig.
Det lönar sig att söka hjälp, om du har något av följande symptom:
sömnlöshet
ingen aptit
vardagen känns tung
du orkar inte arbeta eller träffa människor
fysiska symptom, utan att medicinska orsaker hittas för dessa
ökad alkohol- eller droganvändning
Det är inte ovanligt att söka hjälp för att få stöd med den mentala hälsan.
I Finland lider 20 % av befolkningen av depression i något skede av livet.
Depression(pdf, 110,37 kt)finska _ engelska _ ryska _ franska _ somaliska _ turkiska _ persiska _ arabiska _ kurdiska _ albanska _ vietnamesiska _ burmesiska _ bosniska _ serbiska _ swahili
Var får jag hjälp?
Ofta hjälper det redan att tala om dessa saker med familjen eller vänner. Ibland behövs det även annan hjälp.
Det kan hjälpa att tala med en hälsovårdare (terveydenhoitaja), läkare (lääkäri) eller en psykoterapeut (psykoterapeutti).
Tillsammans kan ni fundera på vilken sorts stöd som skulle passa just dig.
Ofta hjälper terapi, medicinering eller en kombination av båda.
Ibland behövs sjukhusvård.
Sjukhusvården räcker vanligen några veckor.
Målsättningen är att patienten kan återvända hem så fort som möjligt.
Därefter fortsätter vården som öppenvård.r.
Om du har hemkommun i Finland ska du först kontakta din egen hälsostation (terveysasema).
Hälsostationerna har vanligen öppet från måndag till fredag, ungefär kl. 8–16.
Ring hälsostationen genast på morgonen för att boka tid.
Om du behöver hjälp genast ska du tala om det när du ringer.
Läkaren skriver vid behov en remiss till psykiatriska polikliniken (psykiatrian poliklinikka) eller en annan vårdenhet för psykisk hälsa.
Du kan inte gå till polikliniken utan en läkarremiss.
Med läkaren eller psykologen kan du samtala konfidentiellt. De har tystnadsplikt.
De berättar inte om dina saker för andra myndigheter.
Om någon annan hälsovårdsenhet behöver dina uppgifter, ombeds du ge ditt medgivande för överlåtelse av dessa.
På din egen hälsostation får du mer information om hur mentalvårdstjänsterna är ordnade i din hemkommun.
Om du är orolig för en närstående person och tror att han eller hon kan vara i behov av hjälp, kan du rådfråga till exempel hälsovårdaren eller läkaren vid hälsocentralen.
linkkiSocial- och hälsovårdsministeriet:
Mentalvårdstjänsterfinska _ svenska _ engelska _ ryska
Privata mentalvårdstjänster
Du kan också boka tid hos en psykiater eller en psykolog vid en privat läkarstation.
Där får man ibland fortare en tid, men besöket kostar avsevärt mer för kunden.
FPA (Kela) ersätter en del av kostnaderna för besök hos privatläkare om du omfattas av den finländska sjukförsäkringen.
Fråga mer hos FPA.
FPA:s ersättning kan ibland dras av direkt på det belopp som du betalar vid kassan.
Ta med ett intyg över att du omfattas av den finländska sjukförsäkringen.
Du kan också söka ersättning från FPA även i efterhand.
Läs mer om vem som omfattas av den finländska sjukförsäkringen på InfoFinlands sida Den sociala tryggheten i Finland.
Sjukvårdsersättningarfinska _ svenska _ engelska
Privat psykoterapitjänst på Internetfinska _ svenska _ engelska _ ryska _ franska _ spanska _ turkiska _ kinesiska _ tyska _ portugisiska _ norska
_ holländska _ japanska _ italienska
_ danska
Privat läkarstationfinska _ svenska _ engelska
Privat läkarstationfinska _ svenska _ engelska
När hjälpbehovet är brådskande
Om du känner att du behöver hjälp omedelbart kan du kontakta den närmaste jourhavande hälsovårdscentralen eller sjukhusjouren.
Brådskande psykiatrisk sjukvård ges på jourenheter vid psykiatriska sjukhus.
Om din närstående utgör en fara för sig själv eller för andra och inte går med på att träffa en läkare kan du ringa hälstocentralen eller sjukhuset.
Om det behövs hjälp snabbt ska du berätta det vid samtalet.
Nämn också om du är rädd för att din närstående kommer att skada sig själv.
Om din närstående är i mycket dåligt skick och behöver akut psykiatrisk sjukhusvård kan han eller hon intas för vård mot sin vilja.
För detta behövs läkarens remiss för tvångsvård (pakkohoitolähete).
Om någon är i omedelbar livsfara kan du ringa nödnumret 112.
Ring inte nödnumret om situationen inte är akut.
Hjälp telefonledes
Föreningen för mental hälsa i Finland (Suomen Mielenterveysseura) har en kristelefon som ger samtalshjälp för människor i en krissituation.
Du kan även ringa kristelefonen om du är orolig för en närstående person.
Du kan ringa
på finska till numret 01019 5202 må-fre kl. 9–7, på veckoslut och helger kl. 15–7
på engelska och arabiska till numret 040 195 8202 mån., tis., tors. och fre. kl. 11–15 och ons. kl. 18–22.
linkkiFöreningen för mental hälsa i Finland:
Riksomfattande kristelefonfinska _ svenska _ engelska
Barn och unga
Om ditt barn är i en psykiskt påfrestande situation kan du kontakta familjerådgivningen (perheneuvola) i din hemkommun.
På familjerådgivningen kartläggs barnets situation så att barnet får den hjälp som det behöver.
Du kan också boka tid hos barnrådgivningens (lastenneuvola) psykolog eller en läkare på din egen hälsostation.
Om barnet är i skolåldern kan du kontakta skolpsykologen eller skolläkaren.
Mer information om hjälp för barn i problematiska situationer får du på InfoFinlands sida Var hittar jag hjälp när barn eller unga har problem?
Om du är ung kan du berätta om det som bekymrar dig till exempel för skolhälsovårdaren, skolpsykologen eller skolkuratorn.
Du kan också kontakta din egen hälsostation.
Läkaren kan vid behov skriva en remiss till ungdomspsykiatriska polikliniken (nuorisopsykiatrian poliklinikka).
Mer information om hjälp för unga i problematiska situationer får du på InfoFinlands sida Var hittar jag hjälp när barn eller unga har problem?
linkkiMannerheims barnskyddsförbund:
Nätstöd för ungdomar, Nuortennettifinska
linkkiMannerheims Barnskyddsförbund rf:
Stöd för föräldrarfinska
Studerande
I hälsovårdstjänsterna vid läroanstalter ordnas också mentalvårdstjänster för studerande.
Företagshälsovårdens tjänster
Om du har en anställning kan du tala med företagshälsovårdens läkare om sådant som rör den mentala hälsan.
Du kan även ha möjlighet att träffa en psykolog vid företagshälsovården.
Traumatiska upplevelser
Människor som blivit utsatta för traumatiska situationer löper risk att insjukna i posttraumatiskt stressyndrom (traumaperäinen stressihäiriö).
Upplevelser som kan orsaka ett trauma är exempelvis:
förföljelse och diskriminering
fängelse och tortyr
misshandel och våldtäkt
att bevittna våldsamma situationer
krigserfarenheter.
Vid posttraumatiskt stressyndrom väcker olika situationer minnesbilderna från den traumatiska situationen, vilket orsakar kraftig ångest.
I en sådan situation är det viktigt att man skaffar sig hjälp.
Posttraumatiskt stressyndrom påverkar inte bara den som insjuknat utan även dennes närstående.
De flesta som har insjuknat i posttraumatiskt stressyndrom återhämtar sig med rätt behandling.
Rehabiliteringscentret för tortyroffer (Kidutettujen kuntoutuskeskus) hjälper de flyktingar och asylsökande som har blivit utsatta för tortyr i sitt hemland.
Du kan kontakta centret vardagar kl. 8.30–13.30 Telefonnumret är (09) 7750 4584.
Rehabiliteringscentret för tortyrofferfinska _ engelska
Information om posttraumatiskt stressyndromfinska _ engelska _ ryska _ franska _ somaliska _ turkiska _ persiska _ arabiska _ kurdiska _ albanska _ vietnamesiska _ burmesiska _ bosniska _ serbiska _ swahili
Information på olika språk om mental hälsa på webben
På webbsidorna för Föreningen för mental hälsa i Finland hittar du information om
svåra livssituationer
problem med den mentala hälsan
kriser
om hur du kan söka hjälp
om hur du kan återhämta dig.
Informationen finns på finska, engelska, kurdiska, ryska och somaliska.
linkkiFöreningen för Mental Hälsa i Finland:
Information om mental hälsafinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Nödnumret (hätänumero) i Finland är 112.
Du får ringa nödnumret endast i brådskande nödfall där liv, hälsa, egendom eller miljö är i fara.
I nödsituationer får du vård även om du inte har en hemkommun i Finland.
Vårdavgifter kan komma att debiteras av dig i efterhand.
Ring 112 till exempel i följande situationer:
du har råkat ut för en bilolycka (auto-onnettomuus) eller är vittne till en olycka
någon är i livsfara (hengenvaara)
du upptäcker en brand (tulipalo)
du upptäcker ett inbrott (murto)
Ring inte nödnumret om ärendet inte är brådskande.
Du ska inte ringa nödnumret vid vanliga sjukdomsfall.
Du ska inte heller ringa nödnumret om du vill fråga polisen (poliisi) till exempel om ett tillståndsärende.
Onödiga samtal kan orsaka att hjälpen kommer för sent i verkliga nödsituationer.
Du kan straffas för att ha missbrukat nödnumret.
Samtalet besvaras av en utbildad nödcentraloperatör.
Han eller hon ställer dig frågor och bedömer hjälpbehovet.
Därefter larmar han eller hon hjälp.
Operatören berättar också vad du ska göra.
Operatören kopplar inte samtalet vidare, så besvara frågorna noga.
Du kan tala finska eller svenska när du ringer nödnumret.
Du kan också fråga om nödcentraloperatören förstår engelska, med det är inte säkert.
Vid behov bistås nödcentralen av en tolktjänst.
Du kan ringa nödnumret gratis från alla telefoner.
Du behöver inget riktnummer.
Du kan ringa nödnumret utan riktnummer även om du har ett utländskt mobilabonnemang.
Nödnumret 112 fungerar i alla EU-länder.
Om du har installerat den kostnadsfria mobilappen 112 Suomi i din telefon, behöver du inte nödvändigtvis kunna berätta var du befinner dig.
Nödcentraloperatören ser var du är, när du ringer ett nödsamtal via appen.
Du kan ladda ned appen i applikationsbutiken.
När du ringer nödnumret 112:
uppge ditt namn
berätta vad som har hänt
ange exakt adress och kommun
svara på nödcentraloperatörens frågor
följ instruktionerna
avsluta inte samtalet förrän du får lov.
Mer information om nödnumret får du på Nödcentralsverkets (Hätäkeskuslaitos) webbplats.
Om du behöver information om tillståndsärenden som sköts av polisen, fordonsföreskrifter eller hur undersökningen i ett brott som skett tidigare framskrider ska du ringa polisens egna nummer under tjänstetid.
Om du misstänker att någon har förgiftats kan du fråga råd vid Giftinformationscentralen (Myrkytystietokeskus).
Giftinformationscentralens telefontjänst är öppen 24 timmar om dygnet.
Telefonnumret är (09) 471 977.
linkkiNödcentralsverket:
Nödsituationfinska _ svenska _ engelska
linkkiNödcentralsverket:
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
linkkiRöda Kors:
Första hjälpen-anvisningar för olika situationerfinska _ svenska _ engelska
Första hjälpen-anvisningar vid förgiftningfinska _ svenska _ engelska
Graviditet kan också förhindras med spermiedödande medel, till exempel p-skum (emätinvaahto) eller slidpiller (emätinpuikko), men de är inte särskilt effektiva.
Kondom skyddar mot de flesta könssjukdomarna.
Kondomer kan köpas i butiker, bensinstationer, kiosker och apotek. De kan köpas utan recept.
Vissa spermiedödande medel kan köpas receptfritt på apotek.
För hormonella preventivmedel behöver du ett läkarrecept som du får till exempel vid hälsostationen (terveysasema) eller av en privat gynekolog.
Du kan också boka tid vid preventivrådgivningen (ehkäisyneuvonta) antingen ensam eller tillsammans med din partner.
För akutpreventivmedel behövs vanligen inget recept.
P-piller, minipiller, p-plåster och p-ring kan köpas på apoteket med ett läkarrecept.
Kopparspiralen eller hormonspiralen sätts in av en läkare.
Spiralen passar bäst för kvinnor som har fött barn.
Även unga kan boka tid hos läkaren och få ett recept för preventivmedel.
De behöver inte ha föräldrarnas tillstånd.
Du kan diskutera preventivmetoder med skolans hälsovårdare och i vissa kommuner kan skolans hälsovårdare ge dig ett startpaket.
Om du har problem med preventivmedlen eller om du har glömt att använda preventivmedel kan du köpa akut-p-piller (jälkiehkäisypilleri) på apoteket.
Det ska tas så fort efter samlaget som möjligt, senast inom 72 timmar.
Alla som har fyllt 15 år kan köpa ett akut-p-piller receptfritt.
Barn under 15 år behöver ett läkarrecept.
Graviditetspreventionfinska
Även om du inte har värk eller andra symptom, lönar det sig att regelbundet låta undersöka dina tänder.
Tandsjukdomar behandlas på bästa sätt då de upptäcks innan symptom uppkommer.
Mun- och tandhälsan påverkar hälsan i hela din kropps hälsa.
Om du har hemkommun (kotikunta) i Finland kan du utnyttja de offentliga tandvårdstjänsterna.
Mer information finns på InfoFinlands sida Hemkommun i Finland .
I nödfall får du behandling även om du inte har en hemkommun i eller uppehållstillstånd till Finland.
Det är möjligt att vårdutgifterna tas ut av dig i efterskott.
Hälso- och sjukvårdstjänster lämnas på finska och svenska i Finland.
Ofta klarar du dig också på engelska.
Om du inte kan något av dessa språk, ska du fråga om det är möjligt att anlita tolk när du bokar tid till tandvården.
Läs mer på InfoFinlands sida Behöver du en tolk?
När du har bokat tid till tandvård, är det viktigt att komma i tid.
Om du har bokat tid, men inte kan komma, är det väldigt viktigt att du avbokar besöket i tid, vanligen senast dagen innan.
Om du inte kommer och inte har avbokat tiden, måste du betala en ersättning.
linkkiSocial- och hälsovårdsministeriet:
Munhälsafinska _ svenska
Den offentliga tandvården
Kommunerna tillhandahåller tandvård vid hälsostationer (terveysasema) och tandkliniker (hammashoitola).
När du vill boka tid i tandvården ska du ringa tandvårdens tidsbeställning i din hemkommun.
Vårdbehovet bedöms ofta på telefon.
Om du inte behöver brådskande vård kan du tvingas vänta flera månader på en tid.
Intagning för vård måste ske inom sex månader.
När du vill boka tid för akut tandvård ska du ringa tandvårdens jourtidsbeställning (päivystysajanvaraus) i din hemkommun.
Kraftig värk, svullnad eller en olycka är orsaker för att få akut vård.
Brådskande fall sköts så fort som möjligt.
Kvällar och veckoslut är jourmottagningen centraliserad till större vårdenheter.
Om du bor på en liten ort kan du bli tvungen att åka till jourmottagningen i en närliggande stad.
Om du behöver mer krävande vårdåtgärder, som till exempel tandkirurgi, ska du först boka tid hos en tandläkare.
Vid behov skriver tandläkaren en remiss till specialtandvården.
Privata tandvårdstjänster
Du kan också boka tid hos en privat tandläkare.
Privat tandvård är dyrare än offentlig tandvård.
Om du omfattas av den sociala tryggheten i Finland ersätter FPA en del av kostnaderna.
FPA ersätter dock inte till exempel sådan vård som enbart har en kosmetisk effekt.
Mer information hittar du på FPA:s webbplats.
På InfoFinlands sida den sociala tryggheten i Finland får du mer information om vem som omfattas den finländska sjukförsäkringen.
Privat tandvård och ersättningarfinska _ svenska _ engelska
Jämför läkarpriserfinska _ engelska
Barn
Barn får en inbjudan till tandvård med ett brev som skickas hem.
Tandundersökningar ordnas regelbundet för barn.
Offentlig tandvård är gratis för barn under 18 år.
Om du har avlagt examen i något annat land kan du behöva beslut om erkännande av examen för att kunna arbeta eller studera i Finland.
I de flesta situationerna bedömer arbetsgivaren, läroanstalten eller högskolan vilken behörighet och kompetens din utländska examen ger.
Du behöver Utbildningsstyrelsens eller någon annan myndighets beslut om erkännande av examen om du vill arbeta inom ett reglerat yrke eller en uppgift som kräver högskoleexamen på viss nivå.
linkkiUtbildningsstyrelsen:
Erkännande av en examenfinska _ svenska _ engelska
linkkiUtbildningsstyrelsen :
Broschyr om erkännande av examen(pdf, 102,14 kt)finska _ svenska _ engelska _ ryska _ estniska _ franska _ spanska _ kinesiska _ persiska _ arabiska _ portugisiska
linkkiUtbildningsstyrelsen :
Diagram över erkännande av examen(pdf, 410,87 kt)finska _ svenska _ engelska
linkkiUtbildningsstyrelsen:
Servicepriserfinska _ svenska _ engelska
Om du vill fortsätta dina studier i Finland
Högskolor och läroanstalter beslutar om antagning av studerande.
De beslutar också huruvida dina utländska studier och din övriga kompetens kan godkännas som en del av den examen du avlägger i Finland.
Om du har avlagt högskolestudier utomlands och vill fortsätta dina studier i Finland kan du få information och handledning vid högskolornas tjänster för studerande och SIMHE-tjänsterna.
Högskolor som erbjuder SIMHE-tjänsterfinska _ svenska _ engelska
Uppgifter som inte kräver en viss utbildning
Enligt Finlands lag kräver inte alla uppgifter en viss utbildning eller examen på en viss nivå.
Till exempel bedömer arbetsgivare i privatsektorn oftast själv huruvida en utländsk examen ger tillräckliga kvalifikationer för uppgiften.
Jämställande av nivån på en högskolexamen
För uppgifter inom den offentliga sektorn (kommun eller stat) krävs ofta examen på en viss nivå, till exempel en högre högskoleexamen.
Om du har avlagt en högskoleexamen utomlands kan du ansöka om beslut om jämställande av nivån på en högskolexamen vid Utbildningsstyrelsen.
Beslutet är avgiftsbelagt.
När din examensnivå har jämställts med en finländsk högskoleexamen, kan du söka till uppgifter som kräver den nivå på högskoleexamen som du har.
linkkiUtbildningsstyrelsen:
Jämställande av nivån på en högskolexamenfinska _ svenska _ engelska
Reglerade yrken
I Finland är vissa yrken reglerade.
Det betyder att det stadgas i lag vilken utbildning som krävs för dessa yrken.
Sådana uppgifter är till exempel fysioterapeut, läkare, tandläkare, provisor, sjukskötare, advokat, revisor, klasslärare och sotare.
Branschspecifika myndigheter beslutar om rätten att utöva ett reglerat yrke eller använda en yrkesbeteckning.
Till exempel inom social- och hälsovårdsbranschen fattas beslutet av Valvira, och inom undervisningssektorn av Utbildningsstyrelsen.
Beslutet är avgiftsbelagt.
På Utbildningsstyrelsens webbplats hittar du en förteckning över reglerade yrken och de myndigheter som fattar beslut.
linkkiUtbildningsstyrelsen:
Reglerade yrken och ansvariga myndigheterfinska _ svenska _ engelska
Information om erkännande av examen för yrken inom hälsovårdenfinska _ svenska _ engelska
Reglerade yrken och examen från ett annat EU-land
Om
du är medborgare i ett EU-land, EES-land eller Schweiz och du har
förvärvat kvalifikationer för ett yrke som är reglerat i Finland i ett EU-land, EES-land eller Schweiz,
kan du ansöka om erkännande av yrkeskvalifikationer för detta yrke hos den branschspecifika myndigheten.
Om din utbildning skiljer sig mycket från den utbildning som krävs i Finland måste du eventuellt avlägga en anpassningsperiod eller ett lämplighetsprov.
linkkiUtbildningsstyrelsen:
Erkännande av yrkeskvalifikationer som förvärvats i ett EU-landfinska _ svenska _ engelska
linkkiEuropeiska kommissionen:
Information om reglerade yrken i EU-ländernaengelska
Utländsk yrkesexamen
Om du har avlagt en yrkesexamen utomlands kan du ansöka om ett utlåtande om det hos Utbildningsstyrelsen.
I utlåtandet beskrivs examensnivån och innehåll samt för vilka uppgifter examen ger kvalifikationer i det land där du har avlagt examen.
Utlåtandet ger dig dock inte kvalifikationer att utöva ett reglerat yrke i Finland.
linkkiUtbildningsstyrelsen:
Utlåtanden om utländska yrkesexamenfinska _ svenska _ engelska
Översättning av handlingar
Om originalspråket för ditt betyg inte är finska, svenska eller engelska behöver du vanligtvis en officiell översättning av handlingarna som görs av en auktoriserad översättare.
Vissa myndigheter godkänner även handlingar på andra europeiska språk.
Läs noga anvisningarna om ansökning från den branschspecifika myndigheten.
Om du känner att du behöver information eller hjälp i ärenden som rör den sexuella hälsan kan du kontakta din egen hälsostation (terveysasema).
Du kan fråga råd av hälsovårdaren (terveydenhoitaja) eller boka tid hos läkaren (lääkäri).
Till exempel för p-piller behöver du ett recept som endast kan skrivas av en läkare.
Du har rätt att utnyttja tjänsterna vid hälsostationen om du har hemkommun i Finland.
Ungas sexualitetfinska _ engelska
Vuxnas sexualitetfinska _ svenska _ engelska
Sexuell hälsa hos kvinnor
En del läkare inom den offentliga hälsovården gör gynekologiska undersökningar.
Du har rätt att utnyttja de offentliga hälsovårdstjänsterna om du har hemkommun i Finland.
Fråga mer vid din egen hälsostation.
Du kan be om att få tid hos en kvinnlig läkare om du vill.
Du kan också boka tid hos en privat gynekolog. Privatläkares tjänster är avsevärt dyrare för kunden.
I Finland ordnas screeningundersökningar (seulontatutkimus) för kvinnor där man försöker hitta bröstcancer och livmoderhalscancer i ett tidigt skede.
Bröstcancerundersökningen görs för kvinnor i åldern 50–69 år ungefär vartannat år och undersökningen för livmoderhalscancer för kvinnor i åldern 30–60 år med fem års mellanrum.
Om du har hemkommun i Finland.har du rätt att få dessa undersökningar gjorda.
linkkiSocial- och hälsovårdsministeriet:
Screeningsundersökningarfinska _ svenska _ engelska _ ryska
linkkiInstitutet för hälsa och välfärd:
Information om bröstcancerscreeningfinska _ svenska
Anvisning för identifiering av bröstcancer(pdf, 440kt)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ kinesiska _ thai _ rumänska _ samiska
Information om cancerscreeningfinska _ svenska _ engelska
Sexuell hälsa hos män
Om du har hemkommun i Finland kan du boka tid för en urologisk undersökning på din egen hälsostation.
Läkaren kan vid behov skriva en remiss till en specialist på urologiska polikliniken.
Preventivmedel säljs på apoteket.
Kondomer säljs också till exempel i mataffärer.
För hormonella preventivmedel behöver du ett läkarrecept, som du får till exempel från hälsostationen eller av en privat gynekolog.
Du kan också boka tid för preventivrådgivning (ehkäisyneuvonta).
På Väestöliittos webbplats hittar du information om olika preventivmedel.
Graviditetspreventionfinska
Hjälp med att få barn
Om en graviditet inte börjar inom ett år efter att man slutat använda preventivmedel kan saken undersökas.
Ofta kan man få hjälp med att få barn.
Du kan boka tid för en undersökning på din egen hälsostation (terveysasema), hos en gynekolog eller på en privat barnlöshetsklinik (lapsettomuusklinikka).
Det är bra att ni går till kliniken tillsammans.
I undersökningarna utreds orsaken till barnlösheten.
Könssjukdomar
Om du misstänker att du smittats med en könssjukdom kan du boka tid hos läkaren antingen på hälsostationen eller på en privat läkarstation.
I stora städer kan könssjukdomar vårdas på polikliniker för könssjukdomar (sukupuolitautien poliklinikka).
Fråga mer vid din egen hälsostation.
Klamydia och gonorré behandlas med antibiotika.
Virussjukdomar, såsom herpes och kondylom, kan inte botas med läkemedel, men symtomen kan lindras.
Framskridandet av en HIV-infektion kan bromsas med läkemedel.
Det är bra att inleda medicineringen så tidigt som möjligt.
Kondom skyddar mot de flesta könssjukdomarna.
linkkiHivpoint:
Broschyren Information om sexuellt överförda sjukdomar(pdf, 1500kt)finska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
linkkiHivpoint:
Info om HIVfinska _ engelska _ ryska
linkkiHivpoint:
Broschyren Ett gott liv med HIVfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ thai
linkkiHivpoint:
Broschyren HIV i familjen(pdf, 881 kb)finska _ engelska _ ryska
Omskärelse av pojkar
Omskärelse (ympärileikkaus) är alltid ett oåterkalleligt ingrepp.
Om det görs av icke-medicinska orsaker, inkräktar man på en pojkes fysiska integritet.
Omskärelse får endast göras av en legitimerad läkare.
För omskärelse behövs ett skriftligt samtycke av pojkens vårdnadshavare.
Om barnet har två vårdnadshavare, behövs varderas samtycke, i annat fall kan ingreppet inte göras.
Pojken har rätt att vägra att gå med på operationen.
Omskärelse får inte göras utan smärtlindring som ges av läkare, och det ska göras i en steril miljö.
Icke-medicinsk omskärelse omfattas inte av den offentligt finansierade hälsovården, och kan därför inte göras på en offentlig hälsostation, och man måste själv betala det.
Fråga mer om omskärelse på rådgivningen, av läkaren på hälsostationen, skolhälsovårdaren eller skolläkaren.
Omskärelse av flickor
Omskärelse (ympärileikkaus) av flickor är ett brott i Finland. Man kan få ett flera års fängelsestraff för det.
Det är också ett brott att föra en flicka till ett annat land, för att låta henne genomgå omskärelse där.
Om du har omskurits innan du kom till Finland och planerar graviditet, kan du låta operera dig för att få slidmynningen öppnad (avausleikkaus).
Det är lättast om operationen görs innan graviditeten har börjat, men den kan också göras i mitten av graviditeten.
Öppningsoperationen gör förlossningen och undersökningarna under graviditeten lättare.
Operationen görs på sjukhus och återhämtningen tar vanligtvis 1–2 dagar.
Omskärelse av kvinnor och flickorfinska _ engelska _ somaliska _ arabiska
Om ditt barn har hemkommun (kotikunta) i Finland har han eller hon rätt att utnyttja de offentliga hälsovårdstjänsterna.
Läs mer på InfoFinlands sida Hemkommun i Finland.
Om du omfattas av den finländska sjukförsäkringen (sairausvakuutus) kan du teckna en försäkring för ditt barn som täcker en del av kostnaderna för privata hälsovårdstjänster.
När ett barn insjuknar
Om barnet har feber eller annars är sjukt ska det inte tas till dagvården.
Om barnet har hosta eller snuva, men annars mår bra, kan barnet vara i dagvården.
Om ett barn under 10 år insjuknar akut kan barnets mamma eller pappa stanna hemma för att ta hand om barnet.
Vårdledigheten kan vara högst fyra dagar.
I kollektivavtalet bestäms om man får lön för denna tid eller inte.
Om ett barn blir sjukt under skoldagen vårdas han eller hon i skolan.
Vid behov förs barnet till stadens hälsostation.
Om ett sjukt barn behöver läkarhjälp eller uppsöka hälsovårdare ska du kontakta hälsostationen (terveysasema) eller en privat läkarstation i din hemkommun.
Hälsostationerna har öppet från måndag till fredag, vanligen kl. 8–16.
Det är bäst att ringa hälsostationen genast på morgonen när tidsbeställningen öppnar.
Vid tidsbeställningen bedöms vilken slags vård barnet behöver.
Kvällstid och under veckoslut har hälsostationerna stängt.
Då vårdas akuta sjukfall och olycksfall på jourmottagningen (päivystys).
Om barnets sjukdom inte kräver omedelbar vård ska du vänta tills din hälsostation har öppet igen.
Jourmottagningen för barn och unga finns ofta i en separat enhet.
Du kan också boka tid till läkare på en privat hälsostation.
De har ofta öppet också på kvällarna och ibland får man fortare en tid där.
Privata hälsovårdstjänster är dock avsevärt dyrare för kunden än offentliga.
Om du misstänker att ett barn har förgiftats kan du fråga råd vid Giftinformationscentralen (Myrkytystietokeskus).
Giftinformationscentralens telefontjänst är öppen 24 timmar om dygnet. Telefonnumret är (09) 471 977.
Om ett barn är i livsfara eller har hamnat i en olycka ska du ringa nödnumret (hätänumero) 112.
Ambulanser är endast avsedda för allvarliga och brådskande situationer.
Ring inte nödnumret vid vanliga sjukdomsfall.
Om barnet insjuknarfinska _ svenska _ engelska
Sjukvårdsersättningarfinska _ svenska _ engelska
Småbarns hälsa
Hälsotillståndet hos barn under skolåldern följs i barnrådgivningen (lastenneuvola).
Barnrådgivningen följer och stöder den fysiska, psykiska och sociala tillväxten och utvecklingen av barn under skolåldern.
På barnrådgivningen besöker barnen en läkare eller en hälsovårdare.
Familjen till ett barn som är under ett år gammalt kallas till barnrådgivningen minst nio gånger.
Efter det första året kallas man till barnrådgivningen ännu minst sex gånger.
Hälsovårdaren följer barnets utveckling, vaccinerar barnet och ger information om rätt kost.
Hälsovården besöket barnet också hemma direkt efter födseln.
Rådgivningsbyråns tjänster i den egna kommunen är kostnadsfria.
Du kan utnyttja barnrådgivningsbyråns tjänster i din egen kommun om du har hemkommun i Finland.
Mer information finns på InfoFinlands sida Hemkommun i Finland.
Du ska ha med dig kortet på varje besök till rådgivningen.
Hälsovårdaren antecknar uppgifter om barnets hälsa och vaccinationer på kortet.
linkkiSocial- och hälsovårdsministeriet:
Information om rådgivningsbyråernas tjänsterfinska _ svenska _ engelska _ ryska
Skolbarns hälsa
Varje skola har en läkare och en hälsovårdare.
Hälsovårdaren undersöker barnen i skolan.
Hälsovårdaren är på plats i skolan vissa dagar i veckan.
Eleverna kan själva besöka hälsovårdarens mottagning om de har problem.
Vid ett olycksfall i skolan får barnet första hjälpen.
Mer information om skolhälsovården finns på social- och hälsovårdsministeriets (Sosiaali- ja terveysministeriö) webbplats.
linkkiSocial- och hälsovårdsministeriet:
Skolhälsovårdfinska _ svenska
Vaccinationer
I Finland kan barnen vaccineras (rokotus) mot många smittsamma sjukdomar.
Vaccinationerna ges på barnrådgivningen (lastenneuvola) och inom skolhälsovården.
De vaccinationer som ingår i vaccinationsprogrammet är avgiftsfria för familjen.
Vaccinationerna är frivilliga.
De flesta barn i Finland får de vaccinationer som ingår i vaccinationsprogrammet.
Berätta för hälsovårdaren vilka vaccinationer ditt barn har fått innan ni kom till Finland.
Om du vill att ditt barn ska få en vaccination som inte ingår i vaccinationsprogrammet ska du beställa tid till en läkare.
Läkaren kan skriva ett recept på vaccinationen och hälsovårdaren kan vaccinera ditt barn.
Du köper själv vaccinationen på apoteket.
linkkiInstitutet för hälsa och välfärd:
Vaccinationsprogrammet i Finlandfinska _ svenska
Långvarig sjukdom och vård av ett handikappat barn
Om du under en lång tid tar hand om ett sjukt eller handikappat barn under 16 år kan du söka specialvårdpenning (erityishoitoraha) från FPA.
Från FPA kan du även få bidrag för rehabilitering (kuntoutus) av barnet.
Ett barn med en svår sjukdom eller ett handikapp kan även få FPA:s handikappbidrag för barn under 16 år (alle 16-vuotiaan vammaistuki).
FPA:s bidrag är avsedda för personer som omfattas av Den sociala tryggheten i Finland.
Du får mer information om att leva i Finland med ett handikappat barn på InfoFinlands sida Ett handikappat barn.
Specialvårdspenning för barn under 16 årfinska _ svenska _ engelska
Handikappbidrag för barnfinska _ svenska _ engelska
Omskärelse av pojkar
Omskärelse (ympärileikkaus) är alltid ett oåterkalleligt ingrepp.
Om det görs av icke-medicinska orsaker, inkräktar man på en pojkes fysiska integritet.
Omskärelse får endast göras av en legitimerad läkare.
För omskärelse behövs ett skriftligt samtycke av pojkens vårdnadshavare.
Om barnet har två vårdnadshavare, behövs varderas samtycke, i annat fall kan ingreppet inte göras.
Pojken har rätt att vägra att gå med på operationen.
Omskärelse får inte göras utan smärtlindring som ges av läkare, och det ska göras i en steril miljö.
Icke-medicinsk omskärelse omfattas inte av den offentligt finansierade hälsovården, och kan därför inte göras på en offentlig hälsostation, och man måste själv betala det.
Fråga mer om omskärelse på rådgivningen, av läkaren på hälsostationen, skolhälsovårdaren eller skolläkaren.
Omskärelse av flickor
Omskärelse (ympärileikkaus) av flickor är ett brott i Finland. Man kan få ett flera års fängelsestraff för det.
Det är också ett brott att föra en flicka till ett annat land, för att låta henne genomgå omskärelse där.
Omskärelse av kvinnor och flickorfinska _ engelska _ somaliska _ arabiska
Du kan studera i Finland som utbytesstudent eller avlägga hela examen här.
Om du vill hitta arbete i Finland är det viktigt att du studerar finska eller svenska.
I Finland är det ofta svårt att hitta arbete om man inte kan finska eller svenska.
Utbytesstudenter
Du kan komma till Finland som utbytesstudent.
Du kan avlägga utbytesstudier via olika program.
Utbytesstudenter kan få studieplats till exempel via Erasmus, Nordplus, FIRST och Fulbright.
Du kan också studera som utbytesstudent på egen hand.
Om du vill komma till Finland som utbytesstudent ska du ta kontakt med enheten för internationella ärenden eller till exempel studiebyrån i din egen läroanstalt.
Komihåglista för nya studerande
Säkerställ att du har följande när du kommer till Finland för att studera:
uppehållstillstånd
försäkring
pengar
studieplats
bostad
Ansökan för examensstuderande
Du kan söka till en yrkeshögskola eller ett universitet i den gemensamma ansökan till högskolor.
Läs mer på InfoFinlands sida Ansökan till utbildning.
Du hittar mer information om yrkeshögskolor på InfoFinlands sida Yrkeshögskolor.
Läs mer om högskolor på InfoFinlands sida Universitet.
Du kan också avlägga fortsatta studier vid universitet eller yrkeshögskola i Finland.
Läs mer om fortsatta studier på InfoFinlands sidor Universitet och Yrkeshögskolor.
Uppehållstillstånd
När du kommer till Finland för att studera beror behovet av uppehållstillstånd på ditt medborgarskap.
Läs mer på InfoFinlands sida Studerande.
Finansiering av studierna
Utländska studerande får vanligen inget studiestöd.
För att få ett uppehållstillstånd för studerande, ska du kunna visa att din ekonomiska situation ger dig möjlighet att leva i Finland.
Penningunderstöd och stipendier
Utländska studerande kan ansöka om olika penningunderstöd för finländska högskolor.
Alla finländska högskolor har ett eget stipendiesystem för de studerande som kommer från länder utanför EU/EES-området och som har godkänts för att avlägga en kandidat- eller magisterexamen på engelska.
Möjligheten till ett stipendium kan till exempel bero på hur framgångsrik du varit i dina studier.
Stipendiet kan täcka hela läsårsavgiften eller en del av den.
Vissa stipendier kan även täcka andra kostnader.
Ibland krävs att du lyckas tillräckligt bra med dina studier för att du ska få ett stipendium.
Du kan vanligtvis ansöka om ett stipendium samtidigt som du ansöker om en studieplats.
Det finns också särskilda Erasmus Mundus-magisterprogram som har ett eget stipendiesystem.
Utbildningsstyrelsen har stipendieprogram för forskarstuderande som kommer till Finland för att avlägga doktorsexamen.
Studerande från USA kan ansöka om ett Fulbright-stipendium.
Läs mer om stipendier och penningunderstöd på webbplatsen Studyinfinland.fi.
Boende, arbete och försäkring
Det kan vara svårt att hitta en bostad eftersom efterfrågan på bostäder är större än utbudet speciellt i större städer.
Sök en bostad i god tid innan du flyttar till Finland
Du kan hyra en bostad på den öppna marknaden.
Du kan också söka bostad via föreningen Suomen Opiskelija-asunto (Suomen Opiskelija-asunto) (SOA).
Det är dyrt att bo i Finland.
Studentbostäderna är oftast billigare än bostäderna på den öppna marknaden.
Om du arbetar vid sidan av studierna är din arbetstid begränsad.
Vanligen kan du arbeta högst 25 timmar i veckan.
Detta beror dock på vilket land du kommer ifrån.
Läs mer på InfoFinlands sida Studerande.
Du kan också göra ditt slutarbete i något företag eller göra en arbetspraktik.
I dessa har arbetstiden inte begränsats.
Se till att du har försäkringar.
Hur omfattande försäkring du behöver beror på vilket land du kommer ifrån och hur länge dina studier pågår.
Det är mycket viktigt att din försäkring är i kraft hela den tid som du vistas i Finland.
Läs mer på InfoFinlands sida Studerande.
Studier i Finland
Om du inte är medborgare i ett EU-land eller EES-land och inte heller familjemedlem till en medborgare i ett sådant land och du kommer till Finland för att studera i augusti 2017 eller senare, måste du betala terminsavgift för studierna.
Avgiften gäller lägre och högre högskolestudier på engelska.
I Finland kan du studera på finska, svenska och ibland även på engelska.
Högskolorna har vissa utbildningsprogram där undervisningen ges på engelska.
Merparten av studierna är dock på finska eller på svenska.
I Finland finns många aktiva studentorganisationer.
De ordnar verksamhet även för utländska studerande.
I studentorganisationerna lär du dig känna nya människor.
Om du vill hitta en arbetsplats i Finland ska du studera finska eller svenska.
Även om du klarar dig i många dagliga situationer på engelska kräver de flesta arbetsgivare att du kan finska eller svenska.
Läs mer på InfoFinlands sida Finska och svenska språket.
Om inte hinner studera finska vid din egen läroanstalt, finns det kurser i finska vid många andra läroanstalter.
Du kan även studera språket på Internet.
Läs mer på InfoFinlands sida Finska och svenska språket.
Det är också viktigt att du bekantar dig med finländare och arbetslivet i Finland redan under studietiden.
På så sätt hittar du lättare vänner och ett arbete.
Till exempel arbetspraktik (työharjoittelu), hobbyer och organisationer är bra sätt att lära känna det finländska samhället.
Information för utländska studerandeengelska
Information om utbytesprogrammetengelska
När ska jag söka hjälp?
Vem som helst kan behöva hjälp om livssituationen är påfrestande.
Livet kan vara svårt till exempel när man flyttar från ett land till ett annat, har problem på arbetsplatsen, förlorar sin arbetsplats, har problem i familjen, går igenom skilsmässa, förlorar en anhörig, blir sjuk eller när livet förändras på andra sätt.
Också positiva saker, t.ex. att man får barn, kan ändra livet så mycket att man behöver stöd i den nya situationen.
Ibland kan man må dåligt först i efterhand när man redan har lagt den svåra erfarenheten bakom sig och situationen har lugnat ner sig.
Det lönar sig att söka hjälp, om du har något av följande symptom:
sömnlöshet
ingen aptit
vardagen känns tung
du orkar inte arbeta eller träffa människor
fysiska symptom, utan att medicinska orsaker hittas för dessa
ökad alkohol- eller droganvändning
Det är inte ovanligt att söka hjälp för att få stöd med den mentala hälsan.
I Finland lider 20 % av befolkningen av depression i något skede av livet.
Depression(pdf, 110,37 kt)finska _ engelska _ ryska _ franska _ somaliska _ turkiska _ persiska _ arabiska _ kurdiska _ albanska _ vietnamesiska _ burmesiska _ bosniska _ serbiska _ swahili
Var får jag hjälp?
Ofta hjälper det redan att tala om dessa saker med familjen eller vänner. Ibland behövs det även annan hjälp.
Det kan hjälpa att tala med en hälsovårdare (terveydenhoitaja), läkare (lääkäri) eller en psykoterapeut (psykoterapeutti).
Tillsammans kan ni fundera på vilken sorts stöd som skulle passa just dig.
Ofta hjälper terapi, medicinering eller en kombination av båda.
Ibland behövs sjukhusvård.
Sjukhusvården räcker vanligen några veckor.
Målsättningen är att patienten kan återvända hem så fort som möjligt.
Därefter fortsätter vården som öppenvård.r.
Om du har hemkommun i Finland ska du först kontakta din egen hälsostation (terveysasema).
Hälsostationerna har vanligen öppet från måndag till fredag, ungefär kl. 8–16.
Ring hälsostationen genast på morgonen för att boka tid.
Om du behöver hjälp genast ska du tala om det när du ringer.
Läkaren skriver vid behov en remiss till psykiatriska polikliniken (psykiatrian poliklinikka) eller en annan vårdenhet för psykisk hälsa.
Du kan inte gå till polikliniken utan en läkarremiss.
Med läkaren eller psykologen kan du samtala konfidentiellt.
De har tystnadsplikt. De berättar inte om dina saker för andra myndigheter.
Om någon annan hälsovårdsenhet behöver dina uppgifter, ombeds du ge ditt medgivande för överlåtelse av dessa.
På din egen hälsostation får du mer information om hur mentalvårdstjänsterna är ordnade i din hemkommun.
Om du är orolig för en närstående person och tror att han eller hon kan vara i behov av hjälp, kan du rådfråga till exempel hälsovårdaren eller läkaren vid hälsocentralen.
linkkiSocial- och hälsovårdsministeriet:
Mentalvårdstjänsterfinska _ svenska _ engelska _ ryska
Privata mentalvårdstjänster
Du kan också boka tid hos en psykiater eller en psykolog vid en privat läkarstation.
Där får man ibland fortare en tid, men besöket kostar avsevärt mer för kunden.
FPA (Kela) ersätter en del av kostnaderna för besök hos privatläkare om du omfattas av den finländska sjukförsäkringen.
Fråga mer hos FPA.
FPA:s ersättning kan ibland dras av direkt på det belopp som du betalar vid kassan.
Ta med ett intyg över att du omfattas av den finländska sjukförsäkringen.
Du kan också söka ersättning från FPA även i efterhand.
Läs mer om vem som omfattas av den finländska sjukförsäkringen på InfoFinlands sida Den sociala tryggheten i Finland.
Sjukvårdsersättningarfinska _ svenska _ engelska
Privat psykoterapitjänst på Internetfinska _ svenska _ engelska _ ryska _ franska _ spanska _ turkiska _ kinesiska _ tyska _ portugisiska _ norska
_ holländska _ japanska _ italienska
_ danska
Privat läkarstationfinska _ svenska _ engelska
Privat läkarstationfinska _ svenska _ engelska
När hjälpbehovet är brådskande
Om du känner att du behöver hjälp omedelbart kan du kontakta den närmaste jourhavande hälsovårdscentralen eller sjukhusjouren.
Brådskande psykiatrisk sjukvård ges på jourenheter vid psykiatriska sjukhus.
Om din närstående utgör en fara för sig själv eller för andra och inte går med på att träffa en läkare kan du ringa hälstocentralen eller sjukhuset.
Om det behövs hjälp snabbt ska du berätta det vid samtalet.
Nämn också om du är rädd för att din närstående kommer att skada sig själv.
Om din närstående är i mycket dåligt skick och behöver akut psykiatrisk sjukhusvård kan han eller hon intas för vård mot sin vilja.
För detta behövs läkarens remiss för tvångsvård (pakkohoitolähete).
Om någon är i omedelbar livsfara kan du ringa nödnumret 112.
Ring inte nödnumret om situationen inte är akut.
Hjälp telefonledes
Föreningen för mental hälsa i Finland (Suomen Mielenterveysseura) har en kristelefon som ger samtalshjälp för människor i en krissituation.
Du kan även ringa kristelefonen om du är orolig för en närstående person.
Du kan ringa
på finska till numret 01019 5202 må-fre kl. 9–7, på veckoslut och helger kl. 15–7
på engelska och arabiska till numret 040 195 8202 mån., tis., tors. och fre. kl. 11–15 och ons. kl. 18–22.
linkkiFöreningen för mental hälsa i Finland:
Riksomfattande kristelefonfinska _ svenska _ engelska
Barn och unga
Om ditt barn är i en psykiskt påfrestande situation kan du kontakta familjerådgivningen (perheneuvola) i din hemkommun.
På familjerådgivningen kartläggs barnets situation så att barnet får den hjälp som det behöver.
Du kan också boka tid hos barnrådgivningens (lastenneuvola) psykolog eller en läkare på din egen hälsostation.
Om barnet är i skolåldern kan du kontakta skolpsykologen eller skolläkaren.
Mer information om hjälp för barn i problematiska situationer får du på InfoFinlands sida Var hittar jag hjälp när barn eller unga har problem?
Om du är ung kan du berätta om det som bekymrar dig till exempel för skolhälsovårdaren, skolpsykologen eller skolkuratorn.
Du kan också kontakta din egen hälsostation.
Läkaren kan vid behov skriva en remiss till ungdomspsykiatriska polikliniken (nuorisopsykiatrian poliklinikka).
Mer information om hjälp för unga i problematiska situationer får du på InfoFinlands sida Var hittar jag hjälp när barn eller unga har problem?
linkkiMannerheims barnskyddsförbund:
Nätstöd för ungdomar, Nuortennettifinska
linkkiMannerheims Barnskyddsförbund rf:
Stöd för föräldrarfinska
Studerande
I hälsovårdstjänsterna vid läroanstalter ordnas också mentalvårdstjänster för studerande.
Företagshälsovårdens tjänster
Om du har en anställning kan du tala med företagshälsovårdens läkare om sådant som rör den mentala hälsan.
Du kan även ha möjlighet att träffa en psykolog vid företagshälsovården.
Traumatiska upplevelser
Människor som blivit utsatta för traumatiska situationer löper risk att insjukna i posttraumatiskt stressyndrom (traumaperäinen stressihäiriö).
Upplevelser som kan orsaka ett trauma är exempelvis:
förföljelse och diskriminering
fängelse och tortyr
misshandel och våldtäkt
att bevittna våldsamma situationer
krigserfarenheter.
Vid posttraumatiskt stressyndrom väcker olika situationer minnesbilderna från den traumatiska situationen, vilket orsakar kraftig ångest.
I en sådan situation är det viktigt att man skaffar sig hjälp.
Posttraumatiskt stressyndrom påverkar inte bara den som insjuknat utan även dennes närstående.
De flesta som har insjuknat i posttraumatiskt stressyndrom återhämtar sig med rätt behandling.
Rehabiliteringscentret för tortyroffer (Kidutettujen kuntoutuskeskus) hjälper de flyktingar och asylsökande som har blivit utsatta för tortyr i sitt hemland.
Du kan kontakta centret vardagar kl. 8.30–13.30 Telefonnumret är (09) 7750 4584.
Rehabiliteringscentret för tortyrofferfinska _ engelska
Information om posttraumatiskt stressyndromfinska _ engelska _ ryska _ franska _ somaliska _ turkiska _ persiska _ arabiska _ kurdiska _ albanska _ vietnamesiska _ burmesiska _ bosniska _ serbiska _ swahili
Information på olika språk om mental hälsa på webben
På webbsidorna för Föreningen för mental hälsa i Finland hittar du information om
svåra livssituationer
problem med den mentala hälsan
kriser
om hur du kan söka hjälp
om hur du kan återhämta dig.
Informationen finns på finska, engelska, kurdiska, ryska och somaliska.
linkkiFöreningen för Mental Hälsa i Finland:
Information om mental hälsafinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Vilka hälsotjänster kan du använda?
Offentliga hälsovårdstjänster
Privata hälsovårdstjänster
Hälsovård för medborgare i de nordiska länderna
Hälsovård för EU-medborgare
Hälsovård för anställda och företagare
Hälsovård för studerande
Hälsovård för invandrare och asylsökande
Hälsovård för papperslösa
Information på webben
Vilka hälsotjänster kan du använda?
Du kan utnyttja de offentliga hälsovårdstjänsterna i Finland om du har hemkommun (kotikunta) i Finland.
Rätten till hemkommun beror på följande:
från vilket land du kommer till Finland
varför du kommer till Finland (t.ex. arbete, studier)
om du ska bo stadigvarande i Finland eller vistas här tillfälligt
om din vistelse i Finland är tillfällig, beroende på hur länge vistelsen varar.
Om du inte är säker på om du har hemkommun i Finland kan du ta reda på din situation vid magistraten (maistraatti).
Mer information finns på InfoFinlands sida Hemkommun i Finland.
Om du arbetar i Finland, kan du ha rätt till den offentliga hälso- och sjukvården även om du inte har en hemkommun i Finland.
Om du inte har en hemkommun i Finland ska du be FPA utreda din rätt till den offentliga hälso- och sjukvården.
I nödfall får du vård inom den offentliga hälso- och sjukvården fastän du inte har en hemkommun i Finland eller rätt till vård på grund av arbete.
Du kan krävas på vårdkostnaderna i efterhand.
Om du inte har rätt till de offentliga hälsovårdstjänsterna, kan du boka tid på en privat läkarstation.
Privata hälsovårdstjänster är avsevärt dyrare för kunden än de offentliga.
Hälsovårdstjänster ges i Finland på finska och svenska.
Ofta klarar man sig även på engelska.
När du bokar tid till hälsovårdstjänster kan du fråga om möjligheten att använda en tolk (tulkki) om du inte behärskar dessa språk.
Läs mer på InfoFinlands sida Behöver du en tolk?
När du har bokat tid för ett läkarbesök ska du vara punktligt på plats.
Om du har bokat tid för ett läkarbesök men får förhinder är det mycket viktigt att du avbokar besöket i god tid, helst dagen innan.
Om du inte kommer och inte heller har avbokat din tidsbeställning måste du betala en avgift.
Hälsa och rehabiliteringfinska _ svenska _ ryska _ estniska
Sjukvård för utlänningar i Finlandfinska _ svenska _ engelska
Kontaktpunkt för gränsöverskridande hälso- och sjukvårdfinska _ svenska _ engelska
linkkiStödcentralen Hilma för funktionshindrade invandrare :
Handbok med ordlista i hälso- och sjukvård på finska(pdf, 341,02 kt)finska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska
Offentliga hälsovårdstjänster
När du blir sjuk ska du först kontakta din egen hälsostation (terveysasema). Där kan du boka tid hos en allmänläkare eller en hälsovårdare.
Mer information om hälsovårdstjänsterna i olika kommuner hittar du på InfoFinlands sida på de lokala informationssidorna eller på din egen kommuns sida.
Hälsostationens tjänster är relativt förmånliga för klienten eftersom de finansieras med skattemedel.
Hälsostationerna har vanligen öppet från måndag till fredag kl. 310 1671.
Det är klokt att ringa tidsbeställningen genast på morgonen när hälsostationen öppnar.
Om ditt besvär kräver brådskande vård får du en tid snabbt.
Om du inte behöver brådskande vård måste du vänta längre på att få en läkartid.
Vid tidsbeställningen får du veta hur snabbt du kommer att få vård.
Vid tidsbeställningen bedöms även om du behöver vård av läkare eller hälsovårdare.
I Finland kan hälsovårdare ge vård vid flera sjukdomar.
Vid behov kan hälsovårdaren ge remiss till läkare.
Om du har ett FPA-kort (Kela-kortti) ska du ta det med när du besöker hälsovårdsstationen.
Om du behöver en specialist, ska du först boka tid hos en allmänläkare.
Vid behov skriver hälsostationsläkaren en remiss till en specialist.
Specialister finns på vissa hälsostationer, på polikliniker och sjukhus.
Specialsjukvård ges på centralsjukhus och universitetssjukhus.
I Finland gör läkare inom de offentliga hälsovårdstjänsterna inga hembesök.
En del privata läkarstationer erbjuder denna tjänst. Ett hembesök av en privatläkare är dock dyrt.
Om din sjukdom är långvarig och du inte kan arbeta finns det mer information om FPA:s sjukpenning på InfoFinlands sida Stöd när du är sjuk.
Jour inom offentliga hälsovårdstjänster
Hälsostationerna har stängt kvällstid och under veckoslut.
Då vårdas akuta sjukfall på jourmottagningen (päivystys).
Jourmottagningen är avsedd för situationer där man behöver omedelbar vård.
Om din sjukdom inte kräver omedelbar vård ska du beställa tid på din egen hälsostation nästa gång den har öppet.
Jourmottagningen finns ofta i anslutning till sjukhus, i små städer också i en närliggande stad.
Jourmottagningen för barn och unga finns ofta separat.
Fråga mer vid din egen hälsostation under dess öppettider eller leta upp informationen på din hemkommuns webbplats.
Privata hälsovårdstjänster
Kontaktuppgifter till privata läkarstationer hittar du till exempel på internet.
Förmodligen får du en tid snabbare på en privat hälsostation än inom den offentliga hälsovården.
Privata hälsotjänster är avsevärt dyrare för klienten än de offentliga.
Olika läkarstationer erbjuder olika tjänster.
Privata hälsotjänster kan användas av alla, även personer som inte har en hemkommun i Finland.
Om du omfattas av den finländska sjukförsäkringen (sairausvakuutus) ersätter FPA en liten del av kostnaderna för privat sjukvård och tandvård.
Ibland kan också personer som inte omfattas av den finländska sjukförsäkringen ha rätt till ersättning från FPA. Fråga mer hos FPA.
FPA:s ersättning kan ibland dras av direkt på det belopp som du betalar vid kassan.
Du kan också söka ersättning från FPA i efterhand.
Läs mer om sjukförsäkringen i Finland på InfoFinlands sida Den sociala tryggheten i Finland.
Sjukvårdsersättningarfinska _ svenska _ engelska
Jämför läkarpriserfinska _ engelska
Privat läkarstationfinska _ svenska _ engelska
Privat läkarstationfinska _ svenska _ engelska
linkkiAava:
Privat läkarstationfinska _ svenska _ engelska
Hälsovård för medborgare i de nordiska länderna
Om du har en sjukförsäkring i ett annat nordiskt land har du rätt till nödvändig sjukvård i Finland.
Du får vård på samma villkor och till samma kostnad som finländarna.
Ta med dig ett officiellt identitetsbevis när du använder hälsovårdstjänsterna.
Hälsovård för EU-medborgare
Om du har en sjukförsäkring i ett annat EU-land, EES-land eller i Schweiz har du rätt till nödvändig sjukvård i Finland.
För att få vård måste du ha ett europeiskt sjukvårdskort.
Du ska skaffa dig det europeiska sjukvårdskortet i det land där du har din sjukförsäkring.
Det europeiska sjukvårdskortet ger dig rätt till vård om du blir sjuk eller råkar ut för en olycka.
Du får vård även vid en långvarig sjukdom.
Med kortet får du även vård i samband med graviditet och förlossning.
Du får vård till samma kostnad som personer som är stadigvarande bosatta i Finland.
Information om det europeiska sjukvårdskortetfinska _ svenska _ engelska
Hälsovård för anställda och företagare
Om du har kommit till Finland för att arbeta kan du ha rätt att använda de offentliga hälsovårdstjänsterna i Finland.
Detta beror på hurdant och hur långt arbetsavtal du har samt från vilket land du har kommit till Finland.
I Finland är arbetsgivare skyldiga att ordna förebyggande företagshälsovård för sina anställda.
Företagare kan ordna sin egen företagshälsovård om de vill.
Företagare måste alltså inte ordna företagshälsovård för sig.
Företagare måste ändå ordna företagshälsovård för sina anställda.
Företagshälsovården kan ordnas vid den lokala hälsovårdscentralen eller till exempel på en privat läkarcentral.
Mer information får du på InfoFinlands sida Företagshälsovården och på social- och hälsovårdsministeriets webbplats.
linkkiSocial- och hälsovårdsministeriet:
Företagshälsovårdfinska _ svenska _ engelska
Hälsovård för studerande
Om du kommer från ett land som inte är ett EU-land, ett EES-land eller Schweiz till Finland för att studera behöver du vanligtvis ha en täckande sjukförsäkring i ditt hemland för att få uppehållstillstånd i Finland.
Om dina studier beräknas pågå i minst två år får du vanligen en hemkommun i Finland och rätt till de kommunala hälsovårdstjänsterna.
I detta fall räcker det om din sjukförsäkring i första hand täcker läkemedelskostnaderna.
Om du inte är säker på om du har rätt till hemkommun i Finland kan du kontrollera detta vid magistraten.
Du får mer information om hemkommun på InfoFinlands sida Hemkommun i Finland.
Mer information om uppehållstillstånd för studerande och om den sjukförsäkring som krävs för att få uppehållstillstånd får du på Migrationsverkets (Maahanmuuttovirasto) webbplats.
I Finland omfattas högskolestuderande av studerandehälsovården.
Fråga mer vid din egen läroanstalt.
Mer information om studerandehälsovården får du på Studenternas hälsovårdsstiftelses (SHVS) (YTHS) och social- och hälsovårdsministeriets (Sosiaali- ja terveysministeriö) webbplatser.
Information om uppehållstillstånd för studierfinska _ svenska _ engelska
linkkiSHVS:
Hälsovård för högskolestuderandefinska _ svenska _ engelska
linkkiSocial- och hälsovårdsministeriet:
Studerandehälsovårdfinska _ svenska
Hälsovård för invandrare och asylsökande
Om du har kommit till Finland som kvotflykting har du hemkommun i Finland och rätt att utnyttja de offentliga hälsovårdstjänsterna.
Om du är asylsökande och din ansökan inte ännu har behandlats kan du inte registrera dig i magistraten som kommuninvånare och inte heller utnyttja kommunens hälsovårdstjänster.
Fråga mer vid din förläggning.
Om du har fått uppehållstillstånd på grund av behovet av skydd och får rätt till hemkommun i Finland, kan du utnyttja hälsovårdstjänsterna i din egen kommun.
Läs mer om rätten till hemkommun på InfoFinlands sida Hemkommun i Finland.
Hälsovård för papperslösa
Global Clinic är en klinik där du kan få hjälp eller råd av en läkare eller sjukskötare om du vistas i Finland utan uppehållstillstånd.
Global Clinic bedriver verksamhet i följande städer:
Åbo
Uleåborg
Joensuu
Tammerfors
Du kan ringa eller skicka e-post.
En sjukskötare eller läkare besvarar ditt samtal.
Du hittar kontaktinformation på Global Clinic:s hemsidor.
Global Clinic:s tjänster är avgiftsfria för kunderna.
Global Clinic anmäler inte sina kunder till polisen eller andra myndigheter.
Klinikens adress eller öppettider meddelas inte offentligt.
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Information på webben
linkkiTuberkuloosi.fi:
Information om tuberkulosfinska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Din situation avgör hur du kan finansiera dina studier i Finland.
På den här sidan berättar vi om FPA:s stöd till studerande samt om penningunderstöd och stipendier.
Studiestöd
Du kan få FPA:s studiestöd (opintotuki) om du
har det uppehållstillstånd (oleskelulupa) som krävs och
vistas i Finland av någon annan orsak än studier.
Om du flyttar till Finland för att studera kan du inte få studiestöd.
Till exempel utbytesstuderande får inte finskt studiestöd.
Studiestödet består av studiepenning och statsborgen för studielån.
Du kan få studiestöd om
Du studerar i gymnasiet
Du studerar vid en yrkesläroanstalt eller avlägger yrkesinriktade tilläggsstudier
Du studerar vid en högskola.
Du kan få studiepenning om du har fyllt 17 år.
Du måste studera på heltid.
Med heltidsstudier avses att studierna är din huvudsyssla.
Du kan arbeta vid sidan av studierna.
Lönen som du får för ditt arbete kan minska ditt studiestöd.
Du ansöker om studiepenning och statsgaranti för studielån vid FPA.
FPA betalar in studiepenningen på ditt konto månatligen.
På studiepenningens belopp inverkar många omständigheter.
På studiepenningens belopp inverkar bland annat stödmottagarens ålder, om hen bor i sitt eget hem eller hos en förälder, on hen är gift och om hen har minderåriga barn. Kontrollera storleken på din studiepenning på FPA:s webbplats eller vid en FPA-byrå.
Det är inte obligatoriskt att ta studielån.
Du kan högst ta ut ett visst maximibelopp.
Du väljer själv hur mycket studielån du vill ta.
Studielånet är ett lån som finska staten ger garanti för åt studeranden.
Du ansöker om lånet i banken när du har fått FPA:s beslut om statsgaranti.
Du måste betala tillbaka lånet när du har slutfört dina studier.
Du kan få studielån också när du fortbildar dig (täydennyskoulutus) som vuxen.
Dessutom kan du få vuxenutbildningsstöd (aikuiskoulutustuki).
I vissa fall kan du också få bostadstillägg, till exempel om du studerar på en avgiftsbelagd linje vid en folkhögskola och bor på läroanstaltens internat.
Läs mer på FPA:s webbplats.
På InfoFinlands sida Bostadsbidrag finns mer information om FPA:s allmänna bostadsbidrag.
Information om studiestödetfinska _ svenska _ engelska
Information om studiestödetryska _ estniska _ samiska
Information om att ansöka studiestödfinska _ svenska _ engelska
Studiestöd till utländska studerandefinska _ svenska _ engelska
Stöd för skolresor
Du kan få stöd för skolresor (koulumatkatuki) om du bor i Finland och studerar i gymnasiet eller vid en yrkesläroanstalt.
Din skolresa måste vara minst 10 kilometer lång och resekostnaderna måste överstiga 54 euro per månad.
Information om skolresestödetfinska _ svenska _ engelska
Måltidsstöd
Om du studerar vid en högskola får du också måltidsstöd (ateriatuki).
Du kan få måltidsstödet endast i läroanstalternas egna restauranger.
Detta innebär att studeranden betalar mindre för måltiderna än andra som besöker restaurangen.
Du behöver inte ansöka separat om måltidsstödet.
Du behöver bara visa upp ditt studentkort när du betalar för måltiden.
Du har inte rätt till måltidsstöd om du är i Finland endast på arbetspraktik (työharjoittelu) som ingår i en utländsk examen.
Information om måltidsstödetfinska _ svenska _ engelska
Penningunderstöd och stipendier
Utländska studerande kan ansöka om olika penningunderstöd för finländska högskolor.
Alla finländska högskolor har ett eget stipendiesystem för de studerande som kommer från länder utanför EU/EES-området och som har godkänts för att avlägga en kandidat- eller magisterexamen på engelska.
Möjligheten till ett stipendium kan till exempel bero på hur framgångsrik du varit i dina studier.
Stipendiet kan täcka hela läsårsavgiften eller en del av den.
Vissa stipendier kan även täcka andra kostnader.
Ibland krävs att du lyckas tillräckligt bra med dina studier för att du ska få ett stipendium.
Du kan vanligtvis ansöka om ett stipendium samtidigt som du ansöker om en studieplats.
Det finns också särskilda Erasmus Mundus-magisterprogram som har ett eget stipendiesystem.
Utbildningsstyrelsen har stipendieprogram för forskarstuderande som kommer till Finland för att avlägga doktorsexamen.
Studerande från USA kan ansöka om ett Fulbright-stipendium.
Läs mer om stipendier och penningunderstöd på webbplatsen Studyinfinland.fi.
Även om du inte har värk eller andra symptom, lönar det sig att regelbundet låta undersöka dina tänder.
Tandsjukdomar behandlas på bästa sätt då de upptäcks innan symptom uppkommer.
Mun- och tandhälsan påverkar hälsan i hela din kropps hälsa.
Om du har hemkommun (kotikunta) i Finland kan du utnyttja de offentliga tandvårdstjänsterna.
Mer information finns på InfoFinlands sida Hemkommun i Finland .
I nödfall får du behandling även om du inte har en hemkommun i eller uppehållstillstånd till Finland.
Det är möjligt att vårdutgifterna tas ut av dig i efterskott.
Hälso- och sjukvårdstjänster lämnas på finska och svenska i Finland.
Ofta klarar du dig också på engelska.
Om du inte kan något av dessa språk, ska du fråga om det är möjligt att anlita tolk när du bokar tid till tandvården.
Läs mer på InfoFinlands sida Behöver du en tolk?
När du har bokat tid till tandvård, är det viktigt att komma i tid.
Om du har bokat tid, men inte kan komma, är det väldigt viktigt att du avbokar besöket i tid, vanligen senast dagen innan.
Om du inte kommer och inte har avbokat tiden, måste du betala en ersättning.
linkkiSocial- och hälsovårdsministeriet:
Munhälsafinska _ svenska
Den offentliga tandvården
Kommunerna tillhandahåller tandvård vid hälsostationer (terveysasema) och tandkliniker (hammashoitola).
När du vill boka tid i tandvården ska du ringa tandvårdens tidsbeställning i din hemkommun.
Vårdbehovet bedöms ofta på telefon.
Om du inte behöver brådskande vård kan du tvingas vänta flera månader på en tid.
Intagning för vård måste ske inom sex månader.
När du vill boka tid för akut tandvård ska du ringa tandvårdens jourtidsbeställning (päivystysajanvaraus) i din hemkommun.
Kraftig värk, svullnad eller en olycka är orsaker för att få akut vård.
Brådskande fall sköts så fort som möjligt.
Kvällar och veckoslut är jourmottagningen centraliserad till större vårdenheter.
Om du bor på en liten ort kan du bli tvungen att åka till jourmottagningen i en närliggande stad.
Om du behöver mer krävande vårdåtgärder, som till exempel tandkirurgi, ska du först boka tid hos en tandläkare.
Vid behov skriver tandläkaren en remiss till specialtandvården.
Privata tandvårdstjänster
Du kan också boka tid hos en privat tandläkare.
Privat tandvård är dyrare än offentlig tandvård.
Om du omfattas av den sociala tryggheten i Finland ersätter FPA en del av kostnaderna.
FPA ersätter dock inte till exempel sådan vård som enbart har en kosmetisk effekt.
Mer information hittar du på FPA:s webbplats.
På InfoFinlands sida den sociala tryggheten i Finland får du mer information om vem som omfattas den finländska sjukförsäkringen.
Privat tandvård och ersättningarfinska _ svenska _ engelska
Jämför läkarpriserfinska _ engelska
Barn
Barn får en inbjudan till tandvård med ett brev som skickas hem.
Tandundersökningar ordnas regelbundet för barn.
Offentlig tandvård är gratis för barn under 18 år.
Nödnumret (hätänumero) i Finland är 112.
Du får ringa nödnumret endast i brådskande nödfall där liv, hälsa, egendom eller miljö är i fara.
I nödsituationer får du vård även om du inte har en hemkommun i Finland.
Vårdavgifter kan komma att debiteras av dig i efterhand.
Ring 112 till exempel i följande situationer:
du har råkat ut för en bilolycka (auto-onnettomuus) eller är vittne till en olycka
någon är i livsfara (hengenvaara)
du upptäcker en brand (tulipalo)
du upptäcker ett inbrott (murto)
Ring inte nödnumret om ärendet inte är brådskande.
Du ska inte ringa nödnumret vid vanliga sjukdomsfall.
Du ska inte heller ringa nödnumret om du vill fråga polisen (poliisi) till exempel om ett tillståndsärende.
Onödiga samtal kan orsaka att hjälpen kommer för sent i verkliga nödsituationer.
Du kan straffas för att ha missbrukat nödnumret.
Samtalet besvaras av en utbildad nödcentraloperatör.
Han eller hon ställer dig frågor och bedömer hjälpbehovet.
Därefter larmar han eller hon hjälp.
Operatören berättar också vad du ska göra.
Operatören kopplar inte samtalet vidare, så besvara frågorna noga.
Du kan tala finska eller svenska när du ringer nödnumret.
Du kan också fråga om nödcentraloperatören förstår engelska, med det är inte säkert.
Vid behov bistås nödcentralen av en tolktjänst.
Du kan ringa nödnumret gratis från alla telefoner.
Du behöver inget riktnummer.
Du kan ringa nödnumret utan riktnummer även om du har ett utländskt mobilabonnemang.
Nödnumret 112 fungerar i alla EU-länder.
Om du har installerat den kostnadsfria mobilappen 112 Suomi i din telefon, behöver du inte nödvändigtvis kunna berätta var du befinner dig.
Nödcentraloperatören ser var du är, när du ringer ett nödsamtal via appen.
Du kan ladda ned appen i applikationsbutiken.
När du ringer nödnumret 112:
uppge ditt namn
berätta vad som har hänt
ange exakt adress och kommun
svara på nödcentraloperatörens frågor
följ instruktionerna
avsluta inte samtalet förrän du får lov.
Mer information om nödnumret får du på Nödcentralsverkets (Hätäkeskuslaitos) webbplats.
Om du behöver information om tillståndsärenden som sköts av polisen, fordonsföreskrifter eller hur undersökningen i ett brott som skett tidigare framskrider ska du ringa polisens egna nummer under tjänstetid.
Om du misstänker att någon har förgiftats kan du fråga råd vid Giftinformationscentralen (Myrkytystietokeskus).
Giftinformationscentralens telefontjänst är öppen 24 timmar om dygnet.
Telefonnumret är (09) 471 977.
linkkiNödcentralsverket:
Nödsituationfinska _ svenska _ engelska
linkkiNödcentralsverket:
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
linkkiRöda Kors:
Första hjälpen-anvisningar för olika situationerfinska _ svenska _ engelska
Första hjälpen-anvisningar vid förgiftningfinska _ svenska _ engelska
Studierna är inte alltid inriktade på att skaffa ett yrke.
Du kan också ha studier som hobby.
Du kan studera vid flera olika läroanstalter: öppna universitetet (avoin yliopisto) eller öppna yrkeshögskolan (avoin ammattikorkeakoulu), sommaruniversitetet (kesäyliopisto), senioruniversitetet (ikäihmisten yliopisto), medborgarinstitut (kansalaisopisto), arbetarinstitut (työväenopisto) och folkhögskolor (kansanopisto).
Studierna är vanligen avgiftsbelagda.
Många av dessa läroanstalter tillhandahåller undervisning i finska och svenska för invandrare.
Läs mer på InfoFinlands sida Finska och svenska språket.
Du kan även studera flera andra språk, såsom engelska eller franska.
Vid folkhögskolor kan du även avlägga yrkesexamen.
Öppna universitetet och öppna yrkeshögskolan
Öppna universitetet (avoin yliopisto) och öppna yrkeshögskolan (avoin ammattikorkeakoulu) ordnar universitets- och yrkeshögskolekurser.
Vem som helst kan studera vid de öppna högskolorna.
Du kan studera vid öppna högskolor fastän du inte har någon examen.
Du kan studera vid öppna högskolor
om du vill studera som hobby
om du vill bli antagen för studier i ett visst ämne vid en högskola
när du vill utöka din yrkeskunnighet och dina kunskaper
Till de öppna högskolorna ordnas inga inträdesprov.
Du kan anmäla dig till vårens kurser i början av året och till höstens kurser i slutet av sommaren.
Anmäl dig direkt till kurserna.
Du kan välja enskilda kurser eller större studiehelheter.
Vid öppna högskolor är studierna flexibla.
Du kan delta i kurser under dagtid, på kvällar eller på veckoslut.
Du kan också studera på internet.
Studierna vid öppna högskolor är inte heltidsstudier.
Du kan avlägga studier vid öppna högskolan fastän du får arbetslöshetsersättning (työttömyyskorvaus).
Du har nytta av studierna vid öppna högskolan när du studerar vidare.
Om du blir antagen till yrkeshögskolan behöver du inte avlägga de kurser som du redan har avlagt vid öppna yrkeshögskolan.
Om du har studerat vid öppna universitetet och söker till universitetet ansöker du via separat ansökan (erillinen haku).
Information om öppna yrkeshögskolanfinska _ svenska
Information om öppna universitetetfinska _ svenska
Sommaruniversitetet
Kurserna vid sommaruniversitetet (kesäyliopisto) påminner mycket om kurserna vid öppna universitetet.
Man kan studera vid sommaruniversitetet även under andra tider än på sommaren.
Utöver universitetskurser ordnar sommaruniversiteten också annan undervisning, till exempel:
Yrkesinriktad fortbildning (täydennyskoulutus)
Arbetskraftsutbildning (työvoimakoulutus)
Abiturientkurser (abikurssi) för gymnasieelever som förbereder sig för studentskrivningarna
finskakurser för invandrare
Fråga närmare uppgifter om undervisningen vid närmaste sommaruniversitet.
Info om sommaruniversitetfinska _ svenska
Information om sommaruniversitetetfinska _ svenska _ engelska
Senioruniversitetet
Senioruniversitetet (ikäihmisten yliopisto) är avsett för dem som har fyllt 60 år.
Studietillfällena är dock öppna för alla.
Undervisningen vid senioruniversitetet är en del av öppna universitetets verksamhet.
Senioruniversitetet ordnar föreläsningsserier, kurser och studieresor.
Fråga mer om senioruniversitetet i kansliet för närmaste öppna universitet.
Medborgarinstitut och arbetarinstitut
I Finland finns många medborgarinstitut (kansalaisopisto) och arbetarinstitut (työväenopisto).
Vid dem kan du studera bland annat språk, handarbete, idrott, bildkonst och matlagning.
Medborgarinstituten och arbetarinstituten erbjuder hobbystudier.
Vid dem kan man inte avlägga yrkesinriktade studier.
Medborgarinstituten och arbetarinstituten ordnar finskakurser för invandrare.
Fråga närmare uppgifter om kurserna vid närmaste medborgarinstitut eller arbetarinstitut.
Ansökningspraxis varierar.
Vanligen ansöker man till vårens undervisning i början av året och till höstens undervisning på sensommaren.
Fråga om ansökningstiderna vid medborgarinstitutets eller arbetarinstitutets studiebyrå.
Info om medborgarinstituten och arbetarinstitutenfinska _ svenska
Medborgarinstitut i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Folkhögskolor
Folkhögskolorna (kansanopisto) erbjuder både hobbystudier och yrkesinriktad utbildning.
Folkhögskolan kan drivas av en organisation eller också kan de vara självständiga institut.
Vid folkhögskolan kan du utbilda dig till ett yrke.
Vid folkhögskolan kan man till exempel avlägga djurskötarexamen eller massörexamen.
Folkhögskolorna ordnar mycket undervisning för invandrare.
Vid folkhögskolan kan du studera finska eller delta i förberedande utbildning.
Folkhögskolorna ordnar vanligen två olika slags undervisning, kortkurser (lyhytkurssi) och långa utbildningslinjer (pitkä opintolinja).
Kortkurserna är öppna för alla och till dem behöver du inte söka.
Det räcker med att du anmäler dig.
De långa utbildningslinjerna är ofta yrkesinriktade studier.
De pågår vanligen från ett halvår till ett år.
Till de långa utbildningslinjerna måste man söka separat.
Folkhögskolornas ansökningspraxis och ansökningstider varierar.
Fråga mer om antagningen vid folkhögskolans studiebyrå.
Info om folkhögskolorfinska _ svenska
linkkiFinlands folkhögskolförening:
Information om folkhögskolorfinska
linkkiFinlands folkhögskolförening:
Kurser vid folkhögskolor för invandrarefinska
linkkiDövas folkhögskola:
Utbildning för döva invandrarefinska _ svenska _ engelska
På den här sidan finns information om tjänsterna i Rovaniemi.
Du hittar allmän information om arbete och entreprenörskap i Finland på InfoFinlands sida Arbete.
Lapplands arbets- och näringsbyrå
Lapplands arbets- och näringsbyrå
Invandrare får hjälp med jobbsökningen vid Lapplands arbets- och näringsbyrå (TE-byrån).
Kontaktuppgifter:
Valtakatu 16
Öppettiderna för Lapplands TE-byrå
mån kl. 9–16 utan tidsbeställning
tis–fre kl. 9–16, besök hos handläggarna endast med tidsbeställning
Lapplands TE-byrå betjänar kunderna per telefon måndagar, onsdagar, och torsdagar kl. 8–16.15 samt tisdagar och fredagar kl. 9–16.15 på numret 0295 039 501
E-post kan du skicka till adressen: kirjaamo.lappi(at)te-toimisto.fi
Läs mer:
linkkiArbetsministeriet:
Lediga tjänsterfinska
Ainonkatu 1, vån. 2
tfn 040 0377 595
öppettider:
mån–fre kl. 8.00–16.00 (för personligt möte måste du boka tid)
Företagsrådgivare
tfn 0400 187 250
Läs mer:
linkkiFöretags- och näringslivsutveckling i Rovaniemi:
På den här sidan finns information om tjänsterna i Rovaniemi.
Du hittar allmän information om arbete och entreprenörskap i Finland på InfoFinlands sida Arbete.
Lapplands arbets- och näringsbyrå
Lapplands arbets- och näringsbyrå
Invandrare får hjälp med jobbsökningen vid Lapplands arbets- och näringsbyrå (TE-byrån).
Kontaktuppgifter:
Valtakatu 16
Öppettiderna för Lapplands TE-byrå
mån kl. 9–16 utan tidsbeställning
tis–fre kl. 9–16, besök hos handläggarna endast med tidsbeställning
Lapplands TE-byrå betjänar kunderna per telefon måndagar, onsdagar, och torsdagar kl. 8–16.15 samt tisdagar och fredagar kl. 9–16.15 på numret 0295 039 501
E-post kan du skicka till adressen: kirjaamo.lappi(at)te-toimisto.fi
Läs mer:
linkkiArbetsministeriet:
Lediga tjänsterfinska
Ainonkatu 1, vån. 2
tfn 040 0377 595
öppettider:
mån–fre kl. 8.00–16.00 (för personligt möte måste du boka tid)
Företagsrådgivare
tfn 0400 187 250
Läs mer:
linkkiFöretags- och näringslivsutveckling i Rovaniemi:
På den här sidan finns information om tjänsterna i Rovaniemi.
Du hittar allmän information om arbete och entreprenörskap i Finland på InfoFinlands sida Arbete.
Lapplands arbets- och näringsbyrå
Lapplands arbets- och näringsbyrå
Invandrare får hjälp med jobbsökningen vid Lapplands arbets- och näringsbyrå (TE-byrån).
Kontaktuppgifter:
Lapplands arbets- och näringsbyrå
Valtakatu 16
Öppettiderna för Lapplands TE-byrå
mån kl. 9–16 utan tidsbeställning
tis–fre kl. 9–16, besök hos handläggarna endast med tidsbeställning
Lapplands TE-byrå betjänar kunderna per telefon måndagar, onsdagar, och torsdagar kl. 8–16.15 samt tisdagar och fredagar kl. 9–16.15 på numret 0295 039 501
Läs mer:
linkkiArbetsministeriet:
Lediga tjänsterfinska
Ainonkatu 1, vån.
tfn 040 0377 595 öppettider:
mån–fre kl. 8.00–16.00 (för personligt möte måste du boka tid)
tfn 0400 187 250
Läs mer:
linkkiFöretags- och näringslivsutveckling i Rovaniemi:
Om du har hemkommun i Finland kan du utnyttja de offentliga hälsovårdstjänsterna.
När du blir sjuk ska du kontakta hälsostationen (terveysasema) på din ort.
Du får mer information på InfoFinlands sida under rubriken Hälsovårdstjänster i Finland.
Mer information om läkemedel får du på InfoFinlands sida under rubriken Läkemedel.
Information om tjänster som underlättar vardagen för äldre får du på InfoFinlands sida Äldre människor.
Om du vårdar en närstående i hemmet kan du läsa mer på InfoFinlands sida Äldre människor.
Minnet
Orsaken till detta är inte alltid en demenssjukdom. Ibland kan det dock finnas en bakomliggande sjukdom som kan behandlas.
Om du upptäcker att du själv eller en närstående får allt svårare att komma ihåg saker, kan du kontakta hälsostationen i ditt område och boka en tid hos läkaren.
Läkaren diskuterar minnesproblemen med patienten och eventuellt också med dennes närstående och gör ett enkelt minnestest.
Vid behov skriver läkaren en remiss till närmare undersökningar.
linkkiAlzheimer Centralförbundet:
Minnesstörningar och demensfinska _ svenska _ engelska
Man kan insjukna i typ 2-diabetes (diabetes) i vilken ålder som helst men ofta insjuknar man i pensionsåldern.
Symtom på diabetes kan vara trötthet speciellt efter att man ätit, törst, ökat urineringsbehov, depression, retlighet, viktnedgång, benvärk, försämrad syn och ökad infektionskänslighet.
Diabetes kan behandlas med insulin och rätt kost.
Om du misstänker diabetes ska du beställa tid till läkaren på din egen hälsostation eller på en privat läkarstation.
Mer information om diabetes finns på webbplatserna för Institutet för hälsa och välfärd (Terveyden ja hyvinvoinnin laitos) och Diabetesförbundet (Diabetesliitto).
linkkiInstitutet för hälsa och välfärd:
Diabetesfinska _ svenska _ engelska
linkkiDiabetesförbundet:
Fakta om diabetesfinska _ svenska
Synen och hörseln
Många människor får med åldern sämre syn och hörsel.
Låt ögonläkaren undersöka dina ögon regelbundet så att eventuella ögonsjukdomar upptäcks i ett tidigt skede.
Om du upptäcker att din hörsel blivit sämre, boka en tid för en hörselundersökning på hälsostationen i ditt område eller hos en privatläkare.
Efter en preliminär undersökning får du en remiss till fortsatta undersökningar om det behövs.
Läs mer om hjälpmedel för synskadade och hörselskadade på InfoFinlands sida Handikappade personer.
linkkiFinska Hörselförbundet rf:
Åldershörselfinska
Om du har avlagt examen i något annat land kan du behöva beslut om erkännande av examen för att kunna arbeta eller studera i Finland.
I de flesta situationerna bedömer arbetsgivaren, läroanstalten eller högskolan vilken behörighet och kompetens din utländska examen ger.
Du behöver Utbildningsstyrelsens eller någon annan myndighets beslut om erkännande av examen om du vill arbeta inom ett reglerat yrke eller en uppgift som kräver högskoleexamen på viss nivå.
linkkiUtbildningsstyrelsen:
Erkännande av en examenfinska _ svenska _ engelska
linkkiUtbildningsstyrelsen :
Broschyr om erkännande av examen(pdf, 102,14 kt)finska _ svenska _ engelska _ ryska _ estniska _ franska _ spanska _ kinesiska _ persiska _ arabiska
linkkiUtbildningsstyrelsen :
Diagram över erkännande av examen(pdf, 410,87 kt)finska _ svenska _ engelska _ ryska
linkkiUtbildningsstyrelsen:
Servicepriserfinska _ svenska _ engelska
Om du vill fortsätta dina studier i Finland
Högskolor och läroanstalter beslutar om antagning av studerande.
De beslutar också huruvida dina utländska studier och din övriga kompetens kan godkännas som en del av den examen du avlägger i Finland.
Om du har avlagt högskolestudier utomlands och vill fortsätta dina studier i Finland kan du få information och handledning vid högskolornas tjänster för studerande och SIMHE-tjänsterna.
linkkiUtbildningsstyrelsen:
Högskolor som erbjuder SIMHE-tjänsterfinska _ svenska _ engelska
Uppgifter som inte kräver en viss utbildning
Enligt Finlands lag kräver inte alla uppgifter en viss utbildning eller examen på en viss nivå.
Till exempel bedömer arbetsgivare i privatsektorn oftast själv huruvida en utländsk examen ger tillräckliga kvalifikationer för uppgiften.
Jämställande av nivån på en högskolexamen
För uppgifter inom den offentliga sektorn (kommun eller stat) krävs ofta examen på en viss nivå, till exempel en högre högskoleexamen.
Om du har avlagt en högskoleexamen utomlands kan du ansöka om beslut om jämställande av nivån på en högskolexamen vid Utbildningsstyrelsen.
Beslutet är avgiftsbelagt.
När din examensnivå har jämställts med en finländsk högskoleexamen, kan du söka till uppgifter som kräver den nivå på högskoleexamen som du har.
linkkiUtbildningsstyrelsen:
Jämställande av nivån på en högskolexamenfinska _ svenska _ engelska
Reglerade yrken
I Finland är vissa yrken reglerade.
Det betyder att det stadgas i lag vilken utbildning som krävs för dessa yrken.
Sådana uppgifter är till exempel fysioterapeut, läkare, tandläkare, provisor, sjukskötare, advokat, revisor, klasslärare och sotare.
Branschspecifika myndigheter beslutar om rätten att utöva ett reglerat yrke eller använda en yrkesbeteckning.
Till exempel inom social- och hälsovårdsbranschen fattas beslutet av Valvira, och inom undervisningssektorn av Utbildningsstyrelsen.
Beslutet är avgiftsbelagt.
På Utbildningsstyrelsens webbplats hittar du en förteckning över reglerade yrken och de myndigheter som fattar beslut.
linkkiUtbildningsstyrelsen:
Reglerade yrken och ansvariga myndigheterfinska _ svenska _ engelska
Information om erkännande av examen för yrken inom hälsovårdenfinska _ svenska _ engelska
Reglerade yrken och examen från ett annat EU-land
Om
du är medborgare i ett EU-land, EES-land eller Schweiz och du har
förvärvat kvalifikationer för ett yrke som är reglerat i Finland i ett EU-land, EES-land eller Schweiz,
kan du ansöka om erkännande av yrkeskvalifikationer för detta yrke hos den branschspecifika myndigheten.
Om din utbildning skiljer sig mycket från den utbildning som krävs i Finland måste du eventuellt avlägga en anpassningsperiod eller ett lämplighetsprov.
linkkiUtbildningsstyrelsen:
Erkännande av yrkeskvalifikationer som förvärvats i ett EU-landfinska _ svenska _ engelska
linkkiEuropeiska kommissionen:
Information om reglerade yrken i EU-ländernaengelska
Utländsk yrkesexamen
Om du har avlagt en yrkesexamen utomlands kan du ansöka om ett utlåtande om det hos Utbildningsstyrelsen.
I utlåtandet beskrivs examensnivån och innehåll samt för vilka uppgifter examen ger kvalifikationer i det land där du har avlagt examen.
Utlåtandet ger dig dock inte kvalifikationer att utöva ett reglerat yrke i Finland.
linkkiUtbildningsstyrelsen:
Utlåtanden om utländska yrkesexamenfinska _ svenska _ engelska
Översättning av handlingar
Om originalspråket för ditt betyg inte är finska, svenska eller engelska behöver du vanligtvis en officiell översättning av handlingarna som görs av en auktoriserad översättare.
Vissa myndigheter godkänner även handlingar på andra europeiska språk.
Läs noga anvisningarna om ansökning från den branschspecifika myndigheten.
Yrkesinriktad arbetskraftsutbildning hjälper dig att få arbete.
Du kan lära dig nya färdigheter eller till och med ett nytt yrke.
Utbildningen kan också handleda dig i jobbsökningen.
Yrkesinriktad arbetskraftsutbildning är kostnadsfri.
Arbets- och näringsbyrån (TE-toimisto) ordnar den yrkesinriktade arbetskraftsutbildningen.
Du får arbetslöshetsförmån under utbildningstiden.
För vem är yrkesinriktad arbetskraftsutbildning avsedd?
Du kan delta i yrkesinriktad arbetskraftsutbildning, om
du har fyllt 20 år
du är arbetslös eller kommer att bli arbetslös
du har rätt att använda arbets- och näringsbyråns tjänster.
Du har rätt att använda arbets- och näringsbyråns tjänster om du har fått kontinuerligt uppehållstillstånd (A) eller permanent uppehållstillstånd (P).
linkkiArbets- och näringsministeriet:
Yrkesinriktad arbetskraftsutbildningfinska _ svenska _ engelska
Info om arbetskraftsutbildningfinska _ svenska
Hur ansöker jag till yrkesinriktad arbetskraftsutbildning?
Du ansöker till yrkesinriktad arbetskraftsutbildning antingen i arbets- och näringsbyrån eller med en elektronisk blankett på internet.
I ansökningen ska du motivera varför du borde antas till utbildningen.
Överväg din motivering noga.
Motiveringen påverkar antagningen.
Arbets- och näringsbyrån väljer studerandena till den yrkesinriktade arbetskraftsutbildningen.
Vad kan jag studera i yrkesinriktad arbetskraftsutbildning?
Innehållet i yrkesinriktad arbetskraftsutbildning varierar mycket.
Nedan följer några exempel på yrkesinriktad arbetskraftsutbildning:
Du kan lära dig ett nytt yrke eller en ny examensdel.
Du kan studera finska eller svenska.
Du kan få handledning i jobbsökningen.
Du kan få fortbildning eller påbyggnadsutbildning i din egen bransch.
Du kan få handledning i företagande eller företagarutbildning.
Hurdan är den yrkesinriktade arbetskraftsutbildningen?
Arbets- och näringsbyrån köper den yrkesinriktade arbetskraftsutbildningen av olika läroanstalter och företag.
Du studerar alltså inte vid arbets- och näringsbyrån utan vid den läroanstalt som ordnar kursen.
Arbets- och näringsbyrån genomför utbildningar även tillsammans med arbetsgivare.
Vissa läroanstalter ordnar yrkesinriktad arbetskraftsutbildning särskilt för invandrare.
Utbildningen kan vara till exempel studier i finska eller yrkesutbildning.
På vissa kurser kan du skaffa dig behörighet att utöva ditt yrke i Finland.
Till exempel sjukskötare måste avlägga ytterligare studier för att få arbeta som sjukskötare i Finland.
Läs mer på InfoFinlands sida Utländska examina i Finland.
Ekonomiskt stöd under den yrkesinriktade arbetskraftsutbildningen
Under den yrkesinriktade arbetskraftsutbildningen får du samma förmån som när du är arbetslös.
Om du har avtalat om yrkesinriktad arbetskraftsutbildning i din sysselsättningsplan, kan du få förhöjd arbetslöshetsförmån.
Det betyder att du får lite mer pengar i din arbetslöshetsförmån.
Beslut om utbetalning av förhöjningsdelen fattas av den som betalar arbetslöshetsförmånen, alltså arbetslöshetskassan eller FPA.
Du kan även få kostnadsersättning för resekostnader för de dagar som du deltar i utbildningen.
Om den som betalar din arbetslöshetsförmån inte betalar ut kostnadsersättning, kan arbets- och näringsbyrån i vissa fall betala den.
FPA:s kostnadsersättningfinska _ svenska _ engelska
Frivillig utbildning med arbetslöshetsförmån
Du kan även få arbetslöshetsförmån under andra studier om arbets- och näringsbyrån bedömer att du behöver utbildningen.
Arbets- och näringsbyrån skaffar inte utbildningen och väljer inte studeranden till utbildningen såsom i arbetskraftsutbildning.
Du ansöker om studieplats direkt vid läroanstalten.
Du måste avtala om utbildningen med arbets- och näringsbyrån innan du inleder utbildningen.
Du kan få arbetslöshetsförmån under studierna, om
du har anmält dig som arbetssökande vid arbets- och näringsbyrån och din jobbsökning är i kraft
du är minst 25 år gammal
arbets- och näringsbyrån bedömer att utbildningen främjar din yrkeskunnighet eller hjälper dig att få ett jobb
du har avtalat om utbildningen i din sysselsättningsplan med arbets- och näringsbyrån.
För vilka studier kan man få arbetslöshetsförmån?
Med arbetslöshetsförmånen understöds bara heltidsstudier.
Som heltidsstudier räknas följande:
högskoleexamen gymnasiestudier eller
studier, vars omfattning motsvarar heltidsstudier, till exempel fem studiepoäng i månaden eller 25 studietimmar i veckan.
Studierna ska leda till
yrkesinriktade grundexamen, yrkesexamen eller specialyrkesexamen
lägre eller högre högskoleexamen vid universitet eller högskola
avläggande av delar av ovan nämnda examina.
Studierna kan även vara tilläggsutbildning eller påbyggnadsutbildning alternativt studier vid universitet eller yrkeshögskola.
linkkiArbets- och näringsministeriet:
Frivilliga studier med stöd av arbetslöshetsförmånfinska _ svenska _ engelska
Om ditt barn har hemkommun (kotikunta) i Finland har han eller hon rätt att utnyttja de offentliga hälsovårdstjänsterna.
Läs mer på InfoFinlands sida Hemkommun i Finland.
Om du omfattas av den finländska sjukförsäkringen (sairausvakuutus) kan du teckna en försäkring för ditt barn som täcker en del av kostnaderna för privata hälsovårdstjänster.
När ett barn insjuknar
Om barnet har feber eller annars är sjukt ska det inte tas till dagvården.
Om barnet har hosta eller snuva, men annars mår bra, kan barnet vara i dagvården.
Om ett barn under 10 år insjuknar akut kan barnets mamma eller pappa stanna hemma för att ta hand om barnet.
Vårdledigheten kan vara högst fyra dagar.
I kollektivavtalet bestäms om man får lön för denna tid eller inte.
Om ett barn blir sjukt under skoldagen vårdas han eller hon i skolan.
Vid behov förs barnet till stadens hälsostation.
Om ett sjukt barn behöver läkarhjälp eller uppsöka hälsovårdare ska du kontakta hälsostationen (terveysasema) eller en privat läkarstation i din hemkommun.
Hälsostationerna har öppet från måndag till fredag, vanligen kl. 8–16.
Det är bäst att ringa hälsostationen genast på morgonen när tidsbeställningen öppnar.
Vid tidsbeställningen bedöms vilken slags vård barnet behöver.
Kvällstid och under veckoslut har hälsostationerna stängt.
Då vårdas akuta sjukfall och olycksfall på jourmottagningen (päivystys).
Om barnets sjukdom inte kräver omedelbar vård ska du vänta tills din hälsostation har öppet igen.
Jourmottagningen för barn och unga finns ofta i en separat enhet.
Du kan också boka tid till läkare på en privat hälsostation.
De har ofta öppet också på kvällarna och ibland får man fortare en tid där.
Privata hälsovårdstjänster är dock avsevärt dyrare för kunden än offentliga.
Om du misstänker att ett barn har förgiftats kan du fråga råd vid Giftinformationscentralen (Myrkytystietokeskus).
Giftinformationscentralens telefontjänst är öppen 24 timmar om dygnet. Telefonnumret är (09) 471 977.
Om ett barn är i livsfara eller har hamnat i en olycka ska du ringa nödnumret (hätänumero) 112.
Ambulanser är endast avsedda för allvarliga och brådskande situationer.
Ring inte nödnumret vid vanliga sjukdomsfall.
Om barnet insjuknarfinska _ svenska _ engelska
Sjukvårdsersättningarfinska _ svenska _ engelska
Småbarns hälsa
Hälsotillståndet hos barn under skolåldern följs i barnrådgivningen (lastenneuvola).
Barnrådgivningen följer och stöder den fysiska, psykiska och sociala tillväxten och utvecklingen av barn under skolåldern.
På barnrådgivningen besöker barnen en läkare eller en hälsovårdare.
Familjen till ett barn som är under ett år gammalt kallas till barnrådgivningen minst nio gånger.
Efter det första året kallas man till barnrådgivningen ännu minst sex gånger.
Hälsovårdaren följer barnets utveckling, vaccinerar barnet och ger information om rätt kost.
Hälsovården besöket barnet också hemma direkt efter födseln.
Rådgivningsbyråns tjänster i den egna kommunen är kostnadsfria.
Du kan utnyttja barnrådgivningsbyråns tjänster i din egen kommun om du har hemkommun i Finland.
Mer information finns på InfoFinlands sida Hemkommun i Finland.
Du ska ha med dig kortet på varje besök till rådgivningen.
Hälsovårdaren antecknar uppgifter om barnets hälsa och vaccinationer på kortet.
linkkiSocial- och hälsovårdsministeriet:
Information om rådgivningsbyråernas tjänsterfinska _ svenska _ engelska _ ryska
Skolbarns hälsa
Varje skola har en läkare och en hälsovårdare.
Hälsovårdaren undersöker barnen i skolan.
Hälsovårdaren är på plats i skolan vissa dagar i veckan.
Eleverna kan själva besöka hälsovårdarens mottagning om de har problem.
Vid ett olycksfall i skolan får barnet första hjälpen.
Mer information om skolhälsovården finns på social- och hälsovårdsministeriets (Sosiaali- ja terveysministeriö) webbplats.
linkkiSocial- och hälsovårdsministeriet:
Skolhälsovårdfinska _ svenska
Vaccinationer
I Finland kan barnen vaccineras (rokotus) mot många smittsamma sjukdomar.
Vaccinationerna ges på barnrådgivningen (lastenneuvola) och inom skolhälsovården.
De vaccinationer som ingår i vaccinationsprogrammet är avgiftsfria för familjen.
Vaccinationerna är frivilliga.
De flesta barn i Finland får de vaccinationer som ingår i vaccinationsprogrammet.
Berätta för hälsovårdaren vilka vaccinationer ditt barn har fått innan ni kom till Finland.
Om du vill att ditt barn ska få en vaccination som inte ingår i vaccinationsprogrammet ska du beställa tid till en läkare.
Läkaren kan skriva ett recept på vaccinationen och hälsovårdaren kan vaccinera ditt barn.
Du köper själv vaccinationen på apoteket.
linkkiInstitutet för hälsa och välfärd:
Vaccinationsprogrammet i Finlandfinska _ svenska
Långvarig sjukdom och vård av ett handikappat barn
Om du under en lång tid tar hand om ett sjukt eller handikappat barn under 16 år kan du söka specialvårdpenning (erityishoitoraha) från FPA.
Från FPA kan du även få bidrag för rehabilitering (kuntoutus) av barnet.
Ett barn med en svår sjukdom eller ett handikapp kan även få FPA:s handikappbidrag för barn under 16 år (alle 16-vuotiaan vammaistuki).
FPA:s bidrag är avsedda för personer som omfattas av Den sociala tryggheten i Finland.
Du får mer information om att leva i Finland med ett handikappat barn på InfoFinlands sida Ett handikappat barn.
Specialvårdspenning för barn under 16 årfinska _ svenska _ engelska
Handikappbidrag för barnfinska _ svenska _ engelska
Omskärelse av pojkar
Omskärelse (ympärileikkaus) är alltid ett oåterkalleligt ingrepp.
Om det görs av icke-medicinska orsaker, inkräktar man på en pojkes fysiska integritet.
Omskärelse får endast göras av en legitimerad läkare.
För omskärelse behövs ett skriftligt samtycke av pojkens vårdnadshavare.
Om barnet har två vårdnadshavare, behövs varderas samtycke, i annat fall kan ingreppet inte göras.
Pojken har rätt att vägra att gå med på operationen.
Omskärelse får inte göras utan smärtlindring som ges av läkare, och det ska göras i en steril miljö.
Icke-medicinsk omskärelse omfattas inte av den offentligt finansierade hälsovården, och kan därför inte göras på en offentlig hälsostation, och man måste själv betala det.
Fråga mer om omskärelse på rådgivningen, av läkaren på hälsostationen, skolhälsovårdaren eller skolläkaren.
Omskärelse av flickor
Omskärelse (ympärileikkaus) av flickor är ett brott i Finland. Man kan få ett flera års fängelsestraff för det.
Det är också ett brott att föra en flicka till ett annat land, för att låta henne genomgå omskärelse där.
Omskärelse av kvinnor och flickorfinska _ engelska _ somaliska _ arabiska
Du kan studera i Finland som utbytesstudent eller avlägga hela examen här.
Om du vill hitta arbete i Finland är det viktigt att du studerar finska eller svenska.
I Finland är det ofta svårt att hitta arbete om man inte kan finska eller svenska.
Utbytesstudenter
Du kan komma till Finland som utbytesstudent.
Du kan avlägga utbytesstudier via olika program.
Utbytesstudenter kan få studieplats till exempel via Erasmus, Nordplus, FIRST och Fulbright.
Du kan också studera som utbytesstudent på egen hand.
Om du vill komma till Finland som utbytesstudent ska du ta kontakt med enheten för internationella ärenden eller till exempel studiebyrån i din egen läroanstalt.
Komihåglista för nya studerande
Säkerställ att du har följande när du kommer till Finland för att studera:
uppehållstillstånd
försäkring
pengar
studieplats
bostad
Ansökan för examensstuderande
Du kan söka till en yrkeshögskola eller ett universitet i den gemensamma ansökan till högskolor.
Läs mer på InfoFinlands sida Ansökan till utbildning.
Du hittar mer information om yrkeshögskolor på InfoFinlands sida Yrkeshögskolor.
Läs mer om högskolor på InfoFinlands sida Universitet.
Du kan också avlägga fortsatta studier vid universitet eller yrkeshögskola i Finland.
Läs mer om fortsatta studier på InfoFinlands sidor Universitet och Yrkeshögskolor.
Uppehållstillstånd
När du kommer till Finland för att studera beror behovet av uppehållstillstånd på ditt medborgarskap.
Läs mer på InfoFinlands sida Studerande.
Finansiering av studierna
Utländska studerande får vanligen inget studiestöd.
För att få ett uppehållstillstånd för studerande, ska du kunna visa att din ekonomiska situation ger dig möjlighet att leva i Finland.
Penningunderstöd och stipendier
Utländska studerande kan ansöka om olika penningunderstöd för finländska högskolor.
Alla finländska högskolor har ett eget stipendiesystem för de studerande som kommer från länder utanför EU/EES-området och som har godkänts för att avlägga en kandidat- eller magisterexamen på engelska.
Möjligheten till ett stipendium kan till exempel bero på hur framgångsrik du varit i dina studier.
Stipendiet kan täcka hela läsårsavgiften eller en del av den.
Vissa stipendier kan även täcka andra kostnader.
Ibland krävs att du lyckas tillräckligt bra med dina studier för att du ska få ett stipendium.
Du kan vanligtvis ansöka om ett stipendium samtidigt som du ansöker om en studieplats.
Det finns också särskilda Erasmus Mundus-magisterprogram som har ett eget stipendiesystem.
Utbildningsstyrelsen har stipendieprogram för forskarstuderande som kommer till Finland för att avlägga doktorsexamen.
Studerande från USA kan ansöka om ett Fulbright-stipendium.
Läs mer om stipendier och penningunderstöd på webbplatsen Studyinfinland.fi.
Boende, arbete och försäkring
Det kan vara svårt att hitta en bostad eftersom efterfrågan på bostäder är större än utbudet speciellt i större städer.
Sök en bostad i god tid innan du flyttar till Finland
Du kan hyra en bostad på den öppna marknaden.
Du kan också söka bostad via föreningen Suomen Opiskelija-asunto (Suomen Opiskelija-asunto) (SOA).
Det är dyrt att bo i Finland.
Studentbostäderna är oftast billigare än bostäderna på den öppna marknaden.
Om du arbetar vid sidan av studierna är din arbetstid begränsad.
Vanligen kan du arbeta högst 25 timmar i veckan.
Detta beror dock på vilket land du kommer ifrån.
Läs mer på InfoFinlands sida Studerande.
Du kan också göra ditt slutarbete i något företag eller göra en arbetspraktik.
I dessa har arbetstiden inte begränsats.
Se till att du har försäkringar.
Hur omfattande försäkring du behöver beror på vilket land du kommer ifrån och hur länge dina studier pågår.
Det är mycket viktigt att din försäkring är i kraft hela den tid som du vistas i Finland.
Läs mer på InfoFinlands sida Studerande.
Studier i Finland
Om du inte är medborgare i ett EU-land eller EES-land och inte heller familjemedlem till en medborgare i ett sådant land och du kommer till Finland för att studera i augusti 2017 eller senare, måste du betala terminsavgift för studierna.
Avgiften gäller lägre och högre högskolestudier på engelska.
I Finland kan du studera på finska, svenska och ibland även på engelska.
Högskolorna har vissa utbildningsprogram där undervisningen ges på engelska.
Merparten av studierna är dock på finska eller på svenska.
I Finland finns många aktiva studentorganisationer.
De ordnar verksamhet även för utländska studerande.
I studentorganisationerna lär du dig känna nya människor.
Om du vill hitta en arbetsplats i Finland ska du studera finska eller svenska.
Även om du klarar dig i många dagliga situationer på engelska kräver de flesta arbetsgivare att du kan finska eller svenska.
Läs mer på InfoFinlands sida Finska och svenska språket.
Om inte hinner studera finska vid din egen läroanstalt, finns det kurser i finska vid många andra läroanstalter.
Du kan även studera språket på Internet.
Läs mer på InfoFinlands sida Finska och svenska språket.
Det är också viktigt att du bekantar dig med finländare och arbetslivet i Finland redan under studietiden.
På så sätt hittar du lättare vänner och ett arbete.
Till exempel arbetspraktik (työharjoittelu), hobbyer och organisationer är bra sätt att lära känna det finländska samhället.
Information för utländska studerandeengelska
Information om utbytesprogrammetengelska
Gymnasieansökan
Sök till gymnasiet i den gemensamma ansökan till andra stadiet i februari-mars.
Du kan söka till ett gymnasium om du har avlagt lärokursen för den grundläggande utbildningen eller en lärokurs som motsvarar den grundläggande utbildningen.
Fyll ansökan i tjänsten Studieinfo.fi.
Eleverna antas till gymnasiet utifrån vitsorden på avgångsbetyget från grundskolan.
Därtill ordnar vissa gymnasier inträdesprov.
Om du söker till ett vuxengymnasium, kontakta läroanstalten direkt.
Du kan inte söka till ett vuxengymnasium i den gemensamma ansökan.
När du söker till ett vuxengymnasium är inte medeltalet på ditt betyg av betydelse.
Du hittar utbildningar på Studieinfo.fi.
Om du vill förbättra dina kunskaper i finska innan du söker till ett gymnasium, kan du söka till en förberedande gymnasieutbildning
Läs mer på InfoFinlands sida Gymnasieförberedande utbildning.
Ansökan till gymnasium i den gemensamma ansökanfinska _ svenska
Ansökan till yrkesutbildning
Din grundutbildning avgör till hurudan yrkesutbildning du kan söka och på vilket sätt ansökan sker.
Du kan söka till en grundskolebaserad yrkesutbildning om du har avlagt lärokursen för den grundläggande utbildningen eller en lärokurs som motsvarar den grundläggande utbildningen.
Du kan söka till en gymnasiebaserad yrkesutbildning om du har gått färdigt gymnasiet.
Du kan söka till dessa utbildningar i den kontinuerliga ansökan året om eller i den gemensamma ansökan till andra stadiet.
I allmänhet ordnas den gemensamma ansökan i februari-mars.
Fyll ansökan i tjänsten Studieinfo.fi.
Om du redan har avlagt en yrkesexamen eller en högskoleexamen, kan du inte söka till en yrkesutbildning i den gemensamma ansökan.
Då kan du söka till utbildningen i den kontinuerliga ansökan.
Du ska söka till utbildningen i den kontinuerliga ansökan också om du är i arbetslivet och vill byta bransch eller om du vill ansöka till läroavtalsutbildning.
Du kan söka i den kontinuerliga ansökan även i det fall att du inte fick en studieplats i den gemensamma ansökan.
Grunderna för antagning av studeranden beror på utbildningen.
I allmänhet påverkas antagningen av antagningspoängen, som ges bl.a. utifrån dina betyg.
Inträdesprov eller lämplighetsprov ordnas också för många utbildningar.
I vissa branscher ställs krav på hälsotillståndet.
Läroanstalten kan kontrollera att du har tillräckliga språkkunskaper för studierna.
Fråga mer vid den läroanstalt som du ansöker till.
Om du vill ha mera kunskap och färdigheter innan du söker till en yrkesinriktad utbildning, kan du ansöka till VALMA-utbildningen.
Under VALMA-utbildningen kan du även förbättra dina språkkunskaper i finska.
Läs mera på InfoFinlands sida Utbildning som handleder för yrkesutbildning.
Om du behöver särskilt stöd i de yrkesinriktade studierna t.ex. på grund av handikapp eller inlärningssvårigheter ska du ansöka till utbildningen via ansökan till specialundervisning.
Ansökan till yrkesutbildning i den gemensamma ansökanfinska _ svenska
Kontinuerlig ansökan till yrkesutbildning finska _ svenska
Antagningsgrunder till yrkesutbildningfinska _ svenska
Om du har en utländsk examen
Om du har avlagt grundskolan eller gymnasiet utomlands, antas du till en yrkesutbildning enligt prövning.
Vid antagning enligt prövning beaktas
ditt utbildningsbehov
bedömningen av hur bra du kan klara av studierna.
Antagning enligt prövningfinska _ svenska
Ansökan till en yrkesinriktad vuxenutbildning
Du kan söka till en yrkesinriktad vuxenutbildning om du vill avlägga en examen vid sidan om arbetet.
I vuxenutbildningen avlägger du yrkesexamen som fristående examen.
Du kan söka till en yrkesinriktad vuxenutbildning också om du har avlagt en yrkesexamen eller en högskoleexamen.
När du söker till en yrkesinriktad vuxenutbildning, ska du ha en tillräckligt lång arbetserfarenhet.
Du kan inte söka till en yrkesinriktad vuxenutbildning i den gemensamma ansökan.
Ta reda på hur du kan söka till utbildningen i tjänsten Studieinfo.fi eller av läroanstalten.
Ofta är ansökningstiden fortlöpande.
Ansökan till en yrkeshögskola
Du kan söka till en yrkeshögskola för att avlägga en yrkeshögskoleexamen, då du har avlagt t.ex. någon av följande utbildningar:
gymnasiet studentexamen
en yrkesexamen
studentexamen eller en motsvarande examen i ett annat land
Du får närmare uppgifter från tjänsten Studieinfo.fi.
Sök till en yrkeshögskola i den gemensamma ansökan till högskolor.
Den gemensamma ansökan ordnas två gånger per år, på våren och på hösten.
Fyll ansökan i tjänsten Studieinfo.fi.
Grunderna för antagning av studeranden beror på utbildningen.
Ditt betyg, inträdesprovet och din arbetserfarenhet kan påverka antagningen.
Också dina tidigare studier kan spela en roll.
Ansökan till YH-examenfinska _ svenska
Högre yrkeshögskoleexamina
Du kan söka till en YH-examen om du har
en lämplig yrkeshögskoleexamen eller en annan lämplig högskoleexamen och
minst tre års arbetserfarenhet från samma område som din examen och du har inhämtat din arbetserfarenhet efter att du har avlagt examen.
Sök till en YH-examen i den gemensamma ansökan till högskolor på våren eller hösten Till många utbildningar är det möjligt att söka endast på våren.
Fyll i ansökningsblanketten i tjänsten Studieinfo.fi.
Du kan söka till en högre YH-examen på ett främmande språk med en separat ansökan.
Du hittar ansökningsblanketter då du letar efter utbildningar i Studieinfo.fi.
Högre YH-examenfinska _ svenska
Ansökan till universitet
Ansök till ett universitet antingen i den gemensamma ansökan till högskolor eller med en separat ansökan till en viss utbildning.
Du kan söka till många universitetsutbildningar i den gemensamma ansökan till högskolor.
Den ordnas på våren och hösten.
Alternativen är fler på våren.
Den gemensamma ansökan till vissa utbildningar ordnas redan i januari.
Utred i tid när du kan söka.
Fyll ansökan i tjänsten Studieinfo.fi.
Du kan söka till ett universitet om du har avlagt t.ex. någon av följande examina:
en finländsk studentexamen
en minst treårig yrkesinriktad grundexamen
en utländsk examen, som ger möjlighet till universitetsstudier i det land där du avlagt examen
Granska av högskolans studiebyrå att det är möjligt att söka till ett universitet med din examen.
Du får närmare uppgifter också från tjänsten Studieinfo.fi.
När du söker till ett universitet, får du i allmänhet poäng utifrån studentexamen och inträdesprovet.
Det finns skäl att förbereda dig omsorgsfullt för inträdesprovet.
Till vissa utbildningsprogram antas endast en liten del av sökandena.
Vissa inträdesprov omfattar förhandsuppgifter.
Ansökan till universitetfinska _ svenska _ engelska
Separat ansökan
Ansökan till vissa universitetsstudier sker genom en separat ansökan.
Du ska söka med en separat ansökan t.ex.
om du söker till ett magisterprogram
om du flyttar från en högskola till en annan eller
om du har avlagt studier i ett öppet universitet och söker till ett universitet utifrån dessa studier.
Om du söker till ett utbildningsprogram där undervisningsspråket är ett annat än finska eller svenska, beror ansökningssättet på utbildningen.
Det lönar sig att söka till vissa utbildningar på främmande språk i den gemensamma ansökan i januari.
Du hittar närmare information i Studieinfo.fi.
Du kan också fråga direkt av högskolorna.
De separata ansökningarna kan ordnas under olika tidsperioder och ansökningsförfarandena kan avvika från varandra.
Du hittar de separata ansökningarna via tjänsten Studieinfo.fi.
Påbyggnadsexamen
Om du vill avlägga en påbyggnadsexamen vid ett universitet, kontakta universitetet direkt.
Mottagande av studieplats
Läroanstalten meddelar dig att du har antagits för studier med ett brev.
Om du har antagits, meddela så fort som möjligt till läroanstalten att du tar emot studieplatsen.
Brevet innehåller anvisningar om hur du tar emot platsen och hur du anmäler dig.
Om du inte tar emot platsen i tid, förlorar du den.
När du tar emot en studieplats, förbinder du dig att börja studera i läroanstalten.
Du kan söka till många olika läroanstalter i den gemensamma ansökan.
Du kan dock ta emot endast en studieplats.
Vilka hälsotjänster kan du använda?
Offentliga hälsovårdstjänster
Privata hälsovårdstjänster
Hälsovård för medborgare i de nordiska länderna
Hälsovård för EU-medborgare
Hälsovård för anställda och företagare
Hälsovård för studerande
Hälsovård för invandrare och asylsökande
Hälsovård för papperslösa
Information på webben
Vilka hälsotjänster kan du använda?
Du kan utnyttja de offentliga hälsovårdstjänsterna i Finland om du har hemkommun (kotikunta) i Finland.
Rätten till hemkommun beror på följande:
från vilket land du kommer till Finland
varför du kommer till Finland (t.ex. arbete, studier)
om du ska bo stadigvarande i Finland eller vistas här tillfälligt
om din vistelse i Finland är tillfällig, beroende på hur länge vistelsen varar.
Om du inte är säker på om du har hemkommun i Finland kan du ta reda på din situation vid magistraten (maistraatti).
Mer information finns på InfoFinlands sida Hemkommun i Finland.
Om du arbetar i Finland, kan du ha rätt till den offentliga hälso- och sjukvården även om du inte har en hemkommun i Finland.
Om du inte har en hemkommun i Finland ska du be FPA utreda din rätt till den offentliga hälso- och sjukvården.
I nödfall får du vård inom den offentliga hälso- och sjukvården fastän du inte har en hemkommun i Finland eller rätt till vård på grund av arbete.
Du kan krävas på vårdkostnaderna i efterhand.
Om du inte har rätt till de offentliga hälsovårdstjänsterna, kan du boka tid på en privat läkarstation.
Privata hälsovårdstjänster är avsevärt dyrare för kunden än de offentliga.
Hälsovårdstjänster ges i Finland på finska och svenska.
Ofta klarar man sig även på engelska.
När du bokar tid till hälsovårdstjänster kan du fråga om möjligheten att använda en tolk (tulkki) om du inte behärskar dessa språk.
Läs mer på InfoFinlands sida Behöver du en tolk?
När du har bokat tid för ett läkarbesök ska du vara punktligt på plats.
Om du har bokat tid för ett läkarbesök men får förhinder är det mycket viktigt att du avbokar besöket i god tid, helst dagen innan.
Om du inte kommer och inte heller har avbokat din tidsbeställning måste du betala en avgift.
Hälsa och rehabiliteringfinska _ svenska _ ryska _ estniska
Sjukvård för utlänningar i Finlandfinska _ svenska _ engelska
Kontaktpunkt för gränsöverskridande hälso- och sjukvårdfinska _ svenska _ engelska
linkkiStödcentralen Hilma för funktionshindrade invandrare :
Handbok med ordlista i hälso- och sjukvård på finska(pdf, 341,02 kt)finska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska
Offentliga hälsovårdstjänster
När du blir sjuk ska du först kontakta din egen hälsostation (terveysasema). Där kan du boka tid hos en allmänläkare eller en hälsovårdare.
Mer information om hälsovårdstjänsterna i olika kommuner hittar du på InfoFinlands sida på de lokala informationssidorna eller på din egen kommuns sida.
Hälsostationens tjänster är relativt förmånliga för klienten eftersom de finansieras med skattemedel.
Hälsostationerna har vanligen öppet från måndag till fredag kl. 310 1671.
Det är klokt att ringa tidsbeställningen genast på morgonen när hälsostationen öppnar.
Om ditt besvär kräver brådskande vård får du en tid snabbt.
Om du inte behöver brådskande vård måste du vänta längre på att få en läkartid.
Vid tidsbeställningen får du veta hur snabbt du kommer att få vård.
Vid tidsbeställningen bedöms även om du behöver vård av läkare eller hälsovårdare.
I Finland kan hälsovårdare ge vård vid flera sjukdomar.
Vid behov kan hälsovårdaren ge remiss till läkare.
Om du har ett FPA-kort (Kela-kortti) ska du ta det med när du besöker hälsovårdsstationen.
Om du behöver en specialist, ska du först boka tid hos en allmänläkare.
Vid behov skriver hälsostationsläkaren en remiss till en specialist.
Specialister finns på vissa hälsostationer, på polikliniker och sjukhus.
Specialsjukvård ges på centralsjukhus och universitetssjukhus.
I Finland gör läkare inom de offentliga hälsovårdstjänsterna inga hembesök.
En del privata läkarstationer erbjuder denna tjänst. Ett hembesök av en privatläkare är dock dyrt.
Om din sjukdom är långvarig och du inte kan arbeta finns det mer information om FPA:s sjukpenning på InfoFinlands sida Stöd när du är sjuk.
Jour inom offentliga hälsovårdstjänster
Hälsostationerna har stängt kvällstid och under veckoslut.
Då vårdas akuta sjukfall på jourmottagningen (päivystys).
Jourmottagningen är avsedd för situationer där man behöver omedelbar vård.
Om din sjukdom inte kräver omedelbar vård ska du beställa tid på din egen hälsostation nästa gång den har öppet.
Jourmottagningen finns ofta i anslutning till sjukhus, i små städer också i en närliggande stad.
Jourmottagningen för barn och unga finns ofta separat.
Fråga mer vid din egen hälsostation under dess öppettider eller leta upp informationen på din hemkommuns webbplats.
Privata hälsovårdstjänster
Kontaktuppgifter till privata läkarstationer hittar du till exempel på internet.
Förmodligen får du en tid snabbare på en privat hälsostation än inom den offentliga hälsovården.
Privata hälsotjänster är avsevärt dyrare för klienten än de offentliga.
Olika läkarstationer erbjuder olika tjänster.
Privata hälsotjänster kan användas av alla, även personer som inte har en hemkommun i Finland.
Om du omfattas av den finländska sjukförsäkringen (sairausvakuutus) ersätter FPA en liten del av kostnaderna för privat sjukvård och tandvård.
Ibland kan också personer som inte omfattas av den finländska sjukförsäkringen ha rätt till ersättning från FPA.
Fråga mer hos FPA.
FPA:s ersättning kan ibland dras av direkt på det belopp som du betalar vid kassan.
Du kan också söka ersättning från FPA i efterhand.
Läs mer om sjukförsäkringen i Finland på InfoFinlands sida Den sociala tryggheten i Finland.
Sjukvårdsersättningarfinska _ svenska _ engelska
Jämför läkarpriserfinska _ engelska
Privat läkarstationfinska _ svenska _ engelska
Privat läkarstationfinska _ svenska _ engelska
linkkiAava:
Privat läkarstationfinska _ svenska _ engelska
Hälsovård för medborgare i de nordiska länderna
Om du har en sjukförsäkring i ett annat nordiskt land har du rätt till nödvändig sjukvård i Finland.
Du får vård på samma villkor och till samma kostnad som finländarna.
Ta med dig ett officiellt identitetsbevis när du använder hälsovårdstjänsterna.
Hälsovård för EU-medborgare
Om du har en sjukförsäkring i ett annat EU-land, EES-land eller i Schweiz har du rätt till nödvändig sjukvård i Finland.
För att få vård måste du ha ett europeiskt sjukvårdskort.
Du ska skaffa dig det europeiska sjukvårdskortet i det land där du har din sjukförsäkring.
Det europeiska sjukvårdskortet ger dig rätt till vård om du blir sjuk eller råkar ut för en olycka.
Du får vård även vid en långvarig sjukdom.
Med kortet får du även vård i samband med graviditet och förlossning.
Du får vård till samma kostnad som personer som är stadigvarande bosatta i Finland.
Information om det europeiska sjukvårdskortetfinska _ svenska _ engelska
Hälsovård för anställda och företagare
Om du har kommit till Finland för att arbeta kan du ha rätt att använda de offentliga hälsovårdstjänsterna i Finland.
Detta beror på hurdant och hur långt arbetsavtal du har samt från vilket land du har kommit till Finland.
I Finland är arbetsgivare skyldiga att ordna förebyggande företagshälsovård för sina anställda.
Företagare kan ordna sin egen företagshälsovård om de vill.
Företagare måste alltså inte ordna företagshälsovård för sig.
Företagare måste ändå ordna företagshälsovård för sina anställda.
Företagshälsovården kan ordnas vid den lokala hälsovårdscentralen eller till exempel på en privat läkarcentral.
Mer information får du på InfoFinlands sida Företagshälsovården och på social- och hälsovårdsministeriets webbplats.
linkkiSocial- och hälsovårdsministeriet:
Företagshälsovårdfinska _ svenska _ engelska
Hälsovård för studerande
Om du kommer från ett land som inte är ett EU-land, ett EES-land eller Schweiz till Finland för att studera behöver du vanligtvis ha en täckande sjukförsäkring i ditt hemland för att få uppehållstillstånd i Finland.
Om dina studier beräknas pågå i minst två år får du vanligen en hemkommun i Finland och rätt till de kommunala hälsovårdstjänsterna.
I detta fall räcker det om din sjukförsäkring i första hand täcker läkemedelskostnaderna.
Om du inte är säker på om du har rätt till hemkommun i Finland kan du kontrollera detta vid magistraten.
Du får mer information om hemkommun på InfoFinlands sida Hemkommun i Finland.
Mer information om uppehållstillstånd för studerande och om den sjukförsäkring som krävs för att få uppehållstillstånd får du på Migrationsverkets (Maahanmuuttovirasto) webbplats.
I Finland omfattas högskolestuderande av studerandehälsovården.
Fråga mer vid din egen läroanstalt.
Mer information om studerandehälsovården får du på Studenternas hälsovårdsstiftelses (SHVS) (YTHS) och social- och hälsovårdsministeriets (Sosiaali- ja terveysministeriö) webbplatser.
Information om uppehållstillstånd för studierfinska _ svenska _ engelska
linkkiSHVS:
Hälsovård för högskolestuderandefinska _ svenska _ engelska
linkkiSocial- och hälsovårdsministeriet:
Studerandehälsovårdfinska _ svenska
Hälsovård för invandrare och asylsökande
Om du har kommit till Finland som kvotflykting har du hemkommun i Finland och rätt att utnyttja de offentliga hälsovårdstjänsterna.
Om du är asylsökande och din ansökan inte ännu har behandlats kan du inte registrera dig i magistraten som kommuninvånare och inte heller utnyttja kommunens hälsovårdstjänster.
Fråga mer vid din förläggning.
Om du har fått uppehållstillstånd på grund av behovet av skydd och får rätt till hemkommun i Finland, kan du utnyttja hälsovårdstjänsterna i din egen kommun.
Läs mer om rätten till hemkommun på InfoFinlands sida Hemkommun i Finland.
Hälsovård för papperslösa
Global Clinic är en klinik där du kan få hjälp eller råd av en läkare eller sjukskötare om du vistas i Finland utan uppehållstillstånd.
Global Clinic bedriver verksamhet i följande städer:
Åbo
Uleåborg
Joensuu
Tammerfors
Du kan ringa eller skicka e-post.
En sjukskötare eller läkare besvarar ditt samtal.
Du hittar kontaktinformation på Global Clinic:s hemsidor.
Global Clinic:s tjänster är avgiftsfria för kunderna.
Global Clinic anmäler inte sina kunder till polisen eller andra myndigheter.
Klinikens adress eller öppettider meddelas inte offentligt.
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Information på webben
linkkiTuberkuloosi.fi:
Information om tuberkulosfinska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Din situation avgör hur du kan finansiera dina studier i Finland.
På den här sidan berättar vi om FPA:s stöd till studerande samt om penningunderstöd och stipendier.
Studiestöd
Du kan få FPA:s studiestöd (opintotuki) om du
har det uppehållstillstånd (oleskelulupa) som krävs och
vistas i Finland av någon annan orsak än studier.
Om du flyttar till Finland för att studera kan du inte få studiestöd.
Till exempel utbytesstuderande får inte finskt studiestöd.
Studiestödet består av studiepenning och statsborgen för studielån.
Du kan få studiestöd om
Du studerar i gymnasiet
Du studerar vid en yrkesläroanstalt eller avlägger yrkesinriktade tilläggsstudier
Du studerar vid en högskola.
Du kan få studiepenning om du har fyllt 17 år.
Du måste studera på heltid.
Med heltidsstudier avses att studierna är din huvudsyssla.
Du kan arbeta vid sidan av studierna.
Lönen som du får för ditt arbete kan minska ditt studiestöd.
Du ansöker om studiepenning och statsgaranti för studielån vid FPA.
FPA betalar in studiepenningen på ditt konto månatligen.
På studiepenningens belopp inverkar många omständigheter.
På studiepenningens belopp inverkar bland annat stödmottagarens ålder, om hen bor i sitt eget hem eller hos en förälder, on hen är gift och om hen har minderåriga barn. Kontrollera storleken på din studiepenning på FPA:s webbplats eller vid en FPA-byrå.
Det är inte obligatoriskt att ta studielån.
Du kan högst ta ut ett visst maximibelopp.
Du väljer själv hur mycket studielån du vill ta.
Studielånet är ett lån som finska staten ger garanti för åt studeranden.
Du ansöker om lånet i banken när du har fått FPA:s beslut om statsgaranti.
Du måste betala tillbaka lånet när du har slutfört dina studier.
Du kan få studielån också när du fortbildar dig (täydennyskoulutus) som vuxen.
Dessutom kan du få vuxenutbildningsstöd (aikuiskoulutustuki).
I vissa fall kan du också få bostadstillägg, till exempel om du studerar på en avgiftsbelagd linje vid en folkhögskola och bor på läroanstaltens internat.
Läs mer på FPA:s webbplats.
På InfoFinlands sida Bostadsbidrag finns mer information om FPA:s allmänna bostadsbidrag.
Information om studiestödetfinska _ svenska _ engelska
Information om studiestödetryska _ estniska _ samiska
Information om att ansöka studiestödfinska _ svenska _ engelska
Studiestöd till utländska studerandefinska _ svenska _ engelska
Stöd för skolresor
Du kan få stöd för skolresor (koulumatkatuki) om du bor i Finland och studerar i gymnasiet eller vid en yrkesläroanstalt.
Din skolresa måste vara minst 10 kilometer lång och resekostnaderna måste överstiga 54 euro per månad.
Information om skolresestödetfinska _ svenska _ engelska
Måltidsstöd
Om du studerar vid en högskola får du också måltidsstöd (ateriatuki).
Du kan få måltidsstödet endast i läroanstalternas egna restauranger.
Detta innebär att studeranden betalar mindre för måltiderna än andra som besöker restaurangen.
Du behöver inte ansöka separat om måltidsstödet.
Du behöver bara visa upp ditt studentkort när du betalar för måltiden.
Du har inte rätt till måltidsstöd om du är i Finland endast på arbetspraktik (työharjoittelu) som ingår i en utländsk examen.
Information om måltidsstödetfinska _ svenska _ engelska
Penningunderstöd och stipendier
Utländska studerande kan ansöka om olika penningunderstöd för finländska högskolor.
Alla finländska högskolor har ett eget stipendiesystem för de studerande som kommer från länder utanför EU/EES-området och som har godkänts för att avlägga en kandidat- eller magisterexamen på engelska.
Möjligheten till ett stipendium kan till exempel bero på hur framgångsrik du varit i dina studier.
Stipendiet kan täcka hela läsårsavgiften eller en del av den.
Vissa stipendier kan även täcka andra kostnader.
Ibland krävs att du lyckas tillräckligt bra med dina studier för att du ska få ett stipendium.
Du kan vanligtvis ansöka om ett stipendium samtidigt som du ansöker om en studieplats.
Det finns också särskilda Erasmus Mundus-magisterprogram som har ett eget stipendiesystem.
Utbildningsstyrelsen har stipendieprogram för forskarstuderande som kommer till Finland för att avlägga doktorsexamen.
Studerande från USA kan ansöka om ett Fulbright-stipendium.
Läs mer om stipendier och penningunderstöd på webbplatsen Studyinfinland.fi.
I Finland kan man avlägga högskolestudier både vid yrkeshögskolor och vid universitet.
Läs mer om yrkeshögskolan på InfoFinlands sida Yrkeshögskolor.
Ansök om studieplats
Du kan söka till ett universitet om du har avlagt en finländsk studentexamen, en utländsk examen som motsvarar studentexamen eller en yrkesinriktad slutexamen. Sök till ett universitet i den gemensamma ansökan till högskolor.
Läs mer på InfoFinlands sida Ansökan till utbildning.
Gemensam ansökan till universitetfinska _ svenska
Vilka yrken kan studera till?
Vid universitet kan man studera i många olika studieområden.
De som har utexaminerats från en högskola eller ett universitet arbetar i många slags arbetsuppgifter.
En del universitetsstudier leder direkt till ett yrke.
Sådana yrken är till exempel:
lärare
jurist
läkare
skådespelare
diplomingenjör
bildkonstnär
Andra universitetsstudier leder inte till ett visst yrke.
Till exempel studerande vid den samhällsvetenskapliga eller den humanistiska fakulteten utexamineras inte nödvändigtvis till ett yrke.
Dessa människor arbetar till exempel i följande arbetsuppgifter:
forskare
statlig tjänsteman
Studier vid universitet
Vid vissa universitet har olika examen olika namn.
Till exempel är tekniska högskolors motsvarighet till magisterexamen diplomingenjörsexamen (diplomi-insinööri).
När du får en studieplats får du rättighet att avlägga båda examina.
Du kan också avsluta studierna efter lägre högskoleexamen.
Kandidatstudierna pågår ungefär tre år, magisterstudierna ungefär två år.
Hur fort studierna framskrider beror på dig själv.
Du kan också söka till ett separat magisterprogram.
Magisterprogrammet är ett studieprogram som leder till högre högskoleexamen.
För att kunna studera i ett magisterprogram ska du ha avlagt lägre högskoleexamen.
Magisterprogrammen pågår i cirka två år.
Vid dem studerar ofta människor från många olika vetenskapsområden.
Utexaminering från universitetet
När du är klar med dina studier får du antingen kandidatexamen eller magisterexamen.
Om du vill kan du efter magisterexamen söka till fortsatta studier.
Information om högskolestudierfinska _ svenska _ engelska
linkkiFinlands Studentkårers Förbund:
Information om studentkårer i Finlandfinska _ svenska _ engelska
Öppna universitet
De öppna universiteten tillhandahåller universitetskurser.
Vem som helst kan studera vid ett öppet universitet.
Du kan studera vid ett öppet universitet även om du inte har någon examen.
Läs mer på InfoFinlands sida Studier som hobby.
Vetenskaplig fortbildning vid universitet
Vetenskaplig fortbildning vid universitet är examensinriktad fortbildning.
Sådan utbildning förbereder dig till exempel för forskaryrket.
Vid universitetet kan du avlägga licentiatexamen (lisensiaatti) eller doktorsexamen (tohtori).
De flesta studerande som bedriver fortsatta studier avlägger doktorsexamen.
Man kan ansöka till fortsatta studier vid universitet några gånger per år.
Universitet och institutioner har olika ansökningstider.
Kontrollera ansökningstiden vid den institution där du vill bedriva fortsatta studier.
I Finland måste de som bedriver fortsatta studier ofta finansiera studierna själva.
Du kan ansöka om stipendier hos olika stiftelser (säätiö).
Påbyggnadsexamina vid universitetfinska
linkkiStiftelsetjänst:
Information om stiftelser och penningunderstödfinska _ svenska _ engelska
linkkiUtbildningsstyrelsen:
Penningunderstöd för utländska forskarefinska _ engelska
Vägledning i högskolestudier
Vid högskolornas SIMHE-tjänster kan du söka hjälp och information om högskoleutbildning i Finland och om hur du ansöker till högskoleutbildning.
Du kan även få information om andra utbildningsmöjligheter för personer som avlagt högskolestudier.
Du kan få vägledning via SIMHE-tjänsterna om
du har flyttat till Finland
du är intresserad av högskolestudier och
du har avlagt högskolestudier eller högskoleexamen utomlands.
Vägledning kan ges individuellt eller i grupp.
linkkiUtbildningsstyrelsen:
Högskolor som erbjuder SIMHE-tjänsterfinska _ engelska
Högskolor som erbjuder SIMHE-tjänsterfinska _ svenska _ engelska
Nödnumret (hätänumero) i Finland är 112.
Du får ringa nödnumret endast i brådskande nödfall där liv, hälsa, egendom eller miljö är i fara.
I nödsituationer får du vård även om du inte har en hemkommun i Finland.
Vårdavgifter kan komma att debiteras av dig i efterhand.
Ring 112 till exempel i följande situationer:
du har råkat ut för en bilolycka (auto-onnettomuus) eller är vittne till en olycka
någon är i livsfara (hengenvaara)
du upptäcker en brand (tulipalo)
du upptäcker ett inbrott (murto)
Ring inte nödnumret om ärendet inte är brådskande.
Du ska inte ringa nödnumret vid vanliga sjukdomsfall.
Du ska inte heller ringa nödnumret om du vill fråga polisen (poliisi) till exempel om ett tillståndsärende.
Onödiga samtal kan orsaka att hjälpen kommer för sent i verkliga nödsituationer.
Du kan straffas för att ha missbrukat nödnumret.
Samtalet besvaras av en utbildad nödcentraloperatör.
Han eller hon ställer dig frågor och bedömer hjälpbehovet.
Därefter larmar han eller hon hjälp.
Operatören berättar också vad du ska göra.
Operatören kopplar inte samtalet vidare, så besvara frågorna noga.
Du kan tala finska eller svenska när du ringer nödnumret.
Du kan också fråga om nödcentraloperatören förstår engelska, med det är inte säkert.
Vid behov bistås nödcentralen av en tolktjänst.
Du kan ringa nödnumret gratis från alla telefoner.
Du behöver inget riktnummer.
Du kan ringa nödnumret utan riktnummer även om du har ett utländskt mobilabonnemang.
Nödnumret 112 fungerar i alla EU-länder.
Om du har installerat den kostnadsfria mobilappen 112 Suomi i din telefon, behöver du inte nödvändigtvis kunna berätta var du befinner dig.
Nödcentraloperatören ser var du är, när du ringer ett nödsamtal via appen.
Du kan ladda ned appen i applikationsbutiken.
När du ringer nödnumret 112:
uppge ditt namn
berätta vad som har hänt
ange exakt adress och kommun
svara på nödcentraloperatörens frågor
följ instruktionerna
avsluta inte samtalet förrän du får lov.
Mer information om nödnumret får du på Nödcentralsverkets (Hätäkeskuslaitos) webbplats.
Om du behöver information om tillståndsärenden som sköts av polisen, fordonsföreskrifter eller hur undersökningen i ett brott som skett tidigare framskrider ska du ringa polisens egna nummer under tjänstetid.
Om du misstänker att någon har förgiftats kan du fråga råd vid Giftinformationscentralen (Myrkytystietokeskus).
Giftinformationscentralens telefontjänst är öppen 24 timmar om dygnet.
Telefonnumret är (09) 471 977.
linkkiNödcentralsverket:
Nödsituationfinska _ svenska _ engelska
linkkiNödcentralsverket:
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
linkkiRöda Kors:
Första hjälpen-anvisningar för olika situationerfinska _ svenska _ engelska
Första hjälpen-anvisningar vid förgiftningfinska _ svenska _ engelska
Studierna är inte alltid inriktade på att skaffa ett yrke.
Du kan också ha studier som hobby.
Du kan studera vid flera olika läroanstalter: öppna universitetet (avoin yliopisto) eller öppna yrkeshögskolan (avoin ammattikorkeakoulu), sommaruniversitetet (kesäyliopisto), senioruniversitetet (ikäihmisten yliopisto), medborgarinstitut (kansalaisopisto), arbetarinstitut (työväenopisto) och folkhögskolor (kansanopisto).
Studierna är vanligen avgiftsbelagda.
Många av dessa läroanstalter tillhandahåller undervisning i finska och svenska för invandrare.
Läs mer på InfoFinlands sida Finska och svenska språket.
Du kan även studera flera andra språk, såsom engelska eller franska.
Vid folkhögskolor kan du även avlägga yrkesexamen.
Öppna universitetet och öppna yrkeshögskolan
Öppna universitetet (avoin yliopisto) och öppna yrkeshögskolan (avoin ammattikorkeakoulu) ordnar universitets- och yrkeshögskolekurser.
Vem som helst kan studera vid de öppna högskolorna.
Du kan studera vid öppna högskolor fastän du inte har någon examen.
Du kan studera vid öppna högskolor
om du vill studera som hobby
om du vill bli antagen för studier i ett visst ämne vid en högskola
när du vill utöka din yrkeskunnighet och dina kunskaper
Till de öppna högskolorna ordnas inga inträdesprov.
Du kan anmäla dig till vårens kurser i början av året och till höstens kurser i slutet av sommaren.
Anmäl dig direkt till kurserna.
Du kan välja enskilda kurser eller större studiehelheter.
Vid öppna högskolor är studierna flexibla.
Du kan delta i kurser under dagtid, på kvällar eller på veckoslut.
Du kan också studera på internet.
Studierna vid öppna högskolor är inte heltidsstudier.
Du får därför inget studiestöd (opintotuki) och inga studentrabatter när du studerar vid öppna högskolan.
Du kan avlägga studier vid öppna högskolan fastän du får arbetslöshetsersättning (työttömyyskorvaus).
Du har nytta av studierna vid öppna högskolan när du studerar vidare. Om du blir antagen till yrkeshögskolan behöver du inte avlägga de kurser som du redan har avlagt vid öppna yrkeshögskolan.
Om du har studerat vid öppna universitetet och söker till universitetet ansöker du via separat ansökan (erillinen haku).
Information om öppna yrkeshögskolanfinska _ svenska
Information om öppna universitetetfinska _ svenska
Sommaruniversitetet
Kurserna vid sommaruniversitetet (kesäyliopisto) påminner mycket om kurserna vid öppna universitetet.
Man kan studera vid sommaruniversitetet även under andra tider än på sommaren.
Utöver universitetskurser ordnar sommaruniversiteten också annan undervisning, till exempel:
Yrkesinriktad fortbildning (täydennyskoulutus)
Arbetskraftsutbildning (työvoimakoulutus)
Abiturientkurser (abikurssi) för gymnasieelever som förbereder sig för studentskrivningarna
finskakurser för invandrare
Fråga närmare uppgifter om undervisningen vid närmaste sommaruniversitet.
Info om sommaruniversitetfinska _ svenska
Information om sommaruniversitetetfinska _ svenska _ engelska
Senioruniversitetet
Senioruniversitetet (ikäihmisten yliopisto) är avsett för dem som har fyllt 60 år.
Studietillfällena är dock öppna för alla.
Undervisningen vid senioruniversitetet är en del av öppna universitetets verksamhet.
Senioruniversitetet ordnar föreläsningsserier, kurser och studieresor.
Fråga mer om senioruniversitetet i kansliet för närmaste öppna universitet.
Medborgarinstitut och arbetarinstitut
I Finland finns många medborgarinstitut (kansalaisopisto) och arbetarinstitut (työväenopisto).
Vid dem kan du studera bland annat språk, handarbete, idrott, bildkonst och matlagning.
Medborgarinstituten och arbetarinstituten erbjuder hobbystudier.
Vid dem kan man inte avlägga yrkesinriktade studier.
Medborgarinstituten och arbetarinstituten ordnar finskakurser för invandrare.
Fråga närmare uppgifter om kurserna vid närmaste medborgarinstitut eller arbetarinstitut.
Ansökningspraxis varierar.
Vanligen ansöker man till vårens undervisning i början av året och till höstens undervisning på sensommaren.
Fråga om ansökningstiderna vid medborgarinstitutets eller arbetarinstitutets studiebyrå.
Info om medborgarinstituten och arbetarinstitutenfinska _ svenska
Medborgarinstitut i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Folkhögskolor
Folkhögskolorna (kansanopisto) erbjuder både hobbystudier och yrkesinriktad utbildning.
Folkhögskolan kan drivas av en organisation eller också kan de vara självständiga institut.
Vid folkhögskolan kan du utbilda dig till ett yrke.
Vid folkhögskolan kan man till exempel avlägga djurskötarexamen eller massörexamen.
Folkhögskolorna ordnar mycket undervisning för invandrare.
Vid folkhögskolan kan du studera finska eller delta i förberedande utbildning.
Folkhögskolorna ordnar vanligen två olika slags undervisning, kortkurser (lyhytkurssi) och långa utbildningslinjer (pitkä opintolinja).
Kortkurserna är öppna för alla och till dem behöver du inte söka.
Det räcker med att du anmäler dig.
De långa utbildningslinjerna är ofta yrkesinriktade studier.
De pågår vanligen från ett halvår till ett år.
Till de långa utbildningslinjerna måste man söka separat.
Folkhögskolornas ansökningspraxis och ansökningstider varierar.
Fråga mer om antagningen vid folkhögskolans studiebyrå.
Info om folkhögskolorfinska _ svenska
linkkiFinlands folkhögskolförening:
Information om folkhögskolorfinska
linkkiFinlands folkhögskolförening:
Kurser vid folkhögskolor för invandrarefinska
linkkiDövas folkhögskola:
Utbildning för döva invandrarefinska _ svenska _ engelska
Studierna vid en yrkeshögskola (ammattikorkeakoulu) är praktiskt inriktade.
När du utexamineras från en yrkeshögskola får du ofta ett yrke.
Vid yrkeshögskolorna studerar du på finska, svenska eller på engelska.
Vid många yrkeshögskolor finns engelskspråkiga utbildningsprogram.
Ansökan
Du kan söka till en yrkeshögskola då du har avlagt en yrkesskola, gymnasiet eller studentexamen i Finland eller i ett annat land.
Läs mer på InfoFinlands sida Ansökan till utbildning.
Gemensam ansökan till yrkeshögskolorfinska _ svenska
Studier
I yrkeshögskolor kan du studera inom många områden.
Inom parentes anges exempel på yrken som du studera till i olika studieområden:
Naturbruk- och miljöområdet (skogsbruksingenjör, landskapsplanerare)
Den humanistiska och pedagogiska branschen (teckenspråkstolk)
Kulturbranschen (musiker, inredningsarkitekt)
Turism- och kosthållsbranschen (hovmästare, hotellmedarbetare)
Social-, hälso- och idrottsområdet (barnmorska, fysioterapeut, sjuksköterska)
Samhällsvetenskaper, affärsekonomi och förvaltning (försäljningsförhandlare, marknadsföringsassistent)
Teknik och trafik (ingenjör inom bilteknik, maskinmästare i sjöfartsbranschen)
Heltidsstudierna pågår ungefär fyra år.
Studietiden beror på utbildningsprogrammet och din egen studietakt.
Studierna omfattar mycket praktiska övningar.
Studierna omfattar också en arbetspraktik.
Grundläggande information om yrkeshögskolorfinska _ svenska
linkkiUndervisnings- och kulturministeriet:
Förteckning över yrkeshögskolorfinska _ svenska
linkkiSAMOK:
Förbund för studerande vid yrkeshögskolorfinska _ svenska
Förberedande utbildning för invandrare
Yrkeshögskolan kan ordna avgiftsfri utbildning för invandrare med målet att ge den studerande tillräckliga språkkunskaper och andra färdigheter som behövs för att studera vid yrkeshögskolan.
Under studierna tränar studeranden sig i det finska språket, på att läsa saktexter och på sina studiefärdigheter.
Dessutom får studerandena information om utbildningsområdet, arbetsmöjligheter och studier som leder till examen.
Språkkunkapskravet för dem som söker till förberedande utbildning är oftast finskakunskaper på nivån B1 eller B2.
Öppna yrkeshögskolor
De öppna yrkeshögskolorna tillhandahåller yrkeshögskolekurser.
Vem som helst kan studera vid en öppen högskola.
Du kan studera vid en öppen yrkeshögskola även om du inte har någon examen.
Läs mer på InfoFinlands sida Studier som hobby.
Fortsatta studier vid yrkeshögskolor
Om du vill fördjupa dina yrkeskunskaper kan du avlägga högre yrkeshögskoleexamen (ylempi ammattikorkeakoulututkinto).
Den är avsedd för personer som har examen till exempel från en yrkeshögskola och som redan arbetar.
Du kan ansöka till högre yrkeshögskolestudier om du har
någon annan högskoleexamen
minst tre års arbetserfarenhet från en lämplig bransch
Sök till högre yrkeshögskolestudier i den gemensamma ansökan.
Gemensam ansökan ordnas två gånger per år, på hösten och på våren.
Läs mer om den gemensamma ansökan på InfoFinlands sida Ansökan till utbildning.
Du avlägger en högre yrkeshögskoleexamen på ungefär ett eller ett och ett halvt år.
Studiernas omfattning är 60 eller 90 studiepoäng.
Genom högre högskoleexamen kan du fördjupa och utvidga dina kunskaper inom ditt eget yrkesområde.
Till exempel sjukskötare kan avlägga högre yrkeshögskoleexamen inom rehabilitering.
Du kan också välja att avlägga en engelskspråkig examen.
Information om högre yrkeshögskoleexamenfinska _ svenska
Vägledning i högskolestudier
Vid högskolornas SIMHE-tjänster kan du söka hjälp och information om högskoleutbildning i Finland och om hur du ansöker till högskoleutbildning.
Du kan även få information om andra utbildningsmöjligheter för personer som avlagt högskolestudier.
Du kan få vägledning via SIMHE-tjänsterna om
du har flyttat till Finland
du är intresserad av högskolestudier och
du har avlagt högskolestudier eller högskoleexamen utomlands.
Vägledning kan ges individuellt eller i grupp.
Högskolor som erbjuder SIMHE-tjänsterfinska _ svenska _ engelska
linkkiUtbildningsstyrelsen:
Högskolor som erbjuder SIMHE-tjänsterfinska _ engelska
Om du har avlagt en examen utomlands kan du ha nytta av jämställande av examen, erkännande av yrkeskompetens eller av att skaffa dig rätt till yrkesutövning eller en fristående examen.
Erkännande och motsvarighet av examen
Erkännande av examen betyder ett avgörande om vilken behörighet en utländsk examen ger när man söker jobb eller studieplats i Finland.
Erkännande av examen är avgiftsbelagt och söks hos Utbildningsstyrelsen.
När du söker en studieplats krävs inte nödvändigtvis erkännande av examen.
Professionellt erkännande och rätt till yrkesutövning
Personer som söker till uppgifter inom den offentliga sektorn (staten och kommunerna) måste ofta uppfylla vissa behörighetsvillkor beträffande utbildningen.
När någon som studerat utomlands söker till dessa uppgifter behöver han eller hon oftast Utbildningsstyrelsens avgörande om den tjänstebehörighet som hans eller hennes examen ger.
Ett reglerat yrke avser en uppgift som endast kan sökas av personer som har avlagt en viss lagstadgad examen eller vissa studier.
Till reglerade yrken hör både uppdrag inom den offentliga sektorn och yrken för vilka det krävs rätt till yrkesutövning.
Rätt till yrkesutövning krävs till exempel i yrken inom hälsovården och sjöfarten.
Om du har en utländsk examen i något yrke som är reglerat i Finland behöver du ett beslut från någon behörig myndighet innan du kan utöva yrket Finland.
På Utbildningsstyrelsens webbplats finns en förteckning över de reglerade yrkena och de ansvariga myndigheterna.
I den privata sektorn kan arbetsgivaren själv bedöma huruvida den anställdas utländska examen godtas.
I den privata sektorn krävs inget beslut om erkännande, men beslutet kan vara nyttigt då man söker jobb.
Utbildningsstyrelsen ger också expertutlåtanden om utländska yrkesexamina.
Ett sådant utlåtande ger inte tjänstebehörighet i Finland, men det kan ändå vara till hjälp när man ansöker om ett arbete eller en studieplats, eftersom det beskriver innehållet i och nivån på utbildningen som man har avlagt utomlands.
Akademiskt erkännande
Om du vill fortsätta dina studier i Finland kan de studier som du avlagt utomlands tillgodoräknas med hjälp av akademiskt erkännande.
Akademiskt erkännande av examina betyder
att man söker sig till en utbildning på basis av sin utländska utbildning
att de utländska studierna tillgodoräknas som en del av en finländsk examen.
Läroanstalterna beslutar själva om antagningen av studerande och om de tillgodoräknar utländska studier som en del av en examen som avläggs i Finland.
Fråga mer vid den läroanstalt där du vill studera.
linkkiUtbildningsstyrelsen:
Erkännande av en examenfinska _ svenska _ engelska
linkkiUtbildningsstyrelsen :
Broschyr om erkännande av examen(pdf, 102,14 kt)finska _ svenska _ engelska _ ryska _ estniska _ franska _ spanska _ kinesiska _ persiska _ arabiska
linkkiUtbildningsstyrelsen :
Diagram över erkännande av examen(pdf, 410,87 kt)finska _ svenska _ engelska _ ryska
linkkiArbets- och näringsministeriet:
Erkännande av examenfinska _ svenska _ engelska
linkkiUtbildningsstyrelsen:
Reglerade yrkenfinska _ svenska _ engelska
linkkiUtbildningsstyrelsen:
Utlåtanden om utländska yrkesexamenfinska _ svenska _ engelska
Yrkesinriktad arbetskraftsutbildning hjälper dig att få arbete.
Du kan lära dig nya färdigheter eller till och med ett nytt yrke.
Utbildningen kan också handleda dig i jobbsökningen.
Yrkesinriktad arbetskraftsutbildning är kostnadsfri.
Arbets- och näringsbyrån (TE-toimisto) ordnar den yrkesinriktade arbetskraftsutbildningen.
Du får arbetslöshetsförmån under utbildningstiden.
För vem är yrkesinriktad arbetskraftsutbildning avsedd?
Du kan delta i yrkesinriktad arbetskraftsutbildning, om
du har fyllt 20 år
du är arbetslös eller kommer att bli arbetslös
du har rätt att använda arbets- och näringsbyråns tjänster.
Du har rätt att använda arbets- och näringsbyråns tjänster om du har fått kontinuerligt uppehållstillstånd (A) eller permanent uppehållstillstånd (P).
linkkiArbets- och näringsministeriet:
Yrkesinriktad arbetskraftsutbildningfinska _ svenska _ engelska
Info om arbetskraftsutbildningfinska _ svenska
Hur ansöker jag till yrkesinriktad arbetskraftsutbildning?
Du ansöker till yrkesinriktad arbetskraftsutbildning antingen i arbets- och näringsbyrån eller med en elektronisk blankett på internet.
I ansökningen ska du motivera varför du borde antas till utbildningen.
Överväg din motivering noga.
Motiveringen påverkar antagningen.
Arbets- och näringsbyrån väljer studerandena till den yrkesinriktade arbetskraftsutbildningen.
Vad kan jag studera i yrkesinriktad arbetskraftsutbildning?
Innehållet i yrkesinriktad arbetskraftsutbildning varierar mycket.
Nedan följer några exempel på yrkesinriktad arbetskraftsutbildning:
Du kan lära dig ett nytt yrke eller en ny examensdel.
Du kan studera finska eller svenska.
Du kan få handledning i jobbsökningen.
Du kan få fortbildning eller påbyggnadsutbildning i din egen bransch.
Du kan få handledning i företagande eller företagarutbildning.
linkkiArbets- och näringsministeriet:
Arbets- och näringsbyrån köper den yrkesinriktade arbetskraftsutbildningen av olika läroanstalter och företag.
Du studerar alltså inte vid arbets- och näringsbyrån utan vid den läroanstalt som ordnar kursen.
Arbets- och näringsbyrån genomför utbildningar även tillsammans med arbetsgivare.
Vissa läroanstalter ordnar yrkesinriktad arbetskraftsutbildning särskilt för invandrare.
Utbildningen kan vara till exempel studier i finska eller yrkesutbildning.
På vissa kurser kan du skaffa dig behörighet att utöva ditt yrke i Finland.
Till exempel sjukskötare måste avlägga ytterligare studier för att få arbeta som sjukskötare i Finland.
Läs mer på InfoFinlands sida Utländska examina i Finland.
Ekonomiskt stöd under den yrkesinriktade arbetskraftsutbildningen
Under den yrkesinriktade arbetskraftsutbildningen får du samma förmån som när du är arbetslös.
Om du har avtalat om yrkesinriktad arbetskraftsutbildning i din sysselsättningsplan, kan du få förhöjd arbetslöshetsförmån.
Det betyder att du får lite mer pengar i din arbetslöshetsförmån.
Beslut om utbetalning av förhöjningsdelen fattas av den som betalar arbetslöshetsförmånen, alltså arbetslöshetskassan eller FPA.
Du kan även få kostnadsersättning för resekostnader för de dagar som du deltar i utbildningen.
Om den som betalar din arbetslöshetsförmån inte betalar ut kostnadsersättning, kan arbets- och näringsbyrån i vissa fall betala den.
FPA:s kostnadsersättningfinska _ svenska _ engelska
Frivillig utbildning med arbetslöshetsförmån
Du kan även få arbetslöshetsförmån under andra studier om arbets- och näringsbyrån bedömer att du behöver utbildningen.
Arbets- och näringsbyrån skaffar inte utbildningen och väljer inte studeranden till utbildningen såsom i arbetskraftsutbildning.
Du ansöker om studieplats direkt vid läroanstalten.
Du måste avtala om utbildningen med arbets- och näringsbyrån innan du inleder utbildningen.
Du kan få arbetslöshetsförmån under studierna, om
du har anmält dig som arbetssökande vid arbets- och näringsbyrån och din jobbsökning är i kraft
du är minst 25 år gammal
arbets- och näringsbyrån bedömer att utbildningen främjar din yrkeskunnighet eller hjälper dig att få ett jobb
du har avtalat om utbildningen i din sysselsättningsplan med arbets- och näringsbyrån.
För vilka studier kan man få arbetslöshetsförmån?
Med arbetslöshetsförmånen understöds bara heltidsstudier.
Som heltidsstudier räknas följande:
högskoleexamen gymnasiestudier eller
studier, vars omfattning motsvarar heltidsstudier, till exempel fem studiepoäng i månaden eller 25 studietimmar i veckan.
Studierna ska leda till
yrkesinriktade grundexamen, yrkesexamen eller specialyrkesexamen
lägre eller högre högskoleexamen vid universitet eller högskola
avläggande av delar av ovan nämnda examina.
Studierna kan även vara tilläggsutbildning eller påbyggnadsutbildning alternativt studier vid universitet eller yrkeshögskola.
linkkiArbets- och näringsministeriet:
Frivilliga studier med stöd av arbetslöshetsförmånfinska _ svenska _ engelska
Du kan studera i Finland som utbytesstudent eller avlägga hela examen här.
Om du vill hitta arbete i Finland är det viktigt att du studerar finska eller svenska.
I Finland är det ofta svårt att hitta arbete om man inte kan finska eller svenska.
Utbytesstudenter
Du kan komma till Finland som utbytesstudent.
Du kan avlägga utbytesstudier via olika program.
Utbytesstudenter kan få studieplats till exempel via Erasmus, Nordplus, FIRST och Fulbright.
Du kan också studera som utbytesstudent på egen hand.
Om du vill komma till Finland som utbytesstudent ska du ta kontakt med enheten för internationella ärenden eller till exempel studiebyrån i din egen läroanstalt.
Komihåglista för nya studerande
Säkerställ att du har följande när du kommer till Finland för att studera:
uppehållstillstånd
försäkring
pengar
studieplats
bostad
Ansökan för examensstuderande
Du kan söka till en yrkeshögskola eller ett universitet i den gemensamma ansökan till högskolor.
Läs mer på InfoFinlands sida Ansökan till utbildning.
Du hittar mer information om yrkeshögskolor på InfoFinlands sida Yrkeshögskolor.
Läs mer om högskolor på InfoFinlands sida Universitet.
Du kan också avlägga fortsatta studier vid universitet eller yrkeshögskola i Finland.
Läs mer om fortsatta studier på InfoFinlands sidor Universitet och Yrkeshögskolor.
Uppehållstillstånd
När du kommer till Finland för att studera beror behovet av uppehållstillstånd på ditt medborgarskap.
Läs mer på InfoFinlands sida Studerande.
Finansiering av studierna
Utländska studerande får vanligen inget studiestöd.
För att få ett uppehållstillstånd för studerande, ska du kunna visa att din ekonomiska situation ger dig möjlighet att leva i Finland.
Penningunderstöd och stipendier
Utländska studerande kan ansöka om olika penningunderstöd för finländska högskolor.
Alla finländska högskolor har ett eget stipendiesystem för de studerande som kommer från länder utanför EU/EES-området och som har godkänts för att avlägga en kandidat- eller magisterexamen på engelska.
Möjligheten till ett stipendium kan till exempel bero på hur framgångsrik du varit i dina studier.
Stipendiet kan täcka hela läsårsavgiften eller en del av den.
Vissa stipendier kan även täcka andra kostnader.
Ibland krävs att du lyckas tillräckligt bra med dina studier för att du ska få ett stipendium.
Du kan vanligtvis ansöka om ett stipendium samtidigt som du ansöker om en studieplats.
Det finns också särskilda Erasmus Mundus-magisterprogram som har ett eget stipendiesystem.
Utbildningsstyrelsen har stipendieprogram för forskarstuderande som kommer till Finland för att avlägga doktorsexamen.
Studerande från USA kan ansöka om ett Fulbright-stipendium.
Läs mer om stipendier och penningunderstöd på webbplatsen Studyinfinland.fi.
Boende, arbete och försäkring
Det kan vara svårt att hitta en bostad eftersom efterfrågan på bostäder är större än utbudet speciellt i större städer.
Sök en bostad i god tid innan du flyttar till Finland
Du kan hyra en bostad på den öppna marknaden.
Du kan också söka bostad via föreningen Suomen Opiskelija-asunto (Suomen Opiskelija-asunto) (SOA).
Det är dyrt att bo i Finland.
Studentbostäderna är oftast billigare än bostäderna på den öppna marknaden.
Om du arbetar vid sidan av studierna är din arbetstid begränsad.
Vanligen kan du arbeta högst 25 timmar i veckan.
Detta beror dock på vilket land du kommer ifrån.
Läs mer på InfoFinlands sida Studerande.
Du kan också göra ditt slutarbete i något företag eller göra en arbetspraktik.
I dessa har arbetstiden inte begränsats.
Se till att du har försäkringar.
Hur omfattande försäkring du behöver beror på vilket land du kommer ifrån och hur länge dina studier pågår.
Det är mycket viktigt att din försäkring är i kraft hela den tid som du vistas i Finland.
Läs mer på InfoFinlands sida Studerande.
Studier i Finland
Om du inte är medborgare i ett EU-land eller EES-land och inte heller familjemedlem till en medborgare i ett sådant land och du kommer till Finland för att studera i augusti 2017 eller senare, måste du betala terminsavgift för studierna.
Avgiften gäller lägre och högre högskolestudier på engelska.
I Finland kan du studera på finska, svenska och ibland även på engelska.
Högskolorna har vissa utbildningsprogram där undervisningen ges på engelska.
Merparten av studierna är dock på finska eller på svenska.
I Finland finns många aktiva studentorganisationer.
De ordnar verksamhet även för utländska studerande.
I studentorganisationerna lär du dig känna nya människor.
Om du vill hitta en arbetsplats i Finland ska du studera finska eller svenska.
Även om du klarar dig i många dagliga situationer på engelska kräver de flesta arbetsgivare att du kan finska eller svenska.
Läs mer på InfoFinlands sida Finska och svenska språket.
Om inte hinner studera finska vid din egen läroanstalt, finns det kurser i finska vid många andra läroanstalter.
Du kan även studera språket på Internet.
Läs mer på InfoFinlands sida Finska och svenska språket.
Det är också viktigt att du bekantar dig med finländare och arbetslivet i Finland redan under studietiden.
På så sätt hittar du lättare vänner och ett arbete.
Till exempel arbetspraktik (työharjoittelu), hobbyer och organisationer är bra sätt att lära känna det finländska samhället.
Information för utländska studerandeengelska
Information om utbytesprogrammetengelska
Gymnasieansökan
Sök till gymnasiet i den gemensamma ansökan till andra stadiet i februari-mars.
Du kan söka till ett gymnasium om du har avlagt lärokursen för den grundläggande utbildningen eller en lärokurs som motsvarar den grundläggande utbildningen.
Fyll ansökan i tjänsten Studieinfo.fi.
Eleverna antas till gymnasiet utifrån vitsorden på avgångsbetyget från grundskolan.
Därtill ordnar vissa gymnasier inträdesprov.
Om du söker till ett vuxengymnasium, kontakta läroanstalten direkt.
Du kan inte söka till ett vuxengymnasium i den gemensamma ansökan.
När du söker till ett vuxengymnasium är inte medeltalet på ditt betyg av betydelse.
Du hittar utbildningar på Studieinfo.fi.
Om du vill förbättra dina kunskaper i finska innan du söker till ett gymnasium, kan du söka till en förberedande gymnasieutbildning
Läs mer på InfoFinlands sida Gymnasieförberedande utbildning.
Ansökan till gymnasium i den gemensamma ansökanfinska _ svenska
Ansökan till yrkesutbildning
Din grundutbildning avgör till hurudan yrkesutbildning du kan söka och på vilket sätt ansökan sker.
Du kan söka till en grundskolebaserad yrkesutbildning om du har avlagt lärokursen för den grundläggande utbildningen eller en lärokurs som motsvarar den grundläggande utbildningen.
Du kan söka till en gymnasiebaserad yrkesutbildning om du har gått färdigt gymnasiet.
Du kan söka till dessa utbildningar i den kontinuerliga ansökan året om eller i den gemensamma ansökan till andra stadiet.
I allmänhet ordnas den gemensamma ansökan i februari-mars.
Fyll ansökan i tjänsten Studieinfo.fi.
Om du redan har avlagt en yrkesexamen eller en högskoleexamen, kan du inte söka till en yrkesutbildning i den gemensamma ansökan.
Då kan du söka till utbildningen i den kontinuerliga ansökan.
Du ska söka till utbildningen i den kontinuerliga ansökan också om du är i arbetslivet och vill byta bransch eller om du vill ansöka till läroavtalsutbildning.
Du kan söka i den kontinuerliga ansökan även i det fall att du inte fick en studieplats i den gemensamma ansökan.
Grunderna för antagning av studeranden beror på utbildningen.
I allmänhet påverkas antagningen av antagningspoängen, som ges bl.a. utifrån dina betyg.
Inträdesprov eller lämplighetsprov ordnas också för många utbildningar.
I vissa branscher ställs krav på hälsotillståndet.
Läroanstalten kan kontrollera att du har tillräckliga språkkunskaper för studierna.
Fråga mer vid den läroanstalt som du ansöker till.
Om du vill ha mera kunskap och färdigheter innan du söker till en yrkesinriktad utbildning, kan du ansöka till VALMA-utbildningen.
Under VALMA-utbildningen kan du även förbättra dina språkkunskaper i finska.
Läs mera på InfoFinlands sida Utbildning som handleder för yrkesutbildning.
Om du behöver särskilt stöd i de yrkesinriktade studierna t.ex. på grund av handikapp eller inlärningssvårigheter ska du ansöka till utbildningen via ansökan till specialundervisning.
Ansökan till yrkesutbildning i den gemensamma ansökanfinska _ svenska
Kontinuerlig ansökan till yrkesutbildning finska _ svenska
Antagningsgrunder till yrkesutbildningfinska _ svenska
Om du har en utländsk examen
Om du har avlagt grundskolan eller gymnasiet utomlands, antas du till en yrkesutbildning enligt prövning.
Vid antagning enligt prövning beaktas
ditt utbildningsbehov
bedömningen av hur bra du kan klara av studierna.
Antagning enligt prövningfinska _ svenska
Ansökan till en yrkesinriktad vuxenutbildning
Du kan söka till en yrkesinriktad vuxenutbildning om du vill avlägga en examen vid sidan om arbetet.
I vuxenutbildningen avlägger du yrkesexamen som fristående examen.
Du kan söka till en yrkesinriktad vuxenutbildning också om du har avlagt en yrkesexamen eller en högskoleexamen.
När du söker till en yrkesinriktad vuxenutbildning, ska du ha en tillräckligt lång arbetserfarenhet.
Du kan inte söka till en yrkesinriktad vuxenutbildning i den gemensamma ansökan.
Ta reda på hur du kan söka till utbildningen i tjänsten Studieinfo.fi eller av läroanstalten.
Ofta är ansökningstiden fortlöpande.
Ansökan till en yrkeshögskola
Du kan söka till en yrkeshögskola för att avlägga en yrkeshögskoleexamen, då du har avlagt t.ex. någon av följande utbildningar:
gymnasiet
en yrkesexamen
studentexamen eller en motsvarande examen i ett annat land
Du får närmare uppgifter från tjänsten Studieinfo.fi.
Sök till en yrkeshögskola i den gemensamma ansökan till högskolor.
Den gemensamma ansökan ordnas två gånger per år, på våren och på hösten.
Fyll ansökan i tjänsten Studieinfo.fi.
Grunderna för antagning av studeranden beror på utbildningen.
Ditt betyg, inträdesprovet och din arbetserfarenhet kan påverka antagningen.
Också dina tidigare studier kan spela en roll.
Ansökan till YH-examenfinska _ svenska
Högre yrkeshögskoleexamina
Du kan söka till en YH-examen om du har
en lämplig yrkeshögskoleexamen eller en annan lämplig högskoleexamen och
minst tre års arbetserfarenhet från samma område som din examen och du har inhämtat din arbetserfarenhet efter att du har avlagt examen.
Sök till en YH-examen i den gemensamma ansökan till högskolor på våren eller hösten Till många utbildningar är det möjligt att söka endast på våren.
Fyll i ansökningsblanketten i tjänsten Studieinfo.fi.
Du kan söka till en högre YH-examen på ett främmande språk med en separat ansökan.
Du hittar ansökningsblanketter då du letar efter utbildningar i Studieinfo.fi.
Högre YH-examenfinska _ svenska
Ansökan till universitet
Ansök till ett universitet antingen i den gemensamma ansökan till högskolor eller med en separat ansökan till en viss utbildning.
Du kan söka till många universitetsutbildningar i den gemensamma ansökan till högskolor.
Den ordnas på våren och hösten.
Alternativen är fler på våren.
Den gemensamma ansökan till vissa utbildningar ordnas redan i januari.
Utred i tid när du kan söka.
Fyll ansökan i tjänsten Studieinfo.fi.
Du kan söka till ett universitet om du har avlagt t.ex. någon av följande examina:
en finländsk studentexamen
en minst treårig yrkesinriktad grundexamen
en utländsk examen, som ger möjlighet till universitetsstudier i det land där du avlagt examen
Granska av högskolans studiebyrå att det är möjligt att söka till ett universitet med din examen.
Du får närmare uppgifter också från tjänsten Studieinfo.fi.
När du söker till ett universitet, får du i allmänhet poäng utifrån studentexamen och inträdesprovet.
Det finns skäl att förbereda dig omsorgsfullt för inträdesprovet.
Till vissa utbildningsprogram antas endast en liten del av sökandena.
Vissa inträdesprov omfattar förhandsuppgifter.
Ansökan till universitetfinska _ svenska _ engelska
Separat ansökan
Ansökan till vissa universitetsstudier sker genom en separat ansökan.
Du ska söka med en separat ansökan t.ex.
om du söker till ett magisterprogram
om du flyttar från en högskola till en annan eller
om du har avlagt studier i ett öppet universitet och söker till ett universitet utifrån dessa studier.
Om du söker till ett utbildningsprogram där undervisningsspråket är ett annat än finska eller svenska, beror ansökningssättet på utbildningen.
Det lönar sig att söka till vissa utbildningar på främmande språk i den gemensamma ansökan i januari.
Du hittar närmare information i Studieinfo.fi.
Du kan också fråga direkt av högskolorna.
De separata ansökningarna kan ordnas under olika tidsperioder och ansökningsförfarandena kan avvika från varandra.
Du hittar de separata ansökningarna via tjänsten Studieinfo.fi.
Påbyggnadsexamen
Om du vill avlägga en påbyggnadsexamen vid ett universitet, kontakta universitetet direkt.
Mottagande av studieplats
Läroanstalten meddelar dig att du har antagits för studier med ett brev.
Om du har antagits, meddela så fort som möjligt till läroanstalten att du tar emot studieplatsen.
Brevet innehåller anvisningar om hur du tar emot platsen och hur du anmäler dig.
Om du inte tar emot platsen i tid, förlorar du den.
När du tar emot en studieplats, förbinder du dig att börja studera i läroanstalten.
Du kan söka till många olika läroanstalter i den gemensamma ansökan.
Du kan dock ta emot endast en studieplats.
Efter grundskolan (peruskoulu), d.v.s. efter grundstadiet fortsätter studerandena till läroanstalter på andra stadiet (toisen asteen oppilaitos).
Läroanstalter på andra stadiet är gymnasiet och yrkesläroanstalter.
Läs mer om yrkesläroanstalter på InfoFinlands sida Yrkesutbildning.
Gymnasiestudierna är mer teoretiskt inriktade än yrkesutbildning.
Studierna är allmänbildande: fokus ligger speciellt på naturvetenskapliga och humanistiska ämnen.
I vissa gymnasier ges även mycket undervisning i konstämnen.
Vissa gymnasier är specialgymnasier.
De är inriktade på till exempel musik, idrott eller naturvetenskaper.
Specialgymnasierna är mycket populära.
Det kan vara svårt att komma in dit.
Gymnasiet ger förberedande utbildning till exempel för yrkeshögskola och universitet.
Både ungdomar och vuxna kan studera vid gymnasiet.
Ungdomarna studerar vid daggymnasiet (päivälukio) eller distansgymnasiet (etälukio), vuxna studerar ofta vid vuxengymnasiet (aikuislukio).
Information om gymnasiestudierfinska _ svenska
linkkiFörbund för gymnasieelever:
Förbund för gymnasieeleverfinska _ svenska _ engelska
linkkiUtbildningsstyrelsen:
Information om gymnasiestudierfinska _ svenska _ engelska
Att söka till gymnasiet
Sök till gymnasiet i den gemensamma ansökan till andra stadiet.
Om du vill studera vid ett vuxengymnasium ska du ta kontakt direkt med läroanstalten.
Läs mer på InfoFinlands sida Ansökan till utbildning.
Gemensam ansökan till gymnasier och yrkesläroanstalterfinska _ svenska
Att studera vid gymnasiet
Gymnasiestudierna pågår vanligen tre år.
Gymnasiet kan också avläggas på två eller fyra år.
I gymnasiestudierna har du många valmöjligheter.
Utöver de obligatoriska kurserna kan du välja många kurser som passar dig.
I gymnasiet påverkar du själv innehållet i dina studier och din studietakt.
I gymnasiet tas inga terminsavgifter ut.
Utbildningen kostar alltså inget.
Du måste dock själv skaffa gymnasieböckerna.
Böckerna är ofta dyra.
Man kan även köpa gymnasieböckerna begagnade.
Du måste även skaffa dig en bärbar dator.
Om du till exempel har en krävande hobby eller är sjuk en lång tid kan du avlägga gymnasiet som distansstudier.
Fråga mer om distansstudier vid ditt eget gymnasium.
Studentexamen
Gymnasiestudierna siktar till studentexamen (ylioppilastutkinto).
Studentexamen består av prov i olika läroämnen.
Studentskrivningarna (ylioppilaskokeet) skrivs oftast i slutet av studierna.
Modersmålsprovet är ett obligatoriskt prov i studentexamen.
Modersmålsprovet kan skrivas i finska, svenska eller samiska.
Om du inte har finska, svenska eller samiska som modersmål kan du skriva ett prov i finska eller svenska som andra språk.
Utöver modersmålsprovet måste du skriva prov i minst tre andra ämnen.
Om du vill kan du även skriva fler ämnen.
Utöver modersmålsprovet kan du skriva prov i följande andra ämnen:
Det andra inhemska språket (finska eller svenska)
Ett främmande språk: engelska, tyska, ryska, franska, spanska, portugisiska, latin
Matematik
Realämnen (reaali), d.v.s. historia, religion, fysik, kemi, biologi, psykologi, filosofi
Studentskrivningarna ordnas på våren och på hösten.
Om du vill kan du skriva några ämnen på hösten och resten på våren.
Du måste skriva alla prov på högst tre efter varandra följande examenstillfällen.
Info om studentexamenfinska _ svenska
linkkiStudentexamensnämnden:
Information om studentexamenfinska _ svenska _ engelska _ franska _ tyska
Vuxengymnasium
Vuxengymnasiet är i huvudsak avsett för personer som har fyllt 18 år.
Vid vuxengymnasiet är studierna flexibla.
Du kan avlägga hela studentexamen eller bara studera ett ämne.
Undervisningen sker oftast kvällstid.
Många vuxengymnasier erbjuder finskakurser för invandrare.
Fråga om kurserna direkt vid vuxengymnasiet.
Information om vuxengymnasietfinska _ svenska
Din situation avgör hur du kan finansiera dina studier i Finland.
På den här sidan berättar vi om FPA:s stöd till studerande samt om penningunderstöd och stipendier.
Studiestöd
Du kan få FPA:s studiestöd (opintotuki) om du
har det uppehållstillstånd (oleskelulupa) som krävs och
vistas i Finland av någon annan orsak än studier.
Om du flyttar till Finland för att studera kan du inte få studiestöd.
Till exempel utbytesstuderande får inte finskt studiestöd.
Studiestödet består av studiepenning och statsborgen för studielån.
Du kan få studiestöd om
Du studerar i gymnasiet
Du studerar vid en yrkesläroanstalt eller avlägger yrkesinriktade tilläggsstudier
Du studerar vid en högskola.
Du kan få studiepenning om du har fyllt 17 år.
Du måste studera på heltid.
Med heltidsstudier avses att studierna är din huvudsyssla.
Du kan arbeta vid sidan av studierna.
Lönen som du får för ditt arbete kan minska ditt studiestöd.
Du ansöker om studiepenning och statsgaranti för studielån vid FPA.
FPA betalar in studiepenningen på ditt konto månatligen.
På studiepenningens belopp inverkar många omständigheter.
På studiepenningens belopp inverkar bland annat stödmottagarens ålder, om hen bor i sitt eget hem eller hos en förälder, on hen är gift och om hen har minderåriga barn. Kontrollera storleken på din studiepenning på FPA:s webbplats eller vid en FPA-byrå.
Det är inte obligatoriskt att ta studielån.
Du kan högst ta ut ett visst maximibelopp.
Du väljer själv hur mycket studielån du vill ta.
Studielånet är ett lån som finska staten ger garanti för åt studeranden.
Du ansöker om lånet i banken när du har fått FPA:s beslut om statsgaranti.
Du måste betala tillbaka lånet när du har slutfört dina studier.
Du kan få studielån också när du fortbildar dig (täydennyskoulutus) som vuxen.
Dessutom kan du få vuxenutbildningsstöd (aikuiskoulutustuki).
I vissa fall kan du också få bostadstillägg, till exempel om du studerar på en avgiftsbelagd linje vid en folkhögskola och bor på läroanstaltens internat.
Läs mer på FPA:s webbplats.
På InfoFinlands sida Bostadsbidrag finns mer information om FPA:s allmänna bostadsbidrag.
Information om studiestödetfinska _ svenska _ engelska
Information om studiestödetengelska _ ryska _ estniska _ samiska
Information om att ansöka studiestödfinska _ svenska _ engelska
Studiestöd till utländska studerandefinska _ svenska _ engelska
Stöd för skolresor
Du kan få stöd för skolresor (koulumatkatuki) om du bor i Finland och studerar i gymnasiet eller vid en yrkesläroanstalt.
Din skolresa måste vara minst 10 kilometer lång och resekostnaderna måste överstiga 54 euro per månad.
Information om skolresestödetfinska _ svenska _ engelska
Måltidsstöd
Om du studerar vid en högskola får du också måltidsstöd (ateriatuki).
Du kan få måltidsstödet endast i läroanstalternas egna restauranger.
Detta innebär att studeranden betalar mindre för måltiderna än andra som besöker restaurangen.
Du behöver inte ansöka separat om måltidsstödet.
Du behöver bara visa upp ditt studentkort när du betalar för måltiden.
Du har inte rätt till måltidsstöd om du är i Finland endast på arbetspraktik (työharjoittelu) som ingår i en utländsk examen.
Information om måltidsstödetfinska _ svenska _ engelska
Penningunderstöd och stipendier
Utländska studerande kan ansöka om olika penningunderstöd för finländska högskolor.
Alla finländska högskolor har ett eget stipendiesystem för de studerande som kommer från länder utanför EU/EES-området och som har godkänts för att avlägga en kandidat- eller magisterexamen på engelska.
Möjligheten till ett stipendium kan till exempel bero på hur framgångsrik du varit i dina studier.
Stipendiet kan täcka hela läsårsavgiften eller en del av den.
Vissa stipendier kan även täcka andra kostnader.
Ibland krävs att du lyckas tillräckligt bra med dina studier för att du ska få ett stipendium.
Du kan vanligtvis ansöka om ett stipendium samtidigt som du ansöker om en studieplats.
Det finns också särskilda Erasmus Mundus-magisterprogram som har ett eget stipendiesystem.
Utbildningsstyrelsen har stipendieprogram för forskarstuderande som kommer till Finland för att avlägga doktorsexamen.
Studerande från USA kan ansöka om ett Fulbright-stipendium.
Läs mer om stipendier och penningunderstöd på webbplatsen Studyinfinland.fi.
I Finland kan man avlägga högskolestudier både vid yrkeshögskolor och vid universitet.
Läs mer om yrkeshögskolan på InfoFinlands sida Yrkeshögskolor.
Ansök om studieplats
Du kan söka till ett universitet om du har avlagt en finländsk studentexamen, en utländsk examen som motsvarar studentexamen eller en yrkesinriktad slutexamen. Sök till ett universitet i den gemensamma ansökan till högskolor.
Läs mer på InfoFinlands sida Ansökan till utbildning.
Gemensam ansökan till universitetfinska _ svenska
Vilka yrken kan studera till?
Vid universitet kan man studera i många olika studieområden.
De som har utexaminerats från en högskola eller ett universitet arbetar i många slags arbetsuppgifter.
En del universitetsstudier leder direkt till ett yrke.
Sådana yrken är till exempel:
lärare
jurist
läkare
skådespelare
diplomingenjör
bildkonstnär
Andra universitetsstudier leder inte till ett visst yrke.
Till exempel studerande vid den samhällsvetenskapliga eller den humanistiska fakulteten utexamineras inte nödvändigtvis till ett yrke.
Dessa människor arbetar till exempel i följande arbetsuppgifter:
forskare
statlig tjänsteman
Studier vid universitet
Vid vissa universitet har olika examen olika namn.
Till exempel är tekniska högskolors motsvarighet till magisterexamen diplomingenjörsexamen (diplomi-insinööri).
När du får en studieplats får du rättighet att avlägga båda examina.
Du kan också avsluta studierna efter lägre högskoleexamen.
Kandidatstudierna pågår ungefär tre år, magisterstudierna ungefär två år.
Hur fort studierna framskrider beror på dig själv.
Du kan också söka till ett separat magisterprogram.
Magisterprogrammet är ett studieprogram som leder till högre högskoleexamen.
För att kunna studera i ett magisterprogram ska du ha avlagt lägre högskoleexamen.
Magisterprogrammen pågår i cirka två år.
Vid dem studerar ofta människor från många olika vetenskapsområden.
Utexaminering från universitetet
När du är klar med dina studier får du antingen kandidatexamen eller magisterexamen.
Om du vill kan du efter magisterexamen söka till fortsatta studier.
Information om högskolestudierfinska _ svenska _ engelska
linkkiFinlands Studentkårers Förbund:
Information om studentkårer i Finlandfinska _ svenska _ engelska
Öppna universitet
De öppna universiteten tillhandahåller universitetskurser.
Vem som helst kan studera vid ett öppet universitet.
Du kan studera vid ett öppet universitet även om du inte har någon examen.
Läs mer på InfoFinlands sida Studier som hobby.
Vetenskaplig fortbildning vid universitet
Vetenskaplig fortbildning vid universitet är examensinriktad fortbildning.
Sådan utbildning förbereder dig till exempel för forskaryrket.
Vid universitetet kan du avlägga licentiatexamen (lisensiaatti) eller doktorsexamen (tohtori).
De flesta studerande som bedriver fortsatta studier avlägger doktorsexamen.
Man kan ansöka till fortsatta studier vid universitet några gånger per år.
Universitet och institutioner har olika ansökningstider.
Kontrollera ansökningstiden vid den institution där du vill bedriva fortsatta studier.
I Finland måste de som bedriver fortsatta studier ofta finansiera studierna själva.
Du kan ansöka om stipendier hos olika stiftelser (säätiö).
Påbyggnadsexamina vid universitetfinska
linkkiStiftelsetjänst:
Information om stiftelser och penningunderstödfinska _ svenska _ engelska
linkkiCIMO:
Penningunderstöd för utländska forskarefinska _ svenska _ engelska
Vägledning i högskolestudier
Vid högskolornas SIMHE-tjänster kan du söka hjälp och information om högskoleutbildning i Finland och om hur du ansöker till högskoleutbildning.
Du kan även få information om andra utbildningsmöjligheter för personer som avlagt högskolestudier.
Du kan få vägledning via SIMHE-tjänsterna om
du har flyttat till Finland
du är intresserad av högskolestudier och
du har avlagt högskolestudier eller högskoleexamen utomlands.
Vägledning kan ges individuellt eller i grupp.
linkkiUtbildningsstyrelsen:
Högskolor som erbjuder SIMHE-tjänsterfinska _ svenska _ engelska
Utbildning som handleder för grundläggande yrkesutbildning (Ammatilliseen peruskoulutukseen valmentava koulutus) d.v.s. VALMA är avsedd för dem som vill avlägga en grundläggande yrkesutbildning.
Under VALMA-utbildningen får du kunskap och färdigheter som hjälper dig i dina senare yrkesinriktade studier.
Du kan även förbättra din språkkunskap. Du kan också höja dina grundskolebetyg.
VALMA-utbildningen räcker ungefär ett läsår.
Du kan under utbildningen bekanta dig med olika branscher och fundera på vad du vill studera.
Du besöker arbetsplatser och deltar i verkstäder.
I början av utbildningen görs det upp en personlig studieplan för dig.
I den skrivs det in vilka studier du avlägger och hur.
Du får ett betyg för VALMA-utbildningen.
Du får också tilläggspoäng när du ansöker till en yrkesutbildning i den gemensamma ansökan.
VALMA-utbildningen kostar vanligen inget för den studerande.
Information om VALMA-utbildningarfinska _ svenska _ engelska
Ansökan till VALMA-utbildningen
Du kan ansöka till VALMA-utbildningen om du har slutfört grundskolan eller en utbildning som motsvarar grundskolan.
Om läroinrättningen anser att du kan klara av studierna kan du antas som studerande även utan slutbetyg från grundskolan.
Ansök till VALMA-utbildningen efter den egentliga gemensamma ansökan i början av sommaren.
Om du behöver särskilt stöd t.ex. på grund av handikapp ska du ansöka till utbildningen på våren, under ansökan till specialundervisning.
Närmare information om ansökningstiderna hittar du via Studieinfo.fi-tjänsten.
Fyll i ansökningsblanketten i Studieinfo.fi-tjänsten.
Ansökan till VALMA-utbildningfinska _ svenska
Ansökan till specialundervisningfinska _ svenska
Studierna är inte alltid inriktade på att skaffa ett yrke.
Du kan också ha studier som hobby.
Du kan studera vid flera olika läroanstalter: öppna universitetet (avoin yliopisto) eller öppna yrkeshögskolan (avoin ammattikorkeakoulu), sommaruniversitetet (kesäyliopisto), senioruniversitetet (ikäihmisten yliopisto), medborgarinstitut (kansalaisopisto), arbetarinstitut (työväenopisto) och folkhögskolor (kansanopisto).
Studierna är vanligen avgiftsbelagda.
Många av dessa läroanstalter tillhandahåller undervisning i finska och svenska för invandrare.
Läs mer på InfoFinlands sida Finska och svenska språket.
Du kan även studera flera andra språk, såsom engelska eller franska.
Vid folkhögskolor kan du även avlägga yrkesexamen.
Öppna universitetet och öppna yrkeshögskolan
Öppna universitetet (avoin yliopisto) och öppna yrkeshögskolan (avoin ammattikorkeakoulu) ordnar universitets- och yrkeshögskolekurser.
Vem som helst kan studera vid de öppna högskolorna.
Du kan studera vid öppna högskolor fastän du inte har någon examen.
Du kan studera vid öppna högskolor
om du vill studera som hobby
om du vill bli antagen för studier i ett visst ämne vid en högskola
när du vill utöka din yrkeskunnighet och dina kunskaper
Till de öppna högskolorna ordnas inga inträdesprov.
Du kan anmäla dig till vårens kurser i början av året och till höstens kurser i slutet av sommaren.
Anmäl dig direkt till kurserna.
Du kan välja enskilda kurser eller större studiehelheter.
Vid öppna högskolor är studierna flexibla.
Du kan delta i kurser under dagtid, på kvällar eller på veckoslut.
Du kan också studera på internet.
Studierna vid öppna högskolor är inte heltidsstudier.
Du får därför inget studiestöd (opintotuki) och inga studentrabatter när du studerar vid öppna högskolan.
Du kan avlägga studier vid öppna högskolan fastän du får arbetslöshetsersättning (työttömyyskorvaus).
Du har nytta av studierna vid öppna högskolan när du studerar vidare. Om du blir antagen till yrkeshögskolan behöver du inte avlägga de kurser som du redan har avlagt vid öppna yrkeshögskolan.
Om du har studerat vid öppna universitetet och söker till universitetet ansöker du via separat ansökan (erillinen haku).
Information om öppna yrkeshögskolanfinska _ svenska
Information om öppna universitetetfinska _ svenska
Sommaruniversitetet
Kurserna vid sommaruniversitetet (kesäyliopisto) påminner mycket om kurserna vid öppna universitetet.
Man kan studera vid sommaruniversitetet även under andra tider än på sommaren.
Utöver universitetskurser ordnar sommaruniversiteten också annan undervisning, till exempel:
Yrkesinriktad fortbildning (täydennyskoulutus)
Arbetskraftsutbildning (työvoimakoulutus)
Abiturientkurser (abikurssi) för gymnasieelever som förbereder sig för studentskrivningarna
finskakurser för invandrare
Fråga närmare uppgifter om undervisningen vid närmaste sommaruniversitet.
Info om sommaruniversitetfinska _ svenska
Information om sommaruniversitetetfinska _ svenska _ engelska
Senioruniversitetet
Senioruniversitetet (ikäihmisten yliopisto) är avsett för dem som har fyllt 60 år.
Studietillfällena är dock öppna för alla.
Undervisningen vid senioruniversitetet är en del av öppna universitetets verksamhet.
Senioruniversitetet ordnar föreläsningsserier, kurser och studieresor.
Fråga mer om senioruniversitetet i kansliet för närmaste öppna universitet.
Medborgarinstitut och arbetarinstitut
I Finland finns många medborgarinstitut (kansalaisopisto) och arbetarinstitut (työväenopisto).
Vid dem kan du studera bland annat språk, handarbete, idrott, bildkonst och matlagning.
Medborgarinstituten och arbetarinstituten erbjuder hobbystudier.
Vid dem kan man inte avlägga yrkesinriktade studier.
Medborgarinstituten och arbetarinstituten ordnar finskakurser för invandrare.
Fråga närmare uppgifter om kurserna vid närmaste medborgarinstitut eller arbetarinstitut.
Ansökningspraxis varierar.
Vanligen ansöker man till vårens undervisning i början av året och till höstens undervisning på sensommaren.
Fråga om ansökningstiderna vid medborgarinstitutets eller arbetarinstitutets studiebyrå.
Info om medborgarinstituten och arbetarinstitutenfinska _ svenska
Medborgarinstitut i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Folkhögskolor
Folkhögskolorna (kansanopisto) erbjuder både hobbystudier och yrkesinriktad utbildning.
Folkhögskolan kan drivas av en organisation eller också kan de vara självständiga institut.
Vid folkhögskolan kan du utbilda dig till ett yrke.
Vid folkhögskolan kan man till exempel avlägga djurskötarexamen eller massörexamen.
Folkhögskolorna ordnar mycket undervisning för invandrare.
Vid folkhögskolan kan du studera finska eller delta i förberedande utbildning.
Folkhögskolorna ordnar vanligen två olika slags undervisning, kortkurser (lyhytkurssi) och långa utbildningslinjer (pitkä opintolinja).
Kortkurserna är öppna för alla och till dem behöver du inte söka.
Det räcker med att du anmäler dig.
De långa utbildningslinjerna är ofta yrkesinriktade studier.
De pågår vanligen från ett halvår till ett år.
Till de långa utbildningslinjerna måste man söka separat.
Folkhögskolornas ansökningspraxis och ansökningstider varierar.
Fråga mer om antagningen vid folkhögskolans studiebyrå.
Info om folkhögskolorfinska _ svenska
linkkiFinlands folkhögskolförening:
Information om folkhögskolorfinska
linkkiFinlands folkhögskolförening:
Kurser vid folkhögskolor för invandrarefinska
linkkiDövas folkhögskola:
Utbildning för döva invandrarefinska _ svenska _ engelska
Studierna vid en yrkeshögskola (ammattikorkeakoulu) är praktiskt inriktade.
När du utexamineras från en yrkeshögskola får du ofta ett yrke.
Vid yrkeshögskolorna studerar du på finska, svenska eller på engelska.
Vid många yrkeshögskolor finns engelskspråkiga utbildningsprogram.
Ansökan
Du kan söka till en yrkeshögskola då du har avlagt en yrkesskola, gymnasiet eller studentexamen i Finland eller i ett annat land.
Läs mer på InfoFinlands sida Ansökan till utbildning.
Gemensam ansökan till yrkeshögskolorfinska _ svenska
Studier
I yrkeshögskolor kan du studera inom många områden.
Inom parentes anges exempel på yrken som du studera till i olika studieområden:
Naturbruk- och miljöområdet (skogsbruksingenjör, landskapsplanerare)
Den humanistiska och pedagogiska branschen (teckenspråkstolk)
Kulturbranschen (musiker, inredningsarkitekt)
Turism- och kosthållsbranschen (hovmästare, hotellmedarbetare)
Social-, hälso- och idrottsområdet (barnmorska, fysioterapeut, sjuksköterska)
Samhällsvetenskaper, affärsekonomi och förvaltning (försäljningsförhandlare, marknadsföringsassistent)
Teknik och trafik (ingenjör inom bilteknik, maskinmästare i sjöfartsbranschen)
Heltidsstudierna pågår ungefär fyra år.
Studietiden beror på utbildningsprogrammet och din egen studietakt.
Studierna omfattar mycket praktiska övningar.
Studierna omfattar också en arbetspraktik.
Grundläggande information om yrkeshögskolorfinska _ svenska
linkkiUndervisnings- och kulturministeriet:
Förteckning över yrkeshögskolorfinska _ svenska
linkkiSAMOK:
Förbund för studerande vid yrkeshögskolorfinska _ svenska
Förberedande utbildning för invandrare
Yrkeshögskolan kan ordna avgiftsfri utbildning för invandrare med målet att ge den studerande tillräckliga språkkunskaper och andra färdigheter som behövs för att studera vid yrkeshögskolan.
Under studierna tränar studeranden sig i det finska språket, på att läsa saktexter och på sina studiefärdigheter.
Dessutom får studerandena information om utbildningsområdet, arbetsmöjligheter och studier som leder till examen.
Språkkunkapskravet för dem som söker till förberedande utbildning är oftast finskakunskaper på nivån B1 eller B2.
Öppna yrkeshögskolor
De öppna yrkeshögskolorna tillhandahåller yrkeshögskolekurser.
Vem som helst kan studera vid en öppen högskola.
Du kan studera vid en öppen yrkeshögskola även om du inte har någon examen.
Läs mer på InfoFinlands sida Studier som hobby.
Fortsatta studier vid yrkeshögskolor
Om du vill fördjupa dina yrkeskunskaper kan du avlägga högre yrkeshögskoleexamen (ylempi ammattikorkeakoulututkinto).
Den är avsedd för personer som har examen till exempel från en yrkeshögskola och som redan arbetar.
Du kan ansöka till högre yrkeshögskolestudier om du har
någon annan högskoleexamen
minst tre års arbetserfarenhet från en lämplig bransch
Sök till högre yrkeshögskolestudier i den gemensamma ansökan.
Gemensam ansökan ordnas två gånger per år, på hösten och på våren.
Läs mer om den gemensamma ansökan på InfoFinlands sida Ansökan till utbildning.
Du avlägger en högre yrkeshögskoleexamen på ungefär ett eller ett och ett halvt år.
Studiernas omfattning är 60 eller 90 studiepoäng.
Genom högre högskoleexamen kan du fördjupa och utvidga dina kunskaper inom ditt eget yrkesområde.
Till exempel sjukskötare kan avlägga högre yrkeshögskoleexamen inom rehabilitering.
Du kan också välja att avlägga en engelskspråkig examen.
Information om högre yrkeshögskoleexamenfinska _ svenska
Vägledning i högskolestudier
Vid högskolornas SIMHE-tjänster kan du söka hjälp och information om högskoleutbildning i Finland och om hur du ansöker till högskoleutbildning.
Du kan även få information om andra utbildningsmöjligheter för personer som avlagt högskolestudier.
Du kan få vägledning via SIMHE-tjänsterna om
du har flyttat till Finland
du är intresserad av högskolestudier och
du har avlagt högskolestudier eller högskoleexamen utomlands.
Vägledning kan ges individuellt eller i grupp.
linkkiUtbildningsstyrelsen:
Högskolor som erbjuder SIMHE-tjänsterfinska _ svenska _ engelska
Yrkesutbildning ger den studerande behörighet till ett visst yrke.
Därför är utbildningen mycket praktikorienterad.
Du kan söka till en yrkesutbildning när du har avlagt lärokursen för den grundläggande utbildningen.
Även vuxna kan utbilda sig till ett nytt yrke eller komplettera sin kompetens.
Din grundutbildning avgör till hurudan yrkesutbildning du kan söka och på vilket sätt ansökan sker.
Om du har avlagt grundskolans lärokurs kan du ansöka till grundskolebaserad yrkesutbildning (peruskoulupohjainen ammatillinen koulutus).
Om du har avlagt gymnasiet kan du ansöka till gymnasiebaserad yrkesutbildning (lukiopohjainen ammatillinen koulutus).
Om du vill avlägga examen vid sidan av arbetet kan du ansöka till yrkesutbildning för vuxna (ammatillinen aikuiskoulutus).
Läs mer på InfoFinlands sida Ansökan till utbildning.
När du har avlagt yrkesinriktad grundexamen kan du söka dig till fortsatta studier antingen inom yrkesinriktad tilläggsutbildning, vid en yrkeshögskola eller vid ett universitet.
Grundläggande information om yrkesutbildningfinska _ svenska _ engelska
linkkiUtbildningsstyrelsen:
Ytterligare information om yrkesutbildningfinska _ svenska
Gemensam ansökan till gymnasier och yrkesläroanstalterfinska _ svenska
Antagning enligt prövningfinska _ svenska
Utbildningsområden i yrkesutbildningenfinska _ svenska
Förberedande för yrkesutbildning
Utbildning som handleder för grundläggande yrkesutbildning (Ammatilliseen peruskoulutukseen valmentava koulutus) d.v.s. VALMA är avsedd för dem som vill avlägga en grundläggande yrkesutbildning.
Under VALMA-utbildningen får du kunskap och färdigheter som hjälper dig i dina senare yrkesinriktade studier.
Du kan även förbättra din språkkunskap. Du kan också höja dina grundskolebetyg.
VALMA-utbildningen räcker ett läsår.
Läs mera på InfoFinlands sida Utbildning som handleder för yrkesutbildning.
Yrkesinriktad grundexamen
Yrkesutbildning ges av yrkesläroanstalter (ammatillinen oppilaitos), specialyrkesläroanstalter (erityisammattioppilaitos) och av vuxenläroanstalter (aikuisopisto).
Du kan avlägga en yrkesinriktad grundexamen antingen
Inom den grundläggande utbildningen (ungdomar och vuxenstuderande)
Som fristående examen (näyttötutkinto) (vuxenstuderande)
Genom läroavtalsutbildning (oppisopimuskoulutus) (ungdomar och vuxenstuderande)
En yrkesinriktad grundexamen ger dig den grundläggande kompetensen i ett visst yrke.
En grundskolebaserad utbildning varar i cirka tre år.
Du kan också studera vid en yrkesläroanstalt och ett gymnasium samtidigt.
Då kan du avlägga en dubbelexamen (kaksoistutkinto).
Vid yrkesskolorna finns många olika områden som du kan studera.
pedagogiska områden
humanistiska och konstnärliga områden
samhälleliga områden
handel och förvaltning
naturvetenskaper
databehandling och datakommunikation
tekniska områden
jord- och skogsbruksområden
hälso- och välbefinnandeområden
Personlig utvecklingsplan för kunnandet
För varje studerande upprättas en personlig utvecklingsplan för kunnandet (PUK).
I planen nedtecknas vilket kunnande du har förvärvat tidigare och fastställs vilka studier du ska avlägga.
Du kan avlägga studierna i egen takt och påvisa vad du kan i praktiska uppgifter på arbetsplatser.
Utbildningsavtal
Utbildningsavtalet är inlärning i arbetet.
Om du vill skaffa dig praktiska kunskaper på en arbetsplats, är ett utbildningsavtal ett bra alternativ för ett läroavtal.
För utbildningstiden betalas ingen lön.
Utbildningsavtalet kan även kombineras med läroavtal.
Yrkesutbildning efter gymnasiet
Om du har avlagt gymnasiet eller studentexamen, kan du söka till en gymnasiebaserad utbildning.
Då kan du inte söka till en grundskolebaserad yrkesutbildning.
Läs mer på InfoFinlands sida Ansökan till utbildning.
Yrkesutbildning för vuxna
Om du arbetar kan du avlägga en yrkesexamen flexibelt vid sidan om arbetet.
Yrkesutbildning för vuxna omfattar
yrkesinriktade grundexamina
yrkesexamina
specialyrkesexamina.
I utbildningen beaktas din tidigare utbildning och den kunskap som du inhämtat som arbetstagare eller företagare.
Du hittar närmare information om hur du kan söka till en yrkesinriktad vuxenutbildning på InfoFinlands sida Ansökan till utbildning.
Examen vid sidan av arbetet med läroavtal
Läroavtal (oppisopimus) innebär inlärning i arbetet.
Du arbetar på en arbetsplats inom din egen bransch och avlägger examen vid sidan av arbetet.
Genom läroavtalsutbildning kan du avlägga samma examen som vid yrkesläroanstalter.
Yrkesexamen (ammattitutkinto)
Specialyrkesexamen (erityisammattitutkinto)
För att kunna studera genom läroavtal måste du ha en arbetsplats.
Du måste hitta en arbetsgivare som vill anställa dig.
Du kan inte inleda din läroavtalsutbildning om du inte har en arbetsplats.
Arbets- och näringsbyrån (TE-toimisto) kan hjälpa dig att hitta ett jobb.
Läroavtalsplatsen kan också vara din nuvarande arbetsplats.
När du har en arbetsplats ska du kontakta läroavtalsbyrån (oppisopimustoimisto) i din region.
Du kan också kontakta en läroanstalt som tillhandahåller läroavtalsutbildning.
Läroavtalsutbildning ges till exempel vid många vuxenutbildningscentra (aikuiskoulutuskeskus).
Under läroavtalsutbildningen betalar arbetsgivaren dig en lön som motsvarar minst en praktikantlön.
Om din arbetsgivare inte betalar dig lön för den tid som du använder för teoretiska studier har du möjligtvis rätt att ansöka om dagpenning, reseersättning och familjebidrag om du omfattas av Den sociala tryggheten i Finland.
Fråga mer vid din läroanstalt.
Information om läroavtalsutbildningfinska _ svenska
Information om läroavtalsutbildningfinska
Kontaktuppgifter till läroavtalsbyråerfinska
linkkiUtbildningsstyrelsen:
Information om läroavtalsutbildningfinska
Intyg om yrkeskunskap med ett fristående yrkesprov
Du kan påvisa dina yrkeskunskaper med ett fristående yrkesprov.
Då utför du praktiska arbetsuppgifter i verkliga situationer på en arbetsplats.
Utbildningsanordnaren utser två bedömare som bedömer ditt kunnande.
linkkiUtbildningsstyrelsen:
Information om fristående yrkesprovfinska
Yrkesutbildning som anordnas av arbetsgivaren
En del arbetsgivare utbildar människor till arbeten hos dem.
Dessa arbetsgivare ger garanti om en arbetsplats.
Det betyder att den som avlägger utbildningen får en arbetsplats hos arbetsgivaren.
Du får alltså både yrkesutbildning och en arbetsplats.
Till exempel många trafikföretag och VR utbildar de personer som de anställer.
Yrkesinriktad arbetskraftsutbildning hjälper dig att få arbete.
Du kan lära dig nya färdigheter eller till och med ett nytt yrke.
Utbildningen kan också handleda dig i jobbsökningen.
Yrkesinriktad arbetskraftsutbildning är kostnadsfri.
Arbets- och näringsbyrån (TE-toimisto) ordnar den yrkesinriktade arbetskraftsutbildningen.
Du får arbetslöshetsförmån under utbildningstiden.
För vem är yrkesinriktad arbetskraftsutbildning avsedd?
Du kan delta i yrkesinriktad arbetskraftsutbildning, om
du har fyllt 20 år
du är arbetslös eller kommer att bli arbetslös
du har rätt att använda arbets- och näringsbyråns tjänster.
Du har rätt att använda arbets- och näringsbyråns tjänster om du har fått kontinuerligt uppehållstillstånd (A) eller permanent uppehållstillstånd (P).
linkkiArbets- och näringsministeriet:
Yrkesinriktad arbetskraftsutbildningfinska _ svenska _ engelska
Info om arbetskraftsutbildningfinska _ svenska
Hur ansöker jag till yrkesinriktad arbetskraftsutbildning?
Du ansöker till yrkesinriktad arbetskraftsutbildning antingen i arbets- och näringsbyrån eller med en elektronisk blankett på internet.
I ansökningen ska du motivera varför du borde antas till utbildningen.
Överväg din motivering noga.
Motiveringen påverkar antagningen.
Arbets- och näringsbyrån väljer studerandena till den yrkesinriktade arbetskraftsutbildningen.
Vad kan jag studera i yrkesinriktad arbetskraftsutbildning?
Innehållet i yrkesinriktad arbetskraftsutbildning varierar mycket.
Du kan lära dig ett nytt yrke eller en ny examensdel.
Du kan studera finska eller svenska.
Du kan få handledning i jobbsökningen.
Du kan få fortbildning eller påbyggnadsutbildning i din egen bransch.
Du kan få handledning i företagande eller företagarutbildning.
linkkiArbets- och näringsministeriet:
Sök arbetskraftsutbildningarfinska _ svenska
Hurdan är den yrkesinriktade arbetskraftsutbildningen?
Arbets- och näringsbyrån köper den yrkesinriktade arbetskraftsutbildningen av olika läroanstalter och företag.
Du studerar alltså inte vid arbets- och näringsbyrån utan vid den läroanstalt som ordnar kursen.
Arbets- och näringsbyrån genomför utbildningar även tillsammans med arbetsgivare.
Vissa läroanstalter ordnar yrkesinriktad arbetskraftsutbildning särskilt för invandrare.
Utbildningen kan vara till exempel studier i finska eller yrkesutbildning.
På vissa kurser kan du skaffa dig behörighet att utöva ditt yrke i Finland.
Till exempel sjukskötare måste avlägga ytterligare studier för att få arbeta som sjukskötare i Finland.
Läs mer på InfoFinlands sida Utländska examina i Finland.
Ekonomiskt stöd under den yrkesinriktade arbetskraftsutbildningen
Under den yrkesinriktade arbetskraftsutbildningen får du samma förmån som när du är arbetslös.
Om du har avtalat om yrkesinriktad arbetskraftsutbildning i din sysselsättningsplan, kan du få förhöjd arbetslöshetsförmån.
Det betyder att du får lite mer pengar i din arbetslöshetsförmån.
Beslut om utbetalning av förhöjningsdelen fattas av den som betalar arbetslöshetsförmånen, alltså arbetslöshetskassan eller FPA.
Du kan även få kostnadsersättning för resekostnader för de dagar som du deltar i utbildningen.
Om den som betalar din arbetslöshetsförmån inte betalar ut kostnadsersättning, kan arbets- och näringsbyrån i vissa fall betala den.
FPA:s kostnadsersättningfinska _ svenska _ engelska
Frivillig utbildning med arbetslöshetsförmån
Du kan även få arbetslöshetsförmån under andra studier om arbets- och näringsbyrån bedömer att du behöver utbildningen.
Arbets- och näringsbyrån skaffar inte utbildningen och väljer inte studeranden till utbildningen såsom i arbetskraftsutbildning.
Du ansöker om studieplats direkt vid läroanstalten.
Du måste avtala om utbildningen med arbets- och näringsbyrån innan du inleder utbildningen.
Du kan få arbetslöshetsförmån under studierna, om
du har anmält dig som arbetssökande vid arbets- och näringsbyrån och din jobbsökning är i kraft
du är minst 25 år gammal
arbets- och näringsbyrån bedömer att utbildningen främjar din yrkeskunnighet eller hjälper dig att få ett jobb
du har avtalat om utbildningen i din sysselsättningsplan med arbets- och näringsbyrån.
För vilka studier kan man få arbetslöshetsförmån?
Med arbetslöshetsförmånen understöds bara heltidsstudier.
Som heltidsstudier räknas följande:
högskoleexamen gymnasiestudier eller
studier, vars omfattning motsvarar heltidsstudier, till exempel fem studiepoäng i månaden eller 25 studietimmar i veckan.
Studierna ska leda till
yrkesinriktade grundexamen, yrkesexamen eller specialyrkesexamen
lägre eller högre högskoleexamen vid universitet eller högskola
avläggande av delar av ovan nämnda examina.
Studierna kan även vara tilläggsutbildning eller påbyggnadsutbildning alternativt studier vid universitet eller yrkeshögskola.
linkkiArbets- och näringsministeriet:
Frivilliga studier med stöd av arbetslöshetsförmånfinska _ svenska _ engelska
Alla barn som har sitt stadigvarande boende i Finland har läroplikt, vilket innebär att de måste delta i den grundläggande utbildningen.
Läroplikten är lagstadgad.
Läroplikten
börjar det år då barnet fyller 7 år
upphör när grundskolans lärokurs har fullgjorts eller det har förflutit 10 år sedan läroplikten började.
Läroplikten fullgörs vanligtvis i grundskolan.
Grundskolan består av lågstadiet (alakoulu) och högstadiet (yläkoulu).
Lågstadiet omfattar årskurserna 1–6, högstadiet årskurserna 7–9.
Grundskolan är vanligen nioårig: skolan börjar i årskurs 1 och slutar i årskurs 9.
Grundskolan är gratis.
Grundläggande utbildning för invandrarefinska _ svenska
Att börja i skolan
Föräldrarna anmäler sitt barn till skolan.
I början av året skickar staden en anmälan om läroplikt (oppivelvollisuusilmoitus) till hemmen.
I anmälan anges barnets närskola (lähikoulu).
Närskolan är oftast den skola som ligger närmast barnets hem.
Föräldrarna kan också välja en annan skola än närskolan.
Det är ändå inte alltid möjligt att få en plats på en annan skola.
Du kan anmäla ditt barn till skolan i närskolan.
I vissa kommuner kan anmälan göras även på internet.
Anmälningstiden är i början av året, vanligen i januari.
Olika skolor
Barn kan också gå i en skola med en speciell inriktning.
Ibland är dessa skolor privatskolor.
Skolor kan ha till exempel följande inriktningar:
bildkonst
motion
språk
internationalitet (till exempel Europaskolan)
specialpedagogik (till exempel Steinerpedagogik)
I Finland finns några internationella skolor.
I vissa skolor ges undervisningen på något annat språk än finska.
Till exempel i Tyska skolan sker undervisningen på tyska.
Skolor som har andra undervisningsspråk än finska finns i de största städerna.
Även i vanliga grundskolor kan det finnas några klasser där undervisningen sker på ett främmande språk.
linkkiEuropaskolan i Helsingfors:
Europaskolan i Helsingforsfinska _ engelska _ franska
linkkiFörbundet för Steinerpedagogik:
Information om Steinerskolanfinska _ engelska
Skoldagen och studierna
Skolan börjar i augusti och slutar i slutet av maj eller i början av juni.
I juni och juli är det sommarlov.
Längden på skoldagarna varierar i olika årskurser.
På lågstadiet är dagarna kortare än på högstadiet.
Lektionerna är vanligen 45 minuter långa.
Skolveckan består av ungefär 20 lektioner.
Barnen äter en varm måltid i skolan.
Den är gratis.
Om ditt barn har en specialdiet ska du tala om det för läraren.
I grundskolan studerar barnen många obligatoriska ämnen.
I lågstadiets högre klasser och på högstadiet får de även välja tillvalsämnen.
Alla kan få undervisning i den egna religionen eller i livsåskådningskunskap i skolan.
Religionsundervisning måste ordnas när det finns minst tre barn som bekänner en viss religion i kommunen.
I vissa skolor finns det skilda klasser för elever som är duktiga på till exempel musik eller bildkonst.
Oftast söker man separat till dessa klasser.
Invandrare och grundskolan
Barnet eller den unga kan få förberedande undervisning före den grundläggande utbildningen under vilken han eller hon studerar finska (eller svenska) och vissa läroämnen.
Den förberedande undervisningen före grundskolan är avsedd för alla de barn med invandrarbakgrund som inte har tillräckliga kunskaper för att klara sig i undervisningen inom den grundläggande utbildningen.
Den förberedande undervisningen pågår vanligtvis i ett år.
Därefter övergår eleven till en vanlig klass.
Om barnet har ett annat modersmål än finska eller svenska kan kommunen ordna undervisning i barnets eget modersmål.
Då kan barnet även lära sig finska eller svenska som andra språk, som S2-språk (S2-kieli).
Eleven studerar finska (eller svenska) som andra språk om hans eller hennes kunskaper i språket inte är på samma nivå som infödda talares.
Vuxengymnasier ordnar grundläggande utbildning för vuxna invandrare som inte har grundskolans avgångsbetyg från sitt eget land.
Mer information om detta får du vid rådgivningen i din hemkommun eller vid närmaste vuxengymnasium.
Du kan söka kontaktuppgifter tillvuxengymnasier med hjälp av sökmotorer på Internet.
linkkiUndervisnings- och kulturministeriet:
Information om grundundervisningenfinska _ svenska _ engelska
linkkiUtbildningsstyrelsen:
Information om grundundervisningenfinska _ svenska _ engelska
Meddelanden mellan hem och skola
I många kommuner informerar skolan viktiga ärenden i den webbaserade tjänsten Wilma.
Skolan ger barnets föräldrar inloggningsuppgifter till tjänsten.
Via Wilma kan du ha kontakt med barnets lärare och få information om barnets lärande, prov och frånvaron samt händelser i skolan och om skollov.
Om barnet är frånvarande från skolan till exempel på grund av sjukdom ska du meddela skolan om detta på morgonen via Wilma.
Det är viktigt att man regelbundet följer Wilma.
Om du behöver hjälp med att använda Wilma ska du be skolan om en introduktion.
Kervo stad har publicerat anvisningar om användningen av Wilma på olika språk.
Observera att inloggning till Wilma sker på olika adresser i olika städer.
linkkiKervo stad:
Så här använder du Wilma(pdf, 239 kt)finska _ engelska _ ryska _ estniska _ turkiska _ kurdiska _ thai _ vietnamesiska
linkkiVisma:
Stöd för studierna och tionde klassen
Grundskoleelever får stöd i sitt skolarbete.
Studiehandledarna berättar om olika studiemetoder och om fortsatta studier.
De ger också yrkesvägledning.
Studiepsykologer och skolkuratorer hjälper eleverna i problemsituationer.
Läraren kan ge barnet kortvarig stödundervisning.
Barnet får specialundervisning om det har inlärnings- eller koncentrationssvårigheter.
Grupperna i specialundervisningen är mindre än vanliga klasser.
Lärarna håller kontakt med föräldrarna.
De ordnar föräldramöten och berättar för föräldrarna om barnets studier.
Många skolor håller kontakt med föräldrarna med hjälp av webbtjänster.
I skolan ges eventuellt också tilläggsundervisning, på så kallade tionde klasser (kymppiluokka).
Där kan eleverna höja sina vitsord och fundera på vilket studieområde de är intresserade av.
Du kan ansöka till en tionde klass när du har fått ditt avgångsbetyg från grundskolan.
Information om tiondeklassenfinska _ svenska
Gymnasieansökan
Sök till gymnasiet i den gemensamma ansökan till andra stadiet i februari-mars.
Du kan söka till ett gymnasium om du har avlagt lärokursen för den grundläggande utbildningen eller en lärokurs som motsvarar den grundläggande utbildningen.
Fyll ansökan i tjänsten Studieinfo.fi.
Eleverna antas till gymnasiet utifrån vitsorden på avgångsbetyget från grundskolan.
Därtill ordnar vissa gymnasier inträdesprov.
Om du söker till ett vuxengymnasium, kontakta läroanstalten direkt.
Du kan inte söka till ett vuxengymnasium i den gemensamma ansökan.
När du söker till ett vuxengymnasium är inte medeltalet på ditt betyg av betydelse.
Du hittar utbildningar på Studieinfo.fi.
Om du vill förbättra dina kunskaper i finska innan du söker till ett gymnasium, kan du söka till en förberedande gymnasieutbildning
Läs mer på InfoFinlands sida Gymnasieförberedande utbildning.
Ansökan till gymnasium i den gemensamma ansökanfinska _ svenska
Ansökan till yrkesutbildning
Din grundutbildning avgör till hurudan yrkesutbildning du kan söka och på vilket sätt ansökan sker.
Du kan söka till en grundskolebaserad yrkesutbildning om du har avlagt lärokursen för den grundläggande utbildningen eller en lärokurs som motsvarar den grundläggande utbildningen.
Du kan söka till en gymnasiebaserad yrkesutbildning om du har gått färdigt gymnasiet.
Du kan söka till dessa utbildningar i den kontinuerliga ansökan året om eller i den gemensamma ansökan till andra stadiet.
I allmänhet ordnas den gemensamma ansökan i februari-mars och september-oktober.
Fyll ansökan i tjänsten Studieinfo.fi.
Om du redan har avlagt en yrkesexamen eller en högskoleexamen, kan du inte söka till en yrkesutbildning i den gemensamma ansökan.
Då kan du söka direkt till läroverket i den separata ansökningsprocessen som är avsedd för dem som redan avlagt examen.
Du kan även ansöka till yrkesutbildning för vuxna.
Grunderna för antagning av studeranden beror på utbildningen.
I allmänhet påverkas antagningen av antagningspoängen, som ges bl.a. utifrån dina betyg.
Inträdesprov eller lämplighetsprov ordnas också för många utbildningar.
Om ditt modersmål är ett annat än undervisningsspråket, behöver du ett intyg över din språkkunskap.
Det kan exempelvis vara avgångsbetyg från finsk grundskola.
Tjänsten Studieinfo.fi ger dig närmare information om intyg med vilka du kan påvisa din språkkunskap.
Om du inte har intyg över din språkkunskap, får du en inbjudan till ett språkprov.
Om du vill ha mera kunskap och färdigheter innan du söker till en yrkesinriktad utbildning, kan du ansöka till VALMA-utbildningen.
Under VALMA-utbildningen kan du även förbättra dina språkkunskaper i finska.
Läs mera på InfoFinlands sida Utbildning som handleder för yrkesutbildning.
Om du behöver särskilt stöd i de yrkesinriktade studierna t.ex. på grund av handikapp eller inlärningssvårigheter ska du ansöka till utbildningen via ansökan till specialundervisning.
Ansökan till yrkesutbildning i den gemensamma ansökanfinska _ svenska
Kontinuerlig ansökan till yrkesutbildning finska _ svenska
Antagningsgrunder till yrkesutbildningfinska _ svenska
Om du har en utländsk examen
Om du har avlagt grundskolan eller gymnasiet utomlands, antas du till en yrkesutbildning enligt prövning.
Vid antagning enligt prövning beaktas
ditt utbildningsbehov
bedömningen av hur bra du kan klara av studierna.
Antagning enligt prövningfinska _ svenska
Ansökan till en yrkesinriktad vuxenutbildning
Du kan söka till en yrkesinriktad vuxenutbildning om du vill avlägga en examen vid sidan om arbetet.
I vuxenutbildningen avlägger du yrkesexamen som fristående examen.
Du kan söka till en yrkesinriktad vuxenutbildning också om du har avlagt en yrkesexamen eller en högskoleexamen.
När du söker till en yrkesinriktad vuxenutbildning, ska du ha en tillräckligt lång arbetserfarenhet.
Du kan inte söka till en yrkesinriktad vuxenutbildning i den gemensamma ansökan.
Ta reda på hur du kan söka till utbildningen i tjänsten Studieinfo.fi eller av läroanstalten.
Ofta är ansökningstiden fortlöpande.
Ansökan till en yrkeshögskola
Du kan söka till en yrkeshögskola för att avlägga en yrkeshögskoleexamen, då du har avlagt t.ex. någon av följande utbildningar:
gymnasiet
en yrkesexamen
studentexamen eller en motsvarande examen i ett annat land
Du får närmare uppgifter från tjänsten Studieinfo.fi.
Sök till en yrkeshögskola i den gemensamma ansökan till högskolor.
Den gemensamma ansökan ordnas två gånger per år, på våren och på hösten.
Fyll ansökan i tjänsten Studieinfo.fi.
Grunderna för antagning av studeranden beror på utbildningen.
Ditt betyg, inträdesprovet och din arbetserfarenhet kan påverka antagningen.
Också dina tidigare studier kan spela en roll.
Ansökan till YH-examenfinska _ svenska
Högre yrkeshögskoleexamina
Du kan söka till en YH-examen om du har
en lämplig yrkeshögskoleexamen eller en annan lämplig högskoleexamen och
minst tre års arbetserfarenhet från samma område som din examen och du har inhämtat din arbetserfarenhet efter att du har avlagt examen.
Sök till en YH-examen i den gemensamma ansökan till högskolor på våren eller hösten Till många utbildningar är det möjligt att söka endast på våren.
Fyll i ansökningsblanketten i tjänsten Studieinfo.fi.
Du kan söka till en högre YH-examen på ett främmande språk med en separat ansökan.
Du hittar ansökningsblanketter då du letar efter utbildningar i Studieinfo.fi.
Högre YH-examenfinska _ svenska
Ansökan till universitet
Ansök till ett universitet antingen i den gemensamma ansökan till högskolor eller med en separat ansökan till en viss utbildning.
Du kan söka till många universitetsutbildningar i den gemensamma ansökan till högskolor.
Den ordnas på våren och hösten.
Alternativen är fler på våren.
Den gemensamma ansökan till vissa utbildningar ordnas redan i januari.
Utred i tid när du kan söka.
Fyll ansökan i tjänsten Studieinfo.fi.
Du kan söka till ett universitet om du har avlagt t.ex. någon av följande examina:
en finländsk studentexamen
en minst treårig yrkesinriktad grundexamen
en utländsk examen, som ger möjlighet till universitetsstudier i det land där du avlagt examen
Granska av högskolans studiebyrå att det är möjligt att söka till ett universitet med din examen.
Du får närmare uppgifter också från tjänsten Studieinfo.fi.
När du söker till ett universitet, får du i allmänhet poäng utifrån studentexamen och inträdesprovet.
Det finns skäl att förbereda dig omsorgsfullt för inträdesprovet.
Till vissa utbildningsprogram antas endast en liten del av sökandena.
Vissa inträdesprov omfattar förhandsuppgifter.
Ansökan till universitetfinska _ svenska _ engelska
Separat ansökan
Ansökan till vissa universitetsstudier sker genom en separat ansökan.
Du ska söka med en separat ansökan t.ex.
om du söker till ett magisterprogram
om du flyttar från en högskola till en annan eller
om du har avlagt studier i ett öppet universitet och söker till ett universitet utifrån dessa studier.
Om du söker till ett utbildningsprogram där undervisningsspråket är ett annat än finska eller svenska, beror ansökningssättet på utbildningen.
Det lönar sig att söka till vissa utbildningar på främmande språk i den gemensamma ansökan i januari.
Du hittar närmare information i Studieinfo.fi.
Du kan också fråga direkt av högskolorna.
De separata ansökningarna kan ordnas under olika tidsperioder och ansökningsförfarandena kan avvika från varandra.
Du hittar de separata ansökningarna via tjänsten Studieinfo.fi.
Påbyggnadsexamen
Om du vill avlägga en påbyggnadsexamen vid ett universitet, kontakta universitetet direkt.
Mottagande av studieplats
Läroanstalten meddelar dig att du har antagits för studier med ett brev.
Om du har antagits, meddela så fort som möjligt till läroanstalten att du tar emot studieplatsen.
Brevet innehåller anvisningar om hur du tar emot platsen och hur du anmäler dig.
Om du inte tar emot platsen i tid, förlorar du den.
När du tar emot en studieplats, förbinder du dig att börja studera i läroanstalten.
Du kan söka till många olika läroanstalter i den gemensamma ansökan.
Du kan dock ta emot endast en studieplats.
Efter grundskolan (peruskoulu), d.v.s. efter grundstadiet fortsätter studerandena till läroanstalter på andra stadiet (toisen asteen oppilaitos).
Läroanstalter på andra stadiet är gymnasiet och yrkesläroanstalter.
Läs mer om yrkesläroanstalter på InfoFinlands sida Yrkesutbildning.
Gymnasiestudierna är mer teoretiskt inriktade än yrkesutbildning.
Studierna är allmänbildande: fokus ligger speciellt på naturvetenskapliga och humanistiska ämnen.
I vissa gymnasier ges även mycket undervisning i konstämnen.
Vissa gymnasier är specialgymnasier.
De är inriktade på till exempel musik, idrott eller naturvetenskaper.
Specialgymnasierna är mycket populära.
Det kan vara svårt att komma in dit.
Gymnasiet ger förberedande utbildning till exempel för yrkeshögskola och universitet.
Både ungdomar och vuxna kan studera vid gymnasiet.
Ungdomarna studerar vid daggymnasiet (päivälukio) eller distansgymnasiet (etälukio), vuxna studerar ofta vid vuxengymnasiet (aikuislukio).
Information om gymnasiestudierfinska _ svenska
linkkiFörbund för gymnasieelever:
Förbund för gymnasieeleverfinska _ svenska _ engelska
linkkiUtbildningsstyrelsen:
Information om gymnasiestudierfinska _ svenska _ engelska
Att söka till gymnasiet
Sök till gymnasiet i den gemensamma ansökan till andra stadiet.
Om du vill studera vid ett vuxengymnasium ska du ta kontakt direkt med läroanstalten.
Läs mer på InfoFinlands sida Ansökan till utbildning.
Gemensam ansökan till gymnasier och yrkesläroanstalterfinska _ svenska
Att studera vid gymnasiet
Gymnasiestudierna pågår vanligen tre år.
Gymnasiet kan också avläggas på två eller fyra år.
I gymnasiestudierna har du många valmöjligheter.
Utöver de obligatoriska kurserna kan du välja många kurser som passar dig.
I gymnasiet påverkar du själv innehållet i dina studier och din studietakt.
I gymnasiet tas inga terminsavgifter ut.
Utbildningen kostar alltså inget.
Studeranden måste dock själv skaffa gymnasieböckerna.
Böckerna är ofta dyra.
Man kan även köpa gymnasieböckerna begagnade.
Om du till exempel har en krävande hobby eller är sjuk en lång tid kan du avlägga gymnasiet som distansstudier.
Fråga mer om distansstudier vid ditt eget gymnasium.
Studentexamen
Gymnasiestudierna siktar till studentexamen (ylioppilastutkinto).
Studentexamen består av prov i olika läroämnen.
Studentskrivningarna (ylioppilaskokeet) skrivs oftast i slutet av studierna.
Modersmålsprovet är ett obligatoriskt prov i studentexamen.
Modersmålsprovet kan skrivas i finska, svenska eller samiska.
Om du inte har finska, svenska eller samiska som modersmål kan du skriva ett prov i finska eller svenska som andra språk.
Utöver modersmålsprovet måste du skriva prov i minst tre andra ämnen.
Om du vill kan du även skriva fler ämnen.
Utöver modersmålsprovet kan du skriva prov i följande andra ämnen:
Det andra inhemska språket (finska eller svenska)
Ett främmande språk: engelska, tyska, ryska, franska, spanska, portugisiska, latin
Matematik
Realämnen (reaali), d.v.s. historia, religion, fysik, kemi, biologi, psykologi, filosofi
Studentskrivningarna ordnas på våren och på hösten.
Om du vill kan du skriva några ämnen på hösten och resten på våren.
Du måste skriva alla prov på högst tre efter varandra följande examenstillfällen.
Info om studentexamenfinska _ svenska
linkkiStudentexamensnämnden:
Information om studentexamenfinska _ svenska _ engelska _ franska _ tyska
Vuxengymnasium
Vuxengymnasiet är i huvudsak avsett för personer som har fyllt 18 år.
Vid vuxengymnasiet är studierna flexibla.
Du kan avlägga hela studentexamen eller bara studera ett ämne.
Undervisningen sker oftast kvällstid.
Många vuxengymnasier erbjuder finskakurser för invandrare.
Fråga om kurserna direkt vid vuxengymnasiet.
Information om vuxengymnasietfinska _ svenska
linkkiEdu.fi:
Enligt lag ska barn i Finland delta i förskoleundervisning eller motsvarande verksamhet under ett års tid innan läroplikten börjar.
Förskoleundervisningen (esiopetus) förbereder barnen inför grundskolan.
Barnen börjar i förskoleundervisningen vanligen vid sex års ålder och grundskolan vid sju års ålder.
Föräldrarna anmäler sitt barn till förskoleundervisningen vanligtvis i januari eller februari.
Kontrollera tidpunkten i god tid vid skolväsendet (koulutoimi) eller bildningsväsendet (sivistystoimi) i din hemkommun.
Kommunerna ordnar förskoleundervisning.
De kan även köpa förskoleundervisningen till exempel av ett privat daghem.
Förskoleundervisningen är kostnadsfri.
Under dagen får barnet en gratis måltid.
Om barnet bor långt (över 5 km) från undervisningsstället, eller om vägen dit är besvärlig, får barnet gratis skjuts.
Om föräldrarna arbetar eller studerar kan barnet utöver förskoleundervisningen även delta i småbarnspedagogiken.
En dag i förskolan
Förskoledagen är ungefär fyra timmar lång.
Förskolan finns ofta antingen i daghemmets eller skolans lokaler.
I förskolan lär sig barnen bland annat matematik, miljö- och naturkunskap samt konst och kultur.
De lär sig nya saker med lekens hjälp.
Föräldrarna har en viktig roll i förskolan.
De stödjer sitt barns inlärning.
Lärarna utarbetar en egen inlärningsplan för varje barn.
Föräldrarna kan hjälpa ledarna att utarbeta planen.
Språk och kulturer i förskoleundervisningen
Ett barn som har ett annat modersmål än finska eller svenska lär sig finska eller svenska som främmande språk.
Dessutom kan det studera sitt eget modersmål om kommunen ordnar undervisning i det språket.
Barnet kan även få undervisning i den egna religionen eller i livsåskådningskunskap i förskolan.
I förskolan lär sig barnen att uppskatta sitt språk och sin kultur.
De lär sig också att respektera andra människors språk och kulturer.
linkkiUtbildningsstyrelsen:
Information om förskoleundervisningenfinska _ svenska
Förskoleuppgifter på nätetfinska
linkkiUndervisnings- och kulturministeriet:
Information om förskoleundervisningenfinska _ svenska _ engelska
På den här sidan finns information om tjänster för invandrare i Rovaniemi.
Verso Integration av och rådgivning för invandrare
Personer som kommer till Finland som flyktingar kan ta del av integrationsrelaterade socialtjänster vid Rovaniemi stads invandrarbyrå.
I samarbete med berörda myndigheter ansvarar invandrarbyrån för den inledande kartläggningen samt ordnandet av integrationsplan och nödvändiga åtgärder och tjänster.
Kontaktuppgifterna till invandrarbyrån i Rovaniemi är:
Rovaniemi stads invandrarbyrå
Anställda vid invandrarbyrån
Ledande socialarbetare 016-322 3087, 040-731 2557
Socialarbetare 016-322 3088, 040-576 8914
Socialarbetare 016-322 3126, 040-351 6925
Socialhandledare 016-322 3123, 0400-695 037
Socialhandledare 016-322 3125, 040-576 8904
Socialhandledare 016-322 3124, 040-729 8766
Tolkbeställning
p. 050-597 1122
Förmånshandläggare
p. 050-593 0165
Byråarbetare
p. 050-571 5860
Mer information om flytt, uppehållstillstånd och personuppgifter fås från bland annat magistraten, polisen och invandrarbyrån.
Läs mer: Flytta till Rovaniemi
MoniNet, centret för mångkulturell information och verksamhet
MoniNet, som i Rovaniemi upprätthålls av Rovalan Setlementti ry, är ett center för mångkulturell information och verksamhet.
Det betjänar invandrare som är bosatta i Rovaniemi och annorstädes i Lappland.
Mer informtion om MoniNets verksamhet fås via adressen:
MoniNetfinska _ engelska
Samarbetsprojektet Verso
Samarbetsprojektet Verso är ett samarbete mellan Rovaniemi stad och Rovalan Setlementti ry.
Syftet med projektet är att utveckla tjänsteprocesserna för invandrare, avsedda för den inledande tiden direkt efter inflyttningen.
Samarbetsprojektet Versofinska
På den här sidan finns information om tjänster för invandrare i Rovaniemi.
Verso Integration av och rådgivning för invandrare
Personer som kommer till Finland som flyktingar kan ta del av integrationsrelaterade socialtjänster vid Rovaniemi stads invandrarbyrå.
I samarbete med berörda myndigheter ansvarar invandrarbyrån för den inledande kartläggningen samt ordnandet av integrationsplan och nödvändiga åtgärder och tjänster.
Kontaktuppgifterna till invandrarbyrån i Rovaniemi är:
Rovaniemi stads invandrarbyrå
Anställda vid invandrarbyrån
Ledande socialarbetare 016-322 3087, 040-731 2557
Socialarbetare 016-322 3088, 040-576 8914
Socialarbetare 016-322 3126, 040-351 6925
Socialhandledare 016-322 3123, 0400-695 037
Socialhandledare 016-322 3125, 040-576 8904
Socialhandledare 016-322 3124, 040-729 8766
Tolkbeställning
p. 050-597 1122
Förmånshandläggare
p. 050-593 0165
Byråarbetare
p. 050-571 5860
Mer information om flytt, uppehållstillstånd och personuppgifter fås från bland annat magistraten, polisen och invandrarbyrån.
Läs mer: Flytta till Rovaniemi
MoniNet, centret för mångkulturell information och verksamhet
MoniNet, som i Rovaniemi upprätthålls av Rovalan Setlementti ry, är ett center för mångkulturell information och verksamhet.
Det betjänar invandrare som är bosatta i Rovaniemi och annorstädes i Lappland.
Mer informtion om MoniNets verksamhet fås via adressen:
MoniNetfinska _ engelska
Samarbetsprojektet Verso
Samarbetsprojektet Verso är ett samarbete mellan Rovaniemi stad och Rovalan Setlementti ry.
Syftet med projektet är att utveckla tjänsteprocesserna för invandrare, avsedda för den inledande tiden direkt efter inflyttningen.
Samarbetsprojektet Versofinska
Integration av och rådgivning för invandrare
Inledande kartläggning och integrationsplan
Behöver du en tolk eller översättare?
Integration av och rådgivning för invandrare
MoniNet
Kontakta oss om du behöver råd och hjälp i vardagen, vill lära dig finska eller frivilligarbeta, delta i utflykter och evenemang eller utöva fritidsintressen.
MoniNet
Kansankatu 8 (vån. 2)
Tfn 040 559 6564
MoniNet är ett mångkulturellt center som drivs av Rovalan Setlementti ry och ordnar rådgivning och aktiviteter för invandrare.
Syftet med verksamheten är att stödja integrationen av invandrare, främja toleransen och acceptansen av mångfald, öka sysselsättningen, utveckla nya strategier och nätverka med aktörerna i regionen.
MoniNetfinska _ engelska
Välfärds- och servicepunkten Olkkari
Rovaniemi stads välfärds- och servicepunkt ger dig information om stadens tjänster.
Olkkari erbjuder servicehandledning och rådgivning för stadsbor i alla åldrar när det gäller social- och hälsovårdstjänster, kulturella aktiviteter, jobbsökningscoachning, idrottstjänster och organisationsverksamhet.
I samma lokal finns kundtjänsten Osviitta, där du kan köpa resekort till lokaltrafiken.
Köpcentret Rinteenkulma
Tfn 016 322 6800
Välfärds- och servicepunkten Olkkarifinska
Navigatorn
Om du är under 30 år kan du få informations-, rådgivnings- och handledningstjänster på Rovaniemi stads navigator.
Navigatorn ger dig råd om utbildning, arbete, vardagen och livet.
På Navigatorn kan någon i personalen hjälpa dig att reda ut saker och ting.
Navigatorn finska
Integrationsrelaterade socialtjänster
Om du behöver rådgivning och handledning om integration kan du kontakta Rovaniemi stads integrationsrelaterade socialtjänster.
Tjänsten är i första hand avsedd för personer med flyktingbakgrund och deras familjemedlemmar.
Tjänsten kan också användas av andra invandrare som behöver tillfällig rådgivning i specialfrågor som rör integration.
De integrationsrelaterade socialtjänsterna omfattar rådgivning och handledning.
Dessutom görs en inledande kartläggning och integrationsplan för invandrare som inte kan registrera sig som arbetslös arbetssökande.
Socialservicecentret
Invandrarbyrån
Tfn 050 571 5860
Inledande kartläggning och integrationsplan
Invandrare har rätt till en inledande kartläggning.
Den inledande kartläggningen hjälper dig att hitta rätt tjänster i din hemstad.
Utifrån den inledande kartläggningen görs en bedömning av om det även vore bra att göra upp en integrationsplan för dig.
Den inledande kartläggningen och integrationsplanen kan utarbetas tillsammans med dig antingen på Lapplands TE-byrå eller inom Rovaniemi stads socialservice, till exempel inom de integrationsrelaterade socialtjänsterna
eller vuxensocialarbetet.
Lapplands TE-byrå
En anställd vid arbets- och näringsbyrån gör den inledande kartläggningen
och integrationsplanen tillsammans med dig om du anmäler dig till TE-byrån som arbetslös arbetssökande.
Du kan registrera dig som arbetslös arbetssökande elektroniskt
via tjänsten Mina e-tjänster eller per telefon.
När du är arbetslös
kan du ha rätt till integrationsutbildning som ordnas genom TE-byrån.
Om du inte har möjlighet att identifiera dig i Mina e-tjänster eller om du vill uträtta dina ärenden per telefon kan du få information, rådgivning, vägledning och stöd i användningen av nättjänsterna från den nationella telefontjänsten.
Service på finska 0295 025 500
Service på svenska 0295 025 510
Service på engelska 0295 020 713
Service på ryska 0295 020 715
Du måste alltid boka tid till kundtjänsten vid Lapplands TE-byrå i förväg.
I anslutning till TE-byrån finns ett rum där man kan uträtta ärenden på egen hand.
Om det behövs kan du få servicerådgivning om användningen av nättjänsterna.
Lapplands TE-byrå
Servicestället i Rovaniemi
Valtakatu 16
PB 1000
På TE-byråernas webbplats hittar du broschyrer och filmer om registrering som arbetslös arbetssökande, yrkesval, utbildning och utkomstskydd för arbetslösa på flera olika språk.
linkkiTE-tjänster:
Mina e-tjänsterfinska _ svenska
linkkiTE-tjänster:
Information om TE-byråns tjänster för invandrare finska _ svenska _ engelska
linkkiTE-tjänster:
Integrationstjänster för invandrare finska _ svenska _ engelska
Socialservicecentret
Om du är 17–64 år gammal och på grund av din livssituation inte har anmält dig som arbetslös arbetssökande kan personalen på Rovaniemi stads socialservicecenter göra en inledande kartläggning och vid behov även en integrationsplan tillsammans med dig.
Du kan själv be om en inledande kartläggning.
Dessutom kan du få stöd, rådgivning och handledning.
Socialservicecentret
Tjänster för vuxna och personer i arbetsför ålder
Servicerådgivning per telefon
Tfn 016 3222 570.
Vuxensocialarbetefinska
Behöver du en tolk eller översättare?
Om du inte kan finska eller svenska kan du använda en tolk när du uträttar ärenden hos myndigheterna.
I vissa fall får du en tolk genom myndigheten om du meddelar behovet av tolkning i förväg.
I det här fallet är tolkningen avgiftsfri. Tolkning ska alltid begäras i förväg.
Du kan använda en tolk när du vill om du beställer tolken själv och betalar kostnaderna.
Många företag erbjuder tolknings- och översättningstjänster.
Du hittar kontaktuppgifterna till dem till exempel på Finlands översättar- och tolkförbunds webbplats.
linkkiFinlands översättar- och tolkförbund:
Tolknings- och översättningstjänsterfinska _ svenska _ engelska
I Finland kan man avlägga högskolestudier både vid yrkeshögskolor och vid universitet.
Läs mer om yrkeshögskolan på InfoFinlands sida Yrkeshögskolor.
Ansök om studieplats
Du kan söka till ett universitet om du har avlagt en finländsk studentexamen, en utländsk examen som motsvarar studentexamen eller en yrkesinriktad slutexamen. Sök till ett universitet i den gemensamma ansökan till högskolor.
Läs mer på InfoFinlands sida Ansökan till utbildning.
Gemensam ansökan till universitetfinska _ svenska
Vilka yrken kan studera till?
Vid universitet kan man studera i många olika studieområden.
De som har utexaminerats från en högskola eller ett universitet arbetar i många slags arbetsuppgifter.
En del universitetsstudier leder direkt till ett yrke.
Sådana yrken är till exempel:
lärare
jurist
läkare
skådespelare
diplomingenjör
bildkonstnär
Andra universitetsstudier leder inte till ett visst yrke.
Till exempel studerande vid den samhällsvetenskapliga eller den humanistiska fakulteten utexamineras inte nödvändigtvis till ett yrke.
Dessa människor arbetar till exempel i följande arbetsuppgifter:
forskare
statlig tjänsteman
Studier vid universitet
Vid vissa universitet har olika examen olika namn.
Till exempel är tekniska högskolors motsvarighet till magisterexamen diplomingenjörsexamen (diplomi-insinööri).
När du får en studieplats får du rättighet att avlägga båda examina.
Du kan också avsluta studierna efter lägre högskoleexamen.
Kandidatstudierna pågår ungefär tre år, magisterstudierna ungefär två år.
Hur fort studierna framskrider beror på dig själv.
Du kan också söka till ett separat magisterprogram.
Magisterprogrammet är ett studieprogram som leder till högre högskoleexamen.
För att kunna studera i ett magisterprogram ska du ha avlagt lägre högskoleexamen.
Magisterprogrammen pågår i cirka två år.
Vid dem studerar ofta människor från många olika vetenskapsområden.
Utexaminering från universitetet
När du är klar med dina studier får du antingen kandidatexamen eller magisterexamen.
Om du vill kan du efter magisterexamen söka till fortsatta studier.
Information om högskolestudierfinska _ svenska _ engelska
linkkiFinlands Studentkårers Förbund:
Information om studentkårer i Finlandfinska _ svenska _ engelska
Öppna universitet
De öppna universiteten tillhandahåller universitetskurser.
Vem som helst kan studera vid ett öppet universitet.
Du kan studera vid ett öppet universitet även om du inte har någon examen.
Läs mer på InfoFinlands sida Studier som hobby.
Vetenskaplig fortbildning vid universitet
Vetenskaplig fortbildning vid universitet är examensinriktad fortbildning.
Sådan utbildning förbereder dig till exempel för forskaryrket.
Vid universitetet kan du avlägga licentiatexamen (lisensiaatti) eller doktorsexamen (tohtori).
De flesta studerande som bedriver fortsatta studier avlägger doktorsexamen.
Man kan ansöka till fortsatta studier vid universitet några gånger per år.
Universitet och institutioner har olika ansökningstider.
Kontrollera ansökningstiden vid den institution där du vill bedriva fortsatta studier.
I Finland måste de som bedriver fortsatta studier ofta finansiera studierna själva.
Du kan ansöka om stipendier hos olika stiftelser (säätiö).
Påbyggnadsexamina vid universitetfinska
linkkiStiftelsetjänst:
Information om stiftelser och penningunderstödfinska _ svenska _ engelska
linkkiCIMO:
Penningunderstöd för utländska forskarefinska _ svenska _ engelska
Vägledning i högskolestudier
Vid högskolornas SIMHE-tjänster kan du söka hjälp och information om högskoleutbildning i Finland och om hur du ansöker till högskoleutbildning.
Du kan även få information om andra utbildningsmöjligheter för personer som avlagt högskolestudier.
Du kan få vägledning via SIMHE-tjänsterna om
du har flyttat till Finland
du är intresserad av högskolestudier och
du har avlagt högskolestudier eller högskoleexamen utomlands.
Vägledning kan ges individuellt eller i grupp.
linkkiUtbildningsstyrelsen:
Högskolor som erbjuder SIMHE-tjänsterfinska _ svenska _ engelska
Utbildning som handleder för grundläggande yrkesutbildning (Ammatilliseen peruskoulutukseen valmentava koulutus) d.v.s. VALMA är avsedd för dem som vill avlägga en grundläggande yrkesutbildning.
Under VALMA-utbildningen får du kunskap och färdigheter som hjälper dig i dina senare yrkesinriktade studier.
Du kan även förbättra din språkkunskap. Du kan också höja dina grundskolebetyg.
VALMA-utbildningen räcker ungefär ett läsår.
Du kan under utbildningen bekanta dig med olika branscher och fundera på vad du vill studera.
Du besöker arbetsplatser och deltar i verkstäder.
I början av utbildningen görs det upp en personlig studieplan för dig.
I den skrivs det in vilka studier du avlägger och hur.
Du får ett betyg för VALMA-utbildningen.
Du får också tilläggspoäng när du ansöker till en yrkesutbildning i den gemensamma ansökan.
VALMA-utbildningen kostar vanligen inget för den studerande.
Information om VALMA-utbildningarfinska _ svenska _ engelska
Ansökan till VALMA-utbildningen
Du kan ansöka till VALMA-utbildningen om du har slutfört grundskolan eller en utbildning som motsvarar grundskolan.
Om läroinrättningen anser att du kan klara av studierna kan du antas som studerande även utan slutbetyg från grundskolan.
Ansök till VALMA-utbildningen efter den egentliga gemensamma ansökan i början av sommaren.
Om du behöver särskilt stöd t.ex. på grund av handikapp ska du ansöka till utbildningen på våren, under ansökan till specialundervisning.
Närmare information om ansökningstiderna hittar du via Studieinfo.fi-tjänsten.
Fyll i ansökningsblanketten i Studieinfo.fi-tjänsten.
Ansökan till VALMA-utbildningfinska _ svenska
Ansökan till specialundervisningfinska _ svenska
Småbarnspedagogik är avsedd för barn under skolåldern.
I Finland tillhandahåller kommunerna kommunal småbarnspedagogik bland annat i daghem.
Dessutom finns det privata daghem.
Småbarnspedagogik är fostran, undervisning och omsorg som är pedagogiskt planerad och som har noga genomtänkta mål.
Inom småbarnspedagogiken arbetar utbildade lärare i småbarnspedagogik och barnskötare.
Vanligen vårdar någondera av föräldrarna barnet hemma åtminstone under föräldraledigheten (vanhempainvapaa), det vill säga tills barnet är ungefär 9 månader gammalt.
Om du vårdar ditt barn hemma även efter detta har du rätt att vara ledig från ditt arbete för vård av barn tills barnet fyller tre år.
Mer information om ledigheterna får du på InfoFinlands sida Familjeledighet.
Du kan ansöka från Kela om ekonomiskt stöd för hemvård av barn.
Läs mer på InfoFinlands sida Stöd för vård av barn i hemmet.
Kommunal småbarnspedagogik
Om du har din hemkommun i Finland, kan du ansöka om en plats inom den kommunala småbarnspedagogiken för barnet efter föräldraledigheten.
Då är barnet ca nio månader gammalt.
Om du inte har en hemkommun i Finland, räknas du som invånare i den kommun där du vistas.
Om båda föräldrarna arbetar, har barnet rätt till småbarnspedagogik på heltid.
Om den ena föräldern är hemma, beror rätten till småbarnspedagogik på hemkommunen.
I vissa kommuner har barnet rätt till småbarnspedagogik på heltid även då den ena föräldern är hemma.
I vissa kommuner har barnet rätt till 20 timmar småbarnspedagogik per vecka om den ena föräldern är hemma.
Familjen kan ändå söka rätt till småbarnspedagogik på heltid om barnet behöver särskilt stöd till exempel i att lära sig det finska språket eller på grund av att familjen befinner sig i en svår situation.
Du kan ansöka om en plats
på ett daghem (päiväkoti)
På daghemmet är barnen i större gruppen är i gruppfamiljedagvården.
Familjedagvård innebär att skötaren vårdar barnen i sitt eget hem.
Vissa familjedagvårdare vårdar barnen hemma hos de barn som ingår i gruppen.
Ansök om en plats inom den kommunala småbarnspedagogiken från din egen kommun senast fyra månader innan du behöver den.
Man kan få en plats inom två veckor, om föräldrarna får ett arbete eller en studieplats.
Avgiften för småbarnspedagogik (varhaiskasvatusmaksu) beror på
familjens inkomster
familjens storlek och
på hur många timmar per vecka barnet deltar i småbarnspedagogik.
Man får syskonrabatt.
Om familjen inkomster är mycket låga, kan småbarnspedagogiken vara kostnadsfri för familjen.
Fråga mer i din kommuns rådgivningstjänster.
Privat småbarnspedagogik
En plats inom den privata småbarnspedagogiken kan finnas
i ett privat daghem eller i ett gruppfamiljedaghem
i familjedagvård eller
hemma, då familjen anställer en skötare i hemmet
Du kan ansöka om en plats inom småbarnspedagogiken direkt från det privata daghemmet eller gruppfamiljedaghemmet.
Du kan också leta upp en privat familjedagvårdare som vårdar barnen hemma hos sig, eller anställa en skötare i ditt eget hem.
Om du anställer en skötare i ditt hem blir du en arbetsgivare, och du måste uppfylla en arbetsgivares skyldigheter.
Läs mera på InfoFinlands sida Arbetsgivarens rättigheter och skyldigheter.
Familjen kan anställa en skötare i sitt hem även tillsammans med en annan familj.
Kommunen övervakar den privata småbarnspedagogiken.
Priserna för den privata småbarnspedagogiken varierar.
Du kan ändå få stöd för den från FPA.
Då är den inte nödvändigtvis mycket dyrare än den kommunala småbarnspedagogiken.
Stöd för privat dagvård
Om barnet har en hemkommun i Finland, kan du ansöka om Fpa-stöd för privat vård.
Dagvårdsproducenten måste ha kommunens godkännande.
Du kan ansöka om privatvårdsstöd (yksityisen hoidon tuki), om
ditt barn som är under skolåldern är i privat dagvård; eller
barnet har någon annan privat skötare.
Du kan inte ansöka om privatvårdsstöd om skötaren är en medlem i barnets familj eller om barnet och skötaren bor i samma hushåll.
Du kan inte heller ansöka om privatvårdsstöd för den kommunala småbarnspedagogiken.
Stödets storlek beror bland annat på familjens inkomster och kommunen som familjen bor i.
Kela betalar stödet direkt till skötaren eller dagvårdsproducenten.
Man måste betala skatt för privatvårdsstödet.
Stödet betalas inte till utlandet.
Läs mera om privatvårdsstöd på Fpa:s sidor.
Fpa har en telefontjänst för barnfamiljer.
på finska tfn +358 (0)20 692 206
på svenska och engelska tfn +358 (0)20 692 226
På Fpas byråer får du betjäning även på andra språk med hjälp av en tolk.
Stöd för privat vårdfinska _ svenska _ engelska
Vad händer i småbarnspedagogiken?
Till småbarnspedagogiken hör mångsidig verksamhet, till exempel lekar, motion, utevistelse, musik, pyssel och utfärder.
I dagen ingår också en vilostund.
Målsättningen med verksamheten är att främja barnets utveckling och lärande.
Barnet lär sig även sociala färdigheter.
Barnet får stöd i att lära sig det finska eller svenska språket, om hans/hennes modersmål är ett annat språk.
Om barnet behöver, kan hen även få specialundervisning.
Daghemmet är ändå inte en skola.
Barnen studerar inte skolämnen och har inte lektioner.
Barnen äter tre måltider under dagen: frukost, lunch och mellanmål.
Om ditt barn har en specialdiet ska du berätta om det för lärarna i småbarnspedagogiken.
I småbarnspedagogiken beaktas familjens religion eller livsåskådning.
På vissa orter finns det daghem, som fungerar på andra språk än finska eller svenska.
Vanligen börjar daghemsdagen på morgonen och tar slut på eftermiddagen.
Vissa daghem och familjedagvårdare har öppet dygnet runt med anledning av föräldrarnas arbete eller studier.
linkkiFinlands Flyktinghjälp:
Klubbar
Kommunerna, föreningar och församlingar ordnar dagklubbar för barn.
Klubbarna räcker vanligen ett par timmar.
I klubbarna ordnas handledda lekar, sång, pyssel och annat program.
linkkiUndervisnings- och kulturministeriet:
Information om småbarnspedagogikfinska _ svenska _ engelska
Studierna vid en yrkeshögskola (ammattikorkeakoulu) är praktiskt inriktade.
När du utexamineras från en yrkeshögskola får du ofta ett yrke.
Vid yrkeshögskolorna studerar du på finska, svenska eller på engelska.
Vid många yrkeshögskolor finns engelskspråkiga utbildningsprogram.
Ansökan
Du kan söka till en yrkeshögskola då du har avlagt en yrkesskola, gymnasiet eller studentexamen i Finland eller i ett annat land.
Läs mer på InfoFinlands sida Ansökan till utbildning.
Gemensam ansökan till yrkeshögskolorfinska _ svenska
Studier
I yrkeshögskolor kan du studera inom många områden.
Inom parentes anges exempel på yrken som du studera till i olika studieområden:
Naturbruk- och miljöområdet (skogsbruksingenjör, landskapsplanerare)
Den humanistiska och pedagogiska branschen (teckenspråkstolk)
Kulturbranschen (musiker, inredningsarkitekt)
Turism- och kosthållsbranschen (hovmästare, hotellmedarbetare)
Social-, hälso- och idrottsområdet (barnmorska, fysioterapeut, sjuksköterska)
Samhällsvetenskaper, affärsekonomi och förvaltning (försäljningsförhandlare, marknadsföringsassistent)
Teknik och trafik (ingenjör inom bilteknik, maskinmästare i sjöfartsbranschen)
Heltidsstudierna pågår ungefär fyra år.
Studietiden beror på utbildningsprogrammet och din egen studietakt.
Studierna omfattar mycket praktiska övningar.
Studierna omfattar också en arbetspraktik.
Grundläggande information om yrkeshögskolorfinska _ svenska
linkkiUndervisnings- och kulturministeriet:
Förteckning över yrkeshögskolorfinska _ svenska
linkkiSAMOK:
Förbund för studerande vid yrkeshögskolorfinska _ svenska
Förberedande utbildning för invandrare
Yrkeshögskolan kan ordna avgiftsfri utbildning för invandrare med målet att ge den studerande tillräckliga språkkunskaper och andra färdigheter som behövs för att studera vid yrkeshögskolan.
Under studierna tränar studeranden sig i det finska språket, på att läsa saktexter och på sina studiefärdigheter.
Dessutom får studerandena information om utbildningsområdet, arbetsmöjligheter och studier som leder till examen.
Språkkunkapskravet för dem som söker till förberedande utbildning är oftast finskakunskaper på nivån B1 eller B2.
Öppna yrkeshögskolor
De öppna yrkeshögskolorna tillhandahåller yrkeshögskolekurser.
Vem som helst kan studera vid en öppen högskola.
Du kan studera vid en öppen yrkeshögskola även om du inte har någon examen.
Läs mer på InfoFinlands sida Studier som hobby.
Fortsatta studier vid yrkeshögskolor
Om du vill fördjupa dina yrkeskunskaper kan du avlägga högre yrkeshögskoleexamen (ylempi ammattikorkeakoulututkinto).
Den är avsedd för personer som har examen till exempel från en yrkeshögskola och som redan arbetar.
Du kan ansöka till högre yrkeshögskolestudier om du har
någon annan högskoleexamen
minst tre års arbetserfarenhet från en lämplig bransch
Sök till högre yrkeshögskolestudier i den gemensamma ansökan.
Gemensam ansökan ordnas två gånger per år, på hösten och på våren.
Läs mer om den gemensamma ansökan på InfoFinlands sida Ansökan till utbildning.
Du avlägger en högre yrkeshögskoleexamen på ungefär ett eller ett och ett halvt år.
Studiernas omfattning är 60 eller 90 studiepoäng.
Genom högre högskoleexamen kan du fördjupa och utvidga dina kunskaper inom ditt eget yrkesområde.
Till exempel sjukskötare kan avlägga högre yrkeshögskoleexamen inom rehabilitering.
Du kan också välja att avlägga en engelskspråkig examen.
Information om högre yrkeshögskoleexamenfinska _ svenska
Vägledning i högskolestudier
Vid högskolornas SIMHE-tjänster kan du söka hjälp och information om högskoleutbildning i Finland och om hur du ansöker till högskoleutbildning.
Du kan även få information om andra utbildningsmöjligheter för personer som avlagt högskolestudier.
Du kan få vägledning via SIMHE-tjänsterna om
du har flyttat till Finland
du är intresserad av högskolestudier och
du har avlagt högskolestudier eller högskoleexamen utomlands.
Vägledning kan ges individuellt eller i grupp.
linkkiUtbildningsstyrelsen:
Högskolor som erbjuder SIMHE-tjänsterfinska _ svenska _ engelska
Yrkesutbildning ger den studerande behörighet till ett visst yrke.
Därför är utbildningen mycket praktikorienterad.
Du kan söka till en yrkesutbildning när du har avlagt lärokursen för den grundläggande utbildningen.
Även vuxna kan utbilda sig till ett nytt yrke eller komplettera sin kompetens.
Din grundutbildning avgör till hurudan yrkesutbildning du kan söka och på vilket sätt ansökan sker.
Om du har avlagt grundskolans lärokurs kan du ansöka till grundskolebaserad yrkesutbildning (peruskoulupohjainen ammatillinen koulutus).
Om du har avlagt gymnasiet kan du ansöka till gymnasiebaserad yrkesutbildning (lukiopohjainen ammatillinen koulutus).
Om du vill avlägga examen vid sidan av arbetet kan du ansöka till yrkesutbildning för vuxna (ammatillinen aikuiskoulutus).
Läs mer på InfoFinlands sida Ansökan till utbildning.
När du har avlagt yrkesinriktad grundexamen kan du söka dig till fortsatta studier antingen inom yrkesinriktad tilläggsutbildning, vid en yrkeshögskola eller vid ett universitet.
Grundläggande information om yrkesutbildningfinska _ svenska _ engelska
linkkiUtbildningsstyrelsen:
Ytterligare information om yrkesutbildningfinska _ svenska _ engelska
Gemensam ansökan till gymnasier och yrkesläroanstalterfinska _ svenska
Antagning enligt prövningfinska _ svenska
Utbildningsområden i yrkesutbildningenfinska _ svenska
Förberedande för yrkesutbildning
Utbildning som handleder för grundläggande yrkesutbildning (Ammatilliseen peruskoulutukseen valmentava koulutus) d.v.s. VALMA är avsedd för dem som vill avlägga en grundläggande yrkesutbildning.
Under VALMA-utbildningen får du kunskap och färdigheter som hjälper dig i dina senare yrkesinriktade studier.
Du kan även förbättra din språkkunskap. Du kan också höja dina grundskolebetyg.
VALMA-utbildningen räcker ett läsår.
Läs mera på InfoFinlands sida Utbildning som handleder för yrkesutbildning.
Yrkesinriktad grundexamen
Yrkesutbildning ges av yrkesläroanstalter (ammatillinen oppilaitos), specialyrkesläroanstalter (erityisammattioppilaitos) och av vuxenläroanstalter (aikuisopisto).
Du kan avlägga en yrkesinriktad grundexamen antingen
Inom den grundläggande utbildningen (ungdomar och vuxenstuderande)
Som fristående examen (näyttötutkinto) (vuxenstuderande)
Genom läroavtalsutbildning (oppisopimuskoulutus) (ungdomar och vuxenstuderande)
En yrkesinriktad grundexamen ger dig den grundläggande kompetensen i ett visst yrke.
En grundskolebaserad utbildning varar i cirka tre år.
Du kan också studera vid en yrkesläroanstalt och ett gymnasium samtidigt.
Då kan du avlägga en dubbelexamen (kaksoistutkinto).
Vid yrkesskolorna finns många olika områden som du kan studera.
pedagogiska områden
humanistiska och konstnärliga områden
samhälleliga områden
handel och förvaltning
naturvetenskaper
databehandling och datakommunikation
tekniska områden
jord- och skogsbruksområden
hälso- och välbefinnandeområden
Personlig utvecklingsplan för kunnandet
För varje studerande upprättas en personlig utvecklingsplan för kunnandet (PUK).
I planen nedtecknas vilket kunnande du har förvärvat tidigare och fastställs vilka studier du ska avlägga.
Du kan avlägga studierna i egen takt och påvisa vad du kan i praktiska uppgifter på arbetsplatser.
Utbildningsavtal
Utbildningsavtalet är inlärning i arbetet.
Om du vill skaffa dig praktiska kunskaper på en arbetsplats, är ett utbildningsavtal ett bra alternativ för ett läroavtal.
För utbildningstiden betalas ingen lön.
Utbildningsavtalet kan även kombineras med läroavtal.
Yrkesutbildning efter gymnasiet
Om du har avlagt gymnasiet eller studentexamen, kan du söka till en gymnasiebaserad utbildning.
Då kan du inte söka till en grundskolebaserad yrkesutbildning.
Läs mer på InfoFinlands sida Ansökan till utbildning.
Yrkesutbildning för vuxna
Om du arbetar kan du avlägga en yrkesexamen flexibelt vid sidan om arbetet.
Yrkesutbildning för vuxna omfattar
yrkesinriktade grundexamina
yrkesexamina
specialyrkesexamina.
I utbildningen beaktas din tidigare utbildning och den kunskap som du inhämtat som arbetstagare eller företagare.
Du hittar närmare information om hur du kan söka till en yrkesinriktad vuxenutbildning på InfoFinlands sida Ansökan till utbildning.
Examen vid sidan av arbetet med läroavtal
Läroavtal (oppisopimus) innebär inlärning i arbetet.
Du arbetar på en arbetsplats inom din egen bransch och avlägger examen vid sidan av arbetet.
Genom läroavtalsutbildning kan du avlägga samma examen som vid yrkesläroanstalter.
Yrkesexamen (ammattitutkinto)
Specialyrkesexamen (erityisammattitutkinto)
För att kunna studera genom läroavtal måste du ha en arbetsplats.
Du måste hitta en arbetsgivare som vill anställa dig.
Du kan inte inleda din läroavtalsutbildning om du inte har en arbetsplats.
Arbets- och näringsbyrån (TE-toimisto) kan hjälpa dig att hitta ett jobb.
Läroavtalsplatsen kan också vara din nuvarande arbetsplats.
När du har en arbetsplats ska du kontakta läroavtalsbyrån (oppisopimustoimisto) i din region.
Du kan också kontakta en läroanstalt som tillhandahåller läroavtalsutbildning.
Läroavtalsutbildning ges till exempel vid många vuxenutbildningscentra (aikuiskoulutuskeskus).
Under läroavtalsutbildningen betalar arbetsgivaren dig en lön som motsvarar minst en praktikantlön.
Om din arbetsgivare inte betalar dig lön för den tid som du använder för teoretiska studier har du möjligtvis rätt att ansöka om dagpenning, reseersättning och familjebidrag om du omfattas av Den sociala tryggheten i Finland.
Fråga mer vid din läroanstalt.
Information om läroavtalsutbildningfinska _ svenska
Information om läroavtalsutbildningfinska
Kontaktuppgifter till läroavtalsbyråerfinska
linkkiUtbildningsstyrelsen:
Information om läroavtalsutbildningfinska
Bevis för yrkeskunnighet med fristående examen
Fristående examen (näyttötutkinto) är ett sätt att bevisa sin yrkeskunnighet.
Genom fristående examen kan du avlägga
Yrkesexamen (ammattitutkinto)
Yrkesexamen och specialyrkesexamen ger dig behörighet till ett visst yrke.
Dessa examina avläggs alltid genom fristående examen.
Fristående examen är ett lämpligt alternativ också om du har avlagt en yrkesexamen i något annat land och vill jämställa den med en finsk examen.
Om du vill avlägga en fristående examen ska du ta kontakt direkt med läroanstalten.
Fristående examina kan avläggas vid yrkesläroanstalter och vuxenläroanstalter.
För fristående yrkesexamen finns ingen bestämd ansökningstid.
Du avlägga fristående examen vid ett examenstillfälle (tutkintotilanne) där en representant för läroanstalten intygar din yrkeskunnighet.
Sedan får du ett yrkesbevis som bevisar din yrkeskunnighet.
linkkiUtbildningsstyrelsen:
Information om fristående examenfinska _ svenska _ engelska
Yrkesutbildning som anordnas av arbetsgivaren
En del arbetsgivare utbildar människor till arbeten hos dem.
Dessa arbetsgivare ger garanti om en arbetsplats.
Det betyder att den som avlägger utbildningen får en arbetsplats hos arbetsgivaren.
Du får alltså både yrkesutbildning och en arbetsplats.
Till exempel många trafikföretag och VR utbildar de personer som de anställer.
Utbildningen i Finland håller en hög kvalitet.
Skillnaderna i olika skolors studieresultat är små och nästan alla avlägger grundskolan inom den utsatta tiden.
Förskoleundervisning, grundläggande utbildning och utbildning på andra stadiet är kostnadsfria och även därefter är utbildningen till största delen kostnadsfri.
Målet är att alla, oavsett familjens inkomster, ska ha möjlighet att få en högklassig utbildning och växa till aktiva medborgare.
Utbildningssystemet omfattar småbarnspedagogik, förskoleundervisning, grundläggande utbildning, utbildning på andra stadiet och högskoleutbildning.
Vuxenutbildningen är avsedd för vuxna och innehåller många alternativ från grundläggande utbildning till högskoleutbildning.
Småbarnspedagogik
I Finland har barnen rätt till småbarnspedagogik före skolåldern.
Småbarnspedagogiken ordnas i daghem och familjedagvården.
Barnet kan även delta i småbarnspedagogik tillsammans med föräldern i lekparker.
Barnet kan få minst 20 timmar småbarnspedagogik i veckan eller mer om föräldrarna arbetar eller struderar.
Målet är att stödja barnets utveckling och välbefinnande.
Barnet lär sig bland annat sociala färdigheter, att göra saker med händerna och olika kunskaper.
Barnet lär sig också olika färdigheter som hjälper hen att lära sig ytterligare nya saker.
Dagarna innehåller mycket lek och utevistelser.
Om barnet har ett annat modersmål än finska eller svenska, får hen stöd i lärandet av finska eller svenska.
Om barnet behöver, kan hen även få specialundervisning.
I Finland ordnar kommunerna småbarnspedagogiken.
Den finansieras med skattemedel och är därför förmånligare för familjerna.
I Finland finns även privat småbarnspedagogik.
De som arbetar med barnen är utbildade pedagoger inom småbarnsfostran och barnskötare.
Förskoleundervisning
I Finland ska barnen delta i förskoleundervisning under ett års tid innan läroplikten börjar.
Vanligtvis börjar förskoleundervisningen det år då barnet fyller sex år.
Förskoleundervisningen ordnas av kommunerna och är kostnadsfri för familjen.
Förskoleundervisningen ges av pedagoger inom småbarnsfostran som har avlagt universitetsexamen.
Förskoleundervisning ges vanligtvis fyra timmar om dagen från måndag till fredag.
Om föräldrarna arbetar eller studerar kan barnet utöver förskoleundervisningen även delta i småbarnspedagogiken.
Under detta år lär sig barnet kunskaper som hen har nytta av i skolan, till exempel bokstäver.
Barnen undervisas dock inte ännu i läsning.
Om barnet har ett annat modersmål än finska eller svenska, får hen stöd i lärandet av finska eller svenska.
Till dagen hör också lek och utevistelse.
Läs mer på InfoFinlands sida Förskoleundervisning.
Grundläggande utbildning
I Finland börjar den grundläggande utbildningen det år då barnet fyller sju år.
Alla barn som har sitt stadigvarande boende i Finland måste delta i den grundläggande utbildningen.
Grundskolan har nio årskurser.
Läroplikten upphör när barnet har fullgjort hela lärokursen för den grundläggande utbildningen eller det har förflutit tio år sedan läroplikten började.
I Finland reglerar lagstiftningen den grundläggande utbildningen.
Dessutom används nationella läroplansgrunder och lokala läroplaner.
Den grundläggande utbildningen ordnas av kommunerna.
Den finansieras med skattemedel och är därför kostnadsfri för familjerna.
I de lägre årskurserna har man cirka 20 undervisningstimmar i veckan och antalet ökar i de högre årskurserna.
Alla grundskolelärare i Finland har magisterexamen.
Klasslärarna i grundskolan, som undervisar årskurserna 1–6, har läst pedagogik.
Lärarna i årskurserna 7–9 har läst det ämne som de undervisar.
Lärare har stor frihet att planera undervisningen självständigt utifrån den nationella och lokala läroplanen.
På sistone har man i läroplanen betonat bland annat helheter som omfattar flera läroämnen, undersökning av vardagliga fenomen samt data- och kommunikationsteknik.
Barnen har ofta en och samma lärare under de sex första skolåren.
Läraren lär känna eleverna bra och kan utveckla undervisningen så att den passar dem.
Ett viktigt mål är att eleverna lär sig att tänka självständigt och tar eget ansvar för sitt lärande.
Läraren bedömer elevernas framsteg i skolan.
I den grundläggande utbildningen ges alla vitsord av läraren.
Det finns inga egentliga nationella prov.
Däremot följs inlärningsresultaten upp med urvalsbaserade bedömningar.
Dessa ordnas oftast i årskurs nio.
Om barnet eller den unga har flyttat till Finland nyligen, kan hen få förberedande undervisning före den grundläggande utbildningen.
Den förberedande undervisningen varar vanligtvis ett år.
Därefter kan eleven fortfarande läsa finska eller svenska som andraspråk, som S2-språk, om hen behöver stöd med språket.
Vuxna invandrare som inte har grundskolans avgångsbetyg från sitt eget land kan avlägga grundskolan på vuxengymnasiet.
Läs mer om den grundläggande utbildningen på InfoFinlands sida Grundläggande utbildning.
Utbildning på andra stadiet
De vanligaste alternativen efter grundskolan är gymnasium och yrkesutbildning.
Dessa är utbildning på andra stadiet.
Utbildning på andra stadiet är oftast kostnadsfri för studeranden.
Böcker och annat studiematerial måste man dock köpa själv.
Gymnasium
Gymnasiet är en allmänbildande utbildning som inte ger ett yrke.
I gymnasiet läser man samma ämnen som i den grundläggande utbildningen, med undervisningen är mer krävande och studierna mer självständiga.
På slutet avlägger studerandena vanligtvis studentexamen.
Gymnasiet tar 2–4 år, beroende på den studerande.
Efter gymnasiet kan man söka till universitet, yrkeshögskola eller gymnasiebaserad yrkesutbildning.
I de flesta gymnasieskolorna är undervisningsspråket finska eller svenska.
I de stora städerna finns några gymnasieskolor med något annat undervisningsspråk, till exempel engelska eller franska.
Vuxna kan avlägga gymnasiestudier på vuxengymnasiet.
Där kan man avlägga enskilda kurser eller hela gymnasielärokursen och studentexamen.
Undervisningen kan bestå av närundervisning, distansundervisning, webbundervisning och självständiga studier.
Läs mer om gymnasiestudierna på InfoFinlands sida Gymnasium.
Förberedande gymnasieutbildning
På gymnasiet behövs goda språkkunskaper.
Om studeranden har ett annat modersmål än finska eller svenska och saknar tillräckliga språkkunskaper för gymnasiestudierna, kan hen söka till förberedande gymnasieutbildning (LUVA).
Läs mer på InfoFinlands sida Förberedande gymnasieutbildning.
Yrkesutbildning
Yrkesutbildningen är mer praktiknära än gymnasieutbildningen.
En yrkesinriktad grundexamen kan avläggas på ungefär tre år.
Därefter kan man fortsätta studierna och avlägga yrkesexamen eller specialyrkesexamen.
En väsentlig del av studierna är inlärning på arbetsplatsen.
Om man vill, kan man efter yrkesutbildningen fortsätta studierna ända till högskoleutbildning.
Om man redan behärskar de färdigheter som krävs för examen, kan man också avlägga yrkesexamen eller specialyrkesexamen som yrkesprov.
Yrkesexamen kan även avläggas med läroavtal.
Då arbetar studeranden på en arbetsplats inom den egna branschen, får minst samma lön som en praktikant för arbetet och avlägger samtidigt sina studier.
Läs mer på InfoFinlands sida Yrkesutbildning.
Utbildning som handleder för yrkesutbildning
Om du inte har tillräckliga språkkunskaper eller studiefärdigheter för yrkesutbildning, kan du före yrkesutbildningen söka till utbildning som handleder för yrkesutbildning (VALMA).
Läs mer på InfoFinlands sida Utbildning som handleder för yrkesutbildning.
Högskoleutbildning
Efter studierna på andra stadiet kan du gå vidare till högskoleutbildning.
I Finland tillhandahålls högskoleutbildning av yrkeshögskolor och universitet.
Studierna på yrkeshögskola kan vara kostnadsfria eller avgiftsbelagda för studeranden.
Terminsavgift tas ut av personer som inte är medborgare i ett EU-/EES-land eller familjemedlem till en medborgare i ett EU-/EES-land och som avlägger en lägre eller högre högskoleexamen på engelska.
Läs mer på InfoFinlands sida Utländska studerande i Finland.
Yrkeshögskolor
På yrkeshögskolan är undervisningen mer praktiknära än på universitetet.
I undervisningen ingår även inlärning i arbetet.
Yrkeshögskoleexamen kan avläggas på 3,5–4,5 år.
Om man vill fortsätta studierna därefter och avlägga högre yrkeshögskoleexamen, måste man först skaffa sig tre år av arbetserfarenhet från samma område som examen.
Läs mer på InfoFinlands sida Yrkeshögskolor
Undervisningen på universitet är baserad på vetenskaplig forskning.
På universitet kan man avlägga lägre högskoleexamen på cirka tre år och därefter högre högskoleexamen på cirka två år.
Universiteten ordnar undervisning på engelska i vissa utbildningsprogram.
I de flesta utbildningsprogrammen är undervisningsspråket ändå finska eller svenska.
När man har avlagt magisterexamen, kan man ansöka om rätt till fortsatta studier och avlägga licentiat- eller doktorsexamen.
Läs mer på InfoFinlands sida Universitet.
Ansökan till utbildning
På InfoFinlands sida Ansökan till utbildning finns information om hur du ansöker till utbildning på andra stadiet och högskoleutbildning i Finland.
Om du planerar att studera i Finland, läs mer på InfoFinlands sida Utländska studerande i Finland och Studerande.
Andra studiemöjligheter
I Finland finns även många läroanstalter som erbjuder studier som inte leder till examen för människor i alla åldrar.
Största delen av dessa utbildningar är avsedda för vuxna.
Sådana läroanstalter är medborgarinstitut, folkhögskolor, sommaruniversitet, studiecenter och idrottsutbildningscenter.
Studierna är allmänbildande.
Du kan studera till exempel bland annat språk, estetiska ämnen, handarbete och kommunikation.
Oftast betalar den studerande en avgift för studierna.
I vissa situationer kan studierna vid dessa läroanstalter dock vara kostnadsfria.
Om till exempel utbildning i läs- och skrivkunnighet eller någon annan språkutbildning har godkänts till din integrationsplan, tas det inte ut någon avgift för studierna.
Språkutbildning
Om du vill läsa finska eller svenska, läs mer på InfoFinlands sida Finska och svenska språket.
Efter grundskolan (peruskoulu), d.v.s. efter grundstadiet fortsätter studerandena till läroanstalter på andra stadiet (toisen asteen oppilaitos).
Läroanstalter på andra stadiet är gymnasiet och yrkesläroanstalter.
Läs mer om yrkesläroanstalter på InfoFinlands sida Yrkesutbildning.
Gymnasiestudierna är mer teoretiskt inriktade än yrkesutbildning.
Studierna är allmänbildande: fokus ligger speciellt på naturvetenskapliga och humanistiska ämnen.
I vissa gymnasier ges även mycket undervisning i konstämnen.
Vissa gymnasier är specialgymnasier.
De är inriktade på till exempel musik, idrott eller naturvetenskaper.
Specialgymnasierna är mycket populära.
Det kan vara svårt att komma in dit.
Gymnasiet ger förberedande utbildning till exempel för yrkeshögskola och universitet.
Både ungdomar och vuxna kan studera vid gymnasiet.
Ungdomarna studerar vid daggymnasiet (päivälukio) eller distansgymnasiet (etälukio), vuxna studerar ofta vid vuxengymnasiet (aikuislukio).
Information om gymnasiestudierfinska _ svenska
linkkiFörbund för gymnasieelever:
Förbund för gymnasieeleverfinska _ svenska _ engelska
linkkiUtbildningsstyrelsen:
Information om gymnasiestudierfinska _ svenska _ engelska
Att söka till gymnasiet
Sök till gymnasiet i den gemensamma ansökan till andra stadiet.
Om du vill studera vid ett vuxengymnasium ska du ta kontakt direkt med läroanstalten.
Läs mer på InfoFinlands sida Ansökan till utbildning.
Gemensam ansökan till gymnasier och yrkesläroanstalterfinska _ svenska
Att studera vid gymnasiet
Gymnasiestudierna pågår vanligen tre år.
Gymnasiet kan också avläggas på två eller fyra år.
I gymnasiestudierna har du många valmöjligheter.
Utöver de obligatoriska kurserna kan du välja många kurser som passar dig.
I gymnasiet påverkar du själv innehållet i dina studier och din studietakt.
I gymnasiet tas inga terminsavgifter ut.
Utbildningen kostar alltså inget.
Studeranden måste dock själv skaffa gymnasieböckerna.
Böckerna är ofta dyra.
Man kan även köpa gymnasieböckerna begagnade.
Om du till exempel har en krävande hobby eller är sjuk en lång tid kan du avlägga gymnasiet som distansstudier.
Fråga mer om distansstudier vid ditt eget gymnasium.
Studentexamen
Gymnasiestudierna siktar till studentexamen (ylioppilastutkinto).
Studentexamen består av prov i olika läroämnen.
Studentskrivningarna (ylioppilaskokeet) skrivs oftast i slutet av studierna.
Modersmålsprovet är ett obligatoriskt prov i studentexamen.
Modersmålsprovet kan skrivas i finska, svenska eller samiska.
Om du inte har finska, svenska eller samiska som modersmål kan du skriva ett prov i finska eller svenska som andra språk.
Utöver modersmålsprovet måste du skriva prov i minst tre andra ämnen.
Om du vill kan du även skriva fler ämnen.
Utöver modersmålsprovet kan du skriva prov i följande andra ämnen:
Det andra inhemska språket (finska eller svenska)
Ett främmande språk: engelska, tyska, ryska, franska, spanska, portugisiska, latin
Matematik
Realämnen (reaali), d.v.s. historia, religion, fysik, kemi, biologi, psykologi, filosofi
Studentskrivningarna ordnas på våren och på hösten.
Om du vill kan du skriva några ämnen på hösten och resten på våren.
Du måste skriva alla prov på högst tre efter varandra följande examenstillfällen.
Info om studentexamenfinska _ svenska
linkkiStudentexamensnämnden:
Information om studentexamenfinska _ svenska _ engelska _ franska _ tyska
Vuxengymnasium
Vuxengymnasiet är i huvudsak avsett för personer som har fyllt 18 år.
Vid vuxengymnasiet är studierna flexibla.
Du kan avlägga hela studentexamen eller bara studera ett ämne.
Undervisningen sker oftast kvällstid.
Många vuxengymnasier erbjuder finskakurser för invandrare.
Fråga om kurserna direkt vid vuxengymnasiet.
Information om vuxengymnasietfinska _ svenska
linkkiEdu.fi:
Enligt lag ska barn i Finland delta i förskoleundervisning eller motsvarande verksamhet under ett års tid innan läroplikten börjar.
Förskoleundervisningen (esiopetus) förbereder barnen inför grundskolan.
Barnen börjar i förskoleundervisningen vanligen vid sex års ålder och grundskolan vid sju års ålder.
Föräldrarna anmäler sitt barn till förskoleundervisningen vanligtvis i januari eller februari.
Kontrollera tidpunkten i god tid vid skolväsendet (koulutoimi) eller bildningsväsendet (sivistystoimi) i din hemkommun.
Kommunerna ordnar förskoleundervisning.
De kan även köpa förskoleundervisningen till exempel av ett privat daghem.
Förskoleundervisningen är kostnadsfri.
Under dagen får barnet en gratis måltid.
Om barnet bor långt (över 5 km) från undervisningsstället, eller om vägen dit är besvärlig, får barnet gratis skjuts.
Om föräldrarna arbetar eller studerar kan barnet utöver förskoleundervisningen även delta i småbarnspedagogiken.
En dag i förskolan
Förskoledagen är ungefär fyra timmar lång.
Förskolan finns ofta antingen i daghemmets eller skolans lokaler.
I förskolan lär sig barnen bland annat matematik, miljö- och naturkunskap samt konst och kultur.
De lär sig nya saker med lekens hjälp.
Föräldrarna har en viktig roll i förskolan.
De stödjer sitt barns inlärning.
Lärarna utarbetar en egen inlärningsplan för varje barn.
Föräldrarna kan hjälpa ledarna att utarbeta planen.
Språk och kulturer i förskoleundervisningen
Ett barn som har ett annat modersmål än finska eller svenska lär sig finska eller svenska som främmande språk.
Dessutom kan det studera sitt eget modersmål om kommunen ordnar undervisning i det språket.
Barnet kan även få undervisning i den egna religionen eller i livsåskådningskunskap i förskolan.
I förskolan lär sig barnen att uppskatta sitt språk och sin kultur.
De lär sig också att respektera andra människors språk och kulturer.
linkkiUtbildningsstyrelsen:
Information om förskoleundervisningenfinska _ svenska _ engelska
Förskoleuppgifter på nätetfinska
linkkiUndervisnings- och kulturministeriet:
Information om förskoleundervisningenfinska _ svenska _ engelska
Brandsäkerhet
En brandvarnare kan rädda ditt liv.
Om en brand uppstår i din bostad avger brandvarnaren ett högljutt larm och du hinner ut i tid.
Se till att det finns tillräckligt många brandvarnare i ditt hem.
Brandvarnare säljs i varuhus och järnaffärer.
En brandvarnare räcker till 60 kvadratmeter.
Om ditt hem är till exempel 65 kvadratmeter stort behöver du två brandvarnare.
Om ditt hem har fler än en våning måste du räkna ytan separat för varje våning.
Det bör finnas en brandvarnare på varje våning.
Kontrollera regelbundet att brandvarnaren fungerar.
Byt batterier vid behov, gärna en gång per år.
Du ansvarar för brandvarnaren även om du bor i en hyresbostad.
Det finns ofta en bastu i finländska hem.
Även om du inte använder bastun får du aldrig placera något på bastuugnen, eftersom detta kan orsaka en brand.
Torka till exempel inte tvätten ovanför eller i närheten av bastuugnen.
Stäng alltid av en elektrisk bastuugn efter användning.
När du går hemifrån, kom ihåg att kontrollera att spisen och ugnen och till exempel strykjärnet är avstängda.
Det är bra att ha en brandsläckare hemma.
I vissa höghus finns det också en brandsläckare i trappuppgången.
Ta reda på var den närmaste brandsläckaren finns.
Se till att du har en släckningsfilt hemma.
Det är bra att förvara filten till exempel i närheten av spisen.
Lämna inte mat på en het spis utan uppsikt.
Var särskilt försiktig om du lagar mat på natten.
Laga inte mat om du är berusad.
Förvara inte föremål på spisen.
Barn, husdjur eller du själv kan av misstag vrida på spisen.
Då kan sakerna som ligger på spisen fatta eld.
Om fett börjar brinna när du lagar mat, kväv elden med till exempel ett kastrullock eller med en släckningsfilt.
Använd inte vatten.
Kom ihåg att stänga av elapparater efter användning.
Strykjärnet ska också kopplas loss från vägguttaget.
Använd inte elapparater som är i dåligt skick eller vars sladd är trasig.
Om en elapparat börjar brinna, använd inte vatten.
Kväv elden med till exempel en brandsläckare.
Om du har elektriska värmeelement eller värmeaggregat hemma, lägg inte tyger, kläder eller något annat på dem.
Lämna utrymme runt TV:n, mikrovågsugnen, kylskåpet och frysen.
Täck inte över dem.
Det är bra att en gång per år städa bort damm från frysens och kylskåpets bakgaller till exempel med dammsugaren, om möjligt.
Rök inte inomhus.
Lämna inte brinnande ljus utan uppsikt.
Tänd inte ljus i närheten av till exempel gardinerna, ens om du själv är i rummet.
Om en brand uppstår, ring nödnumret 112.
linkkiHelsingfors stads räddningsverk:
Brandsäkerhet i höghusfinska _ svenska _ engelska
linkkiRäddningsbranschens Centralorganisation i Finland:
Information om brandsäkerhetfinska _ svenska _ engelska
linkkiHelsingfors stad, Förortsprojektet:
Mitt hem i ett höghus(pdf, 6,56 MB)finska _ engelska _ ryska _ somaliska _ arabiska
linkkiHelsingfors stads räddningsverk:
Brandsäkerhet i småhusfinska _ svenska _ engelska
Så här undviker du vattenskador
Lämna inte tvättmaskinen eller diskmaskinen på när du går hemifrån.
Kontrollera regelbundet att vattenledningarna i ditt hem inte läcker och att det inte rinner ut vatten från hushållsapparaterna på golvet.
Stäng alltid kranen till tvätt- och diskmaskinen när du inte använder dem.
Det ska finnas ett läckageskydd av plast under kylskåpet, frysen och diskmaskinen.
Skyddet läggs på plats samtidigt som apparaten installeras.
Du får inte installera en diskmaskin själv, utan arbetet måste utföras av en fackman.
Om ett vattenläckage uppstår i ditt hem, försök stänga vattenledningens avstängningsventil.
Om du bor i höghus eller radhus, anmäl läckaget genast till journumret för husets servicebolag.
Om du bor i villa, kontakta en jourhavande rörfirma.
Elarbeten
I Finland är nätspänningen 230 volt.
I Finland utförs egentliga elarbeten endast av personer som är yrkesutbildade inom elbranschen.
Vissa små elarbeten får du utföra själv, om du kan.
Du kan till exempel själv:
byta en säkring
byta lampor
reparera en enfas skarvsladd (spänning 230 V)
hänga upp en lampa i taket med en upphängningsbygel
byta en hel enfas anslutningsledning (spänning 230 V) och stickkontakt i en elapparat, om den gamla gått sönder.
linkkiTukes:
Elarbeten som du får göra självfinska _ svenska _ engelska
Säkerhetslås skyddar mot inbrottstjuvar
Om du har ett säkerhetslås i ditt hem, lås det alltid då du inte är hemma.
Lås inte säkerhetslåset när du är hemma.
Om någon bryter in sig i ditt hem, ring nödnumret 112.
linkkiTukes:
Guiden Ett säkert hem för barnfinska _ svenska _ engelska
Birkalands räddningsverk:
Vad gör jag om det börjar brinna hemma?
Om videon väcker frågor hos dig kan du fråga mer av en expert.
Utbildning som handleder för grundläggande yrkesutbildning (Ammatilliseen peruskoulutukseen valmentava koulutus) d.v.s. VALMA är avsedd för dem som vill avlägga en grundläggande yrkesutbildning.
Under VALMA-utbildningen får du kunskap och färdigheter som hjälper dig i dina senare yrkesinriktade studier.
Du kan även förbättra din språkkunskap. Du kan också höja dina grundskolebetyg.
VALMA-utbildningen räcker ungefär ett läsår.
Du kan under utbildningen bekanta dig med olika branscher och fundera på vad du vill studera.
Du besöker arbetsplatser och deltar i verkstäder.
I början av utbildningen görs det upp en personlig studieplan för dig.
I den skrivs det in vilka studier du avlägger och hur.
Du får ett betyg för VALMA-utbildningen.
Du får också tilläggspoäng när du ansöker till en yrkesutbildning i den gemensamma ansökan.
VALMA-utbildningen kostar vanligen inget för den studerande.
Information om VALMA-utbildningarfinska _ svenska _ engelska
Ansökan till VALMA-utbildningen
Du kan ansöka till VALMA-utbildningen om du har slutfört grundskolan eller en utbildning som motsvarar grundskolan.
Om läroinrättningen anser att du kan klara av studierna kan du antas som studerande även utan slutbetyg från grundskolan.
Ansök till VALMA-utbildningen efter den egentliga gemensamma ansökan i början av sommaren.
Om du behöver särskilt stöd t.ex. på grund av handikapp ska du ansöka till utbildningen på våren, under ansökan till specialundervisning.
Närmare information om ansökningstiderna hittar du via Studieinfo.fi-tjänsten.
Fyll i ansökningsblanketten i Studieinfo.fi-tjänsten.
Ansökan till VALMA-utbildningfinska _ svenska
Ansökan till specialundervisningfinska _ svenska
Småbarnspedagogik är avsedd för barn under skolåldern.
I Finland tillhandahåller kommunerna kommunal småbarnspedagogik bland annat i daghem.
Dessutom finns det privata daghem.
Småbarnspedagogik är fostran, undervisning och omsorg som är pedagogiskt planerad och som har noga genomtänkta mål.
Inom småbarnspedagogiken arbetar utbildade lärare i småbarnspedagogik och barnskötare.
Vanligen vårdar någondera av föräldrarna barnet hemma åtminstone under föräldraledigheten (vanhempainvapaa), det vill säga tills barnet är ungefär 9 månader gammalt.
Om du vårdar ditt barn hemma även efter detta har du rätt att vara ledig från ditt arbete för vård av barn tills barnet fyller tre år.
Mer information om ledigheterna får du på InfoFinlands sida Familjeledighet.
Du kan ansöka från Kela om ekonomiskt stöd för hemvård av barn.
Läs mer på InfoFinlands sida Stöd för vård av barn i hemmet.
Kommunal småbarnspedagogik
Om du har din hemkommun i Finland, kan du ansöka om en plats inom den kommunala småbarnspedagogiken för barnet efter föräldraledigheten.
Då är barnet ca nio månader gammalt.
Om du inte har en hemkommun i Finland, räknas du som invånare i den kommun där du vistas.
Om båda föräldrarna arbetar, har barnet rätt till småbarnspedagogik på heltid.
Om den ena föräldern är hemma, beror rätten till småbarnspedagogik på hemkommunen.
I vissa kommuner har barnet rätt till småbarnspedagogik på heltid även då den ena föräldern är hemma.
I vissa kommuner har barnet rätt till 20 timmar småbarnspedagogik per vecka om den ena föräldern är hemma.
Familjen kan ändå söka rätt till småbarnspedagogik på heltid om barnet behöver särskilt stöd till exempel i att lära sig det finska språket eller på grund av att familjen befinner sig i en svår situation.
Du kan ansöka om en plats
på ett daghem (päiväkoti)
På daghemmet är barnen i större gruppen är i gruppfamiljedagvården.
Familjedagvård innebär att skötaren vårdar barnen i sitt eget hem.
Vissa familjedagvårdare vårdar barnen hemma hos de barn som ingår i gruppen.
Ansök om en plats inom den kommunala småbarnspedagogiken från din egen kommun senast fyra månader innan du behöver den.
Man kan få en plats inom två veckor, om föräldrarna får ett arbete eller en studieplats.
Avgiften för småbarnspedagogik (varhaiskasvatusmaksu) beror på
familjens inkomster
familjens storlek och
på hur många timmar per vecka barnet deltar i småbarnspedagogik.
Man får syskonrabatt.
Om familjen inkomster är mycket låga, kan småbarnspedagogiken vara kostnadsfri för familjen.
Fråga mer i din kommuns rådgivningstjänster.
Privat småbarnspedagogik
En plats inom den privata småbarnspedagogiken kan finnas
i ett privat daghem eller i ett gruppfamiljedaghem
i familjedagvård eller
hemma, då familjen anställer en skötare i hemmet
Du kan ansöka om en plats inom småbarnspedagogiken direkt från det privata daghemmet eller gruppfamiljedaghemmet.
Du kan också leta upp en privat familjedagvårdare som vårdar barnen hemma hos sig, eller anställa en skötare i ditt eget hem.
Om du anställer en skötare i ditt hem blir du en arbetsgivare, och du måste uppfylla en arbetsgivares skyldigheter.
Läs mera på InfoFinlands sida Arbetsgivarens rättigheter och skyldigheter.
Familjen kan anställa en skötare i sitt hem även tillsammans med en annan familj.
Kommunen övervakar den privata småbarnspedagogiken.
Priserna för den privata småbarnspedagogiken varierar.
Du kan ändå få stöd för den från FPA.
Då är den inte nödvändigtvis mycket dyrare än den kommunala småbarnspedagogiken.
Stöd för privat dagvård
Om barnet har en hemkommun i Finland, kan du ansöka om Fpa-stöd för privat vård.
Dagvårdsproducenten måste ha kommunens godkännande.
Du kan ansöka om privatvårdsstöd (yksityisen hoidon tuki), om
ditt barn som är under skolåldern är i privat dagvård; eller
barnet har någon annan privat skötare.
Du kan inte ansöka om privatvårdsstöd om skötaren är en medlem i barnets familj eller om barnet och skötaren bor i samma hushåll.
Du kan inte heller ansöka om privatvårdsstöd för den kommunala småbarnspedagogiken.
Stödets storlek beror bland annat på familjens inkomster och kommunen som familjen bor i.
Kela betalar stödet direkt till skötaren eller dagvårdsproducenten.
Man måste betala skatt för privatvårdsstödet.
Stödet betalas inte till utlandet.
Läs mera om privatvårdsstöd på Fpa:s sidor.
Fpa har en telefontjänst för barnfamiljer.
på finska tfn +358 (0)20 692 206
på svenska och engelska tfn +358 (0)20 692 226
På Fpas byråer får du betjäning även på andra språk med hjälp av en tolk.
Stöd för privat vårdfinska _ svenska _ engelska
Vad händer i småbarnspedagogiken?
Till småbarnspedagogiken hör mångsidig verksamhet, till exempel lekar, motion, utevistelse, musik, pyssel och utfärder.
I dagen ingår också en vilostund.
Målsättningen med verksamheten är att främja barnets utveckling och lärande.
Barnet lär sig även sociala färdigheter.
Barnet får stöd i att lära sig det finska eller svenska språket, om hans/hennes modersmål är ett annat språk.
Om barnet behöver, kan hen även få specialundervisning.
Daghemmet är ändå inte en skola.
Barnen studerar inte skolämnen och har inte lektioner.
Barnen äter tre måltider under dagen: frukost, lunch och mellanmål.
Om ditt barn har en specialdiet ska du berätta om det för lärarna i småbarnspedagogiken.
I småbarnspedagogiken beaktas familjens religion eller livsåskådning.
På vissa orter finns det daghem, som fungerar på andra språk än finska eller svenska.
Vanligen börjar daghemsdagen på morgonen och tar slut på eftermiddagen.
Vissa daghem och familjedagvårdare har öppet dygnet runt med anledning av föräldrarnas arbete eller studier.
linkkiFinlands Flyktinghjälp:
Klubbar
Kommunerna, föreningar och församlingar ordnar dagklubbar för barn.
Klubbarna räcker vanligen ett par timmar.
I klubbarna ordnas handledda lekar, sång, pyssel och annat program.
linkkiUndervisnings- och kulturministeriet:
Information om småbarnspedagogikfinska _ svenska _ engelska
Söka bostad
Att hyra en bostad
Uppsägning av bostad
Att bli av med sin bostad
Konflikter med grannarna
Boendevardag
Fuktproblem
Rådgivningstjänster
Söka bostad
Jag hittar inte en förmånlig hyresbostad.
I de större städerna finns det bara få lediga hyresbostäder.
Bostäderna är dyrare nära stadens centrum.
Därför bor många finländare i ganska små bostäder.
Många bor också långt från centrum eller i en närliggande kommun och pendlar långt till jobbet.
Om du inte hittar en förmånlig bostad där du vill bo, fundera om du kan tänka dig att bo i en mindre bostad eller längre bort från centrum.
På många mindre orter finns det många lediga bostäder och priserna är lägre.
Om du planerar att flytta från en liten ort till en större stad, leta en bostad i förväg.
Läs mer på InfoFinlands sida Hyresbostad.
Jag lämnade en ansökan om en kommunal hyresbostad men jag har inte fått en bostad fastän det har gått tid.
Det finns inte tillräckligt många kommunala bostäder för alla som ansöker om dem.
Det lönar sig att ansöka om bostad på flera ställen.
Följ också utbudet av privata hyresbostäder.
Kom ihåg att uppdatera din ansökan när den är i kraft. Annars löper den ut.
Läs mer på InfoFinlands sida Hyresbostad.
Jag misstänker att jag har blivit diskriminerad när jag letade efter bostad.
Var får jag hjälp?
Enligt lag får hyresvärdar inte diskriminera någon till exempel på grund av etniskt ursprung, religion eller medborgarskap när de väljer hyresgäster.
En privat hyresvärd har dock rätt att själv välja hyresgästen till bostaden och hen behöver inte motivera sitt val.
Om du misstänker att du har blivit diskriminerad kan du fråga om råd till exempel hos diskrimineringsombudsmannens kundtjänst.
Diskrimineringsombudsmannens kundtjänstfinska _ svenska _ engelska
Att hyra en bostad
Måste jag betala ett förmedlingsarvode till bostadsförmedlaren när jag hyr en bostad?
Oftast betalar hyresvärden förmedlingsarvodet.
Du själv betalar förmedlingsarvodet endast om du har ingått ett skriftligt uppdragsavtal med bostadsförmedlaren om att söka en bostad åt dig.
Om du inte har ingått ett skriftligt uppdragsavtal får bostadsförmedlaren inte kräva dig på förmedlingsarvode.
Om hen försöker göra detta kan du polisanmäla hen.
Läs mer på InfoFinlands sida Brott.
Bostadsförmedlaren kräver att jag betalar hen för att få se bostaden.
Måste jag betala?
Du har rätt att se bostaden i förväg och bostadsförmedlaren kan inte kräva att få betalt för detta.
Om du har problem som rör förmedlingsarvodet kan du kontakta Konsumentrådgivningen.
linkkiKonkurrens- och konsumentverket:
Konsumentrådgivningfinska _ svenska _ engelska
Bostadsförmedlaren kräver att jag betalar en reservationsavgift för hyresbostaden.
Måste jag betala?
I Finland tillämpas inga reservationsavgifter för bostäder.
Du ska inte betala någonting förrän du har ett skriftligt hyresavtal för bostaden.
Läs mer om avgifterna för en hyresbostad, till exempel hyresdeposition, på InfoFinlands sida Hyresavtal.
Hyresvärden kräver att jag tecknar en hemförsäkring.
Var får jag en hemförsäkring?
Kan jag säga upp den senare?
Hemförsäkringar säljs av många försäkringsbolag i Finland.
Läs mer på InfoFinlands sida Vardagslivet i Finland.
Det är bra att teckna en hemförsäkring även om det inte krävs i hyresavtalet.
Det är inte tillrådligt att säga upp hemförsäkringen under tiden då du bor i bostaden.
Om du till exempel orsakar en vattenskada måste du själv betala hela renoveringskostnaden.
Fakturan kan uppgå till flera tiotusentals euro.
Vad bör jag beakta innan jag undertecknar hyresavtalet?
Gå och titta på bostaden innan du hyr den.
Kontrollera att bostaden verkligen existerar, alltså att bostaden har samma adress som står på avtalet.
Säkerställ också att bostaden är i det skick som har angetts till dig.
Kontrollera vad hyresavtalet säger till exempel om villkoren för hyresförhållandet och om uppsägningstiden.
Det är också bra att gå igenom bostaden och eventuella fel i bostaden med dess ägare eller hens representant.
Läs mer på InfoFinlands sida Hyresavtal.
När ska jag betala hyresdepositionen?
Betala hyresdepositionen först när du har ett skriftligt hyresavtal.
Hyresvärden kan ange ett konto på vilket du sätter in hyresdepositionen.
Ni kan också öppna ett separat konto för hyresdepositionen på banken.
Läs mer på InfoFinlands sida Hyresavtal.
Hyresvärden föreslog att vi gör ett muntligt hyresavtal.
Är ett muntligt avtal tillräckligt?
Gör hyresavtalet alltid skriftligt.
På så sätt kan du bevisa vad ni kommit överens om, om det skulle uppstå problem.
Förvara hyresavtalet noga.
Det finns brister i hyresbostaden.
Kan hyresvärden i efterhand kräva att jag ersätter för brister som jag inte har orsakat?
Det är bra att skriva upp felen i bostaden tillsammans med hyresvärden när hyresförhållandet inleds.
Du kan även ta fotografier där felen syns.
På så sätt säkerställer du att du inte ställs ansvarig för fel som du inte har orsakat.
Uppsägning av bostad
Jag sade upp min hyresbostad men hyresvärden kräver att jag betalar hyran tills hen hittar en ny hyresgäst.
Måste jag betala?
Om du har ett tills vidare gällande hyresavtal är uppsägningstiden vanligtvis en kalendermånad.
Tiden räknas från slutet av den månad då du säger upp avtalet.
När uppsägningstiden har löpt ut kan hyresvärden inte kräva dig på hyra.
Ett tidsbestämt hyresavtal får inte sägas upp under dess löptid.
Vid behov kan du försöka förhandla om att avsluta hyresavtalet tidigare.
Läs mer på InfoFinlands sida Hyresavtal.
Jag har ett tills vidare gällande hyresavtal.
Jag sade upp avtalet den 2 juni.
Hyresvärden kräver att jag betalar hyra även för juli.
Måste jag betala?
Om inget annat har avtalats i ditt hyresavtal räknas uppsägningstiden enligt lag från slutet av den månad under vilken du säger upp hyresavtalet.
Om du säger upp bostaden den 2 juni, börjar uppsägningstiden den 30 juni och den varar en månad.
Du måste alltså ännu betala hyra för juli.
Läs mer på InfoFinlands sida Hyresavtal.
Att bli av med sin bostad
Jag har inte råd att betala hyran.
Vad kan jag göra?
Kontakta hyresvärden så snart som möjligt och försök förhandla om en förlängning av betalningstiden.
Ta reda på om du kan skjuta upp andra betalningar för att kunna betala hyran.
Kontakta också din bank och ta reda på om banken kan ge dig ett lån så att du kan betala hyran.
Fråga hos FPA om du har rätt till bostadsbidrag eller något annat understöd.
Du kan även be om hjälp och råd vid kommunens skuldrådgivning eller socialverk eller en boenderådgivare vid kommunen eller hyreshusbolaget eller till exempel Garantistiftelsen.
Läs mer på InfoFinlands sida Ekonomiska problem.
Jag måste flytta ut på grund av skilsmässa.
Jag är dessutom rädd att jag kommer att förlora mitt uppehållstillstånd.
Vad kan jag göra?
På InfoFinlands sida Hyresbostad hittar du information om hur du kan söka en ny bostad.
Skilsmässan kan påverka ditt uppehållstillstånd om du har ett tidsbundet uppehållstillstånd på grund av familjeband.
I vissa situationer kan tillståndet dock förlängas om du fortfarande har nära anknytning till Finland, till exempel i form av en arbetsplats.
Läs mer på InfoFinlands sida Kan jag förlora mitt uppehållstillstånd.
Hyresvärden har hotat med att vräka mig från hyresbostaden på grund av högljutt liv.
Om du upprepade gånger bryter mot husets ordningsregler har hyresvärden rätt att häva hyresavtalet.
Försök att enas om saken med hyresvärden innan avtalet hävs.
Du kan också till exempel kontakta grannmedlingscentret Naapuruussovittelun keskus.
Jag var tvungen att flytta ut och jag har inte hittat en ny bostad.
Vad kan jag göra?
I Finland erbjuder kommunerna tjänster för bostadslösa.
Också många organisationer och församlingar hjälper bostadslösa.
Dessa tjänster är avsedda för människor som har en hemkommun i Finland.
Om du blir bostadslös ska du kontakta socialbyrån eller socialstationen i din hemkommun.
Läs mer på InfoFinlands sida Bostadslöshet.
Konflikter med grannarna
Min granne för oljud.
Vad kan jag göra?
Dina grannar får inte föra oljud till exempel på nätterna.
Om din granne ofta och på ett allvarligt sätt bryter mot ordningsreglerna, kan du kontakta disponenten eller hyresvärden.
Min granne klagar ständigt om oljud hos mig.
Hurdana ljud är tillåtna i ett höghus?
Bostadsaktiebolagets ordningsregler anger när det ska vara tyst i huset.
I ett höghus finns ordningsreglerna oftast i trapphuset.
Under de tysta timmarna får man inte vara högljudd, till exempel spela på instrument eller lyssna på musik på hög volym, men normalt liv är tillåtet.
Varifrån kan jag få hjälp vid konflikter med min granne?
Om du och din granne har en konflikt som ni inte klarar av att själva lösa, kan ni be om hjälp vid grannmedlingscentret Naapuruussovittelun keskus eller hos disponenten.
Grannmedling innebär att grannarna diskuterar och en utomstående medlare leder samtalet.
På mötet kan man komma överens om hur situationen ska lösas.
Medlingen är kostnadsfri.
Läs mer på webbplatsen för grannmedlingscentret Naapuruussovittelun keskus.
linkkiCentrum för grannmedling:
Information om grannmedlingfinska _ engelska
Boendevardag
Vad ska jag göra om jag glömmer nyckeln hemma?
I bostadsaktiebolag har fastighetsskötseln eller disponenten oftast kopior på nycklarna och de kan öppna dörren mot en avgift.
I höghus finns ett nummer nära entrédörren som du kan ringa i en sådan situation.
Hur sopsorterar jag rätt?
I Finland sorteras till exempel bioavfall, kartong, glas, metall, farligt avfall och blandavfall.
Läs mer på InfoFinlands sida Avfallshantering och återvinning.
Vad ska jag beakta när jag använder bastun i min bostad?
Du ska aldrig placera något ovanför bastuugnen, använda bastun som förråd eller torka tvätt i bastun, eftersom detta kan orsaka en brand.
Stäng alltid av en elektrisk bastuugn efter användning.
Läs mer på InfoFinlands sida Säkerheten i hemmet.
Vad gör jag när en vattenkran läcker?
Ring fastighetsskötseln som ditt bostadsaktiebolag har avtal med.
Fastighetsskötseln kan göra små reparationer, till exempel reparera en kran eller öppna upp ett avlopp.
Fuktproblem
Jag har fuktproblem eller andra fel i min bostad Vad gör jag?
Kontakta omedelbart fastighetsskötseln, disponenten eller hyresvärden.
Det är viktigt att felen åtgärdas snabbt, innan de förvärras.
När vi lagar mat uppstår det mycket fukt i köket.
Vad kan vi göra?
Om du inte har en mekanisk ventilation i ditt hem ska du öppna fönstren och vädra via dem.
Detta är särskilt viktigt om du upptäcker att det samlas vattenånga eller fukt på fönstren när du lagar mat.
Använd spisfläkten när du lagar mat.
Kontrollera att frånluftsventilerna är öppna.
Om du orsakar skador i bostaden måste du ersätta dem.
Läs mer på InfoFinlands sida Rättigheter och skyldigheter för boende.
Rådgivningstjänster
Var får jag hjälp och råd i boendefrågor?
Det finns många ställen där du kan be om råd i boendefrågor.
Läs mer på InfoFinlands sida Hyresbostad.
Yrkesutbildning ger den studerande behörighet till ett visst yrke.
Därför är utbildningen mycket praktikorienterad.
Du kan söka till en yrkesutbildning när du har avlagt lärokursen för den grundläggande utbildningen.
Även vuxna kan utbilda sig till ett nytt yrke eller komplettera sin kompetens.
Din grundutbildning avgör till hurudan yrkesutbildning du kan söka och på vilket sätt ansökan sker.
Om du har avlagt grundskolans lärokurs kan du ansöka till grundskolebaserad yrkesutbildning (peruskoulupohjainen ammatillinen koulutus).
Om du har avlagt gymnasiet kan du ansöka till gymnasiebaserad yrkesutbildning (lukiopohjainen ammatillinen koulutus).
Om du vill avlägga examen vid sidan av arbetet kan du ansöka till yrkesutbildning för vuxna (ammatillinen aikuiskoulutus).
Läs mer på InfoFinlands sida Ansökan till utbildning.
När du har avlagt yrkesinriktad grundexamen kan du söka dig till fortsatta studier antingen inom yrkesinriktad tilläggsutbildning, vid en yrkeshögskola eller vid ett universitet.
Grundläggande information om yrkesutbildningfinska _ svenska _ engelska
linkkiUtbildningsstyrelsen:
Ytterligare information om yrkesutbildningfinska _ svenska _ engelska
Gemensam ansökan till gymnasier och yrkesläroanstalterfinska _ svenska
Antagning enligt prövningfinska _ svenska
Utbildningsområden i yrkesutbildningenfinska _ svenska
Förberedande för yrkesutbildning
Utbildning som handleder för grundläggande yrkesutbildning (Ammatilliseen peruskoulutukseen valmentava koulutus) d.v.s. VALMA är avsedd för dem som vill avlägga en grundläggande yrkesutbildning.
Under VALMA-utbildningen får du kunskap och färdigheter som hjälper dig i dina senare yrkesinriktade studier.
Du kan även förbättra din språkkunskap. Du kan också höja dina grundskolebetyg.
VALMA-utbildningen räcker ett läsår.
Läs mera på InfoFinlands sida Utbildning som handleder för yrkesutbildning.
Yrkesinriktad grundexamen
Yrkesutbildning ges av yrkesläroanstalter (ammatillinen oppilaitos), specialyrkesläroanstalter (erityisammattioppilaitos) och av vuxenläroanstalter (aikuisopisto).
Du kan avlägga en yrkesinriktad grundexamen antingen
Inom den grundläggande utbildningen (ungdomar och vuxenstuderande)
Som fristående examen (näyttötutkinto) (vuxenstuderande)
Genom läroavtalsutbildning (oppisopimuskoulutus) (ungdomar och vuxenstuderande)
En yrkesinriktad grundexamen ger dig den grundläggande kompetensen i ett visst yrke.
En grundskolebaserad utbildning varar i cirka tre år.
Du kan också studera vid en yrkesläroanstalt och ett gymnasium samtidigt.
Då kan du avlägga en dubbelexamen (kaksoistutkinto).
Vid yrkesskolorna finns många olika områden som du kan studera.
Det humanistiska och pedagogiska området
Det samhällsvetenskapliga, företagsekonomiska och administrativa området
Det naturvetenskapliga området
Teknik och kommunikation
Naturbruk- och miljöområdet
Social-, hälso- och idrottsområdet
turism- och kosthållsbranschen
Säkerhetsbranschen
Personlig utvecklingsplan för kunnandet
För varje studerande upprättas en personlig utvecklingsplan för kunnandet (PUK).
I planen nedtecknas vilket kunnande du har förvärvat tidigare och fastställs vilka studier du ska avlägga.
Du kan avlägga studierna i egen takt och påvisa vad du kan i praktiska uppgifter på arbetsplatser.
Utbildningsavtal
Utbildningsavtalet är inlärning i arbetet.
Om du vill skaffa dig praktiska kunskaper på en arbetsplats, är ett utbildningsavtal ett bra alternativ för ett läroavtal.
För utbildningstiden betalas ingen lön.
Utbildningsavtalet kan även kombineras med läroavtal.
Yrkesutbildning efter gymnasiet
Om du har avlagt gymnasiet eller studentexamen, kan du söka till en gymnasiebaserad utbildning.
Då kan du inte söka till en grundskolebaserad yrkesutbildning.
Läs mer på InfoFinlands sida Ansökan till utbildning.
Yrkesutbildning för vuxna
Om du arbetar kan du avlägga en yrkesexamen flexibelt vid sidan om arbetet.
Yrkesutbildning för vuxna omfattar
yrkesinriktade grundexamina
yrkesexamina
specialyrkesexamina.
I utbildningen beaktas din tidigare utbildning och den kunskap som du inhämtat som arbetstagare eller företagare.
Du hittar närmare information om hur du kan söka till en yrkesinriktad vuxenutbildning på InfoFinlands sida Ansökan till utbildning.
Examen vid sidan av arbetet med läroavtal
Läroavtal (oppisopimus) innebär inlärning i arbetet.
Du arbetar på en arbetsplats inom din egen bransch och avlägger examen vid sidan av arbetet.
Genom läroavtalsutbildning kan du avlägga samma examen som vid yrkesläroanstalter.
Yrkesexamen (ammattitutkinto)
Specialyrkesexamen (erityisammattitutkinto)
För att kunna studera genom läroavtal måste du ha en arbetsplats.
Du måste hitta en arbetsgivare som vill anställa dig.
Du kan inte inleda din läroavtalsutbildning om du inte har en arbetsplats.
Arbets- och näringsbyrån (TE-toimisto) kan hjälpa dig att hitta ett jobb.
Läroavtalsplatsen kan också vara din nuvarande arbetsplats.
När du har en arbetsplats ska du kontakta läroavtalsbyrån (oppisopimustoimisto) i din region.
Du kan också kontakta en läroanstalt som tillhandahåller läroavtalsutbildning.
Läroavtalsutbildning ges till exempel vid många vuxenutbildningscentra (aikuiskoulutuskeskus).
Under läroavtalsutbildningen betalar arbetsgivaren dig en lön som motsvarar minst en praktikantlön.
Om din arbetsgivare inte betalar dig lön för den tid som du använder för teoretiska studier har du möjligtvis rätt att ansöka om dagpenning, reseersättning och familjebidrag om du omfattas av Den sociala tryggheten i Finland.
Fråga mer vid din läroanstalt.
Information om läroavtalsutbildningfinska _ svenska
Information om läroavtalsutbildningfinska
Kontaktuppgifter till läroavtalsbyråerfinska
linkkiUtbildningsstyrelsen:
Information om läroavtalsutbildningfinska
Bevis för yrkeskunnighet med fristående examen
Fristående examen (näyttötutkinto) är ett sätt att bevisa sin yrkeskunnighet.
Genom fristående examen kan du avlägga
Yrkesexamen (ammattitutkinto)
Yrkesexamen och specialyrkesexamen ger dig behörighet till ett visst yrke.
Dessa examina avläggs alltid genom fristående examen.
Fristående examen är ett lämpligt alternativ också om du har avlagt en yrkesexamen i något annat land och vill jämställa den med en finsk examen.
Om du vill avlägga en fristående examen ska du ta kontakt direkt med läroanstalten.
Fristående examina kan avläggas vid yrkesläroanstalter och vuxenläroanstalter.
För fristående yrkesexamen finns ingen bestämd ansökningstid.
Du avlägga fristående examen vid ett examenstillfälle (tutkintotilanne) där en representant för läroanstalten intygar din yrkeskunnighet.
Sedan får du ett yrkesbevis som bevisar din yrkeskunnighet.
linkkiUtbildningsstyrelsen:
Information om fristående examenfinska _ svenska _ engelska
Yrkesutbildning som anordnas av arbetsgivaren
En del arbetsgivare utbildar människor till arbeten hos dem.
Dessa arbetsgivare ger garanti om en arbetsplats.
Det betyder att den som avlägger utbildningen får en arbetsplats hos arbetsgivaren.
Du får alltså både yrkesutbildning och en arbetsplats.
Till exempel många trafikföretag och VR utbildar de personer som de anställer.
Utbildningen i Finland håller en hög kvalitet.
Skillnaderna i olika skolors studieresultat är små och nästan alla avlägger grundskolan inom den utsatta tiden.
Förskoleundervisning, grundläggande utbildning och utbildning på andra stadiet är kostnadsfria och även därefter är utbildningen till största delen kostnadsfri.
Målet är att alla, oavsett familjens inkomster, ska ha möjlighet att få en högklassig utbildning och växa till aktiva medborgare.
Utbildningssystemet omfattar småbarnspedagogik, förskoleundervisning, grundläggande utbildning, utbildning på andra stadiet och högskoleutbildning.
Vuxenutbildningen är avsedd för vuxna och innehåller många alternativ från grundläggande utbildning till högskoleutbildning.
Småbarnspedagogik
I Finland har barnen rätt till småbarnspedagogik före skolåldern.
Småbarnspedagogiken ordnas i daghem och familjedagvården.
Barnet kan även delta i småbarnspedagogik tillsammans med föräldern i lekparker.
Barnet kan få minst 20 timmar småbarnspedagogik i veckan eller mer om föräldrarna arbetar eller struderar.
Målet är att stödja barnets utveckling och välbefinnande.
Barnet lär sig bland annat sociala färdigheter, att göra saker med händerna och olika kunskaper.
Barnet lär sig också olika färdigheter som hjälper hen att lära sig ytterligare nya saker.
Dagarna innehåller mycket lek och utevistelser.
Om barnet har ett annat modersmål än finska eller svenska, får hen stöd i lärandet av finska eller svenska.
Om barnet behöver, kan hen även få specialundervisning.
I Finland ordnar kommunerna småbarnspedagogiken.
Den finansieras med skattemedel och är därför förmånligare för familjerna.
I Finland finns även privat småbarnspedagogik.
De som arbetar med barnen är utbildade pedagoger inom småbarnsfostran och barnskötare.
Förskoleundervisning
I Finland ska barnen delta i förskoleundervisning under ett års tid innan läroplikten börjar.
Vanligtvis börjar förskoleundervisningen det år då barnet fyller sex år.
Förskoleundervisningen ordnas av kommunerna och är kostnadsfri för familjen.
Förskoleundervisningen ges av pedagoger inom småbarnsfostran som har avlagt universitetsexamen.
Förskoleundervisning ges vanligtvis fyra timmar om dagen från måndag till fredag.
Om föräldrarna arbetar eller studerar kan barnet utöver förskoleundervisningen även delta i småbarnspedagogiken.
Under detta år lär sig barnet kunskaper som hen har nytta av i skolan, till exempel bokstäver.
Barnen undervisas dock inte ännu i läsning.
Om barnet har ett annat modersmål än finska eller svenska, får hen stöd i lärandet av finska eller svenska.
Till dagen hör också lek och utevistelse.
Läs mer på InfoFinlands sida Förskoleundervisning.
Grundläggande utbildning
I Finland börjar den grundläggande utbildningen det år då barnet fyller sju år.
Alla barn som har sitt stadigvarande boende i Finland måste delta i den grundläggande utbildningen.
Grundskolan har nio årskurser.
Läroplikten upphör när barnet har fullgjort hela lärokursen för den grundläggande utbildningen eller det har förflutit tio år sedan läroplikten började.
I Finland reglerar lagstiftningen den grundläggande utbildningen.
Dessutom används nationella läroplansgrunder och lokala läroplaner.
Den grundläggande utbildningen ordnas av kommunerna.
Den finansieras med skattemedel och är därför kostnadsfri för familjerna.
I de lägre årskurserna har man cirka 20 undervisningstimmar i veckan och antalet ökar i de högre årskurserna.
Alla grundskolelärare i Finland har magisterexamen.
Klasslärarna i grundskolan, som undervisar årskurserna 1–6, har läst pedagogik.
Lärarna i årskurserna 7–9 har läst det ämne som de undervisar.
Lärare har stor frihet att planera undervisningen självständigt utifrån den nationella och lokala läroplanen.
På sistone har man i läroplanen betonat bland annat helheter som omfattar flera läroämnen, undersökning av vardagliga fenomen samt data- och kommunikationsteknik.
Barnen har ofta en och samma lärare under de sex första skolåren.
Läraren lär känna eleverna bra och kan utveckla undervisningen så att den passar dem.
Ett viktigt mål är att eleverna lär sig att tänka självständigt och tar eget ansvar för sitt lärande.
Läraren bedömer elevernas framsteg i skolan.
I den grundläggande utbildningen ges alla vitsord av läraren.
Det finns inga egentliga nationella prov.
Däremot följs inlärningsresultaten upp med urvalsbaserade bedömningar.
Dessa ordnas oftast i årskurs nio.
Om barnet eller den unga har flyttat till Finland nyligen, kan hen få förberedande undervisning före den grundläggande utbildningen.
Den förberedande undervisningen varar vanligtvis ett år.
Därefter kan eleven fortfarande läsa finska eller svenska som andraspråk, som S2-språk, om hen behöver stöd med språket.
Vuxna invandrare som inte har grundskolans avgångsbetyg från sitt eget land kan avlägga grundskolan på vuxengymnasiet.
Läs mer om den grundläggande utbildningen på InfoFinlands sida Grundläggande utbildning.
Utbildning på andra stadiet
De vanligaste alternativen efter grundskolan är gymnasium och yrkesutbildning.
Dessa är utbildning på andra stadiet.
Utbildning på andra stadiet är oftast kostnadsfri för studeranden.
Böcker och annat studiematerial måste man dock köpa själv.
Gymnasium
Gymnasiet är en allmänbildande utbildning som inte ger ett yrke.
I gymnasiet läser man samma ämnen som i den grundläggande utbildningen, med undervisningen är mer krävande och studierna mer självständiga.
På slutet avlägger studerandena vanligtvis studentexamen.
Gymnasiet tar 2–4 år, beroende på den studerande.
Efter gymnasiet kan man söka till universitet, yrkeshögskola eller gymnasiebaserad yrkesutbildning.
I de flesta gymnasieskolorna är undervisningsspråket finska eller svenska.
I de stora städerna finns några gymnasieskolor med något annat undervisningsspråk, till exempel engelska eller franska.
Vuxna kan avlägga gymnasiestudier på vuxengymnasiet.
Där kan man avlägga enskilda kurser eller hela gymnasielärokursen och studentexamen.
Undervisningen kan bestå av närundervisning, distansundervisning, webbundervisning och självständiga studier.
Läs mer om gymnasiestudierna på InfoFinlands sida Gymnasium.
Förberedande gymnasieutbildning
På gymnasiet behövs goda språkkunskaper.
Om studeranden har ett annat modersmål än finska eller svenska och saknar tillräckliga språkkunskaper för gymnasiestudierna, kan hen söka till förberedande gymnasieutbildning (LUVA).
Läs mer på InfoFinlands sida Förberedande gymnasieutbildning.
Yrkesutbildning
Yrkesutbildningen är mer praktiknära än gymnasieutbildningen.
En yrkesinriktad grundexamen kan avläggas på ungefär tre år.
Därefter kan man fortsätta studierna och avlägga yrkesexamen eller specialyrkesexamen.
En väsentlig del av studierna är inlärning på arbetsplatsen.
Om man vill, kan man efter yrkesutbildningen fortsätta studierna ända till högskoleutbildning.
Om man redan behärskar de färdigheter som krävs för examen, kan man också avlägga yrkesexamen eller specialyrkesexamen som yrkesprov.
Yrkesexamen kan även avläggas med läroavtal.
Då arbetar studeranden på en arbetsplats inom den egna branschen, får minst samma lön som en praktikant för arbetet och avlägger samtidigt sina studier.
Läs mer på InfoFinlands sida Yrkesutbildning.
Utbildning som handleder för yrkesutbildning
Om du inte har tillräckliga språkkunskaper eller studiefärdigheter för yrkesutbildning, kan du före yrkesutbildningen söka till utbildning som handleder för yrkesutbildning (VALMA).
Läs mer på InfoFinlands sida Utbildning som handleder för yrkesutbildning.
Högskoleutbildning
Efter studierna på andra stadiet kan du gå vidare till högskoleutbildning.
I Finland tillhandahålls högskoleutbildning av yrkeshögskolor och universitet.
Studierna på yrkeshögskola kan vara kostnadsfria eller avgiftsbelagda för studeranden.
Terminsavgift tas ut av personer som inte är medborgare i ett EU-/EES-land eller familjemedlem till en medborgare i ett EU-/EES-land och som avlägger en lägre eller högre högskoleexamen på engelska.
Läs mer på InfoFinlands sida Utländska studerande i Finland.
Yrkeshögskolor
På yrkeshögskolan är undervisningen mer praktiknära än på universitetet.
I undervisningen ingår även inlärning i arbetet.
Yrkeshögskoleexamen kan avläggas på 3,5–4,5 år.
Om man vill fortsätta studierna därefter och avlägga högre yrkeshögskoleexamen, måste man först skaffa sig tre år av arbetserfarenhet från samma område som examen.
Läs mer på InfoFinlands sida Yrkeshögskolor
Undervisningen på universitet är baserad på vetenskaplig forskning.
På universitet kan man avlägga lägre högskoleexamen på cirka tre år och därefter högre högskoleexamen på cirka två år.
Universiteten ordnar undervisning på engelska i vissa utbildningsprogram.
I de flesta utbildningsprogrammen är undervisningsspråket ändå finska eller svenska.
När man har avlagt magisterexamen, kan man ansöka om rätt till fortsatta studier och avlägga licentiat- eller doktorsexamen.
Läs mer på InfoFinlands sida Universitet.
Ansökan till utbildning
På InfoFinlands sida Ansökan till utbildning finns information om hur du ansöker till utbildning på andra stadiet och högskoleutbildning i Finland.
Om du planerar att studera i Finland, läs mer på InfoFinlands sida Utländska studerande i Finland och Studerande.
Andra studiemöjligheter
I Finland finns även många läroanstalter som erbjuder studier som inte leder till examen för människor i alla åldrar.
Största delen av dessa utbildningar är avsedda för vuxna.
Sådana läroanstalter är medborgarinstitut, folkhögskolor, sommaruniversitet, studiecenter och idrottsutbildningscenter.
Studierna är allmänbildande.
Du kan studera till exempel bland annat språk, estetiska ämnen, handarbete och kommunikation.
Oftast betalar den studerande en avgift för studierna.
I vissa situationer kan studierna vid dessa läroanstalter dock vara kostnadsfria.
Om till exempel utbildning i läs- och skrivkunnighet eller någon annan språkutbildning har godkänts till din integrationsplan, tas det inte ut någon avgift för studierna.
Språkutbildning
Om du vill läsa finska eller svenska, läs mer på InfoFinlands sida Finska och svenska språket.
På den här sidan har vi sammanställt de viktigaste rättigheter och skyldigheter för boende i Finland.
Du är skyldig
Att följa ordningsreglerna i ditt bostadsaktiebolag om du bor i ett höghus eller ett radhus.
I ordningsreglerna anges vanligtvis till exempel tiderna för när det ska vara tyst i huset.
Ofta innehåller de även anvisningar om användningen av gemensamma utrymmen i huset.
I ett höghus hittar du ordningsreglerna vanligtvis i trapphuset nära entrédörren.
Att se till att även dina gäster följer ordningsreglerna.
Att enbart använda bostaden för det avsedda ändamålet.
Om bostaden är avsedd att användas för boende, kan du inte bo på ett annat ställe och använda bostaden som lokal.
Du har rätt
Att leva ett normalt liv i ditt hem.
Bostadsaktiebolaget kan inte utfärda sådana ordningsregler som står i strid med lagen eller begränsar ett normalt liv i alltför stor omfattning.
Till hemfrid.
Dina grannar får inte störa din hemfrid till exempel genom att föra oljud mitt i natten.
Om en granne ofta bryter mot ordningsreglerna på ett allvarligt sätt, ska du först ta upp saken med grannen.
Om detta inte hjälper, kan du kontakta disponenten eller hyresvärden.
Hemfrid innebär också att du i regel själv får bestämma vem som har tillträde till ditt hem.
Hyresgästens rättigheter och skyldigheter
Du är skyldig
Att betala hyran i tid.
Hyresbeloppet anges i hyresavtalet.
Hyresvärden kan höja hyran i enlighet med vad som anges i hyresavtalet.
Att se till att hyresbostaden hålls i ett gott skick.
Att följa villkoren i hyresavtalet.
Om det till exempel anges i hyresavtalet att det är förbjudet att röka i bostaden, kan du inte röka i ditt hem.
Om hyresavtalet kräver att du har en hemförsäkring, måste du teckna en sådan.
Det är bra att teckna en hemförsäkring även om detta inte krävs i hyresavtalet.
Att fråga om tillstånd hos hyresvärden om du vill göra ändringar i bostaden, till exempel måla en vägg.
Utan tillstånd får du inte göra några ändringar, även om du skulle bekosta renoveringen själv.
Begär tillståndet skriftligt.
Att ersätta hyresvärden för skador som du åsamkar bostaden.
Att meddela hyresvärden om du upptäcker sådana fel i bostaden som hyresvärden ansvarar för.
Hyresvärden ansvarar till exempel för bostadens fasta inredning och ytmaterial.
Att meddela eventuella fel till fastighetsskötseln, till exempel en läckande kran.
Du har rätt
Att bo i hyreslägenheten enligt vad som anges i hyresavtalet.
Hyresvärden får endast beträda bostaden i vissa undantagsfall, till exempel för att övervaka reparationer i bostaden eller visa bostaden för köpare.
Även då måste hen försöka i förväg komma överens om detta med dig.
Att få ett skriftligt meddelande i förväg om hyran höjs.
I meddelandet ska det stå hur mycket och när hyran kommer att höjas och vad som är grunden till höjningen.
Till en uppsägningstid enligt lag.
Att häva hyresavtalet omedelbart om det är skadligt för hälsan att bo i bostaden.
Att hyra ut en del av bostaden till en annan person, om detta inte medför olägenhet för hyresvärden.
Att få ett förhandsmeddelande om reparationer.
Små reparationer ska meddelas 14 dagar i förväg och stora reparationer sex månader i förväg.
Brådskande reparationer kan dock göras utan ett meddelande.
Om det är svårt eller omöjligt att bo i bostaden under reparationerna, har du rätt att säga upp hyresavtalet eller får nedsatt hyra.
Detta måste du emellertid alltid komma överens om med hyresvärden.
Läs mer på InfoFinlands sida Hyresavtal.
Rättigheter och skyldigheter i en ägarbostad
I ett bostadsaktiebolag har du skyldighet att
Betala bolagsvederlag och eventuellt även finansieringsvederlag för bostadsaktiebolagets lån till bostadsaktiebolaget.
Vederlagen används till att sköta bostadsaktiebolaget, till exempel underhålla byggnaderna och gårdsområdet.
Se till att din bostad hålls i gott skick.
I förväg meddela till bostadsaktiebolagets disponent eller styrelse om du ska göra en sådan ändring i din bostad som kan påverka husets bärande konstruktioner, vattenledningar, fuktisolering, elledningar eller ventilationssystem.
Till exempel ska en badrumsrenovering alltid meddelas i förväg.
Genomföra renoveringar på ett sådant sätt att bygganden inte tar skada.
I Finland finns exakta bestämmelser till exempel om hurdant tätskikt ett badrum ska ha.
Meddela bostadsaktiebolaget eller disponenten, i praktiken vanligtvis allra först fastighetsskötseln, om det finns ett sådant fel i din bostad vars åtgärdande åligger bostadsaktiebolaget.
I ett bostadsaktiebolag har du följande rättigheter:
Förvalta den bostad vars aktier du äger.
Du får göra ändringar i din bostad.
Tänk på att renoveringen inte får medföra olägenhet till bostadsaktiebolaget eller de andra aktieägarna.
Hyra ut din bostad eller en del av den till en annan person.
Delta i stämmor och på dem påverka det som händer i bostadsaktiebolaget.
På en stämma kan du rösta om olika saker och kräva att ett ärende tas upp för behandling på stämman.
Bostadsaktiebolaget ska se till att husets konstruktioner, isolering, värmesystem, elledningar, vattenledningar och avlopp samt gårdsområden hålls i gott skick.
På stämman fattas beslut om reparationer gällande dessa.
I vissa bostadsaktiebolag har man beslutat att fördela ansvaret på ett annat sätt.
I detta fall står det i bolagsordningen vem som ansvarar för vad.
Alla barn som har sitt stadigvarande boende i Finland har läroplikt, vilket innebär att de måste delta i den grundläggande utbildningen.
Läroplikten är lagstadgad.
Läroplikten
börjar det år då barnet fyller 7 år
upphör när grundskolans lärokurs har fullgjorts eller det har förflutit 10 år sedan läroplikten började.
Läroplikten fullgörs vanligtvis i grundskolan.
Grundskolan består av lågstadiet (alakoulu) och högstadiet (yläkoulu).
Lågstadiet omfattar årskurserna 1–6, högstadiet årskurserna 7–9.
Grundskolan är vanligen nioårig: skolan börjar i årskurs 1 och slutar i årskurs 9.
Grundskolan är gratis.
Grundläggande utbildning för invandrarefinska _ svenska
Att börja i skolan
Föräldrarna anmäler sitt barn till skolan.
I början av året skickar staden en anmälan om läroplikt (oppivelvollisuusilmoitus) till hemmen.
I anmälan anges barnets närskola (lähikoulu).
Närskolan är oftast den skola som ligger närmast barnets hem.
Föräldrarna kan också välja en annan skola än närskolan.
Det är ändå inte alltid möjligt att få en plats på en annan skola.
Du kan anmäla ditt barn till skolan i närskolan.
I vissa kommuner kan anmälan göras även på internet.
Anmälningstiden är i början av året, vanligen i januari.
Olika skolor
Barn kan också gå i en skola med en speciell inriktning.
Ibland är dessa skolor privatskolor.
Skolor kan ha till exempel följande inriktningar:
bildkonst
motion
språk
internationalitet (till exempel Europaskolan)
specialpedagogik (till exempel Steinerpedagogik)
I Finland finns några internationella skolor.
I vissa skolor ges undervisningen på något annat språk än finska.
Till exempel i Tyska skolan sker undervisningen på tyska.
Skolor som har andra undervisningsspråk än finska finns i de största städerna.
Även i vanliga grundskolor kan det finnas några klasser där undervisningen sker på ett främmande språk.
linkkiEuropaskolan i Helsingfors:
Europaskolan i Helsingforsfinska _ engelska _ franska
linkkiFörbundet för Steinerpedagogik:
Information om Steinerskolanfinska _ engelska
Skoldagen och studierna
Skolan börjar i augusti och slutar i slutet av maj eller i början av juni.
I juni och juli är det sommarlov.
Längden på skoldagarna varierar i olika årskurser.
På lågstadiet är dagarna kortare än på högstadiet.
Lektionerna är vanligen 45 minuter långa.
Skolveckan består av ungefär 20 lektioner.
Barnen äter en varm måltid i skolan.
Den är gratis.
Om ditt barn har en specialdiet ska du tala om det för läraren.
I grundskolan studerar barnen många obligatoriska ämnen.
I lågstadiets högre klasser och på högstadiet får de även välja tillvalsämnen.
Alla kan få undervisning i den egna religionen eller i livsåskådningskunskap i skolan.
Religionsundervisning måste ordnas när det finns minst tre barn som bekänner en viss religion i kommunen.
I vissa skolor finns det skilda klasser för elever som är duktiga på till exempel musik eller bildkonst.
Oftast söker man separat till dessa klasser.
Invandrare och grundskolan
Barnet eller den unga kan få förberedande undervisning före den grundläggande utbildningen under vilken han eller hon studerar finska (eller svenska) och vissa läroämnen.
Den förberedande undervisningen före grundskolan är avsedd för alla de barn med invandrarbakgrund som inte har tillräckliga kunskaper för att klara sig i undervisningen inom den grundläggande utbildningen.
Den förberedande undervisningen pågår vanligtvis i ett år.
Därefter övergår eleven till en vanlig klass.
Om barnet har ett annat modersmål än finska eller svenska kan kommunen ordna undervisning i barnets eget modersmål.
Då kan barnet även lära sig finska eller svenska som andra språk, som S2-språk (S2-kieli).
Eleven studerar finska (eller svenska) som andra språk om hans eller hennes kunskaper i språket inte är på samma nivå som infödda talares.
Vuxengymnasier ordnar grundläggande utbildning för vuxna invandrare som inte har grundskolans avgångsbetyg från sitt eget land.
Mer information om detta får du vid rådgivningen i din hemkommun eller vid närmaste vuxengymnasium.
Du kan söka kontaktuppgifter tillvuxengymnasier med hjälp av sökmotorer på Internet.
linkkiUndervisnings- och kulturministeriet:
Information om grundundervisningenfinska _ svenska _ engelska
linkkiUtbildningsstyrelsen:
Information om grundundervisningenfinska _ svenska _ engelska
Meddelanden mellan hem och skola
I många kommuner informerar skolan viktiga ärenden i den webbaserade tjänsten Wilma.
Skolan ger barnets föräldrar inloggningsuppgifter till tjänsten.
Via Wilma kan du ha kontakt med barnets lärare och få information om barnets lärande, prov och frånvaron samt händelser i skolan och om skollov.
Om barnet är frånvarande från skolan till exempel på grund av sjukdom ska du meddela skolan om detta på morgonen via Wilma.
Det är viktigt att man regelbundet följer Wilma.
Om du behöver hjälp med att använda Wilma ska du be skolan om en introduktion.
Kervo stad har publicerat anvisningar om användningen av Wilma på olika språk.
Observera att inloggning till Wilma sker på olika adresser i olika städer.
linkkiKervo stad:
Så här använder du Wilma(pdf, 239 kt)finska _ engelska _ ryska _ estniska _ turkiska _ kurdiska _ thai _ vietnamesiska
linkkiVisma:
Stöd för studierna och tionde klassen
Grundskoleelever får stöd i sitt skolarbete.
Studiehandledarna berättar om olika studiemetoder och om fortsatta studier.
De ger också yrkesvägledning.
Studiepsykologer och skolkuratorer hjälper eleverna i problemsituationer.
Läraren kan ge barnet kortvarig stödundervisning.
Barnet får specialundervisning om det har inlärnings- eller koncentrationssvårigheter.
Grupperna i specialundervisningen är mindre än vanliga klasser.
Lärarna håller kontakt med föräldrarna.
De ordnar föräldramöten och berättar för föräldrarna om barnets studier.
Många skolor håller kontakt med föräldrarna med hjälp av webbtjänster.
I skolan ges eventuellt också tilläggsundervisning, på så kallade tionde klasser (kymppiluokka).
Där kan eleverna höja sina vitsord och fundera på vilket studieområde de är intresserade av.
Du kan ansöka till en tionde klass när du har fått ditt avgångsbetyg från grundskolan.
Information om tiondeklassenfinska _ svenska
Vanligtvis ska du sortera avfallet hemma innan du gör dig av med det.
Då avfallet sorteras rätt kan man använda materialet för att tillverka nya produkter.
Anvisningarna för sorteringen skiljer sig något från varandra i olika delar av landet.
Anvisningarna finns vanligtvis vid sopbehållarna vid ditt eget hus. Om inte kan du kontakta kommunen eller din hyresvärd.
Kasta inte avfallet ut genom fönstret, i skogen eller på gatan.
Hela saker är inte avfall.
Du kan sälja dem på lopptorg eller på internet eller donera dem till välgörenhet eller återvinningscentraler.
I Finland är det vanligt att köpa använda saker och lätt att hitta använda saker i gott skick.
Hur sorteras avfall?
Sortera avfallet enligt material.
Lägg inte skräp, mat eller kemikaler i avloppet (WC:n).
För alltid farligt avfall till insamlingsställe.
Vid alla hus finns inte alltid samtliga insamlingskärl.
Information om allmänna insamlingsställen finns på adressen kierratys.info.
Du får inte föra ditt eget avfall till insamlingskärl avsedda för ett annat hus.
Du får inte heller lägga avfall från exempelvis ditt företag i sopkärlen avsedda för ditt eget hus.
Insamlingskärl som ofta finns vid husbolaget
Bioavfall (biojäte)
JA: matavfall, även härsken mat, kaffesump, hushållspapper, skal från frukter etc.
Bioavfall komposteras till mylla.
I vissa kommunerer separeras inledningsvis biogas från avfallet för att producera el och värme.
Papper (paperi)
JA: tidningar, reklam, kuvert etc.
NEJ: vått eller mycket smutsigt papper
Av pappret görs dagstidningar eller wc-papper.
Kartong (kartonki)
JA: mjölkförpackningar, papp, papperspåsar, kartongförpackningar
NEJ: våt eller mycket smutsig kartong
Av kartong görs exempelvis papprullar för hushållspapper.
Aluminium i förpackningarna återvinns även.
Glas (lasi)
JA: glasförpackningar (flaskor och matburkar)
NEJ: glasföremål, glaskärl, speglar, porslin
Av glaset tillverkas nya glasförpackningar.
Metall (metalli)
JA: metallföremål och förpackningar som till största delen utgörs av metall
Olika metaller sorteras maskinellt och används för att tillverka nya produkter.
Plast (muovi)
JA: tomma matförpackningar av plast, tomma tvättmedelsflaskor och schampoflaskor, plastpåsar, tomma plastburkar
NEJ: PVC-förpackningar med märkningen 03, förpackningar som innehåller rester av farliga ämnen såsom målarfärg eller kemikalier, plastföremål, leksaker, tandborstar, vattenkannor och så vidare
Av plastförpackningarna tillverkas nya plastprodukter.
Blandavfall (sekajäte) eller övrigt avfall
JA: Allt avfall som du inte kan eller önskar sortera.
NEJ: farligt avfall
Blandavfall bränns vanligtvis vid avfallsverk för att producera el och värme.
Övriga insamlingsställen
Farligt avfall (vaarallinen jäte)
JA: lysrör, energibesparingslampor, kemikalier med ett varningsmärke på förpackningen
VAR: Insamlingsställen för farligt avfall, se kierratys.info
JA: hemmets stora och små batterier, mobiltelefonens batteri
VAR: röda batteriinsamlingslådor i butiker och kiosker
Metallen i batterierna årervinns och de farliga ämnena hanteras på ett säkert sätt.
JA: alla leksaker och utrustning som fungerar med el eller batteri
VAR: små elapparater i butiker som säljer elektronik och större apparater vid insamlingsställen för elskrot, se kierratys.info.
Metall från elapparater (t.ex. guld) återvinns.
Hur kan man minska mängden avfall?
Frys ned mat som blir över.
Förvara maten rätt.
Drick kranvatten, det är gott och säkert i Finland.
Köp endast sådana saker du behöver.
Köp hållbara produkter.
Om du senare vill sälja dem kan du få betalt för dem.
Köp och sälj använda produkter.
Ta hand om dina saker och förvara dem enligt anvisningarna.
Avfallsinsamlingsstationerfinska
linkki4V:
Tips för boende(pdf, 1,5 Mt)finska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
FPA:s bostadsbidrag är avsett för boendekostnader.
FPA:s bostadsbidrag täcker bara en del av boendekostnaderna.
Du kan få bostadsbidrag om du har låga inkomster och bor stadigvarande i Finland.
Med stadigvarande boende i Finland avses att du har ditt egentliga hem i Finland och huvudsakligen också vistas i landet.
För att få bostadsbidrag måste du också du omfattas av den sociala tryggheten i Finland.
Fpa:s stöd för boendet är följande:
allmänt bostadsbidrag
bostadsbidrag för pensionstagare
bostadsunderstöd i samband med militärunderstöd för värnpliktiga och civiltjänstgörare.
Om pengarna inte räcker till för boendekostnaderna fastän du får bostadsbidrag, kan du ansöka om utkomststöd hos FPA.
Läs mer på InfoFinlands sida Ekonomiska problem.
Stöd för boendetfinska _ svenska _ engelska
Fpa:s allmänna bostadsbidrag
Stöd kan betalas till en person eller till ett hushåll (ruokakunta).
Till samma hushåll hör vanligtvis alla som stadigvarande bor i samma bostad.
Vanligen består ett hushåll av ett äkta par, sambor eller en familj.
Också en person kan vara ett hushåll.
Bostadsbidraget beviljas gemensamt för hushållet på basis av en ansökan.
Beakta att om du delar bostad med till exempel en vän och ni har ett gemensamt hyresavtal så anses ni höra till samma hushåll.
Om en av er däremot är huvudhyresgäst och den andra underhyresgäst och ni inte är nära släktingar, anses ni höra till olika hushåll.
Följande kan få allmänt bostadsbidrag
barnfamiljer
studerande
äkta par och registrerade par sambor
ensamboende eller
de som bor i kollektiv.
Hurudana boendekostnader anses skäliga?
Stöd kan beviljas för fast bostad i Finland.
Det är i lagen fastställt vilka boendekostnader om kan anses vara skäliga då stödet beräknas.
Bostaden kan vara:
en hyresbostad
en ägarbostad
en bostadsrättsbostad
en delägarbostad.
Stöd betalas för hyra,vederlag och utgifter för skötseln av bostaden.
Utgifter för skötseln av bostaden är till exempel uppvärmningskostnader och vattenavgifter.
Också en del av räntan på bostadslånet iakttas.
Bostadsbidrag beviljas för skäliga boendekostnader.
I stora städer accepteras högre boendekostnader än på små orter.
Fpa betalar inte alla boendekostnader
En del av boendekostnaderna måste du betala själv.
För detta fastställs en bassjälvrisk.
Bassjälvriskandelens storlek beror på:
hur många vuxna och barn som hör till hushållet
hushållets bruttoinkomster (inkomster före skatt)
Om inkomsterna är mycket låga bortfaller bassjälvrisken.
Då bostadsbidraget kalkyleras avsätts 300 euro per månad av dina förvärvsinkomster.
Detta belopp påverkar inte ditt bostadsbidrag.
Detta kallas förvärvsinkomstavdrag (ansiotulovähennys).
Förvärvsinkomstavdrag görs separat för varje medlem i hushållet.
Bostadsbidrag beviljas endast för skäliga boendekostnader.
Vid fastställande av skäliga boendekostnader beaktas
kommunen där bostaden är belägen
antalet vuxna och barn i hushållets storlek
Om bostaden är större eller dyrare än vad lagen om allmänt bostadsbidrag tillåter växer den andel av boendekostnaderna som du betalar själv.
Det slutliga bostadsbidraget beräknas på följande sätt:
Bassjälvriskandelen dras först bort från boendekostnaderna.
Bostadsbidraget är 80 % av det kvarstående beloppet.
Anmäl ändringar till Fpa
Om dina inkomster, boende- eller familjeförhållanden eller andra omständigheter ändras ska du omgående anmäla ändringen till Fpa.
I Fpa:s beslut anges i detalj vilka omständigheter som bör anmälas.
Allmänt bostadsbidragfinska _ svenska _ engelska
Vad är ett hushållfinska _ svenska _ engelska
Att ansöka om bostadsbidrag
Du ansöker om allmänt bostadsbidrag hos FPA med en ansökan om allmänt bostadsbidrag (AT1).
Du kan också ansöka om bostadsbidraget på internet.
Till din ansökan ska du bifoga:
en kopia av hyresavtalet och en utredning över hyresbeloppet (hyresbostad)
ett intyg på vederlagets belopp och bostadslånet (ägarbostad)
löneverifikat, d.v.s. ett lönebesked som arbetsgivaren gett.
Om du bor i ett kollektiv ska du bifoga ett befullmäktigande av dem som du delar bostad med, d.v.s. en fullmakt att ansöka om bostadsbidrag för alla.
Skicka din ansökan till Fpa:s byrå eller skicka in den på internet.
Fpa betjänar sina kunder på sina byråer, per telefon och post samt via webbtjänsten som finns på FPA:s internetsidor.
När du sköter dina personliga ärenden på en Fpa-byrå ska du ha med dig något identitetsbevis, till exempel pass.
Att ansöka om bostadsbidragfinska _ svenska _ engelska
Enligt lag ska barn i Finland delta i förskoleundervisning eller motsvarande verksamhet under ett års tid innan läroplikten börjar.
Förskoleundervisningen (esiopetus) förbereder barnen inför grundskolan.
Barnen börjar i förskoleundervisningen vanligen vid sex års ålder och grundskolan vid sju års ålder.
Föräldrarna anmäler sitt barn till förskoleundervisningen vanligtvis i januari eller februari.
Kontrollera tidpunkten i god tid vid skolväsendet (koulutoimi) eller bildningsväsendet (sivistystoimi) i din hemkommun.
Kommunerna ordnar förskoleundervisning.
De kan även köpa förskoleundervisningen till exempel av ett privat daghem.
Förskoleundervisningen är kostnadsfri.
Under dagen får barnet en gratis måltid.
Om barnet bor långt (över 5 km) från undervisningsstället, eller om vägen dit är besvärlig, får barnet gratis skjuts.
Om föräldrarna arbetar eller studerar kan barnet utöver förskoleundervisningen även delta i småbarnspedagogiken.
En dag i förskolan
Förskoledagen är ungefär fyra timmar lång.
Förskolan finns ofta antingen i daghemmets eller skolans lokaler.
I förskolan lär sig barnen bland annat matematik, miljö- och naturkunskap samt konst och kultur.
De lär sig nya saker med lekens hjälp.
Föräldrarna har en viktig roll i förskolan.
De stödjer sitt barns inlärning.
Lärarna utarbetar en egen inlärningsplan för varje barn.
Föräldrarna kan hjälpa ledarna att utarbeta planen.
Språk och kulturer i förskoleundervisningen
Ett barn som har ett annat modersmål än finska eller svenska lär sig finska eller svenska som främmande språk.
Dessutom kan det studera sitt eget modersmål om kommunen ordnar undervisning i det språket.
Barnet kan även få undervisning i den egna religionen eller i livsåskådningskunskap i förskolan.
I förskolan lär sig barnen att uppskatta sitt språk och sin kultur.
De lär sig också att respektera andra människors språk och kulturer.
linkkiUtbildningsstyrelsen:
Information om förskoleundervisningenfinska _ svenska _ engelska
Förskoleuppgifter på nätetfinska
linkkiUndervisnings- och kulturministeriet:
Information om förskoleundervisningenfinska _ svenska _ engelska
Brandsäkerhet
En brandvarnare kan rädda ditt liv.
Om en brand uppstår i din bostad avger brandvarnaren ett högljutt larm och du hinner ut i tid.
Se till att det finns tillräckligt många brandvarnare i ditt hem.
Brandvarnare säljs i varuhus och järnaffärer.
En brandvarnare räcker till 60 kvadratmeter.
Om ditt hem är till exempel 65 kvadratmeter stort behöver du två brandvarnare.
Om ditt hem har fler än en våning måste du räkna ytan separat för varje våning.
Det bör finnas en brandvarnare på varje våning.
Kontrollera regelbundet att brandvarnaren fungerar.
Byt batterier vid behov, gärna en gång per år.
Du ansvarar för brandvarnaren även om du bor i en hyresbostad.
Det finns ofta en bastu i finländska hem.
Även om du inte använder bastun får du aldrig placera något på bastuugnen, eftersom detta kan orsaka en brand.
Torka till exempel inte tvätten ovanför eller i närheten av bastuugnen.
Stäng alltid av en elektrisk bastuugn efter användning.
När du går hemifrån, kom ihåg att kontrollera att spisen och ugnen och till exempel strykjärnet är avstängda.
Det är bra att ha en brandsläckare hemma.
I vissa höghus finns det också en brandsläckare i trappuppgången.
Ta reda på var den närmaste brandsläckaren finns.
Se till att du har en släckningsfilt hemma.
Det är bra att förvara filten till exempel i närheten av spisen.
Lämna inte mat på en het spis utan uppsikt.
Var särskilt försiktig om du lagar mat på natten.
Laga inte mat om du är berusad.
Förvara inte föremål på spisen.
Barn, husdjur eller du själv kan av misstag vrida på spisen.
Då kan sakerna som ligger på spisen fatta eld.
Om fett börjar brinna när du lagar mat, kväv elden med till exempel ett kastrullock eller med en släckningsfilt.
Använd inte vatten.
Kom ihåg att stänga av elapparater efter användning.
Strykjärnet ska också kopplas loss från vägguttaget.
Använd inte elapparater som är i dåligt skick eller vars sladd är trasig.
Om en elapparat börjar brinna, använd inte vatten.
Kväv elden med till exempel en brandsläckare.
Om du har elektriska värmeelement eller värmeaggregat hemma, lägg inte tyger, kläder eller något annat på dem.
Lämna utrymme runt TV:n, mikrovågsugnen, kylskåpet och frysen.
Täck inte över dem.
Det är bra att en gång per år städa bort damm från frysens och kylskåpets bakgaller till exempel med dammsugaren, om möjligt.
Rök inte inomhus.
Lämna inte brinnande ljus utan uppsikt.
Tänd inte ljus i närheten av till exempel gardinerna, ens om du själv är i rummet.
Om en brand uppstår, ring nödnumret 112.
linkkiHelsingfors stads räddningsverk:
Brandsäkerhet i höghusfinska _ svenska _ engelska
linkkiRäddningsbranschens Centralorganisation i Finland:
Information om brandsäkerhetfinska _ svenska _ engelska
linkkiHelsingfors stad, Förortsprojektet:
Mitt hem i ett höghus(pdf, 6,56 MB)finska _ engelska _ ryska _ somaliska _ arabiska
linkkiHelsingfors stads räddningsverk:
Brandsäkerhet i småhusfinska _ svenska _ engelska
Så här undviker du vattenskador
Lämna inte tvättmaskinen eller diskmaskinen på när du går hemifrån.
Kontrollera regelbundet att vattenledningarna i ditt hem inte läcker och att det inte rinner ut vatten från hushållsapparaterna på golvet.
Stäng alltid kranen till tvätt- och diskmaskinen när du inte använder dem.
Det ska finnas ett läckageskydd av plast under kylskåpet, frysen och diskmaskinen.
Skyddet läggs på plats samtidigt som apparaten installeras.
Du får inte installera en diskmaskin själv, utan arbetet måste utföras av en fackman.
Om ett vattenläckage uppstår i ditt hem, försök stänga vattenledningens avstängningsventil.
Om du bor i höghus eller radhus, anmäl läckaget genast till journumret för husets servicebolag.
Om du bor i villa, kontakta en jourhavande rörfirma.
Elarbeten
I Finland är nätspänningen 230 volt.
I Finland utförs egentliga elarbeten endast av personer som är yrkesutbildade inom elbranschen.
Vissa små elarbeten får du utföra själv, om du kan.
Du kan till exempel själv:
byta en säkring
byta lampor
reparera en enfas skarvsladd (spänning 230 V)
hänga upp en lampa i taket med en upphängningsbygel
byta en hel enfas anslutningsledning (spänning 230 V) och stickkontakt i en elapparat, om den gamla gått sönder.
linkkiTukes:
Elarbeten som du får göra självfinska _ svenska _ engelska
Säkerhetslås skyddar mot inbrottstjuvar
Om du har ett säkerhetslås i ditt hem, lås det alltid då du inte är hemma.
Lås inte säkerhetslåset när du är hemma.
Om någon bryter in sig i ditt hem, ring nödnumret 112.
linkkiTukes:
Guiden Ett säkert hem för barnfinska _ svenska _ engelska
Birkalands räddningsverk:
Vad gör jag om det börjar brinna hemma?
Om videon väcker frågor hos dig kan du fråga mer av en expert.
Småbarnspedagogik är avsedd för barn under skolåldern.
I Finland tillhandahåller kommunerna kommunal småbarnspedagogik bland annat i daghem.
Dessutom finns det privata daghem.
Småbarnspedagogik är fostran, undervisning och omsorg som är pedagogiskt planerad och som har noga genomtänkta mål.
Inom småbarnspedagogiken arbetar utbildade lärare i småbarnspedagogik och barnskötare.
Vanligen vårdar någondera av föräldrarna barnet hemma åtminstone under föräldraledigheten (vanhempainvapaa), det vill säga tills barnet är ungefär 9 månader gammalt.
Om du vårdar ditt barn hemma även efter detta har du rätt att vara ledig från ditt arbete för vård av barn tills barnet fyller tre år.
Mer information om ledigheterna får du på InfoFinlands sida Familjeledighet.
Du kan ansöka från Kela om ekonomiskt stöd för hemvård av barn.
Läs mer på InfoFinlands sida Stöd för vård av barn i hemmet.
Kommunal småbarnspedagogik
Om du har din hemkommun i Finland, kan du ansöka om en plats inom den kommunala småbarnspedagogiken för barnet efter föräldraledigheten.
Då är barnet ca nio månader gammalt.
Om du inte har en hemkommun i Finland, räknas du som invånare i den kommun där du vistas.
Om båda föräldrarna arbetar, har barnet rätt till småbarnspedagogik på heltid.
Om den ena föräldern är hemma, beror rätten till småbarnspedagogik på hemkommunen.
I vissa kommuner har barnet rätt till småbarnspedagogik på heltid även då den ena föräldern är hemma.
I vissa kommuner har barnet rätt till 20 timmar småbarnspedagogik per vecka om den ena föräldern är hemma.
Familjen kan ändå söka rätt till småbarnspedagogik på heltid om barnet behöver särskilt stöd till exempel i att lära sig det finska språket eller på grund av att familjen befinner sig i en svår situation.
Du kan ansöka om en plats
på ett daghem (päiväkoti)
På daghemmet är barnen i större gruppen är i gruppfamiljedagvården.
Familjedagvård innebär att skötaren vårdar barnen i sitt eget hem.
Vissa familjedagvårdare vårdar barnen hemma hos de barn som ingår i gruppen.
Ansök om en plats inom den kommunala småbarnspedagogiken från din egen kommun senast fyra månader innan du behöver den.
Man kan få en plats inom två veckor, om föräldrarna får ett arbete eller en studieplats.
Avgiften för småbarnspedagogik (varhaiskasvatusmaksu) beror på
familjens inkomster
familjens storlek och
på hur många timmar per vecka barnet deltar i småbarnspedagogik.
Man får syskonrabatt.
Om familjen inkomster är mycket låga, kan småbarnspedagogiken vara kostnadsfri för familjen.
Fråga mer i din kommuns rådgivningstjänster.
Privat småbarnspedagogik
En plats inom den privata småbarnspedagogiken kan finnas
i ett privat daghem eller i ett gruppfamiljedaghem
i familjedagvård eller
hemma, då familjen anställer en skötare i hemmet
Du kan ansöka om en plats inom småbarnspedagogiken direkt från det privata daghemmet eller gruppfamiljedaghemmet.
Du kan också leta upp en privat familjedagvårdare som vårdar barnen hemma hos sig, eller anställa en skötare i ditt eget hem.
Om du anställer en skötare i ditt hem blir du en arbetsgivare, och du måste uppfylla en arbetsgivares skyldigheter.
Läs mera på InfoFinlands sida Arbetsgivarens rättigheter och skyldigheter.
Familjen kan anställa en skötare i sitt hem även tillsammans med en annan familj.
Kommunen övervakar den privata småbarnspedagogiken.
Priserna för den privata småbarnspedagogiken varierar.
Du kan ändå få stöd för den från FPA.
Då är den inte nödvändigtvis mycket dyrare än den kommunala småbarnspedagogiken.
Stöd för privat dagvård
Om barnet har en hemkommun i Finland, kan du ansöka om Fpa-stöd för privat vård.
Dagvårdsproducenten måste ha kommunens godkännande.
Du kan ansöka om privatvårdsstöd (yksityisen hoidon tuki), om
ditt barn som är under skolåldern är i privat dagvård; eller
barnet har någon annan privat skötare.
Du kan inte ansöka om privatvårdsstöd om skötaren är en medlem i barnets familj eller om barnet och skötaren bor i samma hushåll.
Du kan inte heller ansöka om privatvårdsstöd för den kommunala småbarnspedagogiken.
Stödets storlek beror bland annat på familjens inkomster och kommunen som familjen bor i.
Kela betalar stödet direkt till skötaren eller dagvårdsproducenten.
Man måste betala skatt för privatvårdsstödet.
Stödet betalas inte till utlandet.
Läs mera om privatvårdsstöd på Fpa:s sidor.
Fpa har en telefontjänst för barnfamiljer.
på finska tfn +358 (0)20 692 206
på svenska och engelska tfn +358 (0)20 692 226
På Fpas byråer får du betjäning även på andra språk med hjälp av en tolk.
Stöd för privat vårdfinska _ svenska _ engelska
Vad händer i småbarnspedagogiken?
Till småbarnspedagogiken hör mångsidig verksamhet, till exempel lekar, motion, utevistelse, musik, pyssel och utfärder.
I dagen ingår också en vilostund.
Målsättningen med verksamheten är att främja barnets utveckling och lärande.
Barnet lär sig även sociala färdigheter.
Barnet får stöd i att lära sig det finska eller svenska språket, om hans/hennes modersmål är ett annat språk.
Om barnet behöver, kan hen även få specialundervisning.
Daghemmet är ändå inte en skola.
Barnen studerar inte skolämnen och har inte lektioner.
Barnen äter tre måltider under dagen: frukost, lunch och mellanmål.
Om ditt barn har en specialdiet ska du berätta om det för lärarna i småbarnspedagogiken.
I småbarnspedagogiken beaktas familjens religion eller livsåskådning.
På vissa orter finns det daghem, som fungerar på andra språk än finska eller svenska.
Vanligen börjar daghemsdagen på morgonen och tar slut på eftermiddagen.
Vissa daghem och familjedagvårdare har öppet dygnet runt med anledning av föräldrarnas arbete eller studier.
linkkiFinlands Flyktinghjälp:
Klubbar
Kommunerna, föreningar och församlingar ordnar dagklubbar för barn.
Klubbarna räcker vanligen ett par timmar.
I klubbarna ordnas handledda lekar, sång, pyssel och annat program.
linkkiUndervisnings- och kulturministeriet:
Information om småbarnspedagogikfinska _ svenska _ engelska
Söka bostad
Att hyra en bostad
Uppsägning av bostad
Att bli av med sin bostad
Konflikter med grannarna
Boendevardag
Fuktproblem
Rådgivningstjänster
Söka bostad
Jag hittar inte en förmånlig hyresbostad.
I de större städerna finns det bara få lediga hyresbostäder.
Bostäderna är dyrare nära stadens centrum.
Därför bor många finländare i ganska små bostäder.
Många bor också långt från centrum eller i en närliggande kommun och pendlar långt till jobbet.
Om du inte hittar en förmånlig bostad där du vill bo, fundera om du kan tänka dig att bo i en mindre bostad eller längre bort från centrum.
På många mindre orter finns det många lediga bostäder och priserna är lägre.
Om du planerar att flytta från en liten ort till en större stad, leta en bostad i förväg.
Läs mer på InfoFinlands sida Hyresbostad.
Jag lämnade en ansökan om en kommunal hyresbostad men jag har inte fått en bostad fastän det har gått tid.
Det finns inte tillräckligt många kommunala bostäder för alla som ansöker om dem.
Det lönar sig att ansöka om bostad på flera ställen.
Följ också utbudet av privata hyresbostäder.
Kom ihåg att uppdatera din ansökan när den är i kraft. Annars löper den ut.
Läs mer på InfoFinlands sida Hyresbostad.
Jag misstänker att jag har blivit diskriminerad när jag letade efter bostad.
Var får jag hjälp?
Enligt lag får hyresvärdar inte diskriminera någon till exempel på grund av etniskt ursprung, religion eller medborgarskap när de väljer hyresgäster.
En privat hyresvärd har dock rätt att själv välja hyresgästen till bostaden och hen behöver inte motivera sitt val.
Om du misstänker att du har blivit diskriminerad kan du fråga om råd till exempel hos diskrimineringsombudsmannens kundtjänst.
Diskrimineringsombudsmannens kundtjänstfinska _ svenska _ engelska
Att hyra en bostad
Måste jag betala ett förmedlingsarvode till bostadsförmedlaren när jag hyr en bostad?
Oftast betalar hyresvärden förmedlingsarvodet.
Du själv betalar förmedlingsarvodet endast om du har ingått ett skriftligt uppdragsavtal med bostadsförmedlaren om att söka en bostad åt dig.
Om du inte har ingått ett skriftligt uppdragsavtal får bostadsförmedlaren inte kräva dig på förmedlingsarvode.
Om hen försöker göra detta kan du polisanmäla hen.
Läs mer på InfoFinlands sida Brott.
Bostadsförmedlaren kräver att jag betalar hen för att få se bostaden.
Måste jag betala?
Du har rätt att se bostaden i förväg och bostadsförmedlaren kan inte kräva att få betalt för detta.
Om du har problem som rör förmedlingsarvodet kan du kontakta Konsumentrådgivningen.
linkkiKonkurrens- och konsumentverket:
Konsumentrådgivningfinska _ svenska _ engelska
Bostadsförmedlaren kräver att jag betalar en reservationsavgift för hyresbostaden.
Måste jag betala?
I Finland tillämpas inga reservationsavgifter för bostäder.
Du ska inte betala någonting förrän du har ett skriftligt hyresavtal för bostaden.
Läs mer om avgifterna för en hyresbostad, till exempel hyresdeposition, på InfoFinlands sida Hyresavtal.
Hyresvärden kräver att jag tecknar en hemförsäkring.
Var får jag en hemförsäkring?
Kan jag säga upp den senare?
Hemförsäkringar säljs av många försäkringsbolag i Finland.
Läs mer på InfoFinlands sida Vardagslivet i Finland.
Det är bra att teckna en hemförsäkring även om det inte krävs i hyresavtalet.
Det är inte tillrådligt att säga upp hemförsäkringen under tiden då du bor i bostaden.
Om du till exempel orsakar en vattenskada måste du själv betala hela renoveringskostnaden.
Fakturan kan uppgå till flera tiotusentals euro.
Vad bör jag beakta innan jag undertecknar hyresavtalet?
Gå och titta på bostaden innan du hyr den.
Kontrollera att bostaden verkligen existerar, alltså att bostaden har samma adress som står på avtalet.
Säkerställ också att bostaden är i det skick som har angetts till dig.
Kontrollera vad hyresavtalet säger till exempel om villkoren för hyresförhållandet och om uppsägningstiden.
Det är också bra att gå igenom bostaden och eventuella fel i bostaden med dess ägare eller hens representant.
Läs mer på InfoFinlands sida Hyresavtal.
När ska jag betala hyresdepositionen?
Betala hyresdepositionen först när du har ett skriftligt hyresavtal.
Hyresvärden kan ange ett konto på vilket du sätter in hyresdepositionen.
Ni kan också öppna ett separat konto för hyresdepositionen på banken.
Läs mer på InfoFinlands sida Hyresavtal.
Hyresvärden föreslog att vi gör ett muntligt hyresavtal.
Är ett muntligt avtal tillräckligt?
Gör hyresavtalet alltid skriftligt.
På så sätt kan du bevisa vad ni kommit överens om, om det skulle uppstå problem.
Förvara hyresavtalet noga.
Det finns brister i hyresbostaden.
Kan hyresvärden i efterhand kräva att jag ersätter för brister som jag inte har orsakat?
Det är bra att skriva upp felen i bostaden tillsammans med hyresvärden när hyresförhållandet inleds.
Du kan även ta fotografier där felen syns.
På så sätt säkerställer du att du inte ställs ansvarig för fel som du inte har orsakat.
Uppsägning av bostad
Jag sade upp min hyresbostad men hyresvärden kräver att jag betalar hyran tills hen hittar en ny hyresgäst.
Måste jag betala?
Om du har ett tills vidare gällande hyresavtal är uppsägningstiden vanligtvis en kalendermånad.
Tiden räknas från slutet av den månad då du säger upp avtalet.
När uppsägningstiden har löpt ut kan hyresvärden inte kräva dig på hyra.
Ett tidsbestämt hyresavtal får inte sägas upp under dess löptid.
Vid behov kan du försöka förhandla om att avsluta hyresavtalet tidigare.
Läs mer på InfoFinlands sida Hyresavtal.
Jag har ett tills vidare gällande hyresavtal.
Jag sade upp avtalet den 2 juni.
Hyresvärden kräver att jag betalar hyra även för juli.
Måste jag betala?
Om inget annat har avtalats i ditt hyresavtal räknas uppsägningstiden enligt lag från slutet av den månad under vilken du säger upp hyresavtalet.
Om du säger upp bostaden den 2 juni, börjar uppsägningstiden den 30 juni och den varar en månad.
Du måste alltså ännu betala hyra för juli.
Läs mer på InfoFinlands sida Hyresavtal.
Att bli av med sin bostad
Jag har inte råd att betala hyran.
Vad kan jag göra?
Kontakta hyresvärden så snart som möjligt och försök förhandla om en förlängning av betalningstiden.
Ta reda på om du kan skjuta upp andra betalningar för att kunna betala hyran.
Kontakta också din bank och ta reda på om banken kan ge dig ett lån så att du kan betala hyran.
Fråga hos FPA om du har rätt till bostadsbidrag eller något annat understöd.
Du kan även be om hjälp och råd vid kommunens skuldrådgivning eller socialverk eller en boenderådgivare vid kommunen eller hyreshusbolaget eller till exempel Garantistiftelsen.
Läs mer på InfoFinlands sida Ekonomiska problem.
Jag måste flytta ut på grund av skilsmässa.
Jag är dessutom rädd att jag kommer att förlora mitt uppehållstillstånd.
Vad kan jag göra?
På InfoFinlands sida Hyresbostad hittar du information om hur du kan söka en ny bostad.
Skilsmässan kan påverka ditt uppehållstillstånd om du har ett tidsbundet uppehållstillstånd på grund av familjeband.
I vissa situationer kan tillståndet dock förlängas om du fortfarande har nära anknytning till Finland, till exempel i form av en arbetsplats.
Läs mer på InfoFinlands sida Kan jag förlora mitt uppehållstillstånd.
Hyresvärden har hotat med att vräka mig från hyresbostaden på grund av högljutt liv.
Om du upprepade gånger bryter mot husets ordningsregler har hyresvärden rätt att häva hyresavtalet.
Försök att enas om saken med hyresvärden innan avtalet hävs.
Du kan också till exempel kontakta grannmedlingscentret Naapuruussovittelun keskus.
Jag var tvungen att flytta ut och jag har inte hittat en ny bostad.
Vad kan jag göra?
I Finland erbjuder kommunerna tjänster för bostadslösa.
Också många organisationer och församlingar hjälper bostadslösa.
Dessa tjänster är avsedda för människor som har en hemkommun i Finland.
Om du blir bostadslös ska du kontakta socialbyrån eller socialstationen i din hemkommun.
Läs mer på InfoFinlands sida Bostadslöshet.
Konflikter med grannarna
Min granne för oljud.
Vad kan jag göra?
Dina grannar får inte föra oljud till exempel på nätterna.
Om din granne ofta och på ett allvarligt sätt bryter mot ordningsreglerna, kan du kontakta disponenten eller hyresvärden.
Min granne klagar ständigt om oljud hos mig.
Hurdana ljud är tillåtna i ett höghus?
Bostadsaktiebolagets ordningsregler anger när det ska vara tyst i huset.
I ett höghus finns ordningsreglerna oftast i trapphuset.
Under de tysta timmarna får man inte vara högljudd, till exempel spela på instrument eller lyssna på musik på hög volym, men normalt liv är tillåtet.
Varifrån kan jag få hjälp vid konflikter med min granne?
Om du och din granne har en konflikt som ni inte klarar av att själva lösa, kan ni be om hjälp vid grannmedlingscentret Naapuruussovittelun keskus eller hos disponenten.
Grannmedling innebär att grannarna diskuterar och en utomstående medlare leder samtalet.
På mötet kan man komma överens om hur situationen ska lösas.
Medlingen är kostnadsfri.
Läs mer på webbplatsen för grannmedlingscentret Naapuruussovittelun keskus.
linkkiCentrum för grannmedling:
Information om grannmedlingfinska _ engelska
Boendevardag
Vad ska jag göra om jag glömmer nyckeln hemma?
I bostadsaktiebolag har fastighetsskötseln eller disponenten oftast kopior på nycklarna och de kan öppna dörren mot en avgift.
I höghus finns ett nummer nära entrédörren som du kan ringa i en sådan situation.
Hur sopsorterar jag rätt?
I Finland sorteras till exempel bioavfall, kartong, glas, metall, farligt avfall och blandavfall.
Läs mer på InfoFinlands sida Avfallshantering och återvinning.
Vad ska jag beakta när jag använder bastun i min bostad?
Du ska aldrig placera något ovanför bastuugnen, använda bastun som förråd eller torka tvätt i bastun, eftersom detta kan orsaka en brand.
Stäng alltid av en elektrisk bastuugn efter användning.
Läs mer på InfoFinlands sida Säkerheten i hemmet.
Vad gör jag när en vattenkran läcker?
Ring fastighetsskötseln som ditt bostadsaktiebolag har avtal med.
Fastighetsskötseln kan göra små reparationer, till exempel reparera en kran eller öppna upp ett avlopp.
Fuktproblem
Jag har fuktproblem eller andra fel i min bostad Vad gör jag?
Kontakta omedelbart fastighetsskötseln, disponenten eller hyresvärden.
Det är viktigt att felen åtgärdas snabbt, innan de förvärras.
När vi lagar mat uppstår det mycket fukt i köket.
Vad kan vi göra?
Om du inte har en mekanisk ventilation i ditt hem ska du öppna fönstren och vädra via dem.
Detta är särskilt viktigt om du upptäcker att det samlas vattenånga eller fukt på fönstren när du lagar mat.
Använd spisfläkten när du lagar mat.
Kontrollera att frånluftsventilerna är öppna.
Om du orsakar skador i bostaden måste du ersätta dem.
Läs mer på InfoFinlands sida Rättigheter och skyldigheter för boende.
Rådgivningstjänster
Var får jag hjälp och råd i boendefrågor?
Det finns många ställen där du kan be om råd i boendefrågor.
Läs mer på InfoFinlands sida Hyresbostad.
I Finland ordnas stödboende (tukiasuminen) och serviceboende (palveluasuminen) för dem som behöver stöd för att kunna bo självständigt.
Stöd- och serviceboende kan ordnas för
åldringar
handikappade
utvecklingsstörda
människor som återhämtar sig från problem med den mentala hälsan och missbrukarproblem.
Stöd- och serviceboende tillhandahålls av kommuner, organisationer och privata företagare.
Om stöd- eller serviceboende ansöks i hemkommunens socialverk (sosiaalivirasto).
Stödboende
Den som bor i en stödbostad klarar nästan självständigt av de dagliga bestyren.
Stödets omfattning beror på den boendes behov.
Det kan variera allt mellan dagliga till veckovisa hembesök.
En stödbostad kan antingen vara kundens egen ägarbostad, en hyresbostad eller någon annan bostadsform.
Hur länge man bor i stödbostad beror på kundens livssituation och behov.
Avsikten är att kunderna under sin tid i en stödbostad kommer till rätta med sitt liv i den mån att de kan övergå till självständigt boende.
Serviceboende
Serviceboende är en boendeform avsedd för sådana personer som behöver kontinuerlig hjälp men inte är i behov av anstaltsvård.
Serviceboendet omfattar både bostaden och tjänsterna som anknyter till boendet.
Invånaren står själv för boendekostnaderna.
Serviceboende kan ordnas i vanliga bostäder, i ett servicehus, i en servicebostadsgrupp eller i någon annan form.
Invånaren förfogar alltså över en egen bostad och tillgång till tjänster som anknyter till boendet.
Tjänsterna kan vara till exempel hemhjälp, måltidservice, tjänster i anslutning till den personliga hygienen, olika typer av säkerhetstjänster och hälsovårdstjänster.
Kostnader för serviceboende
Kostnaderna för serviceboendet beror på vem som levererar tjänsten.
Serviceboende tillhandahålls såväl av kommuner som av privata företag.
Priserna och tjänsterna varierar mycket.
När du ansöker om serviceboende är det bra att noga reda ut vad det kostar.
Det lönar sig att jämföra kommunalt ägda och privata servicehus.
Den boende betalar boendet och tjänsterna själv om det är möjligt.
Kommunen ska dock säkerställa att invånaren har råd med att bo i ett servicehus om han eller hon är i behov av serviceboende.
Kommunens socialverk kan hjälpa dig med att reda ut de olika boendealternativen.
Åldringar
Åldringar som dagligen behöver utomstående stöd och hjälp har rätt till serviceboende.
De kan själva välja hur mycket hjälp som ska ingå i serviceboendet.
Handikappade personer
Serviceboende ordnas för sådana handikappade personer som på grund av sitt handikapp eller sin sjukdom behöver hjälp för att klara av dagliga sysslor.
På InfoFinlands sida Tjänster för handikappade hittar du information om tjänster för handikappade.
Människor som återhämtar sig från problem med den mentala hälsan och missbrukarproblem
Människor som återhämtar sig från rusmedelsmissbruk eller problem med den mentala hälsan har möjlighet till stödboende.
Stödboendet hjälper dem att lära sig bo på egen hand och föra ett självständigt liv och stödjer dem i återhämtningen.
På InfoFinlands sida Missbruksproblem hittar du information om var du kan få hjälp om du eller en närstående till dig har problem med rusmedel.
linkkiMiljöministeriet:
Information om stöd- och serviceboendefinska _ svenska _ engelska
linkkiSocial- och hälsovårdsministeriet:
Boendetjänsterfinska _ svenska
Utbildningen i Finland håller en hög kvalitet.
Skillnaderna i olika skolors studieresultat är små och nästan alla avlägger grundskolan inom den utsatta tiden.
Förskoleundervisning, grundläggande utbildning och utbildning på andra stadiet är kostnadsfria och även därefter är utbildningen till största delen kostnadsfri.
Målet är att alla, oavsett familjens inkomster, ska ha möjlighet att få en högklassig utbildning och växa till aktiva medborgare.
Utbildningssystemet omfattar småbarnspedagogik, förskoleundervisning, grundläggande utbildning, utbildning på andra stadiet och högskoleutbildning.
Vuxenutbildningen är avsedd för vuxna och innehåller många alternativ från grundläggande utbildning till högskoleutbildning.
Småbarnspedagogik
I Finland har barnen rätt till småbarnspedagogik före skolåldern.
Småbarnspedagogiken ordnas i daghem och familjedagvården.
Barnet kan även delta i småbarnspedagogik tillsammans med föräldern i lekparker.
Barnet kan få minst 20 timmar småbarnspedagogik i veckan eller mer om föräldrarna arbetar eller struderar.
Målet är att stödja barnets utveckling och välbefinnande.
Barnet lär sig bland annat sociala färdigheter, att göra saker med händerna och olika kunskaper.
Barnet lär sig också olika färdigheter som hjälper hen att lära sig ytterligare nya saker.
Dagarna innehåller mycket lek och utevistelser.
Om barnet har ett annat modersmål än finska eller svenska, får hen stöd i lärandet av finska eller svenska.
Om barnet behöver, kan hen även få specialundervisning.
I Finland ordnar kommunerna småbarnspedagogiken.
Den finansieras med skattemedel och är därför förmånligare för familjerna.
I Finland finns även privat småbarnspedagogik.
De som arbetar med barnen är utbildade pedagoger inom småbarnsfostran och barnskötare.
Förskoleundervisning
I Finland ska barnen delta i förskoleundervisning under ett års tid innan läroplikten börjar.
Vanligtvis börjar förskoleundervisningen det år då barnet fyller sex år.
Förskoleundervisningen ordnas av kommunerna och är kostnadsfri för familjen.
Förskoleundervisningen ges av pedagoger inom småbarnsfostran som har avlagt universitetsexamen.
Förskoleundervisning ges vanligtvis fyra timmar om dagen från måndag till fredag.
Om föräldrarna arbetar eller studerar kan barnet utöver förskoleundervisningen även delta i småbarnspedagogiken.
Under detta år lär sig barnet kunskaper som hen har nytta av i skolan, till exempel bokstäver.
Barnen undervisas dock inte ännu i läsning.
Om barnet har ett annat modersmål än finska eller svenska, får hen stöd i lärandet av finska eller svenska.
Till dagen hör också lek och utevistelse.
Läs mer på InfoFinlands sida Förskoleundervisning.
Grundläggande utbildning
I Finland börjar den grundläggande utbildningen det år då barnet fyller sju år.
Alla barn som har sitt stadigvarande boende i Finland måste delta i den grundläggande utbildningen.
Grundskolan har nio årskurser.
Läroplikten upphör när barnet har fullgjort hela lärokursen för den grundläggande utbildningen eller det har förflutit tio år sedan läroplikten började.
I Finland reglerar lagstiftningen den grundläggande utbildningen.
Dessutom används nationella läroplansgrunder och lokala läroplaner.
Den grundläggande utbildningen ordnas av kommunerna.
Den finansieras med skattemedel och är därför kostnadsfri för familjerna.
I de lägre årskurserna har man cirka 20 undervisningstimmar i veckan och antalet ökar i de högre årskurserna.
Alla grundskolelärare i Finland har magisterexamen.
Klasslärarna i grundskolan, som undervisar årskurserna 1–6, har läst pedagogik.
Lärarna i årskurserna 7–9 har läst det ämne som de undervisar.
Lärare har stor frihet att planera undervisningen självständigt utifrån den nationella och lokala läroplanen.
På sistone har man i läroplanen betonat bland annat helheter som omfattar flera läroämnen, undersökning av vardagliga fenomen samt data- och kommunikationsteknik.
Barnen har ofta en och samma lärare under de sex första skolåren.
Läraren lär känna eleverna bra och kan utveckla undervisningen så att den passar dem.
Ett viktigt mål är att eleverna lär sig att tänka självständigt och tar eget ansvar för sitt lärande.
Läraren bedömer elevernas framsteg i skolan.
I den grundläggande utbildningen ges alla vitsord av läraren.
Det finns inga egentliga nationella prov.
Däremot följs inlärningsresultaten upp med urvalsbaserade bedömningar.
Dessa ordnas oftast i årskurs nio.
Om barnet eller den unga har flyttat till Finland nyligen, kan hen få förberedande undervisning före den grundläggande utbildningen.
Den förberedande undervisningen varar vanligtvis ett år.
Därefter kan eleven fortfarande läsa finska eller svenska som andraspråk, som S2-språk, om hen behöver stöd med språket.
Vuxna invandrare som inte har grundskolans avgångsbetyg från sitt eget land kan avlägga grundskolan på vuxengymnasiet.
Läs mer om den grundläggande utbildningen på InfoFinlands sida Grundläggande utbildning.
Utbildning på andra stadiet
De vanligaste alternativen efter grundskolan är gymnasium och yrkesutbildning.
Dessa är utbildning på andra stadiet.
Utbildning på andra stadiet är oftast kostnadsfri för studeranden.
Böcker och annat studiematerial måste man dock köpa själv.
Gymnasium
Gymnasiet är en allmänbildande utbildning som inte ger ett yrke.
I gymnasiet läser man samma ämnen som i den grundläggande utbildningen, med undervisningen är mer krävande och studierna mer självständiga.
På slutet avlägger studerandena vanligtvis studentexamen.
Gymnasiet tar 2–4 år, beroende på den studerande.
Efter gymnasiet kan man söka till universitet, yrkeshögskola eller gymnasiebaserad yrkesutbildning.
I de flesta gymnasieskolorna är undervisningsspråket finska eller svenska.
I de stora städerna finns några gymnasieskolor med något annat undervisningsspråk, till exempel engelska eller franska.
Vuxna kan avlägga gymnasiestudier på vuxengymnasiet.
Där kan man avlägga enskilda kurser eller hela gymnasielärokursen och studentexamen.
Undervisningen kan bestå av närundervisning, distansundervisning, webbundervisning och självständiga studier.
Läs mer om gymnasiestudierna på InfoFinlands sida Gymnasium.
Förberedande gymnasieutbildning
På gymnasiet behövs goda språkkunskaper.
Om studeranden har ett annat modersmål än finska eller svenska och saknar tillräckliga språkkunskaper för gymnasiestudierna, kan hen söka till förberedande gymnasieutbildning (LUVA).
Läs mer på InfoFinlands sida Förberedande gymnasieutbildning.
Yrkesutbildning
Yrkesutbildningen är mer praktiknära än gymnasieutbildningen.
En yrkesinriktad grundexamen kan avläggas på ungefär tre år.
Därefter kan man fortsätta studierna och avlägga yrkesexamen eller specialyrkesexamen.
En väsentlig del av studierna är inlärning på arbetsplatsen.
Om man vill, kan man efter yrkesutbildningen fortsätta studierna ända till högskoleutbildning.
Om man redan behärskar de färdigheter som krävs för examen, kan man också avlägga yrkesexamen eller specialyrkesexamen som yrkesprov.
Yrkesexamen kan även avläggas med läroavtal.
Då arbetar studeranden på en arbetsplats inom den egna branschen, får minst samma lön som en praktikant för arbetet och avlägger samtidigt sina studier.
Läs mer på InfoFinlands sida Yrkesutbildning.
Utbildning som handleder för yrkesutbildning
Om du inte har tillräckliga språkkunskaper eller studiefärdigheter för yrkesutbildning, kan du före yrkesutbildningen söka till utbildning som handleder för yrkesutbildning (VALMA).
Läs mer på InfoFinlands sida Utbildning som handleder för yrkesutbildning.
Högskoleutbildning
Efter studierna på andra stadiet kan du gå vidare till högskoleutbildning.
I Finland tillhandahålls högskoleutbildning av yrkeshögskolor och universitet.
Studierna på yrkeshögskola kan vara kostnadsfria eller avgiftsbelagda för studeranden.
Terminsavgift tas ut av personer som inte är medborgare i ett EU-/EES-land eller familjemedlem till en medborgare i ett EU-/EES-land och som avlägger en lägre eller högre högskoleexamen på engelska.
Läs mer på InfoFinlands sida Utländska studerande i Finland.
Yrkeshögskolor
På yrkeshögskolan är undervisningen mer praktiknära än på universitetet.
I undervisningen ingår även inlärning i arbetet.
Yrkeshögskoleexamen kan avläggas på 3,5–4,5 år.
Om man vill fortsätta studierna därefter och avlägga högre yrkeshögskoleexamen, måste man först skaffa sig tre år av arbetserfarenhet från samma område som examen.
Läs mer på InfoFinlands sida Yrkeshögskolor
Undervisningen på universitet är baserad på vetenskaplig forskning.
På universitet kan man avlägga lägre högskoleexamen på cirka tre år och därefter högre högskoleexamen på cirka två år.
Universiteten ordnar undervisning på engelska i vissa utbildningsprogram.
I de flesta utbildningsprogrammen är undervisningsspråket ändå finska eller svenska.
När man har avlagt magisterexamen, kan man ansöka om rätt till fortsatta studier och avlägga licentiat- eller doktorsexamen.
Läs mer på InfoFinlands sida Universitet.
Ansökan till utbildning
På InfoFinlands sida Ansökan till utbildning finns information om hur du ansöker till utbildning på andra stadiet och högskoleutbildning i Finland.
Om du planerar att studera i Finland, läs mer på InfoFinlands sida Utländska studerande i Finland och Studerande.
Andra studiemöjligheter
I Finland finns även många läroanstalter som erbjuder studier som inte leder till examen för människor i alla åldrar.
Största delen av dessa utbildningar är avsedda för vuxna.
Sådana läroanstalter är medborgarinstitut, folkhögskolor, sommaruniversitet, studiecenter och idrottsutbildningscenter.
Studierna är allmänbildande.
Du kan studera till exempel bland annat språk, estetiska ämnen, handarbete och kommunikation.
Oftast betalar den studerande en avgift för studierna.
I vissa situationer kan studierna vid dessa läroanstalter dock vara kostnadsfria.
Om till exempel utbildning i läs- och skrivkunnighet eller någon annan språkutbildning har godkänts till din integrationsplan, tas det inte ut någon avgift för studierna.
Språkutbildning
Om du vill läsa finska eller svenska, läs mer på InfoFinlands sida Finska och svenska språket.
På den här sidan har vi sammanställt de viktigaste rättigheter och skyldigheter för boende i Finland.
Du är skyldig
Att följa ordningsreglerna i ditt bostadsaktiebolag om du bor i ett höghus eller ett radhus.
I ordningsreglerna anges vanligtvis till exempel tiderna för när det ska vara tyst i huset.
Ofta innehåller de även anvisningar om användningen av gemensamma utrymmen i huset.
I ett höghus hittar du ordningsreglerna vanligtvis i trapphuset nära entrédörren.
Att se till att även dina gäster följer ordningsreglerna.
Att enbart använda bostaden för det avsedda ändamålet.
Om bostaden är avsedd att användas för boende, kan du inte bo på ett annat ställe och använda bostaden som lokal.
Du har rätt
Att leva ett normalt liv i ditt hem.
Bostadsaktiebolaget kan inte utfärda sådana ordningsregler som står i strid med lagen eller begränsar ett normalt liv i alltför stor omfattning.
Till hemfrid.
Dina grannar får inte störa din hemfrid till exempel genom att föra oljud mitt i natten.
Om en granne ofta bryter mot ordningsreglerna på ett allvarligt sätt, ska du först ta upp saken med grannen.
Om detta inte hjälper, kan du kontakta disponenten eller hyresvärden.
Hemfrid innebär också att du i regel själv får bestämma vem som har tillträde till ditt hem.
Hyresgästens rättigheter och skyldigheter
Du är skyldig
Att betala hyran i tid.
Hyresbeloppet anges i hyresavtalet.
Hyresvärden kan höja hyran i enlighet med vad som anges i hyresavtalet.
Att se till att hyresbostaden hålls i ett gott skick.
Att följa villkoren i hyresavtalet.
Om det till exempel anges i hyresavtalet att det är förbjudet att röka i bostaden, kan du inte röka i ditt hem.
Om hyresavtalet kräver att du har en hemförsäkring, måste du teckna en sådan.
Det är bra att teckna en hemförsäkring även om detta inte krävs i hyresavtalet.
Att fråga om tillstånd hos hyresvärden om du vill göra ändringar i bostaden, till exempel måla en vägg.
Utan tillstånd får du inte göra några ändringar, även om du skulle bekosta renoveringen själv.
Begär tillståndet skriftligt.
Att ersätta hyresvärden för skador som du åsamkar bostaden.
Att meddela hyresvärden om du upptäcker sådana fel i bostaden som hyresvärden ansvarar för.
Hyresvärden ansvarar till exempel för bostadens fasta inredning och ytmaterial.
Att meddela eventuella fel till fastighetsskötseln, till exempel en läckande kran.
Du har rätt
Att bo i hyreslägenheten enligt vad som anges i hyresavtalet.
Hyresvärden får endast beträda bostaden i vissa undantagsfall, till exempel för att övervaka reparationer i bostaden eller visa bostaden för köpare.
Även då måste hen försöka i förväg komma överens om detta med dig.
Att få ett skriftligt meddelande i förväg om hyran höjs.
I meddelandet ska det stå hur mycket och när hyran kommer att höjas och vad som är grunden till höjningen.
Till en uppsägningstid enligt lag.
Att häva hyresavtalet omedelbart om det är skadligt för hälsan att bo i bostaden.
Att hyra ut en del av bostaden till en annan person, om detta inte medför olägenhet för hyresvärden.
Att få ett förhandsmeddelande om reparationer.
Små reparationer ska meddelas 14 dagar i förväg och stora reparationer sex månader i förväg.
Brådskande reparationer kan dock göras utan ett meddelande.
Om det är svårt eller omöjligt att bo i bostaden under reparationerna, har du rätt att säga upp hyresavtalet eller får nedsatt hyra.
Detta måste du emellertid alltid komma överens om med hyresvärden.
Läs mer på InfoFinlands sida Hyresavtal.
Rättigheter och skyldigheter i en ägarbostad
I ett bostadsaktiebolag har du skyldighet att
Betala bolagsvederlag och eventuellt även finansieringsvederlag för bostadsaktiebolagets lån till bostadsaktiebolaget.
Vederlagen används till att sköta bostadsaktiebolaget, till exempel underhålla byggnaderna och gårdsområdet.
Se till att din bostad hålls i gott skick.
I förväg meddela till bostadsaktiebolagets disponent eller styrelse om du ska göra en sådan ändring i din bostad som kan påverka husets bärande konstruktioner, vattenledningar, fuktisolering, elledningar eller ventilationssystem.
Till exempel ska en badrumsrenovering alltid meddelas i förväg.
Genomföra renoveringar på ett sådant sätt att bygganden inte tar skada.
I Finland finns exakta bestämmelser till exempel om hurdant tätskikt ett badrum ska ha.
Meddela bostadsaktiebolaget eller disponenten, i praktiken vanligtvis allra först fastighetsskötseln, om det finns ett sådant fel i din bostad vars åtgärdande åligger bostadsaktiebolaget.
I ett bostadsaktiebolag har du följande rättigheter:
Förvalta den bostad vars aktier du äger.
Du får göra ändringar i din bostad.
Tänk på att renoveringen inte får medföra olägenhet till bostadsaktiebolaget eller de andra aktieägarna.
Hyra ut din bostad eller en del av den till en annan person.
Delta i stämmor och på dem påverka det som händer i bostadsaktiebolaget.
På en stämma kan du rösta om olika saker och kräva att ett ärende tas upp för behandling på stämman.
Bostadsaktiebolaget ska se till att husets konstruktioner, isolering, värmesystem, elledningar, vattenledningar och avlopp samt gårdsområden hålls i gott skick.
På stämman fattas beslut om reparationer gällande dessa.
I vissa bostadsaktiebolag har man beslutat att fördela ansvaret på ett annat sätt.
I detta fall står det i bolagsordningen vem som ansvarar för vad.
Om du inte har en stadigvarande bostad, och om du inte officiellt är hyresgäst eller underhyresgäst, är du bostadslös.
I Finland erbjuder kommunerna tjänster för bostadslösa.
Dessa tjänster är avsedda för personer som har hemkommun i Finland.
Om du blir bostadslös, ta då kontakt med socialbyrån eller socialstationen i din hemkommun.
Där får du hjälp när du söker bostad eller tillfällig inkvartering.
En tillfällig inkvartering kan vara ett hem för bostadslösa, ett natthärbärge eller en sådan bostad, som är avsedd för bostadslösa.
Utred din situation tillsammans med socialarbetaren: hur mycket kan du betala i hyra, och kan du få hyresstöd.
Du kan också vända dig till rådgivningstjänsten för invandrare i din kommun.
På InfoFinlands sida Hyresbostad får du information om hur du kan hitta en hyresbostad.
Bostadssituationen varierar mycket mellan olika orter.
Det finns lediga bostäder på till exempel många mindre orter i olika delar av Finland.
Inom huvudstadsregionen kan det vara svårt att hitta en bostad.
Du kan be om råd och hjälp också av Vailla vakinaista asuntoa ry.
Det är en organisation som erbjuder råd, stöd och vägledning i ärenden gällande boende och försöker förbättra de bostadslösas ställning i samhället.
Ohjaamo-verksamheten erbjuder råd och vägledning till unga bostadslösa.
Föreningen för bostadslösafinska _ engelska
Om du inte är stadigvarande bosatt i Finland
Om du inte bor stadigvarande i Finland och blir utan bostad, ta då kontakt med ditt lands beskickning i Finland.
Läs mer på InfoFinlands sida Ambassader i Finland.
Vailla vakinaista asuntoa ry har ett nattcafé, Kalkkers, som erbjuder bostadslösa en varm plats på natten från höst till vår.
Kalkkers håller öppet kl. kl. 22–6.
Det finns inga möjligheter att övernatta på nattcaféet, och det är inte heller drogfritt.
Där är det ingen som frågar om du har uppehållstillstånd.
Nattcaféet finns i Helsingfors på adressen Vasagatan 5, och telefonnumret är 050 443 1068.
På InfoFinlands sida I Finland utan uppehållstillstånd finns det mer information för papperslösa.
Nattcentret Kalkkersfinska
linkkiFlyktingrådgivningen rf:
Information om papperslöshetfinska _ engelska _ franska _ arabiska
Om din bostad har skadats
Om du har en hemförsäkring, och din bostad blir skadad till exempel vid en brand eller till följd av en vattenskada, kontakta då genast ditt försäkringsbolag.
Hemförsäkringen kan eventuellt ersätta hyran för en tillfällig bostad.
Läs mer om kortvarigt boende på InfoFinlands sida Tillfälligt boende.
Om du inte kan betala din hyra
Om du har ekonomiska problem, lönar det sig för dig att alltid först betala hyran och därefter andra räkningar och skulder.
Om du inte kan betala hyran, kontakta då hyresvärden och försök avtala om längre betalningstid.
Läs mer på InfoFinlands sida Ekonomiska problem.
På InfoFinlands sida Bostadsbidrag finns information om det bostadsbidrag som FPA betalar.
På den här sidan finns information om tjänsterna i Rovaniemi.
När du flyttar till ett stadigvarande boende i Rovaniemi ska du registrera dig som invånare i kommunen.
Du kan registrera dig vid magistraten.
Magistratens kontaktuppgifter och närmare anvisningar hittar du på magistratens webbplats.
Registrering av utlänningar i Finland
Adress:
PB 8183
(Statens ämbetshus)
Öppet mån–fre kl. 8–16.15
När du besöker magistraten ska du ta med dig
legitimation (till exempel pass)
uppehållstillstånd och uppehållskort (om du behöver uppehållstillstånd i Finland)
registreringsintyg över uppehållsrätten (om du är medborgare i ett EU-land)
äktenskapsintyg
dina barns födelseattester.
Observera att utländska handlingar ska vara legaliserade.
Registrering av utlänningarfinska _ svenska _ engelska
FPA-kort
tfn 020 435 4810 Öppet mån–fre kl. 9–16
Skattekort, övriga beskattningsärenden
Adress:
tfn 016 367 6000
Mer information om övriga beskattningsärenden: linkkiVerohallinto:
Skattefinska _ svenska _ engelska
På den här sidan finns information om tjänsterna i Rovaniemi.
När du flyttar till ett stadigvarande boende i Rovaniemi ska du registrera dig som invånare i kommunen.
Du kan registrera dig vid magistraten.
Magistratens kontaktuppgifter och närmare anvisningar hittar du på magistratens webbplats.
Registrering av utlänningar i Finland
Adress:
PB 8183
(Statens ämbetshus)
Öppet mån–fre kl. 8–16.15
När du besöker magistraten ska du ta med dig
legitimation (till exempel pass)
uppehållstillstånd och uppehållskort (om du behöver uppehållstillstånd i Finland)
registreringsintyg över uppehållsrätten (om du är medborgare i ett EU-land)
äktenskapsintyg
dina barns födelseattester.
Observera att utländska handlingar ska vara legaliserade.
Registrering av utlänningarfinska _ svenska _ engelska
FPA-kort
tfn 020 435 4810 Öppet mån–fre kl. 9–16
Skattekort, övriga beskattningsärenden
Adress:
tfn 016 367 6000
Mer information om övriga beskattningsärenden: linkkiVerohallinto:
Skattefinska _ svenska _ engelska
På den här sidan finns information om tjänsterna i Rovaniemi.
Annan allmän information i ämnet finns på InfoFinland-sidan Flytta till Finland.
Tillståndsärenden
Registrering som invånare
Den sociala tryggheten i Finland
Tillståndsärenden
Om du vill flytta till Finland måste du ha ett uppehållstillstånd eller så måste du
göra en registrering av EU-medborgares uppehållsrätt. Du kan ansöka om uppehållstillstånd elektroniskt via tjänsten Enter Finland eller genom att besöka Finlands ambassad utomlands eller något av Migrationsverkets serviceställen i Finland.
EU-medborgare ska också registrera sig på Migrationsverket.
Migrationsverket (Migri)
Servicestället i Rovaniemi
Information om uppehållstillståndfinska _ svenska _ engelska
Resedokumentfinska _ svenska _ engelska
linkkiEnterFinland :
Elektronisk ansökanfinska _ svenska _ engelska
Registrering som invånare
När du flyttar till Rovaniemi måste du registrera dig som invånare i kommunen.
Du kan registrera dig på ett av magistratens serviceställen.
Registreringen är viktig, för utan den kommer du inte att ha rätt till exempelvis social trygghet i Finland.
Magistraten i Lappland
Tfn 029 553 9208
Ta med dig följande när du besöker magistraten:
identitetsbevis (till exempel pass)
uppehållstillstånd och uppehållskort (om du behöver uppehållstillstånd i Finland)
registreringsbevis för uppehållsrätt (om du är EU-medborgare)
vigselbevis
födelseattester för barnen
Registrering av utlänningarfinska _ svenska _ engelska
Läs mer Registrering som invånare
Den sociala tryggheten i Finland
Du har rätt till de socialskyddsförmåner som FPA beviljar utifrån boende och arbete.
Du måste alltid lämna in en separat ansökan till FPA om de socialskyddsförmåner som du behöver i din livssituation.
FPA avgör om du har rätt att utnyttja socialskyddsförmånerna på basis av din ansökan.
FPA
Servicestället i Rovaniemi
Kontaktuppgifter till den landsomfattande telefontjänsten finska _ svenska _ engelska
Läs mer Den sociala tryggheten i Finland
Vi svarar på respons på följande språk: finska, svenska och engelska.
Tyvärr kan vi inte svara på respons som är skriven på andra språk.
Du märker väl att vi inte ger råd i hur du ska sköta dina ärenden.
Rådgivningstjänster hittar du på InfoFinlands sida Ring och fråga om råd.
Vi svarar på respons på följande språk: finska, svenska och engelska.
Tyvärr kan vi inte svara på respons som är skriven på andra språk.
Du märker väl att vi inte ger råd i hur du ska sköta dina ärenden.
Rådgivningstjänster hittar du på InfoFinlands sida Ring och fråga om råd.
Vi svarar på respons på följande språk: finska, svenska och engelska.
Tyvärr kan vi inte svara på respons som är skriven på andra språk.
Du märker väl att vi inte ger råd i hur du ska sköta dina ärenden.
Rådgivningstjänster hittar du på InfoFinlands sida Ring och fråga om råd.
Vanligtvis ska du sortera avfallet hemma innan du gör dig av med det.
Då avfallet sorteras rätt kan man använda materialet för att tillverka nya produkter.
Anvisningarna finns vanligtvis vid sopbehållarna vid ditt eget hus.
Om inte kan du kontakta kommunen eller din hyresvärd.
Kasta inte avfallet ut genom fönstret, i skogen eller på gatan.
Hela saker är inte avfall.
Du kan sälja dem på lopptorg eller på internet eller donera dem till välgörenhet eller återvinningscentraler.
I Finland är det vanligt att köpa använda saker och lätt att hitta använda saker i gott skick.
Hur sorteras avfall?
Sortera avfallet enligt material.
Lägg inte skräp, mat eller kemikaler i avloppet (WC:n).
För alltid farligt avfall till insamlingsställe.
Vid alla hus finns inte alltid samtliga insamlingskärl.
Information om allmänna insamlingsställen finns på adressen kierratys.info.
Du får inte föra ditt eget avfall till insamlingskärl avsedda för ett annat hus.
Du får inte heller lägga avfall från exempelvis ditt företag i sopkärlen avsedda för ditt eget hus.
Insamlingskärl som ofta finns vid husbolaget
Bioavfall (biojäte)
JA: matavfall, även härsken mat, kaffesump, hushållspapper, skal från frukter etc.
Bioavfall komposteras till mylla.
I vissa kommunerer separeras inledningsvis biogas från avfallet för att producera el och värme.
Papper (paperi)
JA: tidningar, reklam, kuvert etc.
NEJ: vått eller mycket smutsigt papper
Av pappret görs dagstidningar eller wc-papper.
Kartong (kartonki)
JA: mjölkförpackningar, papp, papperspåsar, kartongförpackningar
NEJ: våt eller mycket smutsig kartong
Av kartong görs exempelvis papprullar för hushållspapper.
Aluminium i förpackningarna återvinns även.
Glas (lasi)
JA: glasförpackningar (flaskor och matburkar)
NEJ: glasföremål, glaskärl, speglar, porslin
Av glaset tillverkas nya glasförpackningar.
Metall (metalli)
JA: metallföremål och förpackningar som till största delen utgörs av metall
Olika metaller sorteras maskinellt och används för att tillverka nya produkter.
Blandavfall (sekajäte) eller övrigt avfall
JA: Allt avfall som du inte kan eller önskar sortera.
NEJ: farligt avfall
Blandavfall bränns vanligtvis vid avfallsverk för att producera el och värme.
Övriga insamlingsställen
Farligt avfall (vaarallinen jäte)
JA: lysrör, energibesparingslampor, kemikalier med ett varningsmärke på förpackningen
VAR: Insamlingsställen för farligt avfall, se kierratys.info
JA: hemmets stora och små batterier, mobiltelefonens batteri
VAR: röda batteriinsamlingslådor i butiker och kiosker
Metallen i batterierna årervinns och de farliga ämnena hanteras på ett säkert sätt.
JA: alla leksaker och utrustning som fungerar med el eller batteri
VAR: små elapparater i butiker som säljer elektronik och större apparater vid insamlingsställen för elskrot, se kierratys.info.
Metall från elapparater (t.ex. guld) återvinns.
JA: påsar, gladpack, askar, emballage och övriga plastförpackningar
NEJ: PVC-plast (kod 03), plastleksaker, plastbehållare, plastsaker
Av plastförpackningar görs nya plastprodukter.
Hur kan man minska mängden avfall?
Frys ned mat som blir över.
Förvara maten rätt.
Drick kranvatten, det är gott och säkert i Finland.
Köp endast sådana saker du behöver.
Köp hållbara produkter.
Om du senare vill sälja dem kan du få betalt för dem.
Köp och sälj använda produkter.
Ta hand om dina saker och förvara dem enligt anvisningarna.
Avfallsinsamlingsstationerfinska
linkki4V:
Tips för boende(pdf, 1,5 Mt)finska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
FPA:s bostadsbidrag är avsett för boendekostnader.
FPA:s bostadsbidrag täcker bara en del av boendekostnaderna.
Du kan få bostadsbidrag om du har låga inkomster och bor stadigvarande i Finland.
Med stadigvarande boende i Finland avses att du har ditt egentliga hem i Finland och huvudsakligen också vistas i landet.
För att få bostadsbidrag måste du också du omfattas av den sociala tryggheten i Finland.
Fpa:s stöd för boendet är följande:
allmänt bostadsbidrag
bostadsbidrag för pensionstagare
bostadsunderstöd i samband med militärunderstöd för värnpliktiga och civiltjänstgörare.
Om pengarna inte räcker till för boendekostnaderna fastän du får bostadsbidrag, kan du ansöka om utkomststöd hos FPA.
Läs mer på InfoFinlands sida Ekonomiska problem.
Stöd för boendetfinska _ svenska _ engelska
Fpa:s allmänna bostadsbidrag
Stöd kan betalas till en person eller till ett hushåll (ruokakunta).
Till samma hushåll hör vanligtvis alla som stadigvarande bor i samma bostad.
Vanligen består ett hushåll av ett äkta par, sambor eller en familj.
Också en person kan vara ett hushåll.
Bostadsbidraget beviljas gemensamt för hushållet på basis av en ansökan.
Beakta att om du delar bostad med till exempel en vän och ni har ett gemensamt hyresavtal så anses ni höra till samma hushåll.
Om en av er däremot är huvudhyresgäst och den andra underhyresgäst och ni inte är nära släktingar, anses ni höra till olika hushåll.
Följande kan få allmänt bostadsbidrag
barnfamiljer
studerande
äkta par och registrerade par
sambor
ensamboende eller
de som bor i kollektiv.
Hurudana boendekostnader anses skäliga?
Stöd kan beviljas för fast bostad i Finland.
Det är i lagen fastställt vilka boendekostnader om kan anses vara skäliga då stödet beräknas.
Bostaden kan vara:
en hyresbostad
en ägarbostad
en bostadsrättsbostad
en delägarbostad.
Stöd betalas för hyra,vederlag och utgifter för skötseln av bostaden.
Utgifter för skötseln av bostaden är till exempel uppvärmningskostnader och vattenavgifter.
Också en del av räntan på bostadslånet iakttas.
Bostadsbidrag beviljas för skäliga boendekostnader.
I stora städer accepteras högre boendekostnader än på små orter.
Fpa betalar inte alla boendekostnader
En del av boendekostnaderna måste du betala själv.
För detta fastställs en bassjälvrisk.
Bassjälvriskandelens storlek beror på:
hur många vuxna och barn som hör till hushållet
hushållets bruttoinkomster (inkomster före skatt)
Om inkomsterna är mycket låga bortfaller bassjälvrisken.
Då bostadsbidraget kalkyleras avsätts 300 euro per månad av dina förvärvsinkomster.
Detta belopp påverkar inte ditt bostadsbidrag.
Detta kallas förvärvsinkomstavdrag (ansiotulovähennys).
Förvärvsinkomstavdrag görs separat för varje medlem i hushållet.
Bostadsbidrag beviljas endast för skäliga boendekostnader.
Vid fastställande av skäliga boendekostnader beaktas
kommunen där bostaden är belägen
antalet vuxna och barn i hushållets storlek
Om bostaden är större eller dyrare än vad lagen om allmänt bostadsbidrag tillåter växer den andel av boendekostnaderna som du betalar själv.
Det slutliga bostadsbidraget beräknas på följande sätt:
Bassjälvriskandelen dras först bort från boendekostnaderna.
Bostadsbidraget är 80 % av det kvarstående beloppet.
Anmäl ändringar till Fpa
Om dina inkomster, boende- eller familjeförhållanden eller andra omständigheter ändras ska du omgående anmäla ändringen till Fpa.
I Fpa:s beslut anges i detalj vilka omständigheter som bör anmälas.
Allmänt bostadsbidragfinska _ svenska _ engelska
Vad är ett hushållfinska _ svenska _ engelska
Att ansöka om bostadsbidrag
Du ansöker om allmänt bostadsbidrag hos FPA med en ansökan om allmänt bostadsbidrag (AT1).
Du kan också ansöka om bostadsbidraget på internet.
Till din ansökan ska du bifoga:
en kopia av hyresavtalet och en utredning över hyresbeloppet (hyresbostad)
ett intyg på vederlagets belopp och bostadslånet (ägarbostad)
löneverifikat, d.v.s. ett lönebesked som arbetsgivaren gett.
Om du bor i ett kollektiv ska du bifoga ett befullmäktigande av dem som du delar bostad med, d.v.s. en fullmakt att ansöka om bostadsbidrag för alla.
Skicka din ansökan till Fpa:s byrå eller skicka in den på internet.
Fpa betjänar sina kunder på sina byråer, per telefon och post samt via webbtjänsten som finns på FPA:s internetsidor.
När du sköter dina personliga ärenden på en Fpa-byrå ska du ha med dig något identitetsbevis, till exempel pass.
Att ansöka om bostadsbidragfinska _ svenska _ engelska
Om du är studerande kan du söka hyresbostäder som är speciellt avsedda för studerande.
Studentbostäder har ofta lägre hyra än vanliga bostäder.
Studentbostäder hyrs ut av studentbostadsstiftelser, universitetens studentkårer, nationer och vissa andra stiftelser.
Dessutom har vissa läroanstalter egna studenthem.
Fråga på din studieort var du kan söka en studentbostad.
Du kan söka bostad direkt när du blivit antagen till studier.
I de största städerna kan det ta flera veckor eller månader innan man får en bostad.
Om du får en studentbostad kan du vanligen bo i den under hela studietiden.
Du måste dock studera på heltid och framskrida i dina studier.
Hyresvärden kan säga upp hyresavtalet om du inte klarar tillräckligt många kurser.
Om du omfattas av den sociala tryggheten i Finland kan du ansöka om bostadsbidrag för boendekostnader hos FPA.
Läs mer om bostadsbidrag på InfoFinlands sida Bostadsbidrag.
Om studierna är den enda orsaken till att du bor i Finland, vistas du tillfälligt i Finland och omfattas därmed inte av den sociala tryggheten.
Om du också har andra orsaker att vistas i Finland, till exempel en arbetsplats, kan du omfattas av den sociala tryggheten i Finland.
Läs mer på InfoFinlands sida Den sociala tryggheten i Finland.
Studentbostäderfinska _ engelska
Information om den sociala tryggheten för studerandefinska _ svenska _ engelska
Brandsäkerhet
En brandvarnare kan rädda ditt liv.
Om en brand uppstår i din bostad avger brandvarnaren ett högljutt larm och du hinner ut i tid.
Se till att det finns tillräckligt många brandvarnare i ditt hem.
Brandvarnare säljs i varuhus och järnaffärer.
En brandvarnare räcker till 60 kvadratmeter.
Om ditt hem är till exempel 65 kvadratmeter stort behöver du två brandvarnare.
Om ditt hem har fler än en våning måste du räkna ytan separat för varje våning.
Det bör finnas en brandvarnare på varje våning.
Kontrollera regelbundet att brandvarnaren fungerar.
Byt batterier vid behov, gärna en gång per år.
Du ansvarar för brandvarnaren även om du bor i en hyresbostad.
Det finns ofta en bastu i finländska hem.
Även om du inte använder bastun får du aldrig placera något på bastuugnen, eftersom detta kan orsaka en brand.
Torka till exempel inte tvätten ovanför eller i närheten av bastuugnen.
Stäng alltid av en elektrisk bastuugn efter användning.
När du går hemifrån, kom ihåg att kontrollera att spisen och ugnen och till exempel strykjärnet är avstängda.
Det är bra att ha en brandsläckare hemma.
I vissa höghus finns det också en brandsläckare i trappuppgången.
Ta reda på var den närmaste brandsläckaren finns.
Se till att du har en släckningsfilt hemma.
Det är bra att förvara filten till exempel i närheten av spisen.
Lämna inte mat på en het spis utan uppsikt.
Var särskilt försiktig om du lagar mat på natten.
Laga inte mat om du är berusad.
Förvara inte föremål på spisen.
Barn, husdjur eller du själv kan av misstag vrida på spisen.
Då kan sakerna som ligger på spisen fatta eld.
Om fett börjar brinna när du lagar mat, kväv elden med till exempel ett kastrullock eller med en släckningsfilt.
Använd inte vatten.
Kom ihåg att stänga av elapparater efter användning.
Strykjärnet ska också kopplas loss från vägguttaget.
Använd inte elapparater som är i dåligt skick eller vars sladd är trasig.
Om en elapparat börjar brinna, använd inte vatten.
Kväv elden med till exempel en brandsläckare.
Om du har elektriska värmeelement eller värmeaggregat hemma, lägg inte tyger, kläder eller något annat på dem.
Lämna utrymme runt TV:n, mikrovågsugnen, kylskåpet och frysen.
Täck inte över dem.
Det är bra att en gång per år städa bort damm från frysens och kylskåpets bakgaller till exempel med dammsugaren, om möjligt.
Rök inte inomhus.
Lämna inte brinnande ljus utan uppsikt.
Tänd inte ljus i närheten av till exempel gardinerna, ens om du själv är i rummet.
Om en brand uppstår, ring nödnumret 112.
linkkiHelsingfors stads räddningsverk:
Brandsäkerhet i höghusfinska _ svenska _ engelska
linkkiRäddningsbranschens Centralorganisation i Finland:
Information om brandsäkerhetfinska _ svenska _ engelska
linkkiHelsingfors stad, Förortsprojektet:
Mitt hem i ett höghus(pdf, 6,56 MB)finska _ engelska _ ryska _ somaliska _ arabiska
linkkiHelsingfors stads räddningsverk:
Brandsäkerhet i småhusfinska _ svenska _ engelska
Så här undviker du vattenskador
Lämna inte tvättmaskinen eller diskmaskinen på när du går hemifrån.
Kontrollera regelbundet att vattenledningarna i ditt hem inte läcker och att det inte rinner ut vatten från hushållsapparaterna på golvet.
Stäng alltid kranen till tvätt- och diskmaskinen när du inte använder dem.
Det ska finnas ett läckageskydd av plast under kylskåpet, frysen och diskmaskinen.
Skyddet läggs på plats samtidigt som apparaten installeras.
Du får inte installera en diskmaskin själv, utan arbetet måste utföras av en fackman.
Om ett vattenläckage uppstår i ditt hem, försök stänga vattenledningens avstängningsventil.
Om du bor i höghus eller radhus, anmäl läckaget genast till journumret för husets servicebolag.
Om du bor i villa, kontakta en jourhavande rörfirma.
Elarbeten
I Finland är nätspänningen 230 volt.
I Finland utförs egentliga elarbeten endast av personer som är yrkesutbildade inom elbranschen.
Vissa små elarbeten får du utföra själv, om du kan.
Du kan till exempel själv:
byta en säkring
byta lampor
reparera en enfas skarvsladd (spänning 230 V)
hänga upp en lampa i taket med en upphängningsbygel
byta en hel enfas anslutningsledning (spänning 230 V) och stickkontakt i en elapparat, om den gamla gått sönder.
linkkiTukes:
Elarbeten som du får göra självfinska
Säkerhetslås skyddar mot inbrottstjuvar
Om du har ett säkerhetslås i ditt hem, lås det alltid då du inte är hemma.
Lås inte säkerhetslåset när du är hemma.
Om någon bryter in sig i ditt hem, ring nödnumret 112.
linkkiTukes:
Guiden Ett säkert hem för barnfinska _ svenska _ engelska
Birkalands räddningsverk:
Vad gör jag om det börjar brinna hemma?
Om videon väcker frågor hos dig kan du fråga mer av en expert.
Söka bostad
Att hyra en bostad
Uppsägning av bostad
Att bli av med sin bostad
Konflikter med grannarna
Boendevardag
Fuktproblem
Rådgivningstjänster
Söka bostad
Jag hittar inte en förmånlig hyresbostad.
I de större städerna finns det bara få lediga hyresbostäder.
Bostäderna är dyrare nära stadens centrum.
Därför bor många finländare i ganska små bostäder.
Många bor också långt från centrum eller i en närliggande kommun och pendlar långt till jobbet.
Om du inte hittar en förmånlig bostad där du vill bo, fundera om du kan tänka dig att bo i en mindre bostad eller längre bort från centrum.
På många mindre orter finns det många lediga bostäder och priserna är lägre.
Om du planerar att flytta från en liten ort till en större stad, leta en bostad i förväg.
Läs mer på InfoFinlands sida Hyresbostad.
Jag lämnade en ansökan om en kommunal hyresbostad men jag har inte fått en bostad fastän det har gått tid.
Det finns inte tillräckligt många kommunala bostäder för alla som ansöker om dem.
Det lönar sig att ansöka om bostad på flera ställen.
Följ också utbudet av privata hyresbostäder.
Kom ihåg att uppdatera din ansökan när den är i kraft. Annars löper den ut.
Läs mer på InfoFinlands sida Hyresbostad.
Jag misstänker att jag har blivit diskriminerad när jag letade efter bostad.
Var får jag hjälp?
Enligt lag får hyresvärdar inte diskriminera någon till exempel på grund av etniskt ursprung, religion eller medborgarskap när de väljer hyresgäster.
En privat hyresvärd har dock rätt att själv välja hyresgästen till bostaden och hen behöver inte motivera sitt val.
Om du misstänker att du har blivit diskriminerad kan du fråga om råd till exempel hos diskrimineringsombudsmannens kundtjänst.
Diskrimineringsombudsmannens kundtjänstfinska _ svenska _ engelska
Att hyra en bostad
Måste jag betala ett förmedlingsarvode till bostadsförmedlaren när jag hyr en bostad?
Oftast betalar hyresvärden förmedlingsarvodet.
Du själv betalar förmedlingsarvodet endast om du har ingått ett skriftligt uppdragsavtal med bostadsförmedlaren om att söka en bostad åt dig.
Om du inte har ingått ett skriftligt uppdragsavtal får bostadsförmedlaren inte kräva dig på förmedlingsarvode.
Om hen försöker göra detta kan du polisanmäla hen.
Läs mer på InfoFinlands sida Brott.
Bostadsförmedlaren kräver att jag betalar hen för att få se bostaden.
Måste jag betala?
Du har rätt att se bostaden i förväg och bostadsförmedlaren kan inte kräva att få betalt för detta.
Om du har problem som rör förmedlingsarvodet kan du kontakta Konsumentrådgivningen.
linkkiKonkurrens- och konsumentverket:
Konsumentrådgivningfinska _ svenska _ engelska
Bostadsförmedlaren kräver att jag betalar en reservationsavgift för hyresbostaden.
Måste jag betala?
I Finland tillämpas inga reservationsavgifter för bostäder.
Du ska inte betala någonting förrän du har ett skriftligt hyresavtal för bostaden.
Läs mer om avgifterna för en hyresbostad, till exempel hyresdeposition, på InfoFinlands sida Hyresavtal.
Hyresvärden kräver att jag tecknar en hemförsäkring.
Var får jag en hemförsäkring?
Kan jag säga upp den senare?
Hemförsäkringar säljs av många försäkringsbolag i Finland.
Läs mer på InfoFinlands sida Vardagslivet i Finland.
Det är bra att teckna en hemförsäkring även om det inte krävs i hyresavtalet.
Det är inte tillrådligt att säga upp hemförsäkringen under tiden då du bor i bostaden.
Om du till exempel orsakar en vattenskada måste du själv betala hela renoveringskostnaden.
Fakturan kan uppgå till flera tiotusentals euro.
Vad bör jag beakta innan jag undertecknar hyresavtalet?
Gå och titta på bostaden innan du hyr den.
Kontrollera att bostaden verkligen existerar, alltså att bostaden har samma adress som står på avtalet.
Säkerställ också att bostaden är i det skick som har angetts till dig.
Kontrollera vad hyresavtalet säger till exempel om villkoren för hyresförhållandet och om uppsägningstiden.
Det är också bra att gå igenom bostaden och eventuella fel i bostaden med dess ägare eller hens representant.
Läs mer på InfoFinlands sida Hyresavtal.
När ska jag betala hyresdepositionen?
Betala hyresdepositionen först när du har ett skriftligt hyresavtal.
Hyresvärden kan ange ett konto på vilket du sätter in hyresdepositionen.
Ni kan också öppna ett separat konto för hyresdepositionen på banken.
Läs mer på InfoFinlands sida Hyresavtal.
Hyresvärden föreslog att vi gör ett muntligt hyresavtal.
Är ett muntligt avtal tillräckligt?
Gör hyresavtalet alltid skriftligt.
På så sätt kan du bevisa vad ni kommit överens om, om det skulle uppstå problem.
Förvara hyresavtalet noga.
Det finns brister i hyresbostaden.
Kan hyresvärden i efterhand kräva att jag ersätter för brister som jag inte har orsakat?
Det är bra att skriva upp felen i bostaden tillsammans med hyresvärden när hyresförhållandet inleds.
Du kan även ta fotografier där felen syns.
På så sätt säkerställer du att du inte ställs ansvarig för fel som du inte har orsakat.
Uppsägning av bostad
Jag sade upp min hyresbostad men hyresvärden kräver att jag betalar hyran tills hen hittar en ny hyresgäst.
Måste jag betala?
Om du har ett tills vidare gällande hyresavtal är uppsägningstiden vanligtvis en kalendermånad.
Tiden räknas från slutet av den månad då du säger upp avtalet.
När uppsägningstiden har löpt ut kan hyresvärden inte kräva dig på hyra.
Ett tidsbestämt hyresavtal får inte sägas upp under dess löptid.
Vid behov kan du försöka förhandla om att avsluta hyresavtalet tidigare.
Läs mer på InfoFinlands sida Hyresavtal.
Jag har ett tills vidare gällande hyresavtal.
Jag sade upp avtalet den 2 juni.
Hyresvärden kräver att jag betalar hyra även för juli.
Måste jag betala?
Om inget annat har avtalats i ditt hyresavtal räknas uppsägningstiden enligt lag från slutet av den månad under vilken du säger upp hyresavtalet.
Om du säger upp bostaden den 2 juni, börjar uppsägningstiden den 30 juni och den varar en månad.
Du måste alltså ännu betala hyra för juli.
Läs mer på InfoFinlands sida Hyresavtal.
Att bli av med sin bostad
Jag har inte råd att betala hyran.
Vad kan jag göra?
Kontakta hyresvärden så snart som möjligt och försök förhandla om en förlängning av betalningstiden.
Ta reda på om du kan skjuta upp andra betalningar för att kunna betala hyran.
Kontakta också din bank och ta reda på om banken kan ge dig ett lån så att du kan betala hyran.
Fråga hos FPA om du har rätt till bostadsbidrag eller något annat understöd.
Du kan även be om hjälp och råd vid kommunens skuldrådgivning eller socialverk eller en boenderådgivare vid kommunen eller hyreshusbolaget eller till exempel Garantistiftelsen.
Läs mer på InfoFinlands sida Ekonomiska problem.
Jag måste flytta ut på grund av skilsmässa.
Jag är dessutom rädd att jag kommer att förlora mitt uppehållstillstånd.
Vad kan jag göra?
På InfoFinlands sida Hyresbostad hittar du information om hur du kan söka en ny bostad.
Skilsmässan kan påverka ditt uppehållstillstånd om du har ett tidsbundet uppehållstillstånd på grund av familjeband.
I vissa situationer kan tillståndet dock förlängas om du fortfarande har nära anknytning till Finland, till exempel i form av en arbetsplats.
Läs mer på InfoFinlands sida Kan jag förlora mitt uppehållstillstånd.
Hyresvärden har hotat med att vräka mig från hyresbostaden på grund av högljutt liv.
Om du upprepade gånger bryter mot husets ordningsregler har hyresvärden rätt att häva hyresavtalet.
Försök att enas om saken med hyresvärden innan avtalet hävs.
Du kan också till exempel kontakta grannmedlingscentret Naapuruussovittelun keskus.
Jag var tvungen att flytta ut och jag har inte hittat en ny bostad.
Vad kan jag göra?
I Finland erbjuder kommunerna tjänster för bostadslösa.
Också många organisationer och församlingar hjälper bostadslösa.
Dessa tjänster är avsedda för människor som har en hemkommun i Finland.
Om du blir bostadslös ska du kontakta socialbyrån eller socialstationen i din hemkommun.
Läs mer på InfoFinlands sida Bostadslöshet.
Konflikter med grannarna
Min granne för oljud.
Vad kan jag göra?
Dina grannar får inte föra oljud till exempel på nätterna.
Om din granne ofta och på ett allvarligt sätt bryter mot ordningsreglerna, kan du kontakta disponenten eller hyresvärden.
Min granne klagar ständigt om oljud hos mig.
Hurdana ljud är tillåtna i ett höghus?
Bostadsaktiebolagets ordningsregler anger när det ska vara tyst i huset.
I ett höghus finns ordningsreglerna oftast i trapphuset.
Under de tysta timmarna får man inte vara högljudd, till exempel spela på instrument eller lyssna på musik på hög volym, men normalt liv är tillåtet.
Varifrån kan jag få hjälp vid konflikter med min granne?
Om du och din granne har en konflikt som ni inte klarar av att själva lösa, kan ni be om hjälp vid grannmedlingscentret Naapuruussovittelun keskus eller hos disponenten.
Grannmedling innebär att grannarna diskuterar och en utomstående medlare leder samtalet.
På mötet kan man komma överens om hur situationen ska lösas.
Medlingen är kostnadsfri.
Läs mer på webbplatsen för grannmedlingscentret Naapuruussovittelun keskus.
linkkiCentrum för grannmedling:
Information om grannmedlingfinska _ engelska
Boendevardag
Vad ska jag göra om jag glömmer nyckeln hemma?
I bostadsaktiebolag har fastighetsskötseln eller disponenten oftast kopior på nycklarna och de kan öppna dörren mot en avgift.
I höghus finns ett nummer nära entrédörren som du kan ringa i en sådan situation.
Hur sopsorterar jag rätt?
I Finland sorteras till exempel bioavfall, kartong, glas, metall, farligt avfall och blandavfall.
Läs mer på InfoFinlands sida Avfallshantering och återvinning.
Vad ska jag beakta när jag använder bastun i min bostad?
Du ska aldrig placera något ovanför bastuugnen, använda bastun som förråd eller torka tvätt i bastun, eftersom detta kan orsaka en brand.
Stäng alltid av en elektrisk bastuugn efter användning.
Läs mer på InfoFinlands sida Säkerheten i hemmet.
Vad gör jag när en vattenkran läcker?
Ring fastighetsskötseln som ditt bostadsaktiebolag har avtal med.
Fastighetsskötseln kan göra små reparationer, till exempel reparera en kran eller öppna upp ett avlopp.
Fuktproblem
Jag har fuktproblem eller andra fel i min bostad Vad gör jag?
Kontakta omedelbart fastighetsskötseln, disponenten eller hyresvärden.
Det är viktigt att felen åtgärdas snabbt, innan de förvärras.
När vi lagar mat uppstår det mycket fukt i köket.
Vad kan vi göra?
Om du inte har en mekanisk ventilation i ditt hem ska du öppna fönstren och vädra via dem.
Detta är särskilt viktigt om du upptäcker att det samlas vattenånga eller fukt på fönstren när du lagar mat.
Använd spisfläkten när du lagar mat.
Kontrollera att frånluftsventilerna är öppna.
Om du orsakar skador i bostaden måste du ersätta dem.
Läs mer på InfoFinlands sida Rättigheter och skyldigheter för boende.
Rådgivningstjänster
Var får jag hjälp och råd i boendefrågor?
Det finns många ställen där du kan be om råd i boendefrågor.
Läs mer på InfoFinlands sida Hyresbostad.
I Finland ordnas stödboende (tukiasuminen) och serviceboende (palveluasuminen) för dem som behöver stöd för att kunna bo självständigt.
Stöd- och serviceboende kan ordnas för
åldringar
handikappade
utvecklingsstörda
människor som återhämtar sig från problem med den mentala hälsan och missbrukarproblem.
Stöd- och serviceboende tillhandahålls av kommuner, organisationer och privata företagare.
Om stöd- eller serviceboende ansöks i hemkommunens socialverk (sosiaalivirasto).
Stödboende
Den som bor i en stödbostad klarar nästan självständigt av de dagliga bestyren.
Stödets omfattning beror på den boendes behov.
Det kan variera allt mellan dagliga till veckovisa hembesök.
En stödbostad kan antingen vara kundens egen ägarbostad, en hyresbostad eller någon annan bostadsform.
Hur länge man bor i stödbostad beror på kundens livssituation och behov.
Avsikten är att kunderna under sin tid i en stödbostad kommer till rätta med sitt liv i den mån att de kan övergå till självständigt boende.
Serviceboende
Serviceboende är en boendeform avsedd för sådana personer som behöver kontinuerlig hjälp men inte är i behov av anstaltsvård.
Serviceboendet omfattar både bostaden och tjänsterna som anknyter till boendet.
Invånaren står själv för boendekostnaderna.
Serviceboende kan ordnas i vanliga bostäder, i ett servicehus, i en servicebostadsgrupp eller i någon annan form.
Invånaren förfogar alltså över en egen bostad och tillgång till tjänster som anknyter till boendet.
Tjänsterna kan vara till exempel hemhjälp, måltidservice, tjänster i anslutning till den personliga hygienen, olika typer av säkerhetstjänster och hälsovårdstjänster.
Kostnader för serviceboende
Kostnaderna för serviceboendet beror på vem som levererar tjänsten.
Serviceboende tillhandahålls såväl av kommuner som av privata företag.
Priserna och tjänsterna varierar mycket.
När du ansöker om serviceboende är det bra att noga reda ut vad det kostar.
Det lönar sig att jämföra kommunalt ägda och privata servicehus.
Den boende betalar boendet och tjänsterna själv om det är möjligt.
Kommunen ska dock säkerställa att invånaren har råd med att bo i ett servicehus om han eller hon är i behov av serviceboende.
Kommunens socialverk kan hjälpa dig med att reda ut de olika boendealternativen.
Åldringar
Åldringar som dagligen behöver utomstående stöd och hjälp har rätt till serviceboende.
De kan själva välja hur mycket hjälp som ska ingå i serviceboendet.
Handikappade personer
Serviceboende ordnas för sådana handikappade personer som på grund av sitt handikapp eller sin sjukdom behöver hjälp för att klara av dagliga sysslor.
På InfoFinlands sida Tjänster för handikappade hittar du information om tjänster för handikappade.
Människor som återhämtar sig från problem med den mentala hälsan och missbrukarproblem
Människor som återhämtar sig från rusmedelsmissbruk eller problem med den mentala hälsan har möjlighet till stödboende.
Stödboendet hjälper dem att lära sig bo på egen hand och föra ett självständigt liv och stödjer dem i återhämtningen.
På InfoFinlands sida Missbruksproblem hittar du information om var du kan få hjälp om du eller en närstående till dig har problem med rusmedel.
linkkiMiljöministeriet:
Information om stöd- och serviceboendefinska _ svenska _ engelska
linkkiSocial- och hälsovårdsministeriet:
Boendetjänsterfinska _ svenska
Möblerade hyresbostäder och lägenhetshotell
Fastighetsförmedlingsbyråer och privatpersoner hyr ut bostäder även för korta perioder.
Boendetiden kan vara från en dag till flera månader.
Oftast är bostäderna som hyrs ut för korta tider färdigt möblerade.
Storleken på hyran varierar beroende på bostadens läge.
Högst är priserna i centralt belägna bostäder.
Det finns även hemlika lägenhetshotell med lägenheter som till exempel kan ha ett eget kök.
Lägenhetshyrorna är vanligen i genomsnitt 100 euro per dygn.
Om du bor i lägenheten en längre tid, till exempel flera veckor, kan priset vara lägre.
linkkiForenom:
Möblerade bostäderfinska _ svenska _ engelska _ ryska
Möblerade bostäderfinska _ engelska
Hotell och vandrarhem
Att bo på hotell är en aning dyrare i Finland än i de flesta andra europeiska länder.
Priset på en hotellnatt varierar också mycket beroende på årstid och hotellets läge.
Ett enkel- eller dubbelrum kostar i genomsnitt 60–100 euro per dygn.
Ett förmånligare alternativ till hotell är att övernatta på ett vandrarhem, men i dessa är servicenivån inte lika hög och man har inte alltid möjlighet att få eget rum.
Priset för en natt är vanligen kring 20–50 euro.
Förmånligast övernattar man i delat rum.
Hotell i Finlandfinska _ svenska _ engelska _ ryska _ kinesiska
Heminkvartering
Du kan också bo som gäst hos vanliga finländare.
Oftast bor man i heminkvartering ett par dygn eller veckor.
Bostadens ägaren bestämmer priset.
Vanligen är detta dock ett lite förmånligare boendealternativ jämfört med ett hotell.
Heminkvarteringengelska _ franska _ spanska _ kinesiska _ tyska _ portugisiska _ italienska
Studentbostäder
Om du kommer till Finland för att studera kan du få en studentbostad där du får bo så länge som dina studier i Finland pågår.
Är du studerande lönar det sig att ansöka om en studentbostad då dessa vanligen är förmånligare än andra hyresbostäder.
Läs mer på InfoFinlands sida Boende för studerande.
Studentbostäderfinska _ engelska
På den här sidan har vi sammanställt de viktigaste rättigheter och skyldigheter för boende i Finland.
Du är skyldig
Att följa ordningsreglerna i ditt bostadsaktiebolag om du bor i ett höghus eller ett radhus.
I ordningsreglerna anges vanligtvis till exempel tiderna för när det ska vara tyst i huset.
Ofta innehåller de även anvisningar om användningen av gemensamma utrymmen i huset.
I ett höghus hittar du ordningsreglerna vanligtvis i trapphuset nära entrédörren.
Att se till att även dina gäster följer ordningsreglerna.
Att enbart använda bostaden för det avsedda ändamålet.
Om bostaden är avsedd att användas för boende, kan du inte bo på ett annat ställe och använda bostaden som lokal.
Du har rätt
Att leva ett normalt liv i ditt hem.
Bostadsaktiebolaget kan inte utfärda sådana ordningsregler som står i strid med lagen eller begränsar ett normalt liv i alltför stor omfattning.
Till hemfrid.
Dina grannar får inte störa din hemfrid till exempel genom att föra oljud mitt i natten.
Om en granne ofta bryter mot ordningsreglerna på ett allvarligt sätt, ska du först ta upp saken med grannen.
Om detta inte hjälper, kan du kontakta disponenten eller hyresvärden.
Hemfrid innebär också att du i regel själv får bestämma vem som har tillträde till ditt hem.
Hyresgästens rättigheter och skyldigheter
Du är skyldig
Att betala hyran i tid.
Hyresbeloppet anges i hyresavtalet.
Hyresvärden kan höja hyran i enlighet med vad som anges i hyresavtalet.
Att se till att hyresbostaden hålls i ett gott skick.
Att följa villkoren i hyresavtalet.
Om det till exempel anges i hyresavtalet att det är förbjudet att röka i bostaden, kan du inte röka i ditt hem.
Om hyresavtalet kräver att du har en hemförsäkring, måste du teckna en sådan.
Det är bra att teckna en hemförsäkring även om detta inte krävs i hyresavtalet.
Att fråga om tillstånd hos hyresvärden om du vill göra ändringar i bostaden, till exempel måla en vägg.
Utan tillstånd får du inte göra några ändringar, även om du skulle bekosta renoveringen själv.
Begär tillståndet skriftligt.
Att ersätta hyresvärden för skador som du åsamkar bostaden.
Att meddela hyresvärden om du upptäcker sådana fel i bostaden som hyresvärden ansvarar för.
Hyresvärden ansvarar till exempel för bostadens fasta inredning och ytmaterial.
Att meddela eventuella fel till fastighetsskötseln, till exempel en läckande kran.
Du har rätt
Att bo i hyreslägenheten enligt vad som anges i hyresavtalet.
Hyresvärden får endast beträda bostaden i vissa undantagsfall, till exempel för att övervaka reparationer i bostaden eller visa bostaden för köpare.
Även då måste hen försöka i förväg komma överens om detta med dig.
Att få ett skriftligt meddelande i förväg om hyran höjs.
I meddelandet ska det stå hur mycket och när hyran kommer att höjas och vad som är grunden till höjningen.
Till en uppsägningstid enligt lag.
Att häva hyresavtalet omedelbart om det är skadligt för hälsan att bo i bostaden.
Att hyra ut en del av bostaden till en annan person, om detta inte medför olägenhet för hyresvärden.
Att få ett förhandsmeddelande om reparationer.
Små reparationer ska meddelas 14 dagar i förväg och stora reparationer sex månader i förväg.
Brådskande reparationer kan dock göras utan ett meddelande.
Om det är svårt eller omöjligt att bo i bostaden under reparationerna, har du rätt att säga upp hyresavtalet eller får nedsatt hyra.
Detta måste du emellertid alltid komma överens om med hyresvärden.
Läs mer på InfoFinlands sida Hyresavtal.
Rättigheter och skyldigheter i en ägarbostad
I ett bostadsaktiebolag har du skyldighet att
Betala bolagsvederlag och eventuellt även finansieringsvederlag för bostadsaktiebolagets lån till bostadsaktiebolaget.
Vederlagen används till att sköta bostadsaktiebolaget, till exempel underhålla byggnaderna och gårdsområdet.
Se till att din bostad hålls i gott skick.
I förväg meddela till bostadsaktiebolagets disponent eller styrelse om du ska göra en sådan ändring i din bostad som kan påverka husets bärande konstruktioner, vattenledningar, fuktisolering, elledningar eller ventilationssystem.
Till exempel ska en badrumsrenovering alltid meddelas i förväg.
Genomföra renoveringar på ett sådant sätt att bygganden inte tar skada.
I Finland finns exakta bestämmelser till exempel om hurdant tätskikt ett badrum ska ha.
Meddela bostadsaktiebolaget eller disponenten, i praktiken vanligtvis allra först fastighetsskötseln, om det finns ett sådant fel i din bostad vars åtgärdande åligger bostadsaktiebolaget.
I ett bostadsaktiebolag har du följande rättigheter:
Förvalta den bostad vars aktier du äger.
Du får göra ändringar i din bostad.
Tänk på att renoveringen inte får medföra olägenhet till bostadsaktiebolaget eller de andra aktieägarna.
Hyra ut din bostad eller en del av den till en annan person.
Delta i stämmor och på dem påverka det som händer i bostadsaktiebolaget.
På en stämma kan du rösta om olika saker och kräva att ett ärende tas upp för behandling på stämman.
Bostadsaktiebolaget ska se till att husets konstruktioner, isolering, värmesystem, elledningar, vattenledningar och avlopp samt gårdsområden hålls i gott skick.
På stämman fattas beslut om reparationer gällande dessa.
I vissa bostadsaktiebolag har man beslutat att fördela ansvaret på ett annat sätt.
I detta fall står det i bolagsordningen vem som ansvarar för vad.
Om du inte har en stadigvarande bostad, och om du inte officiellt är hyresgäst eller underhyresgäst, är du bostadslös.
I Finland erbjuder kommunerna tjänster för bostadslösa.
Dessa tjänster är avsedda för personer som har hemkommun i Finland.
Om du blir bostadslös, ta då kontakt med socialbyrån eller socialstationen i din hemkommun.
Där får du hjälp när du söker bostad eller tillfällig inkvartering.
En tillfällig inkvartering kan vara ett hem för bostadslösa, ett natthärbärge eller en sådan bostad, som är avsedd för bostadslösa.
Utred din situation tillsammans med socialarbetaren: hur mycket kan du betala i hyra, och kan du få hyresstöd.
Du kan också vända dig till rådgivningstjänsten för invandrare i din kommun.
På InfoFinlands sida Hyresbostad får du information om hur du kan hitta en hyresbostad.
Bostadssituationen varierar mycket mellan olika orter.
Det finns lediga bostäder på till exempel många mindre orter i olika delar av Finland.
Inom huvudstadsregionen kan det vara svårt att hitta en bostad.
Du kan be om råd och hjälp också av Vailla vakinaista asuntoa ry.
Det är en organisation som erbjuder råd, stöd och vägledning i ärenden gällande boende och försöker förbättra de bostadslösas ställning i samhället.
Ohjaamo-verksamheten erbjuder råd och vägledning till unga bostadslösa.
Föreningen för bostadslösafinska
Om du inte är stadigvarande bosatt i Finland
Om du inte bor stadigvarande i Finland och blir utan bostad, ta då kontakt med ditt lands beskickning i Finland.
Läs mer på InfoFinlands sida Ambassader i Finland.
Vailla vakinaista asuntoa ry har ett nattcafé, Kalkkers, som erbjuder bostadslösa en varm plats på natten från höst till vår.
Kalkkers håller öppet kl. kl. 22–6.
Det finns inga möjligheter att övernatta på nattcaféet, och det är inte heller drogfritt.
Där är det ingen som frågar om du har uppehållstillstånd.
Nattcaféet finns i Helsingfors på adressen Vasagatan 5, och telefonnumret är 050 443 1068.
På InfoFinlands sida I Finland utan uppehållstillstånd finns det mer information för papperslösa.
Nattcentret Kalkkersfinska
linkkiFlyktingrådgivningen rf:
Information om papperslöshetfinska _ engelska _ franska _ arabiska
Om din bostad har skadats
Om du har en hemförsäkring, och din bostad blir skadad till exempel vid en brand eller till följd av en vattenskada, kontakta då genast ditt försäkringsbolag.
Hemförsäkringen kan eventuellt ersätta hyran för en tillfällig bostad.
Läs mer om kortvarigt boende på InfoFinlands sida Tillfälligt boende.
Om du inte kan betala din hyra
Om du har ekonomiska problem, lönar det sig för dig att alltid först betala hyran och därefter andra räkningar och skulder.
Om du inte kan betala hyran, kontakta då hyresvärden och försök avtala om längre betalningstid.
Läs mer på InfoFinlands sida Ekonomiska problem.
På InfoFinlands sida Bostadsbidrag finns information om det bostadsbidrag som FPA betalar.
En delägarbostad (osaomistusasunto) är ett bra sätt att skaffa en egen bostad om du inte kan köpa dig en egen bostad direkt.
Till en början köper du bara en del av bostaden och bor i bostaden på hyra.
Senare kan du köpa hela bostaden så att den blir helt och hållet din egen.
När du flyttar till en delägarbostad betalar du först ca 10-20 procent av bostadens pris.
Du kan ansöka om ett banklån för detta.
Efter detta bor du i bostaden på hyra och betalar hyra varje månad.
Vanligen är hyrestiden ca 5-12 år.
Du kan samtidigt köpa fler andelar i din bostad om du har kommit överens med byggherren om detta.
Efter hyrestiden köper du bostaden och den blir din egen.
Då har du en vanlig ägarbostad i ett bostadsaktiebolag.
Vissa delägarbostäder byggs med statligt stöd.
Då anger lagstiftningen till exempel hur lång hyrestiden i bostaden är och hur man kan avstå från bostaden.
Det finns även fritt finansierade delägarbostäder (vapaarahoitteinen osaomistusasunto).
Dessa är byggda utan statligt understöd.
Om du köper en fritt finansierad delägarbostad regleras inte hyrestiden eller andra avtalsvillkor i lagen.
Hur får man en delägarbostad?
Samfund och företag som låter bygga delägarbostäder informerar om nya och lediga bostäder.
Du får information om bostäderna även från kommunens bostadsbyrå.
Du kan ansöka om en delägarbostad med en ansökan riktad till bostadens byggherre.
Om delägarbostaden är byggd med statligt stöd kan du få en bostad om
dina inkomster inte är för stora; och
du inte har för stor förmögenhet.
Om du ansöker om en fritt finansierad bostad beaktas inte dina inkomster eller din förmögenhet.
linkkiKonkurrens- och konsumentverket:
Information om att bo i delägarbostadfinska _ svenska _ engelska
linkkiMiljöministeriet:
Information om att bo i delägarbostadfinska _ svenska _ engelska
FPA:s bostadsbidrag är avsett för boendekostnader.
FPA:s bostadsbidrag täcker bara en del av boendekostnaderna.
Du kan få bostadsbidrag om du har låga inkomster och bor stadigvarande i Finland.
Med stadigvarande boende i Finland avses att du har ditt egentliga hem i Finland och huvudsakligen också vistas i landet.
För att få bostadsbidrag måste du också du omfattas av den sociala tryggheten i Finland.
Fpa:s stöd för boendet är följande:
allmänt bostadsbidrag
bostadsbidrag för pensionstagare
bostadsunderstöd i samband med militärunderstöd för värnpliktiga och civiltjänstgörare.
Om pengarna inte räcker till för boendekostnaderna fastän du får bostadsbidrag, kan du ansöka om utkomststöd hos FPA.
Läs mer på InfoFinlands sida Ekonomiska problem.
Stöd för boendetfinska _ svenska _ engelska
Fpa:s allmänna bostadsbidrag
Stöd kan betalas till en person eller till ett hushåll (ruokakunta).
Till samma hushåll hör vanligtvis alla som stadigvarande bor i samma bostad.
Vanligen består ett hushåll av ett äkta par, sambor eller en familj.
Också en person kan vara ett hushåll.
Bostadsbidraget beviljas gemensamt för hushållet på basis av en ansökan.
Beakta att om du delar bostad med till exempel en vän och ni har ett gemensamt hyresavtal så anses ni höra till samma hushåll.
Om en av er däremot är huvudhyresgäst och den andra underhyresgäst och ni inte är nära släktingar, anses ni höra till olika hushåll.
Följande kan få allmänt bostadsbidrag
barnfamiljer
studerande
äkta par och registrerade par sambor
ensamboende eller
de som bor i kollektiv.
Hurudana boendekostnader anses skäliga?
Stöd kan beviljas för fast bostad i Finland.
Det är i lagen fastställt vilka boendekostnader om kan anses vara skäliga då stödet beräknas.
Bostaden kan vara:
en hyresbostad
en ägarbostad
en bostadsrättsbostad
en delägarbostad.
Stöd betalas för hyra,vederlag och utgifter för skötseln av bostaden.
Utgifter för skötseln av bostaden är till exempel uppvärmningskostnader och vattenavgifter.
Också en del av räntan på bostadslånet iakttas.
Bostadsbidrag beviljas för skäliga boendekostnader.
I stora städer accepteras högre boendekostnader än på små orter.
Fpa betalar inte alla boendekostnader
En del av boendekostnaderna måste du betala själv.
För detta fastställs en bassjälvrisk.
Bassjälvriskandelens storlek beror på:
hur många vuxna och barn som hör till hushållet
hushållets bruttoinkomster (inkomster före skatt)
Om inkomsterna är mycket låga bortfaller bassjälvrisken.
Då bostadsbidraget kalkyleras avsätts 300 euro per månad av dina förvärvsinkomster.
Detta belopp påverkar inte ditt bostadsbidrag.
Detta kallas förvärvsinkomstavdrag (ansiotulovähennys).
Förvärvsinkomstavdrag görs separat för varje medlem i hushållet.
Bostadsbidrag beviljas endast för skäliga boendekostnader.
Vid fastställande av skäliga boendekostnader beaktas
kommunen där bostaden är belägen
antalet vuxna och barn i hushållets storlek
Om bostaden är större eller dyrare än vad lagen om allmänt bostadsbidrag tillåter växer den andel av boendekostnaderna som du betalar själv.
Det slutliga bostadsbidraget beräknas på följande sätt:
Bassjälvriskandelen dras först bort från boendekostnaderna.
Bostadsbidraget är 80 % av det kvarstående beloppet.
Anmäl ändringar till Fpa
Om dina inkomster, boende- eller familjeförhållanden eller andra omständigheter ändras ska du omgående anmäla ändringen till Fpa.
I Fpa:s beslut anges i detalj vilka omständigheter som bör anmälas.
Allmänt bostadsbidragfinska _ svenska _ engelska
Vad är ett hushållfinska _ svenska _ engelska
Att ansöka om bostadsbidrag
Du ansöker om allmänt bostadsbidrag hos FPA med en ansökan om allmänt bostadsbidrag (AT1).
Du kan också ansöka om bostadsbidraget på internet.
Till din ansökan ska du bifoga:
en kopia av hyresavtalet och en utredning över hyresbeloppet (hyresbostad)
ett intyg på vederlagets belopp och bostadslånet (ägarbostad)
löneverifikat, d.v.s. ett lönebesked som arbetsgivaren gett.
Om du bor i ett kollektiv ska du bifoga ett befullmäktigande av dem som du delar bostad med, d.v.s. en fullmakt att ansöka om bostadsbidrag för alla.
Skicka din ansökan till Fpa:s byrå eller skicka in den på internet.
Fpa betjänar sina kunder på sina byråer, per telefon och post samt via webbtjänsten som finns på FPA:s internetsidor.
När du sköter dina personliga ärenden på en Fpa-byrå ska du ha med dig något identitetsbevis, till exempel pass.
Att ansöka om bostadsbidragfinska _ svenska _ engelska
Om du är studerande kan du söka hyresbostäder som är speciellt avsedda för studerande.
Studentbostäder har ofta lägre hyra än vanliga bostäder.
Studentbostäder hyrs ut av studentbostadsstiftelser, universitetens studentkårer, nationer och vissa andra stiftelser.
Dessutom har vissa läroanstalter egna studenthem.
Fråga på din studieort var du kan söka en studentbostad.
Du kan söka bostad direkt när du blivit antagen till studier.
I de största städerna kan det ta flera veckor eller månader innan man får en bostad.
Om du får en studentbostad kan du vanligen bo i den under hela studietiden.
Du måste dock studera på heltid och framskrida i dina studier.
Hyresvärden kan säga upp hyresavtalet om du inte klarar tillräckligt många kurser.
Om du omfattas av den sociala tryggheten i Finland kan du ansöka om bostadsbidrag för boendekostnader hos FPA.
Läs mer om bostadsbidrag på InfoFinlands sida Bostadsbidrag.
Om studierna är den enda orsaken till att du bor i Finland, vistas du tillfälligt i Finland och omfattas därmed inte av den sociala tryggheten.
Om du också har andra orsaker att vistas i Finland, till exempel en arbetsplats, kan du omfattas av den sociala tryggheten i Finland.
Läs mer på InfoFinlands sida Den sociala tryggheten i Finland.
Studentbostäderfinska _ engelska
Information om den sociala tryggheten för studerandefinska _ svenska _ engelska
Du får bo i en bostadsrättsbostad om du först betalar bostadsrättsavgiften (asumisoikeusmaksu).
Avgiften är ca 15 procent av bostadens pris.
Om du inte har pengar till bostadsrättsavgiften kan du ansöka om lån från banken.
Du kan dra av låneräntan i beskattningen.
Därefter betalar du varje månad en bestämd summa det vill säga bruksvederlag (käyttövastike).
Bruksvederlagets storlek beror på bostaden och orten.
Bruksvederlaget får inte vara större än hyran för bostäder av samma typ på samma område.
Om dina inkomster är små kan du ansöka om bostadsbidrag för bruksvederlaget.
Läs mera på InfoFinlands sida Bostadsbidrag.
Man kan inte köpa en bostadsrättsbostad.
Varför bostadsrättsbostad?
Bostadsrättsbostäder är inte förknippade med ekonomiska risker.
Därför är det en tryggare boendeform än en ägarbostad.
Du behöver inget stort lån för en bostadsrättsbostad.
När du vill flytta behöver du inte sälja bostaden.
Du kan bo i bostadsrättsbostaden så länge du vill.
Husets ägare kan inte säga upp bostadsrättskontraktet.
En bostadsrättsbostad är alltså mer bestående än en hyresbostad.
Du kan också låta bostadsrätten gå i arv.
Den boendes skyldigheter
Om du har en bostadsrättsbostad måste du själv vara fast bosatt i den.
Du kan hyra ut bostaden till någon annan under högst två år.
Du behöver dock tillstånd till detta av husets ägare.
Vem kan få en bostadsrättsbostad?
Om bostadsrättsbostaden inte har byggts med statsstöd kan husets ägare välja boende själv.
Om bostaden är byggd med statsstöd, kan du ansöka om
du har fyllt 18 år;
du inte har en ägarbostad på samma område; och
du inte har råd att skaffa en ägarbostad på samma område.
Din egendom beaktas ändå inte om du är över 55 år gammal eller flyttar från en bostadsrättsbostad till en annan bostadsrättsbostad.
Ibland kan det utöver dessa förekomma övriga villkor.
Hur ansöker man om en bostadsrättsbostad?
Det finns bostadsrättsbostäder i de största kommunerna.
Om du vill ha en bostadsrättsbostad, hämta först ett könummer på kommunens bostadsbyrå.
Du kan skaffa könummer i flera olika kommuner.
Könumret kostar ingenting.
Även om du har ett nummer behöver du inte ansöka om en bostad.
Välj sedan det hus där du vill ha en bostadsrättsbostad.
Anmäl dig till husets ägare.
Berätta också hurdan bostad du letar efter.
Du kan ansöka om bostadsrättsbostad i många olika hus.
Du kan bli tvungen att vänta länge på en bostad.
Bostadsrättsavtal
Då du får en bostad ska du göra ett skriftligt bostadsrättsavtal (asumisoikeussopimus) med husets ägare.
I bostadsrättsavtalet fastställs storleken på bostadsrättsavgiften, bruksvederlaget och övriga eventuella villkor.
Du kan flytta in i bostadsrättsbostaden när du har gjort bostadsrättskontraktet och betalat bostadsrättsavgiften.
När du flyttar ut
Om du vill flytta ut ur bostaden måste du göra en avträdelseanmälan (luopumisilmoitus) till husets ägare.
Du får bostadsrättsavgiften tillbaka, när du har avträtt bostaden.
linkkiKonkurrens- och konsumentverket:
Information om att bo i bostadsrättsbostadfinska _ svenska _ engelska
linkkiMiljöministeriet:
Att ansöka om en bostadsrättsbostadfinska _ svenska _ engelska
linkkiMiljöministeriet:
Information om att bo i bostadsrättsbostadfinska _ svenska _ engelska
Oy:
Bostadsrättsbostäderfinska
Bostadsrättsbostäderfinska
Bostadsrättsbostäderfinska
Bostadsrättsbostäderfinska
En ägarbostad är ofta på lång sikt förmånligare än en hyresbostad.
Största delen av finländarna bor ägarbostäder.
Det finns också andra alternativ än ägarbostad och hyresbostad.
Läs mer på InfoFinlands sidor Bostadsrättsbostad och Delägarbostad.
Bostadsaktie och fastighet
Då du köper en bostad, köper du antingen en bostadsaktie (asunto-osake) eller en fastighet (kiinteistö).
Höghuslägenheter och radhuslägenheter är bostadsaktier.
De finns i hus som ägs av ett bostadsaktiebolag.
Då du köper ett egnahemshus köper du en fastighet.
Fastigheten utgörs vanligen av egnahemshuset och dess tomt.
Hur hittar jag en ägarbostad?
När du letar efter en bostad är det bra att räkna med att det tar till och med flera månader.
Bostäder säljs av privatpersoner, fastighetsförmedlingar och byggherrar.
Bland annat på internet och i dagstidningar finns det annonser för bostäder som är till salu.
När du hittar en bostad som intresserar dig kan du komma överens med försäljaren om en visning av bostaden.
Ibland finns det i annonsen en utsatt tid då bostaden visas.
I så fall behöver du inte avtala en tid.
linkkiEtuovi.com:
Sökning av ägarbostäderfinska _ engelska
Sökning av ägarbostäderfinska
linkkiKonkurrens- och konsumentverket:
Information om att köpa en bostadfinska _ svenska _ engelska
Utred bostadens skick och andra frågor
Ta reda på allt som berör bostaden när du har hittat en bostad du tycker om.
Särskilt lönar det sig att utreda bostadens skick grundligt.
Om du tänker köpa en bostadsaktie, ta då även reda på vilka renoveringar bostadsaktiebolaget planerar och vad de kostar.
Till exempel ett stambyte kan kosta bostadsägaren många tiotusentals euro.
Säljarens och köparens ansvar vid bostadsköp
Den som säljer bostaden är ansvarig för fel i bostaden ännu under någon tid efter att bostaden har sålts.
Den som säljer en bostadsaktie är vanligen ansvarig för fel under två år.
För den som säljer en fastighet varar ansvaret fem år.
Enligt lagen måste den som säljer bostaden berätta om de fel som han/hon känner till innan försäljningen av bostaden.
Om det står klart att försäljaren har känt till fel i bostaden utan att berätta om detta för köparen, kan säljaren tvingas ersätta köparen för felet.
Granska om det finns fel i bostaden innan du köper en bostad.
Du kan inte efteråt kräva ersättning för fel, om
felet kan upptäckas vid granskning av bostaden; eller
du har känt till det innan köpet.
Det kan också finnas dolda fel i bostaden.
De är fel som ingen känner till.
Dolda fel är ofta till exempel fuktproblem.
Säljaren måste betala ut en ersättning till köparen ifall det i bostaden finns ett allvarligt fel, som skulle ha påverkat bostadsköpet ifall man känt till det.
Bostadslån
Vanligen betalar man bostaden med ett bostadslån (asuntolaina).
Vem som helst kan ansöka om ett bostadslån hos banken.
För att du ska kunna få ett bostadslån måste du ha tillräckliga inkomster för att betala tillbaka lånet utan problem.
På bankernas webbsidor finns det låneräknare.
Med hjälp av dem kan du på förhand uppskatta om du kan betala tillbaka lånet.
Om du inte är säker på huruvida banken ger dig ett lån lönar det sig att gå till banken och förhandla om lånet i god tid innan du köper bostaden.
Lånet återbetalas det vill säga amorteras en gång i månaden.
Dessutom måste man betala ränta (korko) för lånet till banken.
Du kan be om låneerbjudanden från flera banker och jämföra dem.
Olika lån har olika villkor.
Då du funderar på vilket lån du ska välja bör du beakta
hur stor ränta lånet har
hur stor summa du betalar tillbaka per månad
hur många år du återbetalar lånet
Märk väl att om räntorna stiger så stiger även lånekostnaderna.
Då stiger den månatliga avgiften eller också förlängs lånetiden.
Du kan dra av en del av räntan på bostadslånet i beskattningen.
linkkiKonkurrens- och konsumentverket:
Information om bostadslånfinska _ svenska _ engelska
Säkerhet och borgen för bostadslån
För ett bostadslån behövs det vanligen en säkerhet (vakuus).
Bostaden som du köper täcker en del av säkerheten, vanligen ca 70 procent.
Utöver detta behöver du en säkerhet för resten av lånesumman.
Du kan ordna säkerheten till exempel så att
Statsborgen kan utgöra högst 20 procent av lånet och högst 50 000 euro.
du ber en släktning eller vän gå i borgen för ditt lån.
Om du inte själv kan betala tillbaka lånet, blir borgensmannen tvungen att betala den summan som han eller hon gått i borgen för.
Du behöver ändå inte borgensmän för ditt lån om du har sparat ihop en del av bostadens pris på förhand, eller om du har annan egendom som duger som säkerhet för lånet.
linkkiMiljöministeriet:
Information om statsborgen för bostadslånfinska _ svenska _ engelska
Stöd vid bostadsköp
Staten beviljar räntestöd (korkotuki) för bostadslån.
Räntestöd beviljas för unga som skaffar sin första ägarbostad.
Det beviljas även för dem som köper eller bygger ett egnahemshus.
Läs mera på miljöministeriets sidor.
linkkiMiljöministeriet:
Information om räntestödetfinska _ svenska _ engelska
Överlåtelseskatt
När du köper en bostad måste du också betala överlåtelseskatt (varainsiirtovero).
Om du köper en bostadsaktie är överlåtelseskatten 2 procent av bostadens skuldfria pris.
Om du köper en fastighet är skatten 4 procent av bostadens skuldfria pris.
Du behöver ändå inte betala överlåtelseskatt om alla följande villkor uppfylls:
du är 18–39 år gammal
du har inte tidigare ägt en bostad i Finland eller något annat land
du äger minst 50 % av bostaden
du är själv fast bosatt i bostaden
linkkiSkatteförvaltningen:
Befrielse från överlåtelseskatt på första bostadfinska _ svenska _ engelska
Köpeanbud
När du är säker på att du vill och kan köpa en bostad kan du göra ett köpeanbud på bostaden.
Det lönar sig att göra ett skriftligt anbud.
Anbudet kan vara t.ex. 5-10 procent lägre än priset som säljaren har bett om för bostaden.
Säljaren kanske ändå inte vill sälja bostaden billigare.
Köpeanbudet är bindande.
Det betyder att du inte kan ta tillbaka anbudet.
Om du tar tillbaka köpeanbudet kan du bli tvungen att betala säljaren böter eller en handpenning.
Denna summa är vanligen några procent av bostadens pris.
Information om priser på sålda bostäderfinska _ svenska
Bostadsköp
Om säljaren av bostaden godtar köpeanbudet görs bostadsköpet upp i köparens bank.
Vanligen närvarar köparen och säljaren av bostaden samt bostadsförmedlaren, om en förmedlare har använts.
Köpebrevet är ett kontrakt där t.ex. bostadens pris, bostadens storlek, bostadens skick och datumet då köparen får tillgång till bostaden finns inskrivet.
Vanligen görs köpebrevet upp av banken eller bostadsförmedlaren.
Köparen har rätt att läsa köpebrevet före dagen då köpet genomförs.
Banken lånar bolånepengarna åt köparen, och summan flyttas över på säljarens konto.
Handpenning
Handpenningen (käsiraha) är en avgift, som betalas för bostaden på förhand.
Köparen kan betala handpenningen åt säljaren i det skedet då köpet förbereds.
Handpenningen är vanligen ca tre procent av bostadens pris.
Om du inte kan betala handpenningen av dina egna besparingar kan du låna summan av banken som en del av bostadslånet.
Kostnader för ägarbostad
På boendekostnaderna inverkar
bostadslånets storlek
bostadens storlek
bostadens skick
bostadens läge.
Bostadsaktie
Om du äger en bostadsaktie betalar du vanligen
ränta och amorteringar på bostadslånet
finansieringsvederlag (rahoitusvastike), om bostadsaktiebolaget har skulder
el och vatten
eventuella reparationsarbeten
Fastighet
Om du äger en fastighet betalar du vanligen
ränta och amorteringar på bostadslånet
fastighetsskatt (kiinteistövero)
el och vatten
värme
sophämtning
eventuella reparationsarbeten
Hushållsavfall
I Finland ska hushållsavfall sorteras i olika sopkärl.
Läs mer på InfoFinlands sida Avfallshantering och återvinning.
I Finland ordnas stödboende (tukiasuminen) och serviceboende (palveluasuminen) för dem som behöver stöd för att kunna bo självständigt.
Stöd- och serviceboende kan ordnas för
åldringar
handikappade
utvecklingsstörda
människor som återhämtar sig från problem med den mentala hälsan och missbrukarproblem.
Stöd- och serviceboende tillhandahålls av kommuner, organisationer och privata företagare.
Om stöd- eller serviceboende ansöks i hemkommunens socialverk (sosiaalivirasto).
Stödboende
Den som bor i en stödbostad klarar nästan självständigt av de dagliga bestyren.
Stödets omfattning beror på den boendes behov.
Det kan variera allt mellan dagliga till veckovisa hembesök.
En stödbostad kan antingen vara kundens egen ägarbostad, en hyresbostad eller någon annan bostadsform.
Hur länge man bor i stödbostad beror på kundens livssituation och behov.
Avsikten är att kunderna under sin tid i en stödbostad kommer till rätta med sitt liv i den mån att de kan övergå till självständigt boende.
Serviceboende
Serviceboende är en boendeform avsedd för sådana personer som behöver kontinuerlig hjälp men inte är i behov av anstaltsvård.
Serviceboendet omfattar både bostaden och tjänsterna som anknyter till boendet.
Invånaren står själv för boendekostnaderna.
Serviceboende kan ordnas i vanliga bostäder, i ett servicehus, i en servicebostadsgrupp eller i någon annan form.
Invånaren förfogar alltså över en egen bostad och tillgång till tjänster som anknyter till boendet.
Tjänsterna kan vara till exempel hemhjälp, måltidservice, tjänster i anslutning till den personliga hygienen, olika typer av säkerhetstjänster och hälsovårdstjänster.
Kostnader för serviceboende
Kostnaderna för serviceboendet beror på vem som levererar tjänsten.
Serviceboende tillhandahålls såväl av kommuner som av privata företag.
Priserna och tjänsterna varierar mycket.
När du ansöker om serviceboende är det bra att noga reda ut vad det kostar.
Det lönar sig att jämföra kommunalt ägda och privata servicehus.
Den boende betalar boendet och tjänsterna själv om det är möjligt.
Kommunen ska dock säkerställa att invånaren har råd med att bo i ett servicehus om han eller hon är i behov av serviceboende.
Kommunens socialverk kan hjälpa dig med att reda ut de olika boendealternativen.
Åldringar
Åldringar som dagligen behöver utomstående stöd och hjälp har rätt till serviceboende.
De kan själva välja hur mycket hjälp som ska ingå i serviceboendet.
Handikappade personer
Serviceboende ordnas för sådana handikappade personer som på grund av sitt handikapp eller sin sjukdom behöver hjälp för att klara av dagliga sysslor.
På InfoFinlands sida Tjänster för handikappade hittar du information om tjänster för handikappade.
Människor som återhämtar sig från problem med den mentala hälsan och missbrukarproblem
Människor som återhämtar sig från rusmedelsmissbruk eller problem med den mentala hälsan har möjlighet till stödboende.
Stödboendet hjälper dem att lära sig bo på egen hand och föra ett självständigt liv och stödjer dem i återhämtningen.
På InfoFinlands sida Missbruksproblem hittar du information om var du kan få hjälp om du eller en närstående till dig har problem med rusmedel.
linkkiMiljöministeriet:
Information om stöd- och serviceboendefinska _ svenska _ engelska
linkkiSocial- och hälsovårdsministeriet:
Boendetjänsterfinska _ svenska
Möblerade hyresbostäder och lägenhetshotell
Fastighetsförmedlingsbyråer och privatpersoner hyr ut bostäder även för korta perioder.
Boendetiden kan vara från en dag till flera månader.
Oftast är bostäderna som hyrs ut för korta tider färdigt möblerade.
Storleken på hyran varierar beroende på bostadens läge.
Högst är priserna i centralt belägna bostäder.
Det finns även hemlika lägenhetshotell med lägenheter som till exempel kan ha ett eget kök.
Lägenhetshyrorna är vanligen i genomsnitt 100 euro per dygn.
Om du bor i lägenheten en längre tid, till exempel flera veckor, kan priset vara lägre.
linkkiForenom:
Möblerade bostäderfinska _ svenska _ engelska _ ryska
Möblerade bostäderfinska _ engelska
Hotell och vandrarhem
Att bo på hotell är en aning dyrare i Finland än i de flesta andra europeiska länder.
Priset på en hotellnatt varierar också mycket beroende på årstid och hotellets läge.
Ett enkel- eller dubbelrum kostar i genomsnitt 60–100 euro per dygn.
Ett förmånligare alternativ till hotell är att övernatta på ett vandrarhem, men i dessa är servicenivån inte lika hög och man har inte alltid möjlighet att få eget rum.
Priset för en natt är vanligen kring 20–50 euro.
Förmånligast övernattar man i delat rum.
Hotell i Finlandfinska _ svenska _ engelska _ ryska _ kinesiska
Heminkvartering
Du kan också bo som gäst hos vanliga finländare.
Oftast bor man i heminkvartering ett par dygn eller veckor.
Bostadens ägaren bestämmer priset.
Vanligen är detta dock ett lite förmånligare boendealternativ jämfört med ett hotell.
Heminkvarteringengelska _ franska _ spanska _ kinesiska _ tyska _ portugisiska _ italienska
Studentbostäder
Om du kommer till Finland för att studera kan du få en studentbostad där du får bo så länge som dina studier i Finland pågår.
Är du studerande lönar det sig att ansöka om en studentbostad då dessa vanligen är förmånligare än andra hyresbostäder.
Läs mer på InfoFinlands sida Boende för studerande.
Studentbostäderfinska _ engelska
Ett hyresavtal kan vara
ett hyresavtal som gäller tillsvidare eller
ett tidsbestämt hyresavtal.
Ett hyresavtal som gäller tillsvidare (Toistaiseksi voimassa oleva vuokrasopimus) fortsätter fram till dess att hyresgästen eller hyresvärden säger upp avtalet.
Om du på förhand inte vet hur länge du kommer att bo i bostaden, är ett sådant avtal ett bra alternativ.
Ett tidsbestämt avtal (Määräaikainen vuokrasopimus) innebär att hyresvärden och hyresgästen från början kommer överens om när avtalet upphör.
Ett tidsbestämt hyresavtal upphör automatiskt utan uppsägning på den dag som antecknats i avtalet.
Om du fortfarande vill bo i bostaden efter detta behöver du ett nytt hyresavtal.
Det är inte möjligt att säga upp ett tidsbestämt avtal under dess giltighetstid.
Detta gäller för såväl hyresgästen som för hyresvärden.
Om du på förhand vet att du behöver bostaden enbart för en viss tid, är ett tidsbestämt hyresavtal ett bra alternativ.
Betalning av hyra
Hyra betalas vanligen en gång per månad.
Hyran ska betalas senast på förfallodatumet.
Förfallodagen har antecknats i hyresavtalet.
Betala hyran som en girering till hyresvärdens konto.
Du kan inte betala hyran med ett kreditkort.
Hyresgaranti
När du ingår ett hyresavtal i Finland, ska du nästan alltid betala en hyresgaranti.
Detta innebär att du på förhand betalar ett penningbelopp som motsvarar några månaders hyra till hyresvärden.
Vanligen motsvarar garantin beloppet på två månaders hyra.
Den kan högst uppgå till beloppet på tre månaders hyra.
Betala hyresgarantin senast på det datum som överenskommits i hyresavtalet.
I allmänhet får du nycklarna till bostaden när du betalat hyresgarantin.
När hyresavtalet upphör utförs en slutsyn i bostaden.
Hyresgarantin betalas tillbaka till dig i sin helhet om du
skött bostaden omsorgsfullt och
betalat alla avgifter som överenskommits med hyresvärden.
Om du söndrat bostaden eller inte betalat hela hyran, får du inte tillbaka hyresgarantin i sin helhet.
Hyresgarantin kan inte användas för att betala hyran för de sista månaderna.
Övriga avgifter
Reservera pengar för andra avgifter än hyran.
Vatten
Ofta ska du betala en vattenavgift för bostaden.
Betala vattenavgiften till hyresvärdens eller husbolagets konto på samma gång som du betalar hyra.
Beloppet på vattenavgiften beror ofta på det antal personer som bor i bostaden.
Om det finns en vattenmätare i bostaden, fastställs vattenavgiften enligt vattenkonsumtionen.
El
Ofta ska du själv ingå ett elavtal.
Du ingår ett elavtal genom att ringa ett elbolag och uppge ditt namn och din nya adress.
Om du vill hitta det förmånligaste priset, kan du jämföra olika elbolags priser.
Uppvärmning
Om bostaden har centralvärme, ingår uppvärmningen i allmänhet i hyran.
Om bostaden har oljevärme eller elvärme, ska avgiften ibland betalas separat.
Bastu, tvättstuga och bilplats
Det kostar i allmänhet att använda husbolagets bastu, tvättstuga och bilplatser.
I allmänhet ska dessa avgifter betalas direkt till husbolaget.
Avgifter i egnahemshus
Om du bor på hyra i ett egnahemshus, ska du ofta betala för uppvärmningen och avfallshanteringen.
Uppsägning av hyresavtal
Med uppsägningstid avses den tid som avtalet är i kraft efter att det sagts upp.
Uppsägningstiden gäller hyresavtal som gäller tillsvidare.
Uppsägningstiden för hyresgäster är en kalendermånad.
Du bör beakta hur uppsägningstiden räknas.
Uppsägningstiden börjar i allmänhet först från slutet av den månad då avtalet sägs upp.
Om du vill flytta ut från bostaden t.ex. 1.12, lönar det sig att säga upp bostaden senast 31.10.
Annars måste du betala hyra också för december månad.
Ge alltid ett skriftligt uppsägningsmeddelande.
Du måste kunna bevisa att du gett hyresvärden ett meddelande.
Hyresvärdens uppsägningstid beror på hur länge hyresavtalet varit i kraft.
Om avtalet varit i kraft i kortare tid än ett år, är uppsägningstiden tre månader.
Om avtalet varit i kraft i över ett år, är uppsägningstiden sex månader.
Ett tidsbestämt hyresavtal kan inte sägas upp mitt i avtalsperioden.
Underuthyrning
Med underuthyrning avses att hyresgästen hyr ut en del av bostaden till en annan person.
Hyresgästen har rätt att göra detta, om bostadens egentliga hyresvärd godkänner detta.
Innan du flyttar in som underhyresgäst ska du säkerställa att hyresgästen har rätt att ta en underhyresgäst.
Du är underhyresgäst också när du hyrt endast en del av en bostad och bostadsägaren själv bor i samma bostad.
Uppsägningstiden för en underhyresgäst är kortare än för en hyresgäst.
Uthyrning i andra hand
Med uthyrning i andra hand avses att hyresgästen hyr ut hela bostaden till en annan person.
Ett tillstånd av hyresvärden behövs alltid för detta.
Uppsägningsvillkoren är de samma som för hyresgäster.
Mallar för hyresavtalfinska
Guiden God hyressed(pdf, 546 kB)finska _ svenska _ engelska
Om du inte har en stadigvarande bostad, och om du inte officiellt är hyresgäst eller underhyresgäst, är du bostadslös.
I Finland erbjuder kommunerna tjänster för bostadslösa.
Dessa tjänster är avsedda för personer som har hemkommun i Finland.
Om du blir bostadslös, ta då kontakt med socialbyrån eller socialstationen i din hemkommun.
Där får du hjälp när du söker bostad eller tillfällig inkvartering.
En tillfällig inkvartering kan vara ett hem för bostadslösa, ett natthärbärge eller en sådan bostad, som är avsedd för bostadslösa.
Utred din situation tillsammans med socialarbetaren: hur mycket kan du betala i hyra, och kan du få hyresstöd.
Du kan också vända dig till rådgivningstjänsten för invandrare i din kommun.
På InfoFinlands sida Hyresbostad får du information om hur du kan hitta en hyresbostad.
Bostadssituationen varierar mycket mellan olika orter.
Det finns lediga bostäder på till exempel många mindre orter i olika delar av Finland.
Inom huvudstadsregionen kan det vara svårt att hitta en bostad.
Du kan be om råd och hjälp också av Vailla vakinaista asuntoa ry.
Det är en organisation som erbjuder råd, stöd och vägledning i ärenden gällande boende och försöker förbättra de bostadslösas ställning i samhället.
Ohjaamo-verksamheten erbjuder råd och vägledning till unga bostadslösa.
Föreningen för bostadslösafinska
Om du inte är stadigvarande bosatt i Finland
Om du inte bor stadigvarande i Finland och blir utan bostad, ta då kontakt med ditt lands beskickning i Finland.
Läs mer på InfoFinlands sida Ambassader i Finland.
Vailla vakinaista asuntoa ry har ett nattcafé, Kalkkers, som erbjuder bostadslösa en varm plats på natten från höst till vår.
Kalkkers håller öppet kl. kl. 22–6.
Det finns inga möjligheter att övernatta på nattcaféet, och det är inte heller drogfritt.
Där är det ingen som frågar om du har uppehållstillstånd.
Nattcaféet finns i Helsingfors på adressen Vasagatan 5, och telefonnumret är 050 443 1068.
På InfoFinlands sida I Finland utan uppehållstillstånd finns det mer information för papperslösa.
Nattcentret Kalkkersfinska
linkkiFlyktingrådgivningen rf:
Information om papperslöshetfinska _ engelska _ franska _ arabiska
Om din bostad har skadats
Om du har en hemförsäkring, och din bostad blir skadad till exempel vid en brand eller till följd av en vattenskada, kontakta då genast ditt försäkringsbolag.
Hemförsäkringen kan eventuellt ersätta hyran för en tillfällig bostad.
Läs mer om kortvarigt boende på InfoFinlands sida Tillfälligt boende.
Om du inte kan betala din hyra
Om du har ekonomiska problem, lönar det sig för dig att alltid först betala hyran och därefter andra räkningar och skulder.
Om du inte kan betala hyran, kontakta då hyresvärden och försök avtala om längre betalningstid.
Läs mer på InfoFinlands sida Ekonomiska problem.
På InfoFinlands sida Bostadsbidrag finns information om det bostadsbidrag som FPA betalar.
En delägarbostad (osaomistusasunto) är ett bra sätt att skaffa en egen bostad om du inte kan köpa dig en egen bostad direkt.
Till en början köper du bara en del av bostaden och bor i bostaden på hyra.
Senare kan du köpa hela bostaden så att den blir helt och hållet din egen.
När du flyttar till en delägarbostad betalar du först ca 10-20 procent av bostadens pris.
Du kan ansöka om ett banklån för detta.
Efter detta bor du i bostaden på hyra och betalar hyra varje månad.
Vanligen är hyrestiden ca 5-12 år.
Du kan samtidigt köpa fler andelar i din bostad om du har kommit överens med byggherren om detta.
Efter hyrestiden köper du bostaden och den blir din egen.
Då har du en vanlig ägarbostad i ett bostadsaktiebolag.
Vissa delägarbostäder byggs med statligt stöd.
Då anger lagstiftningen till exempel hur lång hyrestiden i bostaden är och hur man kan avstå från bostaden.
Det finns även fritt finansierade delägarbostäder (vapaarahoitteinen osaomistusasunto).
Dessa är byggda utan statligt understöd.
Om du köper en fritt finansierad delägarbostad regleras inte hyrestiden eller andra avtalsvillkor i lagen.
Hur får man en delägarbostad?
Samfund och företag som låter bygga delägarbostäder informerar om nya och lediga bostäder.
Du får information om bostäderna även från kommunens bostadsbyrå.
Du kan ansöka om en delägarbostad med en ansökan riktad till bostadens byggherre.
Om delägarbostaden är byggd med statligt stöd kan du få en bostad om
dina inkomster inte är för stora; och
du inte har för stor förmögenhet.
Om du ansöker om en fritt finansierad bostad beaktas inte dina inkomster eller din förmögenhet.
linkkiKonkurrens- och konsumentverket:
Information om att bo i delägarbostadfinska _ svenska _ engelska
linkkiMiljöministeriet:
Information om att bo i delägarbostadfinska _ svenska _ engelska
I Finland bor många människor i hyresbostäder.
Det som är bra med en hyresbostad är att det är lätt att byta bostad, eftersom du inte behöver sälja och köpa bostaden.
Men å andra sidan kan hyresvärden bestämma sig för att säga upp hyresavtalet, om han eller hon har en godtagbar anledning.
Då måste du flytta från hyresbostaden, även om du inte vill det.
På InfoFinlands sida Hyresavtal finns viktig information om uppsägning av hyresbostad, betalning av hyran, hyresdeposition och andra utgifter i en hyresbostad.
I större städer är det ofta svårare att hitta en lämplig hyresbostad. Även hyran är högre.
Reservera tillräckligt med tid för att hitta en bostad.
En del områden är väldigt populära. I sådana områden hyrs bostäderna ut mycket snabbt.
När du har hittat en lämplig bostad bör du snabbt bestämma dig om du vill ha den.
Då hyrsvärden väljer hyresgäst får han eller hon enligt lagen inte diskriminera någon exempelvis på grund av etniskt ursprung, religion eller nationalitet.
Läs mer på InfoFinlands sida Diskriminering och rasism.
Hur skaffar jag en hyresbostad?
När du letar efter en hyresbostad kan du leta efter annonser till exempel på internet.
Skriv in sökordet ”hyresbostad”.
Du kan även titta i lokaltidningarna.
Sökning av hyresbostäderfinska _ engelska
Sökning av hyresbostäderfinska
Privata hyresbostäder
Man får oftast en privat hyresbostad snabbare än en kommunal hyresbostad. Hyran för en privat bostad är ofta högre.
Du behöver inte anlita en bostadsmäklare för att söka bostad.
Du kan själv söka information om lediga bostäder.
Då behöver du inte heller betala mäklararvode (välityspalkkio).
Du kan söka privata hyresbostäder på internet och i lokaltidningar.
Du kan även publicera en egen annons.
Om du vill hyra en privat hyresbostad ska du kontakta den som hyr ut bostaden.
Kom överens om när du kan gå och titta på bostaden. En bostadsvisning ordnas oftast för alla intresserade på samma gång.
Samtidigt får du en ansökningsblankett.
Fyll i den om du vill flytta in i bostaden.
Om du vill att en mäklare söker en lämplig hyresbostad åt dig, ska du ingå ett skriftligt uppdragsavtal (toimeksiantosopimus) med mäklaren.
Du måste då betala mäklararvode till mäklaren.
Avtala om arvodet skriftligen på förhand.
Arvodet kan till exempel vara lika stort som en månads hyra.
Jämför olika mäklarbyråers priser på förhand.
När du hyr en privat bostad ska du göra ett hyresavtal med hyresvärden.
Läs mera på InfoFinlands sida Hyresavtal.
Priser på icke subventionerade hyresbostäderengelska
Kommunernas hyresbostäder
Även kommunerna äger hyresbostäder. De är ofta förmånligare än andra hyresbostäder.
Du kan söka boende i en hyresbostad som staten stödjer, om du har något av följande:
Finskt medborgarskap;
registrerat uppehållstillstånd;
uppehållskort;
uppehållstillstånd som är giltigt i minst ett år; eller
uppehållstillstånd för studerande.
Om du vill ansöka om en kommunal hyresbostad fyller du i ansökningsblanketten på bostadskontoret i din kommun.
Ofta kan du även fylla i och skicka blanketten på kommunens webbsida.
I en del kommuner är hyresbostäderna så populära att man kan vara tvungen att stå i kö mycket länge.
Köerna till bostäderna kan vara långa till exempel i huvudstadsregionen (Helsingfors, Esbo och Vanda), men det finns lediga bostäder på mindre orter runt om i Finland.
När hyresgästerna väljs beaktas
inkomster
egendom
behovet av bostad.
I Finland finns även många allmännyttiga samfund som har förmånliga hyresbostäder.
Priser på hyresbostäder med statliga stödengelska
Studentbostäder
Om du är studerande kan du söka en hyresbostad som är avsedd särskild för studerande. Studentbostäderna har oftast en lägre hyra än andra bostäder.
Läs mer på InfoFinlands sida Boende för studerande.
Bostadsansökan och bilagor
När du lämnar in en bostadsansökan kan du behöva också andra dokument som bilagor till ansökan.
Dessa beror på varifrån du söker bostaden.
senaste löneintyg
kopia på beskattningsbeslutet där din egendom framgår
intyg över lån
kopia på uppehållstillstånd eller pass om du inte är EU-medborgare.
Ofta granskas även den bostadssökandes kredituppgifter.
linkkiKonkurrens- och konsumentverket:
Att hyra en bostadfinska _ svenska _ engelska
Information för hyresgästenfinska _ svenska _ engelska
linkkiMiljöministeriet:
Information om hyresboendefinska _ svenska _ engelska
linkkiKonsumentförbundet ry:
Hyreshandboken(pdf, 1,11 MB)finska _ svenska _ ryska _ franska _ somaliska _ arabiska
Hyresbostadens utrustning
I utrustningen i en hyresbostad ingår nästan alltid köksskåpen, kylskåpet och spisen.
Även klädskåp och skåp i hallen ingår vanligtvis.
Duschen, vattenkranarna och toalettstolen hör alltid till utrustningen.
Hyresbostäder är vanligtvis inte möblerade.
Det händer dock att lägenheter hyrs ut med möbler.
Vilka möbler som ingår varierar.
Kontrollera alltid med hyresvärden vilka möbler som ingår.
Hushållsavfall
I Finland ska hushållsavfall sorteras i olika sopkärl.
Läs mer på InfoFinlands sida Avfallshantering och återvinning.
Rådgivningstjänster
Vill du söka råd om att hyra en bostad?
Finlands Konsumentförbund erbjuder råd och handledning både för hyresgäster och hyresvärder.
Finlands Konsumentförbunds rådgivningstjänst:
tfn 010 8022 40
tis-fre kl. 10–12 och tis kl. 17–19
Du kan ringa till tjänsten och endast betala lokalsamtalsavgift överallt i Finland.
Du kan fråga råd på tjänsten även på nätet genom att fylla i en blankett. Du får svar per e-post.
Även Marthaförbundet och Finlands flyktinghjälp erbjuder bostadsrådgivning åt invandrare.
linkkiKonsumentförbundet:
Boenderådgivningfinska
linkkiFlyktinghjälp:
Flyktinghjälpens regionkontorfinska
linkkiMarthaförbundet:
Kontaktuppgifter till Marthaförbundetfinska _ engelska
Om du är studerande kan du söka hyresbostäder som är speciellt avsedda för studerande.
Studentbostäder har ofta lägre hyra än vanliga bostäder.
Studentbostäder hyrs ut av studentbostadsstiftelser, universitetens studentkårer, nationer och vissa andra stiftelser.
Dessutom har vissa läroanstalter egna studenthem.
Fråga på din studieort var du kan söka en studentbostad.
Du kan söka bostad direkt när du blivit antagen till studier.
I de största städerna kan det ta flera veckor eller månader innan man får en bostad.
Om du får en studentbostad kan du vanligen bo i den under hela studietiden.
Du måste dock studera på heltid och framskrida i dina studier.
Hyresvärden kan säga upp hyresavtalet om du inte klarar tillräckligt många kurser.
Om du omfattas av den sociala tryggheten i Finland kan du ansöka om bostadsbidrag för boendekostnader hos FPA.
Läs mer om bostadsbidrag på InfoFinlands sida Bostadsbidrag.
Om studierna är den enda orsaken till att du bor i Finland, vistas du tillfälligt i Finland och omfattas därmed inte av den sociala tryggheten.
Om du också har andra orsaker att vistas i Finland, till exempel en arbetsplats, kan du omfattas av den sociala tryggheten i Finland.
Läs mer på InfoFinlands sida Den sociala tryggheten i Finland.
Studentbostäderfinska _ engelska
Information om den sociala tryggheten för studerandefinska _ svenska _ engelska
Du får bo i en bostadsrättsbostad om du först betalar bostadsrättsavgiften (asumisoikeusmaksu).
Avgiften är ca 15 procent av bostadens pris.
Om du inte har pengar till bostadsrättsavgiften kan du ansöka om lån från banken.
Du kan dra av låneräntan i beskattningen.
Därefter betalar du varje månad en bestämd summa det vill säga bruksvederlag (käyttövastike).
Bruksvederlagets storlek beror på bostaden och orten.
Bruksvederlaget får inte vara större än hyran för bostäder av samma typ på samma område.
Om dina inkomster är små kan du ansöka om bostadsbidrag för bruksvederlaget.
Läs mera på InfoFinlands sida Bostadsbidrag.
Man kan inte köpa en bostadsrättsbostad.
Varför bostadsrättsbostad?
Bostadsrättsbostäder är inte förknippade med ekonomiska risker.
Därför är det en tryggare boendeform än en ägarbostad.
Du behöver inget stort lån för en bostadsrättsbostad.
När du vill flytta behöver du inte sälja bostaden.
Du kan bo i bostadsrättsbostaden så länge du vill.
Husets ägare kan inte säga upp bostadsrättskontraktet.
En bostadsrättsbostad är alltså mer bestående än en hyresbostad.
Du kan också låta bostadsrätten gå i arv.
Den boendes skyldigheter
Om du har en bostadsrättsbostad måste du själv vara fast bosatt i den.
Du kan hyra ut bostaden till någon annan under högst två år.
Du behöver dock tillstånd till detta av husets ägare.
Vem kan få en bostadsrättsbostad?
Om bostadsrättsbostaden inte har byggts med statsstöd kan husets ägare välja boende själv.
Om bostaden är byggd med statsstöd, kan du ansöka om
du har fyllt 18 år;
du inte har en ägarbostad på samma område; och
du inte har råd att skaffa en ägarbostad på samma område.
Din egendom beaktas ändå inte om du är över 55 år gammal eller flyttar från en bostadsrättsbostad till en annan bostadsrättsbostad.
Ibland kan det utöver dessa förekomma övriga villkor.
Hur ansöker man om en bostadsrättsbostad?
Det finns bostadsrättsbostäder i de största kommunerna.
Om du vill ha en bostadsrättsbostad, hämta först ett könummer på kommunens bostadsbyrå.
Du kan skaffa könummer i flera olika kommuner.
Könumret kostar ingenting.
Även om du har ett nummer behöver du inte ansöka om en bostad.
Välj sedan det hus där du vill ha en bostadsrättsbostad.
Anmäl dig till husets ägare.
Berätta också hurdan bostad du letar efter.
Du kan ansöka om bostadsrättsbostad i många olika hus.
Du kan bli tvungen att vänta länge på en bostad.
Bostadsrättsavtal
Då du får en bostad ska du göra ett skriftligt bostadsrättsavtal (asumisoikeussopimus) med husets ägare.
I bostadsrättsavtalet fastställs storleken på bostadsrättsavgiften, bruksvederlaget och övriga eventuella villkor.
Du kan flytta in i bostadsrättsbostaden när du har gjort bostadsrättskontraktet och betalat bostadsrättsavgiften.
När du flyttar ut
Om du vill flytta ut ur bostaden måste du göra en avträdelseanmälan (luopumisilmoitus) till husets ägare.
Du får bostadsrättsavgiften tillbaka, när du har avträtt bostaden.
linkkiKonkurrens- och konsumentverket:
Information om att bo i bostadsrättsbostadfinska _ svenska _ engelska
linkkiMiljöministeriet:
Att ansöka om en bostadsrättsbostadfinska _ svenska _ engelska
linkkiMiljöministeriet:
Information om att bo i bostadsrättsbostadfinska _ svenska _ engelska
Oy:
Bostadsrättsbostäderfinska
Bostadsrättsbostäderfinska
Bostadsrättsbostäderfinska
Bostadsrättsbostäderfinska
Checklista för dig som flyttar
När du flyttar i Finland från en bostad till en annan:
Kom ihåg att göra flyttanmälan (muuttoilmoitus).
Du kan göra flyttanmälan högst en månad före flyttningsdagen, men den bör göras senast en vecka efter att du har flyttat.
Flyttanmälan ska alltid göras till magistraten (maistraatti).
Du kan göra flyttanmälan
på nätet
telefonledes på finska på numret 0295 535 535 eller på svenska på numret 0295 535 536 eller
på en blankett som du får på posten eller hos magistraten.
Om du bor i höghus eller radhus ska du alltid också komma ihåg att meddela husets disponent (isännöitsijä) att du flyttar.
Meddela din nya adress till alla instanser som skickar dig post.
Vissa organisationer och företag får din nya adress direkt från befolkningsregistret.
Du har ändå själv ansvaret för att dina fakturor skickas till rätt adress och betalas i tid.
Om du bor i en hyresbostad ska du komma ihåg att säga upp din gamla bostad i tid.
Det är bäst att göra uppsägningen skriftligt.
Kontrollera hur lång uppsägningstid du har för bostaden.
Vanligen är den en kalendermånad.
Läs mer på InfoFinlands sida Hyresavtal.
Om du har barn ska du se till att skaffa dem nya dagvårds- och skolplatser.
Du måste meddela daghemmet och skolan när barnen slutar där.
Samtidigt är det bra att anmäla barnen till det nya daghemmet eller den nya skolan.
Kom ihåg att skaffa eventuell flytthjälp i tid.
Bland annat vid månadsskift och på veckoslut är flyttfirmorna alltid upptagna.
Avtala med din tjänsteleverantör om överföringen av din internetanslutning i god tid så att det inte blir ett avbrott i servicen.
Säg upp ditt gamla elavtal innan du flyttar och gör upp ett nytt.
Det lönar sig att jämföra olika elbolags priser så att du hittar det förmånligaste.
Du får ett elavtal genom att ringa upp elbolaget och meddela ditt namn och din nya adress.
Om du flyttar till ett egnahemshus ska du också komma ihåg att teckna andra avtal, såsom avtal om vattenförsörjning och avfallshantering.
Om huset värms upp med olja ska du komma ihåg att kontrollera oljemängden.
Kontrollera om dina nuvarande försäkringar, som hemförsäkringen, är tillräckliga även för den nya bostaden.
Om du till exempel flyttar från höghus till egnahemshus behöver du förmodligen en annorlunda försäkring.
Städa den gamla bostaden innan du flyttar och töm vinden, källarförrådet och garaget på saker.
Om du bor i en hyresbostad ska du ge ägaren eller disponenten alla nycklar till den gamla bostaden.
linkkiFörbundet för ungdomsbostäder:
Ordlista om boendefinska
Flyttanmälanfinska _ svenska _ engelska
linkkiEnergimarknadsverket:
Jämför elpriserfinska
Flyttjänsterfinska _ engelska
Flyttjänsterfinska _ engelska _ ryska
Flyttjänsterfinska _ svenska _ engelska
När du flyttar till Finland
Om du vill ha information om praktiska frågor i anslutning till att du flyttar till Finland, läs mer på sidan Komihåglista för dig som flyttar till Finland.
Om du nyligen har flyttat till Finland, måste du registrera dig som invånare.
Lär mer på InfoFinlands sida Registrering som invånare.
Flytta från Finland
Planerar du att flytta från Finland till ett annat land?
Läs mer på InfoFinlands sida Flytta från Finland.
En ägarbostad är ofta på lång sikt förmånligare än en hyresbostad.
Största delen av finländarna bor ägarbostäder.
Det finns också andra alternativ än ägarbostad och hyresbostad.
Läs mer på InfoFinlands sidor Bostadsrättsbostad och Delägarbostad.
Bostadsaktie och fastighet
Då du köper en bostad, köper du antingen en bostadsaktie (asunto-osake) eller en fastighet (kiinteistö).
Höghuslägenheter och radhuslägenheter är bostadsaktier.
De finns i hus som ägs av ett bostadsaktiebolag.
Då du köper ett egnahemshus köper du en fastighet.
Fastigheten utgörs vanligen av egnahemshuset och dess tomt.
Hur hittar jag en ägarbostad?
När du letar efter en bostad är det bra att räkna med att det tar till och med flera månader.
Bostäder säljs av privatpersoner, fastighetsförmedlingar och byggherrar.
Bland annat på internet och i dagstidningar finns det annonser för bostäder som är till salu.
När du hittar en bostad som intresserar dig kan du komma överens med försäljaren om en visning av bostaden.
Ibland finns det i annonsen en utsatt tid då bostaden visas.
I så fall behöver du inte avtala en tid.
linkkiEtuovi.com:
Sökning av ägarbostäderfinska _ engelska
Sökning av ägarbostäderfinska
linkkiKonkurrens- och konsumentverket:
Information om att köpa en bostadfinska _ svenska _ engelska
Utred bostadens skick och andra frågor
Ta reda på allt som berör bostaden när du har hittat en bostad du tycker om.
Särskilt lönar det sig att utreda bostadens skick grundligt.
Om du tänker köpa en bostadsaktie, ta då även reda på vilka renoveringar bostadsaktiebolaget planerar och vad de kostar.
Till exempel ett stambyte kan kosta bostadsägaren många tiotusentals euro.
Säljarens och köparens ansvar vid bostadsköp
Den som säljer bostaden är ansvarig för fel i bostaden ännu under någon tid efter att bostaden har sålts.
Den som säljer en bostadsaktie är vanligen ansvarig för fel under två år.
För den som säljer en fastighet varar ansvaret fem år.
Enligt lagen måste den som säljer bostaden berätta om de fel som han/hon känner till innan försäljningen av bostaden.
Om det står klart att försäljaren har känt till fel i bostaden utan att berätta om detta för köparen, kan säljaren tvingas ersätta köparen för felet.
Granska om det finns fel i bostaden innan du köper en bostad.
Du kan inte efteråt kräva ersättning för fel, om
felet kan upptäckas vid granskning av bostaden; eller
du har känt till det innan köpet.
Det kan också finnas dolda fel i bostaden.
De är fel som ingen känner till.
Dolda fel är ofta till exempel fuktproblem.
Säljaren måste betala ut en ersättning till köparen ifall det i bostaden finns ett allvarligt fel, som skulle ha påverkat bostadsköpet ifall man känt till det.
Bostadslån
Vanligen betalar man bostaden med ett bostadslån (asuntolaina).
Vem som helst kan ansöka om ett bostadslån hos banken.
För att du ska kunna få ett bostadslån måste du ha tillräckliga inkomster för att betala tillbaka lånet utan problem.
På bankernas webbsidor finns det låneräknare.
Med hjälp av dem kan du på förhand uppskatta om du kan betala tillbaka lånet.
Om du inte är säker på huruvida banken ger dig ett lån lönar det sig att gå till banken och förhandla om lånet i god tid innan du köper bostaden.
Lånet återbetalas det vill säga amorteras en gång i månaden.
Dessutom måste man betala ränta (korko) för lånet till banken.
Du kan be om låneerbjudanden från flera banker och jämföra dem.
Olika lån har olika villkor.
Då du funderar på vilket lån du ska välja bör du beakta
hur stor ränta lånet har
hur stor summa du betalar tillbaka per månad
hur många år du återbetalar lånet
Märk väl att om räntorna stiger så stiger även lånekostnaderna.
Då stiger den månatliga avgiften eller också förlängs lånetiden.
Du kan dra av en del av räntan på bostadslånet i beskattningen.
linkkiKonkurrens- och konsumentverket:
Information om bostadslånfinska _ svenska _ engelska
Säkerhet och borgen för bostadslån
För ett bostadslån behövs det vanligen en säkerhet (vakuus).
Bostaden som du köper täcker en del av säkerheten, vanligen ca 70 procent.
Utöver detta behöver du en säkerhet för resten av lånesumman.
Du kan ordna säkerheten till exempel så att
Statsborgen kan utgöra högst 20 procent av lånet och högst 50 000 euro.
du ber en släktning eller vän gå i borgen för ditt lån.
Om du inte själv kan betala tillbaka lånet, blir borgensmannen tvungen att betala den summan som han eller hon gått i borgen för.
Du behöver ändå inte borgensmän för ditt lån om du har sparat ihop en del av bostadens pris på förhand, eller om du har annan egendom som duger som säkerhet för lånet.
linkkiMiljöministeriet:
Information om statsborgen för bostadslånfinska _ svenska _ engelska
Stöd vid bostadsköp
Staten beviljar räntestöd (korkotuki) för bostadslån.
Räntestöd beviljas för unga som skaffar sin första ägarbostad.
Det beviljas även för dem som köper eller bygger ett egnahemshus.
Läs mera på miljöministeriets sidor.
linkkiMiljöministeriet:
Information om räntestödetfinska _ svenska _ engelska
Överlåtelseskatt
När du köper en bostad måste du också betala överlåtelseskatt (varainsiirtovero).
Om du köper en bostadsaktie är överlåtelseskatten 2 procent av bostadens skuldfria pris.
Om du köper en fastighet är skatten 4 procent av bostadens skuldfria pris.
Du behöver ändå inte betala överlåtelseskatt om alla följande villkor uppfylls:
du är 18–39 år gammal
du har inte tidigare ägt en bostad i Finland eller något annat land
du äger minst 50 % av bostaden
du är själv fast bosatt i bostaden
linkkiSkatteförvaltningen:
Befrielse från överlåtelseskatt på första bostadfinska _ svenska _ engelska
Köpeanbud
När du är säker på att du vill och kan köpa en bostad kan du göra ett köpeanbud på bostaden.
Det lönar sig att göra ett skriftligt anbud.
Anbudet kan vara t.ex. 5-10 procent lägre än priset som säljaren har bett om för bostaden.
Säljaren kanske ändå inte vill sälja bostaden billigare.
Köpeanbudet är bindande.
Det betyder att du inte kan ta tillbaka anbudet.
Om du tar tillbaka köpeanbudet kan du bli tvungen att betala säljaren böter eller en handpenning.
Denna summa är vanligen några procent av bostadens pris.
Information om priser på sålda bostäderfinska _ svenska
Bostadsköp
Om säljaren av bostaden godtar köpeanbudet görs bostadsköpet upp i köparens bank.
Vanligen närvarar köparen och säljaren av bostaden samt bostadsförmedlaren, om en förmedlare har använts.
Köpebrevet är ett kontrakt där t.ex. bostadens pris, bostadens storlek, bostadens skick och datumet då köparen får tillgång till bostaden finns inskrivet.
Vanligen görs köpebrevet upp av banken eller bostadsförmedlaren.
Köparen har rätt att läsa köpebrevet före dagen då köpet genomförs.
Banken lånar bolånepengarna åt köparen, och summan flyttas över på säljarens konto.
Handpenning
Handpenningen (käsiraha) är en avgift, som betalas för bostaden på förhand.
Köparen kan betala handpenningen åt säljaren i det skedet då köpet förbereds.
Handpenningen är vanligen ca tre procent av bostadens pris.
Om du inte kan betala handpenningen av dina egna besparingar kan du låna summan av banken som en del av bostadslånet.
Kostnader för ägarbostad
På boendekostnaderna inverkar
bostadslånets storlek
bostadens storlek
bostadens skick
bostadens läge.
Bostadsaktie
Om du äger en bostadsaktie betalar du vanligen
ränta och amorteringar på bostadslånet
finansieringsvederlag (rahoitusvastike), om bostadsaktiebolaget har skulder
el och vatten
eventuella reparationsarbeten
Fastighet
Om du äger en fastighet betalar du vanligen
ränta och amorteringar på bostadslånet
fastighetsskatt (kiinteistövero)
el och vatten
värme
sophämtning
eventuella reparationsarbeten
Hushållsavfall
I Finland ska hushållsavfall sorteras i olika sopkärl.
Läs mer på InfoFinlands sida Avfallshantering och återvinning.
God morgon!
God dag!
God kväll!
God natt!
Välkommen!
Tack.
Var så god.
Förlåt.
Jag älskar dig.
Hur står det till?
Hejdå.
Adjö.
Jag förstår inte, kan du upprepa?
Jag talar inte finska.
Jag talar bara lite finska.
Talar du engelska/svenska?
Jag är lärare / ingenjör / studerande.
Vad är ditt telefonnummer / din e-postadress?
Var finns det en affär / ett apotek / en skola / ett daghem / en busstation / en metrostation?
Möblerade hyresbostäder och lägenhetshotell
Fastighetsförmedlingsbyråer och privatpersoner hyr ut bostäder även för korta perioder.
Boendetiden kan vara från en dag till flera månader.
Oftast är bostäderna som hyrs ut för korta tider färdigt möblerade.
Storleken på hyran varierar beroende på bostadens läge.
Högst är priserna i centralt belägna bostäder.
Det finns även hemlika lägenhetshotell med lägenheter som till exempel kan ha ett eget kök.
Lägenhetshyrorna är vanligen i genomsnitt 100 euro per dygn.
Om du bor i lägenheten en längre tid, till exempel flera veckor, kan priset vara lägre.
linkkiForenom:
Möblerade bostäderfinska _ svenska _ engelska _ ryska
Möblerade bostäderfinska _ engelska
Hotell och vandrarhem
Att bo på hotell är en aning dyrare i Finland än i de flesta andra europeiska länder.
Priset på en hotellnatt varierar också mycket beroende på årstid och hotellets läge.
Ett enkel- eller dubbelrum kostar i genomsnitt 60–100 euro per dygn.
Ett förmånligare alternativ till hotell är att övernatta på ett vandrarhem, men i dessa är servicenivån inte lika hög och man har inte alltid möjlighet att få eget rum.
Priset för en natt är vanligen kring 20–50 euro.
Förmånligast övernattar man i delat rum.
Hotell i Finlandfinska _ svenska _ engelska _ ryska _ kinesiska
Heminkvartering
Du kan också bo som gäst hos vanliga finländare.
Oftast bor man i heminkvartering ett par dygn eller veckor.
Bostadens ägaren bestämmer priset.
Vanligen är detta dock ett lite förmånligare boendealternativ jämfört med ett hotell.
Heminkvarteringengelska _ franska _ spanska _ kinesiska _ tyska _ portugisiska _ italienska
Studentbostäder
Om du kommer till Finland för att studera kan du få en studentbostad där du får bo så länge som dina studier i Finland pågår.
Är du studerande lönar det sig att ansöka om en studentbostad då dessa vanligen är förmånligare än andra hyresbostäder.
Läs mer på InfoFinlands sida Boende för studerande.
Studentbostäderfinska _ engelska
Ett hyresavtal kan vara
ett hyresavtal som gäller tillsvidare eller
ett tidsbestämt hyresavtal.
Ett hyresavtal som gäller tillsvidare (Toistaiseksi voimassa oleva vuokrasopimus) fortsätter fram till dess att hyresgästen eller hyresvärden säger upp avtalet.
Om du på förhand inte vet hur länge du kommer att bo i bostaden, är ett sådant avtal ett bra alternativ.
Ett tidsbestämt avtal (Määräaikainen vuokrasopimus) innebär att hyresvärden och hyresgästen från början kommer överens om när avtalet upphör.
Ett tidsbestämt hyresavtal upphör automatiskt utan uppsägning på den dag som antecknats i avtalet.
Om du fortfarande vill bo i bostaden efter detta behöver du ett nytt hyresavtal.
Det är inte möjligt att säga upp ett tidsbestämt avtal under dess giltighetstid.
Detta gäller för såväl hyresgästen som för hyresvärden.
Om du på förhand vet att du behöver bostaden enbart för en viss tid, är ett tidsbestämt hyresavtal ett bra alternativ.
Betalning av hyra
Hyra betalas vanligen en gång per månad.
Hyran ska betalas senast på förfallodatumet.
Förfallodagen har antecknats i hyresavtalet.
Betala hyran som en girering till hyresvärdens konto.
Du kan inte betala hyran med ett kreditkort.
Hyresgaranti
När du ingår ett hyresavtal i Finland, ska du nästan alltid betala en hyresgaranti.
Detta innebär att du på förhand betalar ett penningbelopp som motsvarar några månaders hyra till hyresvärden.
Vanligen motsvarar garantin beloppet på två månaders hyra.
Den kan högst uppgå till beloppet på tre månaders hyra.
Betala hyresgarantin senast på det datum som överenskommits i hyresavtalet.
I allmänhet får du nycklarna till bostaden när du betalat hyresgarantin.
När hyresavtalet upphör utförs en slutsyn i bostaden.
Hyresgarantin betalas tillbaka till dig i sin helhet om du
skött bostaden omsorgsfullt och
betalat alla avgifter som överenskommits med hyresvärden.
Om du söndrat bostaden eller inte betalat hela hyran, får du inte tillbaka hyresgarantin i sin helhet.
Hyresgarantin kan inte användas för att betala hyran för de sista månaderna.
Övriga avgifter
Reservera pengar för andra avgifter än hyran.
Vatten
Ofta ska du betala en vattenavgift för bostaden.
Betala vattenavgiften till hyresvärdens eller husbolagets konto på samma gång som du betalar hyra.
Beloppet på vattenavgiften beror ofta på det antal personer som bor i bostaden.
Om det finns en vattenmätare i bostaden, fastställs vattenavgiften enligt vattenkonsumtionen.
El
Ofta ska du själv ingå ett elavtal.
Du ingår ett elavtal genom att ringa ett elbolag och uppge ditt namn och din nya adress.
Om du vill hitta det förmånligaste priset, kan du jämföra olika elbolags priser.
Uppvärmning
Om bostaden har centralvärme, ingår uppvärmningen i allmänhet i hyran.
Om bostaden har oljevärme eller elvärme, ska avgiften ibland betalas separat.
Bastu, tvättstuga och bilplats
Det kostar i allmänhet att använda husbolagets bastu, tvättstuga och bilplatser.
I allmänhet ska dessa avgifter betalas direkt till husbolaget.
Avgifter i egnahemshus
Om du bor på hyra i ett egnahemshus, ska du ofta betala för uppvärmningen och avfallshanteringen.
Uppsägning av hyresavtal
Med uppsägningstid avses den tid som avtalet är i kraft efter att det sagts upp.
Uppsägningstiden gäller hyresavtal som gäller tillsvidare.
Uppsägningstiden för hyresgäster är en kalendermånad.
Du bör beakta hur uppsägningstiden räknas.
Uppsägningstiden börjar i allmänhet först från slutet av den månad då avtalet sägs upp.
Om du vill flytta ut från bostaden t.ex. 1.12, lönar det sig att säga upp bostaden senast 31.10.
Annars måste du betala hyra också för december månad.
Ge alltid ett skriftligt uppsägningsmeddelande.
Du måste kunna bevisa att du gett hyresvärden ett meddelande.
Hyresvärdens uppsägningstid beror på hur länge hyresavtalet varit i kraft.
Om avtalet varit i kraft i kortare tid än ett år, är uppsägningstiden tre månader.
Om avtalet varit i kraft i över ett år, är uppsägningstiden sex månader.
Ett tidsbestämt hyresavtal kan inte sägas upp mitt i avtalsperioden.
Underuthyrning
Med underuthyrning avses att hyresgästen hyr ut en del av bostaden till en annan person.
Hyresgästen har rätt att göra detta, om bostadens egentliga hyresvärd godkänner detta.
Innan du flyttar in som underhyresgäst ska du säkerställa att hyresgästen har rätt att ta en underhyresgäst.
Du är underhyresgäst också när du hyrt endast en del av en bostad och bostadsägaren själv bor i samma bostad.
Uppsägningstiden för en underhyresgäst är kortare än för en hyresgäst.
Uthyrning i andra hand
Med uthyrning i andra hand avses att hyresgästen hyr ut hela bostaden till en annan person.
Ett tillstånd av hyresvärden behövs alltid för detta.
Uppsägningsvillkoren är de samma som för hyresgäster.
Mallar för hyresavtalfinska
Guiden God hyressed(pdf, 546 kB)finska _ svenska _ engelska
Finland är ett tvåspråkigt land
Finland har två officiella språk, finska och svenska.
Båda språken har långa traditioner i Finland.
Ungefär 90 procent av finländarna har finska som modersmål och ungefär fem procent av finländarna har svenska som modersmål.
När du uträttar ärenden med statliga myndigheter, till exempel vid arbets- och näringsbyrån (työ- ja elinkeinotoimisto), kan du använda endera språket.
Svenska talas mest på Finlands väst- och sydkust.
På somliga orter är svenskan vanligare än finskan.
Kontrollera vilket som är det vanligaste språket på din ort.
Kommunerna kan vara antingen enspråkiga eller tvåspråkiga.
I tvåspråkiga kommuner kan du använda antingen finska eller svenska när du uträttar ärenden med anställda inom kommunen, till exempel på socialbyrån (sosiaalitoimisto).
På vissa arbetsplatser måste man kunna både finska och svenska.
I skolorna i Finland lär man sig både finska och svenska.
Elever som har finska som modersmål lär sig svenska i skolan.
Elever som har svenska som modersmål lär sig finska i skolan.
Om ett invandrarbarn går i en skola där undervisningsspråket är finska studerar barnet också svenska som främmande språk tillsammans med de finskspråkiga eleverna.
Hurdant är det finska språket?
Finskan är ett finsk-ugriskt språk.
Besläktade språk är till exempel estniska och ungerska.
Finskan har många böjningsformer, till exempel kasusformer av nomen, personformer av verb och tempusformer.
Finskan har färre prepositioner än till exempel de indoeuropeiska språken.
Finskan har också en del postpositioner.
Ordföljden är friare än i många andra språk.
Finskan har även många lånord från till exempel svenska, tyska, ryska och engelska.
Finskans uttal är mycket regelbundet.
Betoningen ligger alltid på den första stavelsen.
I Finland är det vanligt att dua.
Ibland kan det vara artigt att nia.
Till exempel kunder och äldre människor nias ofta.
Hurdant är det svenska språket?
Svenskan är ett indoeuropeiskt språk som tillhör de nordeuropeiska germanska språken.
Besläktade språk är till exempel norska, danska och tyska.
I svenskan finns också många lånord från till exempel franskan.
I svenskan böjs verben i olika tempus.
Substantiven kategoriseras i två genus.
Adjektiven böjs efter dessa genus.
I svenskan är det vanligt med prepositioner och ordföljden är mycket regelbunden.
Den svenska som talas i Finland kallas finlandssvenska.
Den uttalas lite annorlunda än den svenska som talas i Sverige.
Svenskans uttal är relativt regelbundet.
Inhemska minoritetsspråk
Förutom finska och svenska talas även andra inhemska språk i Finland.
De samiska språken tillhör urspråken i Finland.
I Finlands talas tre olika varieteter av samiska.
De är finsk-ugriska språk.
Finsk romani hör till de indoeuropeiska språken.
I Finland finns också ett eget teckenspråk.
Mer information om dessa språk får du på webbplatsen för Forskningscentralen för de inhemska språken.
Information om språklagenfinska _ svenska _ engelska
linkkiKommuner.net:
Svenskspråkiga och tvåspråkiga kommunerfinska _ svenska
linkkiInstitutet för de inhemska språken:
Information om finska språketfinska _ svenska
linkkiInstitutet för de inhemska språken:
Information om svenska språketfinska _ svenska
linkkiInstitutet för de inhemska språken:
Information om de samiska språkenfinska _ svenska
linkkiInstitutet för de inhemska språken:
Information om finska romanifinska
linkkiInstitutet för de inhemska språken:
Information om det finska teckenspråketfinska _ svenska
Ordbok i det finska teckenspråketfinska
En delägarbostad (osaomistusasunto) är ett bra sätt att skaffa en egen bostad om du inte kan köpa dig en egen bostad direkt.
Till en början köper du bara en del av bostaden och bor i bostaden på hyra.
Senare kan du köpa hela bostaden så att den blir helt och hållet din egen.
När du flyttar till en delägarbostad betalar du först ca 10-20 procent av bostadens pris.
Du kan ansöka om ett banklån för detta.
Efter detta bor du i bostaden på hyra och betalar hyra varje månad.
Vanligen är hyrestiden ca 5-12 år.
Du kan samtidigt köpa fler andelar i din bostad om du har kommit överens med byggherren om detta.
Efter hyrestiden köper du bostaden och den blir din egen.
Då har du en vanlig ägarbostad i ett bostadsaktiebolag.
Vissa delägarbostäder byggs med statligt stöd.
Då anger lagstiftningen till exempel hur lång hyrestiden i bostaden är och hur man kan avstå från bostaden.
Det finns även fritt finansierade delägarbostäder (vapaarahoitteinen osaomistusasunto).
Dessa är byggda utan statligt understöd.
Om du köper en fritt finansierad delägarbostad regleras inte hyrestiden eller andra avtalsvillkor i lagen.
Hur får man en delägarbostad?
Samfund och företag som låter bygga delägarbostäder informerar om nya och lediga bostäder.
Du får information om bostäderna även från kommunens bostadsbyrå.
Du kan ansöka om en delägarbostad med en ansökan riktad till bostadens byggherre.
Om delägarbostaden är byggd med statligt stöd kan du få en bostad om
dina inkomster inte är för stora; och
du inte har för stor förmögenhet.
Om du ansöker om en fritt finansierad bostad beaktas inte dina inkomster eller din förmögenhet.
linkkiKonkurrens- och konsumentverket:
Information om att bo i delägarbostadfinska _ svenska _ engelska
linkkiMiljöministeriet:
Information om att bo i delägarbostadfinska _ svenska _ engelska
I Finland bor många människor i hyresbostäder.
Det som är bra med en hyresbostad är att det är lätt att byta bostad, eftersom du inte behöver sälja och köpa bostaden.
Men å andra sidan kan hyresvärden bestämma sig för att säga upp hyresavtalet, om han eller hon har en godtagbar anledning.
Då måste du flytta från hyresbostaden, även om du inte vill det.
På InfoFinlands sida Hyresavtal finns viktig information om uppsägning av hyresbostad, betalning av hyran, hyresdeposition och andra utgifter i en hyresbostad.
I större städer är det ofta svårare att hitta en lämplig hyresbostad. Även hyran är högre.
Reservera tillräckligt med tid för att hitta en bostad.
En del områden är väldigt populära. I sådana områden hyrs bostäderna ut mycket snabbt.
När du har hittat en lämplig bostad bör du snabbt bestämma dig om du vill ha den.
Då hyrsvärden väljer hyresgäst får han eller hon enligt lagen inte diskriminera någon exempelvis på grund av etniskt ursprung, religion eller nationalitet.
Läs mer på InfoFinlands sida Diskriminering och rasism.
Hur skaffar jag en hyresbostad?
När du letar efter en hyresbostad kan du leta efter annonser till exempel på internet.
Skriv in sökordet ”hyresbostad”.
Du kan även titta i lokaltidningarna.
Sökning av hyresbostäderfinska _ engelska
Sökning av hyresbostäderfinska
Privata hyresbostäder
Man får oftast en privat hyresbostad snabbare än en kommunal hyresbostad. Hyran för en privat bostad är ofta högre.
Du behöver inte anlita en bostadsmäklare för att söka bostad.
Du kan själv söka information om lediga bostäder.
Då behöver du inte heller betala mäklararvode (välityspalkkio).
Du kan söka privata hyresbostäder på internet och i lokaltidningar.
Du kan även publicera en egen annons.
Om du vill hyra en privat hyresbostad ska du kontakta den som hyr ut bostaden.
Kom överens om när du kan gå och titta på bostaden. En bostadsvisning ordnas oftast för alla intresserade på samma gång.
Samtidigt får du en ansökningsblankett.
Fyll i den om du vill flytta in i bostaden.
Om du vill att en mäklare söker en lämplig hyresbostad åt dig, ska du ingå ett skriftligt uppdragsavtal (toimeksiantosopimus) med mäklaren.
Du måste då betala mäklararvode till mäklaren.
Avtala om arvodet skriftligen på förhand.
Arvodet kan till exempel vara lika stort som en månads hyra.
Jämför olika mäklarbyråers priser på förhand.
När du hyr en privat bostad ska du göra ett hyresavtal med hyresvärden.
Läs mera på InfoFinlands sida Hyresavtal.
Priser på icke subventionerade hyresbostäderengelska
Kommunernas hyresbostäder
Även kommunerna äger hyresbostäder. De är ofta förmånligare än andra hyresbostäder.
Du kan söka boende i en hyresbostad som staten stödjer, om du har något av följande:
Finskt medborgarskap;
registrerat uppehållstillstånd;
uppehållskort;
uppehållstillstånd som är giltigt i minst ett år; eller
uppehållstillstånd för studerande.
Om du vill ansöka om en kommunal hyresbostad fyller du i ansökningsblanketten på bostadskontoret i din kommun.
Ofta kan du även fylla i och skicka blanketten på kommunens webbsida.
I en del kommuner är hyresbostäderna så populära att man kan vara tvungen att stå i kö mycket länge.
Köerna till bostäderna kan vara långa till exempel i huvudstadsregionen (Helsingfors, Esbo och Vanda), men det finns lediga bostäder på mindre orter runt om i Finland.
När hyresgästerna väljs beaktas
inkomster
egendom
behovet av bostad.
I Finland finns även många allmännyttiga samfund som har förmånliga hyresbostäder.
Priser på hyresbostäder med statliga stödengelska
Studentbostäder
Om du är studerande kan du söka en hyresbostad som är avsedd särskild för studerande.
Läs mer på InfoFinlands sida Boende för studerande.
Bostadsansökan och bilagor
När du lämnar in en bostadsansökan kan du behöva också andra dokument som bilagor till ansökan.
Dessa beror på varifrån du söker bostaden.
senaste löneintyg
kopia på beskattningsbeslutet där din egendom framgår
intyg över lån
kopia på uppehållstillstånd eller pass om du inte är EU-medborgare.
Ofta granskas även den bostadssökandes kredituppgifter.
linkkiKonkurrens- och konsumentverket:
Att hyra en bostadfinska _ svenska _ engelska
Information för hyresgästenfinska _ svenska _ engelska
linkkiMiljöministeriet:
Information om hyresboendefinska _ svenska _ engelska
linkkiKonsumentförbundet ry:
Hyreshandboken(pdf, 1,11 MB)finska _ svenska _ ryska _ franska _ somaliska _ arabiska
Hyresbostadens utrustning
I utrustningen i en hyresbostad ingår nästan alltid köksskåpen, kylskåpet och spisen.
Även klädskåp och skåp i hallen ingår vanligtvis.
Duschen, vattenkranarna och toalettstolen hör alltid till utrustningen.
Hyresbostäder är vanligtvis inte möblerade.
Det händer dock att lägenheter hyrs ut med möbler.
Vilka möbler som ingår varierar.
Kontrollera alltid med hyresvärden vilka möbler som ingår.
Hushållsavfall
I Finland ska hushållsavfall sorteras i olika sopkärl.
Läs mer på InfoFinlands sida Avfallshantering och återvinning.
Rådgivningstjänster
Vill du söka råd om att hyra en bostad?
Finlands Konsumentförbund erbjuder råd och handledning både för hyresgäster och hyresvärder.
Finlands Konsumentförbunds rådgivningstjänst:
tfn 010 8022 40
tis-fre kl. 10–12 och tis kl. 17–19
Du kan ringa till tjänsten och endast betala lokalsamtalsavgift överallt i Finland.
Du kan fråga råd på tjänsten även på nätet genom att fylla i en blankett. Du får svar per e-post.
Även Marthaförbundet och Finlands flyktinghjälp erbjuder bostadsrådgivning åt invandrare.
linkkiKonsumentförbundet:
Boenderådgivningfinska
linkkiFlyktinghjälp:
Flyktinghjälpens regionkontorfinska
linkkiMarthaförbundet:
Kontaktuppgifter till Marthaförbundetfinska _ engelska
Tvåspråkiga kommuner i Finland
Finland har två officiella språk, finska och svenska.
Finska är modersmålet för cirka 90 procent av finländarna.
Svenska är modersmålet för cirka 5 procent av finländarna.
Svenska talas mest på Finlands väst- och sydkust.
Svenskan som talas i Finland är finlandssvenska.
Uttalet skiljer sig något från svenskan i Sverige.
Om du vill ansöka om finskt medborgarskap behöver du ett intyg över tillräckliga kunskaper i finska eller svenska.
Läs mer på InfoFinlands sida Officiellt intyg över språkkunskaper.
Du kan använda svenska med statliga myndigheter, till exempel FPA eller TE-byrån.
Ange ditt kontaktspråk till magistraten när du registrerar dig som invånare.
Du kan även ändra kontaktspråket senare.
Kommunerna i Finland kan vara antingen enspråkiga eller tvåspråkiga.
De flesta kommunerna i Finland är finskspråkiga.
Tvåspråkiga kommuner finns på väst- och sydkusten.
Om din hemkommun är tvåspråkig, kan du använda svenska även inom de kommunala tjänsterna, till exempel på hälsostationen.
linkkiKommuner.net:
Svenskspråkiga och tvåspråkiga kommunerfinska _ svenska
Integration på svenska kan vara ett bra alternativ för dig till exempel om:
Du bor i ett område med många svensktalande.
Du har svenskspråkiga familjemedlemmar eller släktingar.
Du kan lite svenska redan.
Det kan vara fördelaktigt att kunna svenska när du söker jobb.
Tänk ändå på att kunskaper i finska krävs på de flesta arbetsplatserna.
Även om du väljer integrationsutbildning på svenska lönar det sig för dig att i något skede även lära dig finska.
I en del kommuner kan du delta i integrationsutbildning på svenska.
Om du inte blir antagen till integrationsutbildning på svenska kan du i vissa fall få stöd för frivilliga studier i svenska, om detta överenskommits i din integrations- eller sysselsättningsplan.
Fråga om integration på svenska när din inledande kartläggning och integrationsplan görs.
Enligt lag har du rätt att välja antingen finska eller svenska som integrationsspråk.
linkkiArbets- och näringsministeriet:
Information om integration på svenskafinska _ svenska
Språkstudier som arbetskraftsutbildning
Om du är kund vid arbets- och näringsbyrån kan du också studera svenska som arbetskraftsutbildning.
Arbetskraftsutbildningen är avsedd för arbetslösa arbetssökande.
Läs på InfoFinlands sida Arbets- och näringsbyråns tjänster vad som krävs för att du ska kunna bli kund hos arbets- och näringsbyrån.
Arbetskraftsutbildningen är kostnadsfri för dig.
Fråga mer om kurser i svenska vid din egen arbets- och näringsbyrå.
Barndagvård och utbildning för barn
I Finland ges dagvård, förskoleundervisning och grundläggande utbildning vanligtvis på finska eller svenska.
Om du vill att ditt barn ska börja i svenskspråkig dagvård, förskola eller skola, fråga om möjligheterna i din hemkommun.
Vissa kommuner ordnar förberedande undervisning före den grundläggande utbildningen för elever som ännu inte har tillräckligt bra språkkunskaper för den vanliga undervisningen.
Fråga i din hemkommun om förberedande undervisning ordnas på svenska i kommunen.
Om barnet har något annat modersmål än finska eller svenska, kan kommunen ordna undervisning i barnets eget modersmål för barnet.
Om barnet går i en svensk skola kan hen läsa svenska som andra språk.
Läs mer om barndagvård, förskoleundervisning och grundläggande utbildning på InfoFinlands sida Det finländska utbildningssystemet.
Gymnasium och yrkesläroanstalt
Efter grundskolan kan du studera på gymnasiet eller en yrkesläroanstalt.
Svenskspråkiga yrkesläroanstalter och gymnasieskolor finns i svenskspråkiga och tvåspråkiga kommuner och i en del finskspråkiga kommuner.
Vissa yrkesläroanstalter och gymnasieskolor ordnar förberedande utbildning före studierna.
I den förberedande utbildningen får du sådana kunskaper och färdigheter som du behöver i dina fortsatta studier.
Du kan också förbättra dina språkkunskaper.
Du kan söka svenskspråkig yrkes- och gymnasieutbildning samt förberedande utbildning före dessa via tjänsten Opintopolku.fi.
Läs mer på InfoFinlands sida: Efter grundskolan.
Grundläggande information om yrkesutbildningfinska _ svenska _ engelska
Information om gymnasiestudierfinska _ svenska
Högskoleutbildning
I Finland finns svenskspråkiga yrkeshögskolor och universitet.
Dessutom finns det några tvåspråkiga universitet där du kan läsa på svenska.
Du kan söka svenskspråkiga högskoleutbildningar via tjänsten Opintopolku.fi.
Information om högskolestudierfinska _ svenska _ engelska
Var kan jag läsa svenska?
Du kan läsa svenska till exempel vid medborgarinstitut, arbetarinstitut och sommaruniversitet.
Fråga om studier i svenska hos utbildningsväsendet i din hemkommun, studievägledarna vid läroanstalter eller rådgivningstjänsterna för invandrare.
Läs mer på InfoFinlands sida: Studier som hobby.
Svenska på internet
Appar
Du kan lära dig svenska med hjälp av appar som du kan ladda ned i din telefon eller surfplatta.
Sök appar för svenska i din appbutik (t.ex. Google Play och App Store) med sökorden ”learn Swedish”, ”Swedish language”, ”lär dig svenska” eller ”svenska”.
En del appar kostar pengar.
Övningar och kurser på internet
På internet hittar du kurser i det svenska språket på olika nivåer.
På internet kan du till exempel göra övningar och spela spel, lära dig grammatik och vokabulär samt läsa texter.
linkkiYle:
Övningar för allmänna språkexaminafinska
Svenska på internetfinska _ svenska _ engelska
linkkiYle.fi:
Övningar och kurser på internetfinska
linkkiBab.la:
Flerspråkiga ordböckerfinska _ svenska _ engelska
Du får bo i en bostadsrättsbostad om du först betalar bostadsrättsavgiften (asumisoikeusmaksu).
Avgiften är ca 15 procent av bostadens pris.
Om du inte har pengar till bostadsrättsavgiften kan du ansöka om lån från banken.
Du kan dra av låneräntan i beskattningen.
Därefter betalar du varje månad en bestämd summa det vill säga bruksvederlag (käyttövastike).
Bruksvederlagets storlek beror på bostaden och orten.
Bruksvederlaget får inte vara större än hyran för bostäder av samma typ på samma område.
Om dina inkomster är små kan du ansöka om bostadsbidrag för bruksvederlaget.
Läs mera på InfoFinlands sida Bostadsbidrag.
Man kan inte köpa en bostadsrättsbostad.
Varför bostadsrättsbostad?
Bostadsrättsbostäder är inte förknippade med ekonomiska risker.
Därför är det en tryggare boendeform än en ägarbostad.
Du behöver inget stort lån för en bostadsrättsbostad.
När du vill flytta behöver du inte sälja bostaden.
Du kan bo i bostadsrättsbostaden så länge du vill.
Husets ägare kan inte säga upp bostadsrättskontraktet.
En bostadsrättsbostad är alltså mer bestående än en hyresbostad.
Du kan också låta bostadsrätten gå i arv.
Den boendes skyldigheter
Om du har en bostadsrättsbostad måste du själv vara fast bosatt i den.
Du kan hyra ut bostaden till någon annan under högst två år.
Du behöver dock tillstånd till detta av husets ägare.
Vem kan få en bostadsrättsbostad?
Om bostadsrättsbostaden inte har byggts med statsstöd kan husets ägare välja boende själv.
Om bostaden är byggd med statsstöd, kan du ansöka om
du har fyllt 18 år;
du inte har en ägarbostad på samma område; och
du inte har råd att skaffa en ägarbostad på samma område.
Din egendom beaktas ändå inte om du är över 55 år gammal eller flyttar från en bostadsrättsbostad till en annan bostadsrättsbostad.
Ibland kan det utöver dessa förekomma övriga villkor.
Hur ansöker man om en bostadsrättsbostad?
Det finns bostadsrättsbostäder i de största kommunerna.
Om du vill ha en bostadsrättsbostad, hämta först ett könummer på kommunens bostadsbyrå.
Du kan skaffa könummer i flera olika kommuner.
Könumret kostar ingenting.
Även om du har ett nummer behöver du inte ansöka om en bostad.
Välj sedan det hus där du vill ha en bostadsrättsbostad.
Anmäl dig till husets ägare.
Berätta också hurdan bostad du letar efter.
Du kan ansöka om bostadsrättsbostad i många olika hus.
Du kan bli tvungen att vänta länge på en bostad.
Bostadsrättsavtal
Då du får en bostad ska du göra ett skriftligt bostadsrättsavtal (asumisoikeussopimus) med husets ägare.
I bostadsrättsavtalet fastställs storleken på bostadsrättsavgiften, bruksvederlaget och övriga eventuella villkor.
Du kan flytta in i bostadsrättsbostaden när du har gjort bostadsrättskontraktet och betalat bostadsrättsavgiften.
När du flyttar ut
Om du vill flytta ut ur bostaden måste du göra en avträdelseanmälan (luopumisilmoitus) till husets ägare.
Du får bostadsrättsavgiften tillbaka, när du har avträtt bostaden.
linkkiKonkurrens- och konsumentverket:
Information om att bo i bostadsrättsbostadfinska _ svenska _ engelska
linkkiMiljöministeriet:
Att ansöka om en bostadsrättsbostadfinska _ svenska _ engelska
linkkiMiljöministeriet:
Information om att bo i bostadsrättsbostadfinska _ svenska _ engelska
Oy:
Bostadsrättsbostäderfinska
Bostadsrättsbostäderfinska
Bostadsrättsbostäderfinska
Bostadsrättsbostäderfinska
Checklista för dig som flyttar
När du flyttar i Finland från en bostad till en annan:
Kom ihåg att göra flyttanmälan (muuttoilmoitus).
Du kan göra flyttanmälan högst en månad före flyttningsdagen, men den bör göras senast en vecka efter att du har flyttat.
Flyttanmälan ska alltid göras till magistraten (maistraatti).
Du kan göra flyttanmälan
på nätet
telefonledes på finska på numret 0295 535 535 eller på svenska på numret 0295 535 536 eller
på en blankett som du får på posten eller hos magistraten.
Om du bor i höghus eller radhus ska du alltid också komma ihåg att meddela husets disponent (isännöitsijä) att du flyttar.
Meddela din nya adress till alla instanser som skickar dig post.
Vissa organisationer och företag får din nya adress direkt från befolkningsregistret.
Du har ändå själv ansvaret för att dina fakturor skickas till rätt adress och betalas i tid.
Om du bor i en hyresbostad ska du komma ihåg att säga upp din gamla bostad i tid.
Det är bäst att göra uppsägningen skriftligt.
Kontrollera hur lång uppsägningstid du har för bostaden.
Vanligen är den en kalendermånad.
Läs mer på InfoFinlands sida Hyresavtal.
Om du har barn ska du se till att skaffa dem nya dagvårds- och skolplatser.
Du måste meddela daghemmet och skolan när barnen slutar där.
Samtidigt är det bra att anmäla barnen till det nya daghemmet eller den nya skolan.
Kom ihåg att skaffa eventuell flytthjälp i tid.
Bland annat vid månadsskift och på veckoslut är flyttfirmorna alltid upptagna.
Avtala med din tjänsteleverantör om överföringen av din internetanslutning i god tid så att det inte blir ett avbrott i servicen.
Säg upp ditt gamla elavtal innan du flyttar och gör upp ett nytt.
Det lönar sig att jämföra olika elbolags priser så att du hittar det förmånligaste.
Du får ett elavtal genom att ringa upp elbolaget och meddela ditt namn och din nya adress.
Om du flyttar till ett egnahemshus ska du också komma ihåg att teckna andra avtal, såsom avtal om vattenförsörjning och avfallshantering.
Om huset värms upp med olja ska du komma ihåg att kontrollera oljemängden.
Kontrollera om dina nuvarande försäkringar, som hemförsäkringen, är tillräckliga även för den nya bostaden.
Om du till exempel flyttar från höghus till egnahemshus behöver du förmodligen en annorlunda försäkring.
Städa den gamla bostaden innan du flyttar och töm vinden, källarförrådet och garaget på saker.
Om du bor i en hyresbostad ska du ge ägaren eller disponenten alla nycklar till den gamla bostaden.
linkkiFörbundet för ungdomsbostäder:
Ordlista om boendefinska
Flyttanmälanfinska _ svenska _ engelska
linkkiEnergimarknadsverket:
Jämför elpriserfinska
Flyttjänsterfinska _ engelska
Flyttjänsterfinska _ engelska _ ryska
Flyttjänsterfinska _ svenska _ engelska
När du flyttar till Finland
Om du vill ha information om praktiska frågor i anslutning till att du flyttar till Finland, läs mer på sidan Komihåglista för dig som flyttar till Finland.
Om du nyligen har flyttat till Finland, måste du registrera dig som invånare.
Lär mer på InfoFinlands sida Registrering som invånare.
Flytta från Finland
Planerar du att flytta från Finland till ett annat land?
Läs mer på InfoFinlands sida Flytta från Finland.
Om du vill ansöka om finskt medborgarskap behöver du ett officiellt intyg över dina kunskaper i finska eller svenska.
Du kan behöva intyget också när du söker ett jobb eller en studieplats.
Du kan påvisa dina språkkunskaper:
med en allmän språkexamen (yleinen kielitutkinto)
med vitsordet i finska eller svenska på ditt avgångsbetyg (päättötodistus).
Allmän språkexamen
Allmän språkexamen, ASE, är ett språktest för vuxna.
Med en allmän språkexamen kan du påvisa dina kunskaper i finska eller svenska.
Examen är avgiftsbelagd.
När du avlagt examen får du ett intyg som anger nivån på dina språkkunskaper.
Språkexamen finns på tre olika nivåer: grundnivån, mellannivån och högsta nivån.
Varje examensnivå består av två färdighetsnivåer, vilka det alltså finns sammanlagt sex av.
Grundnivån är avsedd för personer som kan använda språket i vardagliga sammanhang.
Deras färdighetsnivå är 1–2.
Medelnivån är avsedd för personer som kan språket relativt väl. Deras färdighetsnivå är 3–4.
Den högsta nivån är avsedd för personer som kan språket mycket väl. Deras färdighetsnivå är 5–6.
Närmare beskrivningar av de olika färdighetsnivåerna finns på Utbildningsstyrelsens webbplats.
Om du vill ansöka om finskt medborgarskap (kansalaisuus) kan du påvisa att du har tillräckliga kunskaper i finska eller svenska genom att avlägga den muntliga och skriftliga delen av en allmän språkexamen minst på nivå 3.
Språkexamenstillfället pågår 3–6 timmar.
Uppgifternas ämnesområden rör det vardagliga livet såsom fritid, utbildning och vanliga situationer på arbetet.
I examen ingår olika uppgifter där följande färdigheter krävs:
textförståelse
skriftliga färdigheter
grammatik och vokabulär
talförståelse
Du kan avlägga examen på olika orter i Finland.
Mer information om anmälan får du på Utbildningsstyrelsens (Opetushallitus) webbplats.
Examina kategoriseras på en annan skala än kurserna.
Om du har slutfört en språkkurs som kategoriserats enligt den europeiska referensramen motsvarar kursen nivån på den allmänna språkexamen ungefär enligt följande tabell:
A1 – ASE 1
A2 – ASE 2
B1 – ASE 3
B2 – ASE 4
C1 – ASE 5
C2 – ASE 6
Innan du anmäler dig till examen ska du göra dig förtrogen med kraven på de olika examensnivåerna.
Du kan även fråga din lärare i finska.
Mer information om den allmänna språkexamen får du på Utbildningsstyrelsens webbplats.
linkkiUtbildningsstyrelsen:
Allmänna språkexaminafinska _ svenska _ engelska
linkkiUtbildningsstyrelsen:
Färdighetsnivåerna i allmänna språkexamina(pdf, 100 KB)finska _ svenska _ engelska
linkkiUtbildningsstyrelsen:
Att anmäla sig till en allmän språkexamen och examensavgifterfinska _ svenska _ engelska
Statsförvaltningens språkexamen om kunskaper i finska och svenska
Om du vill arbeta inom den offentliga förvaltningen behöver du vanligtvis ett intyg över dina kunskaper i finska eller svenska.
Du kan påvisa dina kunskaper i finska eller svenska med statsförvaltningens språkexamen.
Fråga din arbetsgivare hurdana språkkunskapskrav som gäller på den arbetsplats som du vill söka.
Språkexamen finns på tre olika nivåer: för nöjaktiga, goda och utmärkta språkkunskaper.
Det beror på din arbets- eller studieplats vilken examensnivå du måste avlägga.
För finskt medborgarskap behöver du ett intyg för åtminstone nöjaktiga språkkunskaper.
Du kan avlägga examen för nöjaktiga eller goda språkkunskaper olika orter i Finland.
På Utbildningsstyrelsens webbplats hittar du en förteckning över de städer där examen kan avläggas.
Examen på utmärkt nivå kan endast avläggas i Helsingfors.
Examen omfattar olika tester. I dem ska du läsa och lyssna på texter och svara på frågor.
Därtill finns det intervjuer, diskussioner och skriftliga uppgifter.
Du kan ersätta statsförvaltningens språkexamen med vissa andra studier.
Till exempel motsvarar statsförvaltningens språkexamen som gäller goda språkkunskaper ett mognadsprov (kypsyysnäyte) som du har avlagt på finska eller svenska vid universitetet.
Mer information får du på Utbildningsstyrelsens webbplats.
linkkiUtbildningsstyrelsen:
Statsförvaltningens språkexaminafinska _ svenska
linkkiUtbildningsstyrelsen:
Mottagare av statsförvaltningens språkexamina, finska språketfinska _ svenska
linkkiUtbildningsstyrelsen:
Mottagare av statsförvaltningens språkexamina, svenska språketfinska _ svenska
Intyg över språkkunskaper på basis av studier
Om du vill ansöka om finskt medborgarskap kan du påvisa dina kunskaper i finska eller svenska även med något av följande intyg:
avgångsbetyg från grundskolan med ett godkänt vitsord i finska eller svenska som modersmål eller som andra språk
avgångsbetyg från gymnasiet med ett godkänt vitsord i finska eller svenska som modersmål eller som andra språk
studentexamen på finska eller svenska med ett godkänt vitsord i finska eller svenska som modersmål eller som andra språk
intyg på yrkesinriktad grundexamen som du har avlagt på finska eller svenska
intyg på yrkesexamen som du har avlagt på finska eller svenska
intyg på studier i tjänstemannafinska eller -svenska som du har avlagt vid universitet eller högskola
intyg på mognadsprov som du har avlagt på finska eller svenska för universitetsexamen eller yrkeshögskoleexamen
Mer information får du på Migrationsverkets (Maahanmuuttovirasto) webbplats.
linkkiUtbildningsstyrelsen:
Språkkunskaper och finskt medborgarskapfinska _ svenska _ engelska
En ägarbostad är ofta på lång sikt förmånligare än en hyresbostad.
Största delen av finländarna bor ägarbostäder.
Det finns också andra alternativ än ägarbostad och hyresbostad.
Läs mer på InfoFinlands sidor Bostadsrättsbostad och Delägarbostad.
Bostadsaktie och fastighet
Då du köper en bostad, köper du antingen en bostadsaktie (asunto-osake) eller en fastighet (kiinteistö).
Höghuslägenheter och radhuslägenheter är bostadsaktier.
De finns i hus som ägs av ett bostadsaktiebolag.
Då du köper ett egnahemshus köper du en fastighet.
Fastigheten utgörs vanligen av egnahemshuset och dess tomt.
Hur hittar jag en ägarbostad?
När du letar efter en bostad är det bra att räkna med att det tar till och med flera månader.
Bostäder säljs av privatpersoner, fastighetsförmedlingar och byggherrar.
Bland annat på internet och i dagstidningar finns det annonser för bostäder som är till salu.
När du hittar en bostad som intresserar dig kan du komma överens med försäljaren om en visning av bostaden.
Ibland finns det i annonsen en utsatt tid då bostaden visas.
I så fall behöver du inte avtala en tid.
linkkiEtuovi.com:
Sökning av ägarbostäderfinska _ engelska
Sökning av ägarbostäderfinska
linkkiKonkurrens- och konsumentverket:
Information om att köpa en bostadfinska _ svenska _ engelska
Utred bostadens skick och andra frågor
Ta reda på allt som berör bostaden när du har hittat en bostad du tycker om.
Särskilt lönar det sig att utreda bostadens skick grundligt.
Om du tänker köpa en bostadsaktie, ta då även reda på vilka renoveringar bostadsaktiebolaget planerar och vad de kostar.
Till exempel ett stambyte kan kosta bostadsägaren många tiotusentals euro.
Säljarens och köparens ansvar vid bostadsköp
Den som säljer bostaden är ansvarig för fel i bostaden ännu under någon tid efter att bostaden har sålts.
Den som säljer en bostadsaktie är vanligen ansvarig för fel under två år.
För den som säljer en fastighet varar ansvaret fem år.
Enligt lagen måste den som säljer bostaden berätta om de fel som han/hon känner till innan försäljningen av bostaden.
Om det står klart att försäljaren har känt till fel i bostaden utan att berätta om detta för köparen, kan säljaren tvingas ersätta köparen för felet.
Granska om det finns fel i bostaden innan du köper en bostad.
Du kan inte efteråt kräva ersättning för fel, om
felet kan upptäckas vid granskning av bostaden; eller
du har känt till det innan köpet.
Det kan också finnas dolda fel i bostaden.
De är fel som ingen känner till.
Dolda fel är ofta till exempel fuktproblem.
Säljaren måste betala ut en ersättning till köparen ifall det i bostaden finns ett allvarligt fel, som skulle ha påverkat bostadsköpet ifall man känt till det.
Bostadslån
Vanligen betalar man bostaden med ett bostadslån (asuntolaina).
Vem som helst kan ansöka om ett bostadslån hos banken.
För att du ska kunna få ett bostadslån måste du ha tillräckliga inkomster för att betala tillbaka lånet utan problem.
På bankernas webbsidor finns det låneräknare.
Med hjälp av dem kan du på förhand uppskatta om du kan betala tillbaka lånet.
Om du inte är säker på huruvida banken ger dig ett lån lönar det sig att gå till banken och förhandla om lånet i god tid innan du köper bostaden.
Lånet återbetalas det vill säga amorteras en gång i månaden.
Dessutom måste man betala ränta (korko) för lånet till banken.
Du kan be om låneerbjudanden från flera banker och jämföra dem.
Olika lån har olika villkor.
Då du funderar på vilket lån du ska välja bör du beakta
hur stor ränta lånet har
hur stor summa du betalar tillbaka per månad
hur många år du återbetalar lånet
Märk väl att om räntorna stiger så stiger även lånekostnaderna.
Då stiger den månatliga avgiften eller också förlängs lånetiden.
Du kan dra av en del av räntan på bostadslånet i beskattningen.
linkkiKonkurrens- och konsumentverket:
Information om bostadslånfinska _ svenska _ engelska
Säkerhet och borgen för bostadslån
För ett bostadslån behövs det vanligen en säkerhet (vakuus).
Bostaden som du köper täcker en del av säkerheten, vanligen ca 70 procent.
Utöver detta behöver du en säkerhet för resten av lånesumman.
Du kan ordna säkerheten till exempel så att
Statsborgen kan utgöra högst 20 procent av lånet och högst 50 000 euro.
du ber en släktning eller vän gå i borgen för ditt lån.
Om du inte själv kan betala tillbaka lånet, blir borgensmannen tvungen att betala den summan som han eller hon gått i borgen för.
Du behöver ändå inte borgensmän för ditt lån om du har sparat ihop en del av bostadens pris på förhand, eller om du har annan egendom som duger som säkerhet för lånet.
linkkiMiljöministeriet:
Information om statsborgen för bostadslånfinska _ svenska _ engelska
Stöd vid bostadsköp
Staten beviljar räntestöd (korkotuki) för bostadslån.
Räntestöd beviljas för unga som skaffar sin första ägarbostad.
Det beviljas även för dem som köper eller bygger ett egnahemshus.
Läs mera på miljöministeriets sidor.
linkkiMiljöministeriet:
Information om räntestödetfinska _ svenska _ engelska
Överlåtelseskatt
När du köper en bostad måste du också betala överlåtelseskatt (varainsiirtovero).
Om du köper en bostadsaktie är överlåtelseskatten 2 procent av bostadens skuldfria pris.
Om du köper en fastighet är skatten 4 procent av bostadens skuldfria pris.
Du behöver ändå inte betala överlåtelseskatt om alla följande villkor uppfylls:
du är 18–39 år gammal
du har inte tidigare ägt en bostad i Finland eller något annat land
du äger minst 50 % av bostaden
du är själv fast bosatt i bostaden
linkkiSkatteförvaltningen:
Befrielse från överlåtelseskatt på första bostadfinska _ svenska _ engelska
Köpeanbud
När du är säker på att du vill och kan köpa en bostad kan du göra ett köpeanbud på bostaden.
Det lönar sig att göra ett skriftligt anbud.
Anbudet kan vara t.ex. 5-10 procent lägre än priset som säljaren har bett om för bostaden.
Säljaren kanske ändå inte vill sälja bostaden billigare.
Köpeanbudet är bindande.
Det betyder att du inte kan ta tillbaka anbudet.
Om du tar tillbaka köpeanbudet kan du bli tvungen att betala säljaren böter eller en handpenning.
Denna summa är vanligen några procent av bostadens pris.
Information om priser på sålda bostäderfinska _ svenska
Bostadsköp
Om säljaren av bostaden godtar köpeanbudet görs bostadsköpet upp i köparens bank.
Vanligen närvarar köparen och säljaren av bostaden samt bostadsförmedlaren, om en förmedlare har använts.
Köpebrevet är ett kontrakt där t.ex. bostadens pris, bostadens storlek, bostadens skick och datumet då köparen får tillgång till bostaden finns inskrivet.
Vanligen görs köpebrevet upp av banken eller bostadsförmedlaren.
Köparen har rätt att läsa köpebrevet före dagen då köpet genomförs.
Banken lånar bolånepengarna åt köparen, och summan flyttas över på säljarens konto.
Handpenning
Handpenningen (käsiraha) är en avgift, som betalas för bostaden på förhand.
Köparen kan betala handpenningen åt säljaren i det skedet då köpet förbereds.
Handpenningen är vanligen ca tre procent av bostadens pris.
Om du inte kan betala handpenningen av dina egna besparingar kan du låna summan av banken som en del av bostadslånet.
Kostnader för ägarbostad
På boendekostnaderna inverkar
bostadslånets storlek
bostadens storlek
bostadens skick
bostadens läge.
Bostadsaktie
Om du äger en bostadsaktie betalar du vanligen
ränta och amorteringar på bostadslånet
finansieringsvederlag (rahoitusvastike), om bostadsaktiebolaget har skulder
el och vatten
eventuella reparationsarbeten
Fastighet
Om du äger en fastighet betalar du vanligen
ränta och amorteringar på bostadslånet
fastighetsskatt (kiinteistövero)
el och vatten
värme
sophämtning
eventuella reparationsarbeten
Hushållsavfall
I Finland ska hushållsavfall sorteras i olika sopkärl.
Läs mer på InfoFinlands sida Avfallshantering och återvinning.
God morgon!
God dag!
God kväll!
God natt!
Välkommen!
Tack.
Var så god.
Förlåt.
Jag älskar dig.
Hur står det till?
Hejdå.
Adjö.
Jag förstår inte, kan du upprepa?
Jag talar inte finska.
Jag talar bara lite finska.
Talar du engelska/svenska?
Jag är lärare / ingenjör / studerande.
Vad är ditt telefonnummer / din e-postadress?
Var finns det en affär / ett apotek / en skola / ett daghem / en busstation / en metrostation?
På nätet hittar du finskakurser på många olika nivåer.
På nätet kan du till exempel göra övningar, spela spel, lära dig grammatik och vokabulär och läsa texter.
De flesta webbkurser är på finska eller svenska, men det finns även andra alternativ:
Nybörjarnivån
linkkiYle:
Nybörjarkurs i finska, Easyfinnishfinska
Nybörjarkurs i finska "A Taste of Finnish"engelska
linkkiTammerfors yrkeshögskola:
Nybörjarkurs i finska, Uunofinska
Nybörjarkurs i finska, Tavataan taasengelska _ franska _ tyska _ bulgariska
Nybörjarkurs i finskafinska _ svenska _ engelska _ arabiska
linkkiWordDive:
Nybörjarkurs i finskafinska _ svenska _ engelska _ ryska _ kinesiska _ tyska
Inledningskurs i finskaengelska
Tilläggsövningar till läroboken Hyvin meneefinska
Mångsidiga övningar i finska språketfinska
Ordspel för nybörjareengelska _ franska _ japanska
Applikationen Suomipassi med flera stödspråkfinska _ engelska
Grundnivån
linkkiYle:
Övningar för allmänna språkexaminafinska
Webbkurs med många hjälpspråksvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ portugisiska
Vokabulärövningarfinska
linkkiYle:
Läromaterial från TV-serien Supisuomeafinska
linkkiUtbildningsstyrelsen:
Finska i arbetslivetfinska
Mångsidiga övningar i finska språketfinska
Lär dig finska med hjälp av filmerfinska _ engelska _ persiska _ arabiska
Självständiga språkanvändare
linkkiYle:
Nyheter på klarspråkfinska
Information om olika ämnen på klarspråkfinska
Nyheter på lättläst finskafinska
linkkiUtbildningsstyrelsen:
linkkiUtbildningsstyrelsen:
Finska i arbetslivetfinska
Avancerade språkanvändare
Lyssna på finska dialekterfinska
linkkiWordDive:
Finskans grammatikfinska _ svenska _ engelska _ ryska _ spanska _ tyska _ japanska
Finskans grammatikengelska
Finskans grammatikengelska
Verbböjningengelska
linkkiInstitutet för de inhemska språken:
Grammatiken Iso suomen kielioppi på nätetfinska
Information om finska språketengelska
Ordböcker på nätet
Flerspråkiga ordböckerfinska
linkkiBab.la:
Flerspråkiga ordböckerfinska _ svenska _ engelska
Ett hyresavtal kan vara
ett hyresavtal som gäller tillsvidare eller
ett tidsbestämt hyresavtal.
Ett hyresavtal som gäller tillsvidare (Toistaiseksi voimassa oleva vuokrasopimus) fortsätter fram till dess att hyresgästen eller hyresvärden säger upp avtalet.
Om du på förhand inte vet hur länge du kommer att bo i bostaden, är ett sådant avtal ett bra alternativ.
Ett tidsbestämt avtal (Määräaikainen vuokrasopimus) innebär att hyresvärden och hyresgästen från början kommer överens om när avtalet upphör.
Ett tidsbestämt hyresavtal upphör automatiskt utan uppsägning på den dag som antecknats i avtalet.
Om du fortfarande vill bo i bostaden efter detta behöver du ett nytt hyresavtal.
Det är inte möjligt att säga upp ett tidsbestämt avtal under dess giltighetstid.
Detta gäller för såväl hyresgästen som för hyresvärden.
Om du på förhand vet att du behöver bostaden enbart för en viss tid, är ett tidsbestämt hyresavtal ett bra alternativ.
Betalning av hyra
Hyra betalas vanligen en gång per månad.
Hyran ska betalas senast på förfallodatumet.
Förfallodagen har antecknats i hyresavtalet.
Betala hyran som en girering till hyresvärdens konto.
Du kan inte betala hyran med ett kreditkort.
Hyresgaranti
När du ingår ett hyresavtal i Finland, ska du nästan alltid betala en hyresgaranti.
Detta innebär att du på förhand betalar ett penningbelopp som motsvarar några månaders hyra till hyresvärden.
Vanligen motsvarar garantin beloppet på två månaders hyra.
Den kan högst uppgå till beloppet på tre månaders hyra.
Betala hyresgarantin senast på det datum som överenskommits i hyresavtalet.
I allmänhet får du nycklarna till bostaden när du betalat hyresgarantin.
När hyresavtalet upphör utförs en slutsyn i bostaden.
Hyresgarantin betalas tillbaka till dig i sin helhet om du
skött bostaden omsorgsfullt och
betalat alla avgifter som överenskommits med hyresvärden.
Om du söndrat bostaden eller inte betalat hela hyran, får du inte tillbaka hyresgarantin i sin helhet.
Hyresgarantin kan inte användas för att betala hyran för de sista månaderna.
Övriga avgifter
Reservera pengar för andra avgifter än hyran.
Vatten
Ofta ska du betala en vattenavgift för bostaden.
Betala vattenavgiften till hyresvärdens eller husbolagets konto på samma gång som du betalar hyra.
Beloppet på vattenavgiften beror ofta på det antal personer som bor i bostaden.
Om det finns en vattenmätare i bostaden, fastställs vattenavgiften enligt vattenkonsumtionen.
El
Ofta ska du själv ingå ett elavtal.
Du ingår ett elavtal genom att ringa ett elbolag och uppge ditt namn och din nya adress.
Om du vill hitta det förmånligaste priset, kan du jämföra olika elbolags priser.
Uppvärmning
Om bostaden har centralvärme, ingår uppvärmningen i allmänhet i hyran.
Om bostaden har oljevärme eller elvärme, ska avgiften ibland betalas separat.
Bastu, tvättstuga och bilplats
Det kostar i allmänhet att använda husbolagets bastu, tvättstuga och bilplatser.
I allmänhet ska dessa avgifter betalas direkt till husbolaget.
Avgifter i egnahemshus
Om du bor på hyra i ett egnahemshus, ska du ofta betala för uppvärmningen och avfallshanteringen.
Uppsägning av hyresavtal
Med uppsägningstid avses den tid som avtalet är i kraft efter att det sagts upp.
Uppsägningstiden gäller hyresavtal som gäller tillsvidare.
Uppsägningstiden för hyresgäster är en kalendermånad.
Du bör beakta hur uppsägningstiden räknas.
Uppsägningstiden börjar i allmänhet först från slutet av den månad då avtalet sägs upp.
Om du vill flytta ut från bostaden t.ex. 1.12, lönar det sig att säga upp bostaden senast 31.10.
Annars måste du betala hyra också för december månad.
Ge alltid ett skriftligt uppsägningsmeddelande.
Du måste kunna bevisa att du gett hyresvärden ett meddelande.
Hyresvärdens uppsägningstid beror på hur länge hyresavtalet varit i kraft.
Om avtalet varit i kraft i kortare tid än ett år, är uppsägningstiden tre månader.
Om avtalet varit i kraft i över ett år, är uppsägningstiden sex månader.
Ett tidsbestämt hyresavtal kan inte sägas upp mitt i avtalsperioden.
Underuthyrning
Med underuthyrning avses att hyresgästen hyr ut en del av bostaden till en annan person.
Hyresgästen har rätt att göra detta, om bostadens egentliga hyresvärd godkänner detta.
Innan du flyttar in som underhyresgäst ska du säkerställa att hyresgästen har rätt att ta en underhyresgäst.
Du är underhyresgäst också när du hyrt endast en del av en bostad och bostadsägaren själv bor i samma bostad.
Uppsägningstiden för en underhyresgäst är kortare än för en hyresgäst.
Uthyrning i andra hand
Med uthyrning i andra hand avses att hyresgästen hyr ut hela bostaden till en annan person.
Ett tillstånd av hyresvärden behövs alltid för detta.
Uppsägningsvillkoren är de samma som för hyresgäster.
Mallar för hyresavtalfinska
Guiden God hyressed(pdf, 546 kB)finska _ svenska _ engelska
Finland är ett tvåspråkigt land
Finland har två officiella språk, finska och svenska.
Båda språken har långa traditioner i Finland.
Ungefär 90 procent av finländarna har finska som modersmål och ungefär fem procent av finländarna har svenska som modersmål.
När du uträttar ärenden med statliga myndigheter, till exempel vid arbets- och näringsbyrån (työ- ja elinkeinotoimisto), kan du använda endera språket.
Svenska talas mest på Finlands väst- och sydkust.
På somliga orter är svenskan vanligare än finskan.
Kontrollera vilket som är det vanligaste språket på din ort.
Kommunerna kan vara antingen enspråkiga eller tvåspråkiga.
I tvåspråkiga kommuner kan du använda antingen finska eller svenska när du uträttar ärenden med anställda inom kommunen, till exempel på socialbyrån (sosiaalitoimisto).
På vissa arbetsplatser måste man kunna både finska och svenska.
I skolorna i Finland lär man sig både finska och svenska.
Elever som har finska som modersmål lär sig svenska i skolan.
Elever som har svenska som modersmål lär sig finska i skolan.
Om ett invandrarbarn går i en skola där undervisningsspråket är finska studerar barnet också svenska som främmande språk tillsammans med de finskspråkiga eleverna.
Hurdant är det finska språket?
Finskan är ett finsk-ugriskt språk.
Besläktade språk är till exempel estniska och ungerska.
Finskan har många böjningsformer, till exempel kasusformer av nomen, personformer av verb och tempusformer.
Finskan har färre prepositioner än till exempel de indoeuropeiska språken.
Finskan har också en del postpositioner.
Ordföljden är friare än i många andra språk.
Finskan har även många lånord från till exempel svenska, tyska, ryska och engelska.
Finskans uttal är mycket regelbundet.
Betoningen ligger alltid på den första stavelsen.
I Finland är det vanligt att dua.
Ibland kan det vara artigt att nia.
Till exempel kunder och äldre människor nias ofta.
Hurdant är det svenska språket?
Svenskan är ett indoeuropeiskt språk som tillhör de nordeuropeiska germanska språken.
Besläktade språk är till exempel norska, danska och tyska.
I svenskan finns också många lånord från till exempel franskan.
I svenskan böjs verben i olika tempus.
Substantiven kategoriseras i två genus.
Adjektiven böjs efter dessa genus.
I svenskan är det vanligt med prepositioner och ordföljden är mycket regelbunden.
Den svenska som talas i Finland kallas finlandssvenska.
Den uttalas lite annorlunda än den svenska som talas i Sverige.
Svenskans uttal är relativt regelbundet.
Inhemska minoritetsspråk
Förutom finska och svenska talas även andra inhemska språk i Finland.
De samiska språken tillhör urspråken i Finland.
I Finlands talas tre olika varieteter av samiska.
De är finsk-ugriska språk.
Finsk romani hör till de indoeuropeiska språken.
I Finland finns också ett eget teckenspråk.
Mer information om dessa språk får du på webbplatsen för Forskningscentralen för de inhemska språken.
Information om språklagenfinska _ svenska _ engelska
linkkiKommuner.net:
Svenskspråkiga och tvåspråkiga kommunerfinska _ svenska
linkkiInstitutet för de inhemska språken:
Information om finska språketfinska _ svenska
linkkiInstitutet för de inhemska språken:
Information om svenska språketfinska _ svenska
linkkiInstitutet för de inhemska språken:
Information om de samiska språkenfinska _ svenska
linkkiInstitutet för de inhemska språken:
Information om finska romanifinska
linkkiInstitutet för de inhemska språken:
Information om det finska teckenspråketfinska _ svenska
Ordbok i det finska teckenspråketfinska
I Finland beskrivs språkkursernas nivåer på olika sätt.
Ofta använder man bedömningsskalan enligt den gemensamma europeiska referensramen (GER).
(Eurooppalainen viitekehys EVK) Denna skala omfattar följande nivåer:
nivåerna A1 och A2: grundläggande språkkunskaper (peruskielitaito)
nivåerna B1 och B2: en självständig språkanvändares språkkunskaper (itsenäisen kielenkäyttäjän kielitaito)
nivåerna C1 och C2: en avancerad språkanvändares språkkunskaper (taitavan kielenkäyttäjän kielitaito)
Dessa nivåer delas ytterligare in i undernivåer.
Till exempel omfattar nivå A1 kurserna A1.1, A1.2 och A1.3 och nivå A2 kurserna A2.1 och A2.2.
Mer information om hurdana kunskaper de olika nivåerna avser i praktiken får du på Utbildningsstyrelsens (Opetushallitus) webbplats.
Du kan också fråga direkt vid läroanstalterna.
I InfoFinland under rubriken Officiellt intyg över språkkunskaper får du information om hur du kan jämföra kursernas nivåer med nivån på den allmänna språkexamen (yleinen kielitutkinto).
linkkiUtbildningsstyrelsen:
Skala för beskrivning av språkkunskapsnivåer(pdf, 119,85 kb)finska _ svenska
linkkiEuropass.eu:
Utvärdera nivån på din språkkunskapfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
I Finland bor många människor i hyresbostäder.
Det som är bra med en hyresbostad är att det är lätt att byta bostad, eftersom du inte behöver sälja och köpa bostaden.
Men å andra sidan kan hyresvärden bestämma sig för att säga upp hyresavtalet, om han eller hon har en godtagbar anledning.
Då måste du flytta från hyresbostaden, även om du inte vill det.
På InfoFinlands sida Hyresavtal finns viktig information om uppsägning av hyresbostad, betalning av hyran, hyresdeposition och andra utgifter i en hyresbostad.
I större städer är det ofta svårare att hitta en lämplig hyresbostad. Även hyran är högre.
Reservera tillräckligt med tid för att hitta en bostad.
En del områden är väldigt populära. I sådana områden hyrs bostäderna ut mycket snabbt.
När du har hittat en lämplig bostad bör du snabbt bestämma dig om du vill ha den.
Då hyrsvärden väljer hyresgäst får han eller hon enligt lagen inte diskriminera någon exempelvis på grund av etniskt ursprung, religion eller nationalitet.
Läs mer på InfoFinlands sida Diskriminering och rasism.
Hur skaffar jag en hyresbostad?
När du letar efter en hyresbostad kan du leta efter annonser till exempel på internet.
Skriv in sökordet ”hyresbostad”.
Du kan även titta i lokaltidningarna.
Sökning av hyresbostäderfinska _ engelska
Sökning av hyresbostäderfinska
Privata hyresbostäder
Man får oftast en privat hyresbostad snabbare än en kommunal hyresbostad. Hyran för en privat bostad är ofta högre.
Du behöver inte anlita en bostadsmäklare för att söka bostad.
Du kan själv söka information om lediga bostäder.
Då behöver du inte heller betala mäklararvode (välityspalkkio).
Du kan söka privata hyresbostäder på internet och i lokaltidningar.
Du kan även publicera en egen annons.
Om du vill hyra en privat hyresbostad ska du kontakta den som hyr ut bostaden. Kom överens om när du kan gå och titta på bostaden.
En bostadsvisning ordnas oftast för alla intresserade på samma gång.
Samtidigt får du en ansökningsblankett.
Fyll i den om du vill flytta in i bostaden.
Om du vill att en mäklare söker en lämplig hyresbostad åt dig, ska du ingå ett skriftligt uppdragsavtal (toimeksiantosopimus) med mäklaren.
Du måste då betala mäklararvode till mäklaren.
Avtala om arvodet skriftligen på förhand.
Arvodet kan till exempel vara lika stort som en månads hyra.
Jämför olika mäklarbyråers priser på förhand.
När du hyr en privat bostad ska du göra ett hyresavtal med hyresvärden.
Läs mera på InfoFinlands sida Hyresavtal.
Priser på icke subventionerade hyresbostäderengelska
Kommunernas hyresbostäder
Även kommunerna äger hyresbostäder. De är ofta förmånligare än andra hyresbostäder.
Du kan söka boende i en hyresbostad som staten stödjer, om du har något av följande:
Finskt medborgarskap;
registrerat uppehållstillstånd;
uppehållskort;
uppehållstillstånd som är giltigt i minst ett år; eller
uppehållstillstånd för studerande.
Om du vill ansöka om en kommunal hyresbostad fyller du i ansökningsblanketten på bostadskontoret i din kommun.
Ofta kan du även fylla i och skicka blanketten på kommunens webbsida.
I en del kommuner är hyresbostäderna så populära att man kan vara tvungen att stå i kö mycket länge.
Köerna till bostäderna kan vara långa till exempel i huvudstadsregionen (Helsingfors, Esbo och Vanda), men det finns lediga bostäder på mindre orter runt om i Finland.
När hyresgästerna väljs beaktas
inkomster
egendom
behovet av bostad.
I Finland finns även många allmännyttiga samfund som har förmånliga hyresbostäder.
Priser på hyresbostäder med statliga stödengelska
Studentbostäder
Om du är studerande kan du söka en hyresbostad som är avsedd särskild för studerande.
Läs mer på InfoFinlands sida Boende för studerande.
Bostadsansökan och bilagor
När du lämnar in en bostadsansökan kan du behöva också andra dokument som bilagor till ansökan.
Dessa beror på varifrån du söker bostaden.
senaste löneintyg
kopia på beskattningsbeslutet där din egendom framgår
intyg över lån
kopia på uppehållstillstånd eller pass om du inte är EU-medborgare.
Ofta granskas även den bostadssökandes kredituppgifter.
linkkiKonkurrens- och konsumentverket:
Att hyra en bostadfinska _ svenska _ engelska
Information för hyresgästenfinska _ svenska _ engelska
linkkiMiljöministeriet:
Information om hyresboendefinska _ svenska _ engelska
linkkiKonsumentförbundet ry:
Hyreshandboken(pdf, 1,11 MB)finska _ svenska _ ryska _ franska _ somaliska _ arabiska
Hyresbostadens utrustning
I utrustningen i en hyresbostad ingår nästan alltid köksskåpen, kylskåpet och spisen.
Även klädskåp och skåp i hallen ingår vanligtvis.
Duschen, vattenkranarna och toalettstolen hör alltid till utrustningen.
Hyresbostäder är vanligtvis inte möblerade.
Det händer dock att lägenheter hyrs ut med möbler.
Vilka möbler som ingår varierar.
Kontrollera alltid med hyresvärden vilka möbler som ingår.
Hushållsavfall
I Finland ska hushållsavfall sorteras i olika sopkärl.
Läs mer på InfoFinlands sida Avfallshantering och återvinning.
Rådgivningstjänster
Vill du söka råd om att hyra en bostad?
Finlands Konsumentförbund erbjuder råd och handledning både för hyresgäster och hyresvärder.
Finlands Konsumentförbunds rådgivningstjänst:
tfn 010 8022 40
tis-fre kl. 10–12 och tis kl. 17–19
Du kan ringa till tjänsten och endast betala lokalsamtalsavgift överallt i Finland.
Du kan fråga råd på tjänsten även på nätet genom att fylla i en blankett. Du får svar per e-post.
Även Marthaförbundet och Finlands flyktinghjälp erbjuder bostadsrådgivning åt invandrare.
linkkiKonsumentförbundet:
Boenderådgivningfinska
linkkiFlyktinghjälp:
Flyktinghjälpens regionkontorfinska
linkkiMarthaförbundet:
Kontaktuppgifter till Marthaförbundetfinska _ engelska
Tvåspråkiga kommuner i Finland
Finland har två officiella språk, finska och svenska.
Finska är modersmålet för cirka 90 procent av finländarna.
Svenska är modersmålet för cirka 5 procent av finländarna.
Svenska talas mest på Finlands väst- och sydkust.
Svenskan som talas i Finland är finlandssvenska.
Uttalet skiljer sig något från svenskan i Sverige.
Om du vill ansöka om finskt medborgarskap behöver du ett intyg över tillräckliga kunskaper i finska eller svenska.
Läs mer på InfoFinlands sida Officiellt intyg över språkkunskaper.
Du kan använda svenska med statliga myndigheter, till exempel FPA eller TE-byrån.
Ange ditt kontaktspråk till magistraten när du registrerar dig som invånare.
Du kan även ändra kontaktspråket senare.
Kommunerna i Finland kan vara antingen enspråkiga eller tvåspråkiga.
De flesta kommunerna i Finland är finskspråkiga.
Tvåspråkiga kommuner finns på väst- och sydkusten.
Om din hemkommun är tvåspråkig, kan du använda svenska även inom de kommunala tjänsterna, till exempel på hälsostationen.
linkkiKommuner.net:
Svenskspråkiga och tvåspråkiga kommunerfinska _ svenska
Integration på svenska kan vara ett bra alternativ för dig till exempel om:
Du bor i ett område med många svensktalande.
Du har svenskspråkiga familjemedlemmar eller släktingar.
Du kan lite svenska redan.
Det kan vara fördelaktigt att kunna svenska när du söker jobb.
Tänk ändå på att kunskaper i finska krävs på de flesta arbetsplatserna.
Även om du väljer integrationsutbildning på svenska lönar det sig för dig att i något skede även lära dig finska.
I en del kommuner kan du delta i integrationsutbildning på svenska.
Om du inte blir antagen till integrationsutbildning på svenska kan du i vissa fall få stöd för frivilliga studier i svenska, om detta överenskommits i din integrations- eller sysselsättningsplan.
Fråga om integration på svenska när din inledande kartläggning och integrationsplan görs.
Enligt lag har du rätt att välja antingen finska eller svenska som integrationsspråk.
linkkiArbets- och näringsministeriet:
Information om integration på svenskafinska _ svenska
Språkstudier som arbetskraftsutbildning
Om du är kund vid arbets- och näringsbyrån kan du också studera svenska som arbetskraftsutbildning.
Arbetskraftsutbildningen är avsedd för arbetslösa arbetssökande.
Läs på InfoFinlands sida Arbets- och näringsbyråns tjänster vad som krävs för att du ska kunna bli kund hos arbets- och näringsbyrån.
Arbetskraftsutbildningen är kostnadsfri för dig.
Fråga mer om kurser i svenska vid din egen arbets- och näringsbyrå.
Barndagvård och utbildning för barn
I Finland ges dagvård, förskoleundervisning och grundläggande utbildning vanligtvis på finska eller svenska.
Om du vill att ditt barn ska börja i svenskspråkig dagvård, förskola eller skola, fråga om möjligheterna i din hemkommun.
Vissa kommuner ordnar förberedande undervisning före den grundläggande utbildningen för elever som ännu inte har tillräckligt bra språkkunskaper för den vanliga undervisningen.
Fråga i din hemkommun om förberedande undervisning ordnas på svenska i kommunen.
Om barnet har något annat modersmål än finska eller svenska, kan kommunen ordna undervisning i barnets eget modersmål för barnet.
Om barnet går i en svensk skola kan hen läsa svenska som andra språk.
Läs mer om barndagvård, förskoleundervisning och grundläggande utbildning på InfoFinlands sida Det finländska utbildningssystemet.
Gymnasium och yrkesläroanstalt
Efter grundskolan kan du studera på gymnasiet eller en yrkesläroanstalt.
Svenskspråkiga yrkesläroanstalter och gymnasieskolor finns i svenskspråkiga och tvåspråkiga kommuner och i en del finskspråkiga kommuner.
Vissa yrkesläroanstalter och gymnasieskolor ordnar förberedande utbildning före studierna.
I den förberedande utbildningen får du sådana kunskaper och färdigheter som du behöver i dina fortsatta studier.
Du kan också förbättra dina språkkunskaper.
Du kan söka svenskspråkig yrkes- och gymnasieutbildning samt förberedande utbildning före dessa via tjänsten Opintopolku.fi.
Läs mer på InfoFinlands sida: Efter grundskolan.
Grundläggande information om yrkesutbildningfinska _ svenska _ engelska
Information om gymnasiestudierfinska _ svenska
Högskoleutbildning
I Finland finns svenskspråkiga yrkeshögskolor och universitet.
Dessutom finns det några tvåspråkiga universitet där du kan läsa på svenska.
Du kan söka svenskspråkiga högskoleutbildningar via tjänsten Opintopolku.fi.
Läs mer om högskoleutbildning på InfoFinlands sida: Högskoleutbildning.
Information om högskolestudierfinska _ svenska _ engelska
Var kan jag läsa svenska?
Du kan läsa svenska till exempel vid medborgarinstitut, arbetarinstitut och sommaruniversitet.
Fråga om studier i svenska hos utbildningsväsendet i din hemkommun, studievägledarna vid läroanstalter eller rådgivningstjänsterna för invandrare.
Läs mer på InfoFinlands sida: Studier som hobby.
Svenska på internet
Appar
Du kan lära dig svenska med hjälp av appar som du kan ladda ned i din telefon eller surfplatta.
Sök appar för svenska i din appbutik (t.ex. Google Play och App Store) med sökorden ”learn Swedish”, ”Swedish language”, ”lär dig svenska” eller ”svenska”.
En del appar kostar pengar.
Övningar och kurser på internet
På internet hittar du kurser i det svenska språket på olika nivåer.
På internet kan du till exempel göra övningar och spela spel, lära dig grammatik och vokabulär samt läsa texter.
linkkiYle:
Övningar för allmänna språkexaminafinska
Svenska på internetfinska _ svenska _ engelska
linkkiYle.fi:
Övningar och kurser på internetfinska
linkkiBab.la:
Flerspråkiga ordböckerfinska _ svenska _ engelska
I Finland finns många möjligheter att studera finska.
Olika kurser ordnas för både barn och vuxna.
Undervisning i finska för vuxna
Du hittar information om kurser i finska till exempel hos medborgarinstitut, arbetarinstitut, universitet och sommaruniversitet.
Fråga mer vid rådgivningstjänsterna för invandrare, utbildningsväsendet i din hemkommun eller studievägledarna vid lokala läroanstalter.
På vissa orter har informationen om kurserna samlats på ett och samma ställe.
Till exempel finns det information om kurserna i finska språket i Helsingfors, Tammerfors och Åbo i tjänsten Finnishcourses.fi.
Vid läroanstalterna börjar kurserna vanligtvis i augusti eller september och i januari.
Språkkurserna är ofta fullsatta.
Därför är det viktigt att anmäla sig till kursen i god tid.
Medborgarinstitut i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Kurser i finska och svenska språketfinska _ engelska _ ryska
Språkstudier i anslutning till annan utbildning
Du kan studera finska också i arbetskraftsutbildning och i förberedande utbildning före yrkesutbildning (VALMA) eller förberedande gymnasieutbildning (LUVA).
Om du är kund vid arbets- och näringsbyrån kan du få plats på en kurs i finska via arbets- och näringsbyrån.
Hurdan språkundervisning du behöver bedöms på arbets- och näringsbyrån i samband med att du får en integrations- eller sysselsättningsplan.
Du kan studera finska som arbetskraftsutbildning.
Arbetskraftsutbildning är i huvudsak utbildning avsedd för arbetslösa arbetssökande.
Utbildningen är kostnadsfri för deltagarna.
Fråga om kurserna i finska på din egen arbets- och näringsbyrå.
linkkiArbets- och näringsministeriet:
Kontaktuppgifter till TE-byråerfinska _ svenska
linkkiArbets- och näringsministeriet:
Utbildning i finska och svenska språketfinska _ svenska _ engelska
Finska på arbetsplatsen
Vissa arbetsgivare ordnar finskundervisning för sina arbetstagare.
Fråga din arbetsgivare om du kan studera finska på din arbetsplats.
Arbetsgivaren kan ansöka om stöd för arbetstagarnas finskundervisning via arbets- och näringslivstjänsterna.
linkkiTE-tjänster:
Finska på arbetsplatsenfinska _ svenska _ engelska
Undervisning i finska för barn
Barn lär sig nya språk snabbt, även om det kan kännas svårt i början.
Finskundervisning ges på daghem, i förskola och skola.
Undervisningen kallas finska som andra språk eller S2-undervisning.
Barnet eller den unga kan även delta i förberedande undervisning.
Den är avsedd för de elever som ännu inte har särskilt bra kunskaper i finska.
Under den förberedande undervisningen studerar barnet eller den unga finska och några läroämnen.
Den förberedande undervisningen är avsedd för 7–16-åringar.
Undervisningen varar vanligtvis ett år.
Därefter flyttas eleven till en vanlig klass.
linkkiUtbildningsstyrelsen:
Finska som andra språk i den grundläggande undervisningenfinska _ svenska
Checklista för dig som flyttar
När du flyttar i Finland från en bostad till en annan:
Kom ihåg att göra flyttanmälan (muuttoilmoitus).
Du kan göra flyttanmälan högst en månad före flyttningsdagen, men den bör göras senast en vecka efter att du har flyttat.
Flyttanmälan ska alltid göras till magistraten (maistraatti).
Du kan göra flyttanmälan
på nätet
telefonledes på finska på numret 0295 535 535 eller på svenska på numret 0295 535 536 eller
på en blankett som du får på posten eller hos magistraten.
Om du bor i höghus eller radhus ska du alltid också komma ihåg att meddela husets disponent (isännöitsijä) att du flyttar.
Meddela din nya adress till alla instanser som skickar dig post.
Vissa organisationer och företag får din nya adress direkt från befolkningsregistret.
Du har ändå själv ansvaret för att dina fakturor skickas till rätt adress och betalas i tid.
Om du bor i en hyresbostad ska du komma ihåg att säga upp din gamla bostad i tid.
Det är bäst att göra uppsägningen skriftligt.
Kontrollera hur lång uppsägningstid du har för bostaden.
Vanligen är den en kalendermånad.
Läs mer på InfoFinlands sida Hyresavtal.
Om du har barn ska du se till att skaffa dem nya dagvårds- och skolplatser.
Du måste meddela daghemmet och skolan när barnen slutar där.
Samtidigt är det bra att anmäla barnen till det nya daghemmet eller den nya skolan.
Kom ihåg att skaffa eventuell flytthjälp i tid.
Bland annat vid månadsskift och på veckoslut är flyttfirmorna alltid upptagna.
Avtala med din tjänsteleverantör om överföringen av din internetanslutning i god tid så att det inte blir ett avbrott i servicen.
Säg upp ditt gamla elavtal innan du flyttar och gör upp ett nytt.
Det lönar sig att jämföra olika elbolags priser så att du hittar det förmånligaste.
Du får ett elavtal genom att ringa upp elbolaget och meddela ditt namn och din nya adress.
Om du flyttar till ett egnahemshus ska du också komma ihåg att teckna andra avtal, såsom avtal om vattenförsörjning och avfallshantering.
Om huset värms upp med olja ska du komma ihåg att kontrollera oljemängden.
Kontrollera om dina nuvarande försäkringar, som hemförsäkringen, är tillräckliga även för den nya bostaden.
Om du till exempel flyttar från höghus till egnahemshus behöver du förmodligen en annorlunda försäkring.
Städa den gamla bostaden innan du flyttar och töm vinden, källarförrådet och garaget på saker.
Om du bor i en hyresbostad ska du ge ägaren eller disponenten alla nycklar till den gamla bostaden.
linkkiFörbundet för ungdomsbostäder:
Ordlista om boendefinska
Flyttanmälanfinska _ svenska _ engelska
linkkiEnergimarknadsverket:
Jämför elpriserfinska
Flyttjänsterfinska _ engelska
Flyttjänsterfinska _ engelska _ ryska
Flyttjänsterfinska _ svenska _ engelska
När du flyttar till Finland
Om du vill ha information om praktiska frågor i anslutning till att du flyttar till Finland, läs mer på sidan Komihåglista för dig som flyttar till Finland.
Om du nyligen har flyttat till Finland, måste du registrera dig som invånare.
Lär mer på InfoFinlands sida Registrering som invånare.
Flytta från Finland
Planerar du att flytta från Finland till ett annat land?
Läs mer på InfoFinlands sida Flytta från Finland.
Om du vill ansöka om finskt medborgarskap behöver du ett officiellt intyg över dina kunskaper i finska eller svenska.
Du kan behöva intyget också när du söker ett jobb eller en studieplats.
Du kan påvisa dina språkkunskaper:
med en allmän språkexamen (yleinen kielitutkinto)
med vitsordet i finska eller svenska på ditt avgångsbetyg (päättötodistus).
Allmän språkexamen
Allmän språkexamen, ASE, är ett språktest för vuxna.
Med en allmän språkexamen kan du påvisa dina kunskaper i finska eller svenska.
Examen är avgiftsbelagd.
När du avlagt examen får du ett intyg som anger nivån på dina språkkunskaper.
Språkexamen finns på tre olika nivåer: grundnivån, mellannivån och högsta nivån.
Varje examensnivå består av två färdighetsnivåer, vilka det alltså finns sammanlagt sex av.
Grundnivån är avsedd för personer som kan använda språket i vardagliga sammanhang.
Deras färdighetsnivå är 1–2.
Medelnivån är avsedd för personer som kan språket relativt väl. Deras färdighetsnivå är 3–4.
Den högsta nivån är avsedd för personer som kan språket mycket väl. Deras färdighetsnivå är 5–6.
Närmare beskrivningar av de olika färdighetsnivåerna finns på Utbildningsstyrelsens webbplats.
Om du vill ansöka om finskt medborgarskap (kansalaisuus) kan du påvisa att du har tillräckliga kunskaper i finska eller svenska genom att avlägga den muntliga och skriftliga delen av en allmän språkexamen minst på nivå 3.
Språkexamenstillfället pågår 3–6 timmar.
Uppgifternas ämnesområden rör det vardagliga livet såsom fritid, utbildning och vanliga situationer på arbetet.
I examen ingår olika uppgifter där följande färdigheter krävs:
textförståelse
skriftliga färdigheter
grammatik och vokabulär
talförståelse
Du kan avlägga examen på olika orter i Finland.
Mer information om anmälan får du på Utbildningsstyrelsens (Opetushallitus) webbplats.
Examina kategoriseras på en annan skala än kurserna.
Om du har slutfört en språkkurs som kategoriserats enligt den europeiska referensramen motsvarar kursen nivån på den allmänna språkexamen ungefär enligt följande tabell:
A1 – ASE 1
A2 – ASE 2
B1 – ASE 3
B2 – ASE 4
C1 – ASE 5
C2 – ASE 6
Innan du anmäler dig till examen ska du göra dig förtrogen med kraven på de olika examensnivåerna.
Du kan även fråga din lärare i finska.
Mer information om den allmänna språkexamen får du på Utbildningsstyrelsens webbplats.
linkkiUtbildningsstyrelsen:
Allmänna språkexaminafinska _ svenska _ engelska
linkkiUtbildningsstyrelsen:
Färdighetsnivåerna i allmänna språkexaminafinska _ svenska _ engelska
linkkiUtbildningsstyrelsen:
Att anmäla sig till en allmän språkexamen och examensavgifterfinska _ svenska _ engelska
Statsförvaltningens språkexamen om kunskaper i finska och svenska
Om du vill arbeta inom den offentliga förvaltningen behöver du vanligtvis ett intyg över dina kunskaper i finska eller svenska.
Du kan påvisa dina kunskaper i finska eller svenska med statsförvaltningens språkexamen.
Fråga din arbetsgivare hurdana språkkunskapskrav som gäller på den arbetsplats som du vill söka.
Språkexamen finns på tre olika nivåer: för nöjaktiga, goda och utmärkta språkkunskaper.
Det beror på din arbets- eller studieplats vilken examensnivå du måste avlägga.
För finskt medborgarskap behöver du ett intyg för åtminstone nöjaktiga språkkunskaper.
Du kan avlägga examen för nöjaktiga eller goda språkkunskaper olika orter i Finland.
På Utbildningsstyrelsens webbplats hittar du en förteckning över de städer där examen kan avläggas.
Examen på utmärkt nivå kan endast avläggas i Helsingfors.
Examen omfattar olika tester. I dem ska du läsa och lyssna på texter och svara på frågor.
Därtill finns det intervjuer, diskussioner och skriftliga uppgifter.
Du kan ersätta statsförvaltningens språkexamen med vissa andra studier.
Till exempel motsvarar statsförvaltningens språkexamen som gäller goda språkkunskaper ett mognadsprov (kypsyysnäyte) som du har avlagt på finska eller svenska vid universitetet.
Mer information får du på Utbildningsstyrelsens webbplats.
linkkiUtbildningsstyrelsen:
Statsförvaltningens språkexaminafinska _ svenska
linkkiUtbildningsstyrelsen:
Färdighetsnivåerna i statsförvaltningens språkexaminafinska _ svenska
linkkiUtbildningsstyrelsen:
Mottagare av statsförvaltningens språkexamina, finska språketfinska _ svenska
linkkiUtbildningsstyrelsen:
Mottagare av statsförvaltningens språkexamina, svenska språketfinska _ svenska
Intyg över språkkunskaper på basis av studier
Om du vill ansöka om finskt medborgarskap kan du påvisa dina kunskaper i finska eller svenska även med något av följande intyg:
avgångsbetyg från grundskolan med ett godkänt vitsord i finska eller svenska som modersmål eller som andra språk
avgångsbetyg från gymnasiet med ett godkänt vitsord i finska eller svenska som modersmål eller som andra språk
studentexamen på finska eller svenska med ett godkänt vitsord i finska eller svenska som modersmål eller som andra språk
intyg på yrkesinriktad grundexamen som du har avlagt på finska eller svenska
intyg på yrkesexamen som du har avlagt på finska eller svenska
intyg på studier i tjänstemannafinska eller -svenska som du har avlagt vid universitet eller högskola
intyg på mognadsprov som du har avlagt på finska eller svenska för universitetsexamen eller yrkeshögskoleexamen
Mer information får du på Migrationsverkets (Maahanmuuttovirasto) webbplats.
linkkiUtbildningsstyrelsen:
Språkkunskaper och finskt medborgarskapfinska _ svenska _ engelska
Ungefär 90 procent av finländarna har finska som modersmål.
Ungefär fem procent av finländarna har svenska som modersmål.
När du funderar på om det är finska eller svenska som du borde lära dig ska du beakta vilket språk som talas på din hemort och i din näromgivning.
Om du vill ansöka om finskt medborgarskap måste du kunna finska, svenska eller i det finska teckenspråket.
När du ansöker om medborgarskap, bifoga ett intyg över dina språkkunskaper.
Läs mer om språkkunskapskraven på InfoFinlands sida Officiellt intyg över språkkunskaper.
På de flesta arbetsplatser är det nödvändigt att kunna finska.
Om du vill studera i Finland behöver du sannolikt kunna finska.
Det kan vara bra att lära sig finska eller svenska trots att du inte tänker bo en lång tid i landet.
Även om finländarna i allmänhet behärskar engelska relativt väl har du ändå mycket nytta av att kunna finska eller svenska.
När du behärskar språket är det lättare för dig att trivas i landet och anpassa dig till livet i Finland.
Du har lättare att sköta dina ärenden med myndigheter, följa nyheter, få nya bekantskaper och vänner.
Du lär dig språket bäst om du vågar använda det.
Du behöver inte alltid förstå allting, det räcker med att du förstår det viktigaste.
Dra dig alltså inte för situationer där du har möjlighet att tala finska eller svenska.
Information om språklagenfinska _ svenska _ engelska
linkkiKommuner.net:
Svenskspråkiga och tvåspråkiga kommunerfinska _ svenska
God morgon!
God dag!
God kväll!
God natt!
Välkommen!
Tack.
Var så god.
Förlåt.
Jag älskar dig.
Hur står det till?
Hejdå.
Adjö.
Jag förstår inte, kan du upprepa?
Jag talar inte finska.
Jag talar bara lite finska.
Talar du engelska/svenska?
Jag är lärare / ingenjör / studerande.
Vad är ditt telefonnummer / din e-postadress?
Var finns det en affär / ett apotek / en skola / ett daghem / en busstation / en metrostation?
På nätet hittar du finskakurser på många olika nivåer.
På nätet kan du till exempel göra övningar, spela spel, lära dig grammatik och vokabulär och läsa texter.
De flesta webbkurser är på finska eller svenska, men det finns även andra alternativ:
Nybörjarnivån
linkkiYle:
Nybörjarkurs i finska, Easyfinnishfinska
Nybörjarkurs i finska "A Taste of Finnish"engelska
linkkiTammerfors yrkeshögskola:
Nybörjarkurs i finska, Uunofinska
Nybörjarkurs i finska, Tavataan taasengelska _ franska _ tyska _ bulgariska
Nybörjarkurs i finskafinska _ svenska _ engelska _ arabiska
linkkiWordDive:
Nybörjarkurs i finskafinska _ svenska _ engelska _ ryska _ kinesiska _ tyska
Inledningskurs i finskaengelska
Tilläggsövningar till läroboken Hyvin meneefinska
Mångsidiga övningar i finska språketfinska
Ordspel för nybörjareengelska _ franska _ japanska
Applikationen Suomipassi med flera stödspråkfinska _ engelska
Grundnivån
linkkiYle:
Övningar för allmänna språkexaminafinska
Webbkurs med många hjälpspråksvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ portugisiska
linkkiEdu.fi:
Vardagsfinska: videoinspelning med intervjuerfinska
Vokabulärövningarfinska
linkkiYle:
Läromaterial från TV-serien Supisuomeafinska
linkkiUtbildningsstyrelsen:
Finska i arbetslivetfinska
Mångsidiga övningar i finska språketfinska
Lär dig finska med hjälp av filmerfinska _ engelska _ persiska _ arabiska
Självständiga språkanvändare
linkkiYle:
Nyheter på klarspråkfinska
Information om olika ämnen på klarspråkfinska
Nyheter på lättläst finskafinska
linkkiUtbildningsstyrelsen:
linkkiUtbildningsstyrelsen:
Finska i arbetslivetfinska
Avancerade språkanvändare
Lyssna på finska dialekterfinska
linkkiWordDive:
Finskans grammatikfinska _ svenska _ engelska _ ryska _ spanska _ tyska _ japanska
Finskans grammatikengelska
Finskans grammatikengelska
Verbböjningengelska
linkkiInstitutet för de inhemska språken:
Grammatiken Iso suomen kielioppi på nätetfinska
Information om finska språketengelska
Ordböcker på nätet
Flerspråkiga ordböckerfinska
linkkiBab.la:
Flerspråkiga ordböckerfinska _ svenska _ engelska
Intern kommunikation på arbetsplatsen
Vanligen informerar man om kommande händelser och ändringar på arbetsplatsen vid möten.
Om man deltar i möten kan man påverka, föreslå ändringar och utveckla sitt eget arbete.
På varje arbetsplats finns också andra kanaler för den interna kommunikationen, såsom anslagstavlor, e-post eller de anställdas postfack.
Följ informationen på arbetsplatsen.
Pauser
I arbetsavtalet står det ofta hur långa pauser som ingår i arbetsdagen och tidpunkten för dessa.
Vanligen har man en kort kaffepaus på förmiddagen, en lunchpaus mitt på dagen och en kaffepaus till på eftermiddagen.
Längden på lunchpausen varierar mellan olika arbetsplatser.
Fråga din chef hur långa pauser du har.
Arbetsplatsbespisningen är ordnad på olika sätt på olika arbetsplatser: vissa arbetsplatser har en egen personalmatsal, på andra ställen tar de anställda med sig maten hemifrån.
På vissa arbetsplatser kan man köpa förmånliga lunchsedlar som man kan använda på matställen i närheten av arbetsplatsen.
Under lunchen arbetar man vanligtvis inte.
Att sköta egna ärenden under arbetsdagen
På arbetstid får man inte sköta sina privata angelägenheter, utan detta måste göras utanför arbetstiden.
Antalet arbetstimmar som står i arbetsavtalet är bindande och det avtalade antalet arbetstimmar ska fullgöras.
Under pauserna kan du till exempel ringa viktiga samtal.
Du kan också ansöka om oavlönad ledighet om din situation kräver att du är frånvarande en längre tid.
Om du av någon anledning inte till exempel lyckas få en läkartid utanför arbetstiden, ska du komma överens med din chef om att du är borta och hur du ersätter din frånvaro.
Företagshälsovården kan du besöka under arbetstid.
Utbildning som rör arbetet
Även om arbetstagaren har sådan utbildning som krävs för yrket redan när anställningen inleds, uppmuntrar många arbetsgivare sina anställda att skaffa sig mer utbildning.
Ofta kan du utbilda dig på arbetstid och arbetsgivaren kan betala för utbildningen.
De flesta arbetsgivare värdesätter att den anställda vill utveckla sig i sitt arbete och inhämta nya kunskaper.
Vanligen ger man inte varandra presenter på arbetsplatserna.
På viktiga bemärkelsedagar (födelsedagar, äktenskap, pensionering) uppmärksammar arbetskamraterna och arbetsgivaren festföremålet med en liten present eller en blombukett.
Arbetstid och semester
En normal arbetsdag är vanligtvis åtta timmar.
Arbetstagaren kan även komma överens om någon annan tid med arbetsgivaren.
I Finland gör arbetstagare vanligtvis inte mycket övertid.
Man arbetar de timmar som står i anställningsavtalet.
I Finland börjar semesterperioden i början av maj.
Antalet intjänade semesterdagar beror på anställningstiden i år och när anställningen har börjat.
Utöver den betalda semesterna kan du ansöka om obetald ledighet.
Jämfört med många andra länder har arbetstagare i Finland långa semestrar.
Arbetshälsa och rekreation
På många arbetsplatser vill man stödja de anställdas arbetsmotivation och -trivsel med olika rekreationsdagar och fester på arbetsplatsen. Arbetsgivaren kan också erbjuda sina anställda olika hobbymöjligheter vid sidan av arbetet.
Årliga helger
Vissa dagar är allmänna lediga dagar i Finland.
Till dem hör följande:
nyårsdagen 1.1
trettondagen 6.1
påsk: tidpunkten varierar, i mars-april
första maj 1.5
midsommarafton: i juni, alltid en fredag
självständighetsdagen 6.12
juldagen 25.12
annandag jul 26.12
Läs mer om dessa dagar på sidan Finländska helgdagar.
På vissa arbetsplatser, till exempel sjukhus, arbetar man även under helgerna.
För arbetet under helgerna betalas högre lön.
Kontrollera ersättningen i ditt kollektivavtal.
Finland är ett tvåspråkigt land
Finland har två officiella språk, finska och svenska.
Båda språken har långa traditioner i Finland.
Ungefär 90 procent av finländarna har finska som modersmål och ungefär fem procent av finländarna har svenska som modersmål.
När du uträttar ärenden med statliga myndigheter, till exempel vid arbets- och näringsbyrån (työ- ja elinkeinotoimisto), kan du använda endera språket.
Svenska talas mest på Finlands väst- och sydkust.
På somliga orter är svenskan vanligare än finskan.
Kontrollera vilket som är det vanligaste språket på din ort.
Kommunerna kan vara antingen enspråkiga eller tvåspråkiga.
I tvåspråkiga kommuner kan du använda antingen finska eller svenska när du uträttar ärenden med anställda inom kommunen, till exempel på socialbyrån (sosiaalitoimisto).
På vissa arbetsplatser måste man kunna både finska och svenska.
I skolorna i Finland lär man sig både finska och svenska.
Elever som har finska som modersmål lär sig svenska i skolan.
Elever som har svenska som modersmål lär sig finska i skolan.
Om ett invandrarbarn går i en skola där undervisningsspråket är finska studerar barnet också svenska som främmande språk tillsammans med de finskspråkiga eleverna.
Hurdant är det finska språket?
Finskan är ett finsk-ugriskt språk.
Besläktade språk är till exempel estniska och ungerska.
Finskan har många böjningsformer, till exempel kasusformer av nomen, personformer av verb och tempusformer.
Finskan har färre prepositioner än till exempel de indoeuropeiska språken.
Finskan har också en del postpositioner.
Ordföljden är friare än i många andra språk.
Finskan har även många lånord från till exempel svenska, tyska, ryska och engelska.
Finskans uttal är mycket regelbundet.
Betoningen ligger alltid på den första stavelsen.
I Finland är det vanligt att dua.
Ibland kan det vara artigt att nia.
Till exempel kunder och äldre människor nias ofta.
Hurdant är det svenska språket?
Svenskan är ett indoeuropeiskt språk som tillhör de nordeuropeiska germanska språken.
Besläktade språk är till exempel norska, danska och tyska.
I svenskan finns också många lånord från till exempel franskan.
I svenskan böjs verben i olika tempus.
Substantiven kategoriseras i två genus.
Adjektiven böjs efter dessa genus.
I svenskan är det vanligt med prepositioner och ordföljden är mycket regelbunden.
Den svenska som talas i Finland kallas finlandssvenska.
Den uttalas lite annorlunda än den svenska som talas i Sverige.
Svenskans uttal är relativt regelbundet.
Inhemska minoritetsspråk
Förutom finska och svenska talas även andra inhemska språk i Finland.
De samiska språken tillhör urspråken i Finland.
I Finlands talas tre olika varieteter av samiska.
De är finsk-ugriska språk.
Finsk romani hör till de indoeuropeiska språken.
I Finland finns också ett eget teckenspråk.
Mer information om dessa språk får du på webbplatsen för Forskningscentralen för de inhemska språken.
Information om språklagenfinska _ svenska _ engelska
linkkiKommuner.net:
Svenskspråkiga och tvåspråkiga kommunerfinska _ svenska
linkkiInstitutet för de inhemska språken:
Information om finska språketfinska _ svenska
linkkiInstitutet för de inhemska språken:
Information om svenska språketfinska _ svenska
linkkiInstitutet för de inhemska språken:
Information om de samiska språkenfinska _ svenska
linkkiInstitutet för de inhemska språken:
Information om finska romanifinska
linkkiInstitutet för de inhemska språken:
Information om det finska teckenspråketfinska _ svenska
Ordbok i det finska teckenspråketfinska
I Finland beskrivs språkkursernas nivåer på olika sätt.
Ofta använder man bedömningsskalan enligt den gemensamma europeiska referensramen (GER).
(Eurooppalainen viitekehys EVK) Denna skala omfattar följande nivåer:
nivåerna A1 och A2: grundläggande språkkunskaper (peruskielitaito)
nivåerna B1 och B2: en självständig språkanvändares språkkunskaper (itsenäisen kielenkäyttäjän kielitaito)
nivåerna C1 och C2: en avancerad språkanvändares språkkunskaper (taitavan kielenkäyttäjän kielitaito)
Dessa nivåer delas ytterligare in i undernivåer.
Till exempel omfattar nivå A1 kurserna A1.1, A1.2 och A1.3 och nivå A2 kurserna A2.1 och A2.2.
Mer information om hurdana kunskaper de olika nivåerna avser i praktiken får du på Utbildningsstyrelsens (Opetushallitus) webbplats.
Du kan också fråga direkt vid läroanstalterna.
I InfoFinland under rubriken Officiellt intyg över språkkunskaper får du information om hur du kan jämföra kursernas nivåer med nivån på den allmänna språkexamen (yleinen kielitutkinto).
linkkiUtbildningsstyrelsen:
Skala för beskrivning av språkkunskapsnivåer(pdf, 119,85 kb)finska
linkkiEuropass.eu:
Utvärdera nivån på din språkkunskapfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
I Finland värdesätts ärlighet, punktlighet och jämställdhet.
Det syns överallt i den finländska kulturen, även i arbetslivet.
På den här sidan finns mer information om den finländska arbetskulturen.
Lagar och avtal i arbetslivet
Arbetslivet i Finland styrs av många regler som arbetstagaren och arbetsgivaren måste följa.
I lagstiftningen och kollektivavtalen fastställs till exempel minimilöner, arbetstider, semester, lön under sjukskrivning och uppsägningsvillkor.
Ibland kan arbetsgivaren be arbetstagaren arbeta övertid.
Enligt lag ska arbetsgivaren betala högre lön för övertid.
Du kan även få ersättningen i form av ledighet.
Du har rätt att vägra övertidsarbete.
Information om arbetstagarnas rättigheter och skyldigheter i Finland hittar du på InfoFinlands sida Arbetstagarens rättigheter och skyldigheter.
linkkiFFC:
Arbetslivet i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ kinesiska _ arabiska
Lär dig finska eller svenska
Du kan utveckla dina språkkunskaper på kurser eller i arbetet.
Dra dig inte för att prata finska eller svenska med dina kollegor.
Läs mer om språkstudier i InfoFinlands avsnitt Finska och svenska språket.
Jämlikhet och jämställdhet i arbetslivet
Enligt finsk lag är alla slags diskriminering på arbetsplatserna förbjuden.
Arbetsgivaren ska se till att jämlikhet och jämställdhet mellan könen förverkligas på arbetsplatsen.
Läs mer på InfoFinlands sida Jämlikhet och jämställdhet i arbetslivet.
Eget initiativtagande och ansvar
På en finländsk arbetsplats övervakar chefen inte de anställdas arbete hela tiden.
Arbetstagarna tillfrågas om sina åsikter och åsikterna beaktas i planeringen av arbetet.
Man kommer överens om utförandet av arbetet på gemensamma möten och alla håller fast vid det man kommit överens om.
Chefen ger den anställda arbetsuppgifter och förväntar sig att den anställda själv fattar beslut om detaljerna i arbetets utförande.
Om den anställda inte kan eller förmår utföra arbetsuppgiften som anvisats, går han eller hon själv till andra anställda eller chefen för att be om råd.
Pålitlighet och att hålla tidtabeller
I den finländska arbetskulturen är det viktigt att hålla fast vid överenskommelser.
När man har beslutat något tillsammans förväntar sig både de anställda och arbetsgivaren att alla gör det man kommit överens om.
I Finland är det också viktigt att man håller fast vid tider.
Man kommer punktligt till arbetet på den avtalade tiden.
Klockan 8.00 betyder prick klockan 8.00, inte klockan 8.10.
Det är oartigt att komma för sent eftersom de andra då tvingas vänta på den som är försenad.
Om du vet att du kommer att bli sen till arbetet ska du tala om det för din chef.
På många arbetsplatser har man flexibel arbetstid och man kan komma till arbetet till exempel mellan klockan 7 och 9 och gå hem mellan klockan 15 och 17.
Om man har flexibel arbetstid ska den anställda själv se till att han eller hon arbetar den tid som avtalats.
Kommunikationsstil
Finländarna är ofta rakt på sak och frispråkighet upplevs inte som något oartigt.
Rättframhet är också vanligt i arbetslivet.
Om man till exempel inte har tillräckligt med tid för att göra en arbetsuppgift, är det bra att säga det uppriktigt till chefen.
På möten och vid diskussioner är det vanligt att man går rakt på sak genast efter att man hälsat på varandra.
I den finländska arbetskulturen tilltalar man varandra på ett mycket informellt sätt.
På de flesta arbetsplatserna duar alla varandra oberoende av sin ställning.
Religionens påverkan på arbetslivet
Många finländare är kristna men inte speciellt religiösa.
I den finländska kulturen följs dock fortfarande många kristna seder.
I arbetslivet syns religionens inflytande i de många lediga dagarna som anställda får.
Under de kristna helgerna, såsom på jul och påsk, har man lagstadgade lediga dagar.
Läs mer om högtidsdagarna på InfoFinlands sida Finländska helgdagar.
Religiösa seder eller ritualer hör inte hemma på den finländska arbetsplatsen.
På vissa arbetsplatser har man ordnat en plats för bön om de anställda framfört önskemål om det.
Sådan praxis är dock ovanlig på arbetsplatser.
Om en anställd till exempel vill hålla en bönestund under arbetsdagen ska detta göras under de avtalade pauserna.
Yttre religiösa symboler, såsom huvuddukar, är tillåtna i Finland, men de klädregler som gäller på arbetsplatserna måste följas.
Orsaken till detta är arbetssäkerhets- och hygienföreskrifter som anknyter till arbetsuppgifterna.
Du kan läsa mer om värderingar och seder i det finländska samhället på sidan Finländska seder.
Tvåspråkiga kommuner i Finland
Finland har två officiella språk, finska och svenska.
Finska är modersmålet för cirka 90 procent av finländarna.
Svenska är modersmålet för cirka 5 procent av finländarna.
Svenska talas mest på Finlands väst- och sydkust.
Svenskan som talas i Finland är finlandssvenska.
Uttalet skiljer sig något från svenskan i Sverige.
Om du vill ansöka om finskt medborgarskap behöver du ett intyg över tillräckliga kunskaper i finska eller svenska.
Läs mer på InfoFinlands sida Officiellt intyg över språkkunskaper.
Du kan använda svenska med statliga myndigheter, till exempel FPA eller TE-byrån.
Ange ditt kontaktspråk till magistraten när du registrerar dig som invånare.
Du kan även ändra kontaktspråket senare.
Kommunerna i Finland kan vara antingen enspråkiga eller tvåspråkiga.
De flesta kommunerna i Finland är finskspråkiga.
Tvåspråkiga kommuner finns på väst- och sydkusten.
Om din hemkommun är tvåspråkig, kan du använda svenska även inom de kommunala tjänsterna, till exempel på hälsostationen.
linkkiKommuner.net:
Svenskspråkiga och tvåspråkiga kommunerfinska _ svenska
Integration på svenska kan vara ett bra alternativ för dig till exempel om:
Du bor i ett område med många svensktalande.
Du har svenskspråkiga familjemedlemmar eller släktingar.
Du kan lite svenska redan.
Det kan vara fördelaktigt att kunna svenska när du söker jobb.
Tänk ändå på att kunskaper i finska krävs på de flesta arbetsplatserna.
Även om du väljer integrationsutbildning på svenska lönar det sig för dig att i något skede även lära dig finska.
I en del kommuner kan du delta i integrationsutbildning på svenska.
Om du inte blir antagen till integrationsutbildning på svenska kan du i vissa fall få stöd för frivilliga studier i svenska, om detta överenskommits i din integrations- eller sysselsättningsplan.
Fråga om integration på svenska när din inledande kartläggning och integrationsplan görs.
Enligt lag har du rätt att välja antingen finska eller svenska som integrationsspråk.
linkkiArbets- och näringsministeriet:
Information om integration på svenskafinska _ svenska
Språkstudier som arbetskraftsutbildning
Om du är kund vid arbets- och näringsbyrån kan du också studera svenska som arbetskraftsutbildning.
Arbetskraftsutbildningen är avsedd för arbetslösa arbetssökande.
Läs på InfoFinlands sida Arbets- och näringsbyråns tjänster vad som krävs för att du ska kunna bli kund hos arbets- och näringsbyrån.
Arbetskraftsutbildningen är kostnadsfri för dig.
Fråga mer om kurser i svenska vid din egen arbets- och näringsbyrå.
Barndagvård och utbildning för barn
I Finland ges dagvård, förskoleundervisning och grundläggande utbildning vanligtvis på finska eller svenska.
Om du vill att ditt barn ska börja i svenskspråkig dagvård, förskola eller skola, fråga om möjligheterna i din hemkommun.
Vissa kommuner ordnar förberedande undervisning före den grundläggande utbildningen för elever som ännu inte har tillräckligt bra språkkunskaper för den vanliga undervisningen.
Fråga i din hemkommun om förberedande undervisning ordnas på svenska i kommunen.
Om barnet har något annat modersmål än finska eller svenska, kan kommunen ordna undervisning i barnets eget modersmål för barnet.
Om barnet går i en svensk skola kan hen läsa svenska som andra språk.
Läs mer om barndagvård, förskoleundervisning och grundläggande utbildning på InfoFinlands sida Utbildning för barn.
Gymnasium och yrkesläroanstalt
Efter grundskolan kan du studera på gymnasiet eller en yrkesläroanstalt.
Svenskspråkiga yrkesläroanstalter och gymnasieskolor finns i svenskspråkiga och tvåspråkiga kommuner och i en del finskspråkiga kommuner.
Vissa yrkesläroanstalter och gymnasieskolor ordnar förberedande utbildning före studierna.
I den förberedande utbildningen får du sådana kunskaper och färdigheter som du behöver i dina fortsatta studier.
Du kan också förbättra dina språkkunskaper.
Du kan söka svenskspråkig yrkes- och gymnasieutbildning samt förberedande utbildning före dessa via tjänsten Opintopolku.fi.
Läs mer på InfoFinlands sida: Efter grundskolan.
Grundläggande information om yrkesutbildningfinska _ svenska _ engelska
Information om gymnasiestudierfinska _ svenska
Högskoleutbildning
I Finland finns svenskspråkiga yrkeshögskolor och universitet.
Dessutom finns det några tvåspråkiga universitet där du kan läsa på svenska.
Du kan söka svenskspråkiga högskoleutbildningar via tjänsten Opintopolku.fi.
Läs mer om högskoleutbildning på InfoFinlands sida: Högskoleutbildning.
Information om högskolestudierfinska _ svenska _ engelska
Var kan jag läsa svenska?
Du kan läsa svenska till exempel vid medborgarinstitut, arbetarinstitut och sommaruniversitet.
Fråga om studier i svenska hos utbildningsväsendet i din hemkommun, studievägledarna vid läroanstalter eller rådgivningstjänsterna för invandrare.
Läs mer på InfoFinlands sida: Studier som hobby.
Svenska på internet
Appar
Du kan lära dig svenska med hjälp av appar som du kan ladda ned i din telefon eller surfplatta.
Sök appar för svenska i din appbutik (t.ex. Google Play och App Store) med sökorden ”learn Swedish”, ”Swedish language”, ”lär dig svenska” eller ”svenska”.
En del appar kostar pengar.
Övningar och kurser på internet
På internet hittar du kurser i det svenska språket på olika nivåer.
På internet kan du till exempel göra övningar och spela spel, lära dig grammatik och vokabulär samt läsa texter.
linkkiYle:
Övningar för allmänna språkexaminafinska
Svenska på internetfinska _ svenska _ engelska
linkkiYle.fi:
Övningar och kurser på internetfinska
linkkiBab.la:
Flerspråkiga ordböckerfinska _ svenska _ engelska
I Finland finns många möjligheter att studera finska.
Olika kurser ordnas för både barn och vuxna.
Undervisning i finska för vuxna
Du hittar information om kurser i finska till exempel hos medborgarinstitut, arbetarinstitut, universitet och sommaruniversitet.
Fråga mer vid rådgivningstjänsterna för invandrare, utbildningsväsendet i din hemkommun eller studievägledarna vid lokala läroanstalter.
På vissa orter har informationen om kurserna samlats på ett och samma ställe.
Till exempel finns det information om kurserna i finska språket i Helsingfors, Tammerfors och Åbo i tjänsten Finnishcourses.fi.
Vid läroanstalterna börjar kurserna vanligtvis i augusti eller september och i januari.
Språkkurserna är ofta fullsatta.
Därför är det viktigt att anmäla sig till kursen i god tid.
Medborgarinstitut i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Kurser i finska och svenska språketfinska _ engelska _ ryska
Språkstudier i anslutning till annan utbildning
Du kan studera finska också i arbetskraftsutbildning och i förberedande utbildning före yrkesutbildning (VALMA) eller förberedande gymnasieutbildning (LUVA).
Om du är kund vid arbets- och näringsbyrån kan du få plats på en kurs i finska via arbets- och näringsbyrån.
Hurdan språkundervisning du behöver bedöms på arbets- och näringsbyrån i samband med att du får en integrations- eller sysselsättningsplan.
Du kan studera finska som arbetskraftsutbildning.
Arbetskraftsutbildning är i huvudsak utbildning avsedd för arbetslösa arbetssökande.
Utbildningen är kostnadsfri för deltagarna.
Fråga om kurserna i finska på din egen arbets- och näringsbyrå.
linkkiArbets- och näringsministeriet:
Kontaktuppgifter till TE-byråerfinska _ svenska
linkkiArbets- och näringsministeriet:
Utbildning i finska och svenska språketfinska _ svenska _ engelska
Finska på arbetsplatsen
Vissa arbetsgivare ordnar finskundervisning för sina arbetstagare.
Fråga din arbetsgivare om du kan studera finska på din arbetsplats.
Arbetsgivaren kan ansöka om stöd för arbetstagarnas finskundervisning via arbets- och näringslivstjänsterna.
linkkiTE-tjänster:
Finska på arbetsplatsenfinska _ svenska _ engelska
Undervisning i finska för barn
Barn lär sig nya språk snabbt, även om det kan kännas svårt i början.
Finskundervisning ges på daghem, i förskola och skola.
Undervisningen kallas finska som andra språk eller S2-undervisning.
Barnet eller den unga kan även delta i förberedande undervisning.
Den är avsedd för de elever som ännu inte har särskilt bra kunskaper i finska.
Under den förberedande undervisningen studerar barnet eller den unga finska och några läroämnen.
Den förberedande undervisningen är avsedd för 7–16-åringar.
Undervisningen varar vanligtvis ett år.
Därefter flyttas eleven till en vanlig klass.
linkkiEdu.fi:
Finska som andra språk i den grundläggande undervisningenfinska
I Finland finns två pensionssystem som kompletterar varandra:
Arbetspensionen intjänas med det egna lönearbetet och företagandet.
Arbetsgivaren är skyldig att teckna pensionsförsäkring åt alla sina anställda och betala försäkringspremierna.
Privatföretagare sköter sina premier själva.
Folkpensionen och garantipensionen är avsedda för de pensionärer som inte får arbetspension eller vars pension är mycket liten.
Båda pensionssystemen omfattar ålderspension och invalidpension.
Du kan få folkpension när du har fyllt 65 år.
Ditt födelseår avgör i vilken ålder du kan få arbetspension.
Kontrollera din pensionsålder på ditt arbetspensionsutdrag eller hos din arbetspensionsanstalt.
Om man är arbetsoförmögen kan man få invalidpension före ålderspensionen.
Om man vill kan man också arbeta när man är pensionerad.
Om du är i ålderspension påverkar din arbetsinkomst inte pensionens storlek.
I Finland betalas skatt på pensionerna.
Arbetsgivarna och arbetstagarna finansierar pensionsskyddet tillsammans.
Arbetsgivaren drar av arbetstagarens andel från lönen och betalar den och sin egen andel av försäkringspremierna till pensionsanstalten.
Arbetspensionens belopp beror på hur länge du har arbetat och hur stor lön du har haft.
Arbetspensionsförsäkringsbolag, pensionskassor och -stiftelser har hand om arbetspensionsförsäkringarna.
Pensionsskyddscentralen sköter centraliserat frågor som rör pensionsskyddet.
linkkiPensionsskyddscentralen:
Arbetspensionfinska _ svenska _ engelska
Kontrollera på arbetspensionsutdraget hur stor pension du tjänat in
Din pensionsanstalt skickar regelbundet ett arbetspensionsutdrag till dig.
På arbetspensionsutdraget finns en uppskattning av din intjänade pension.
Du kan också beställa ett arbetspensionsutdrag från din pensionsanstalt eller Pensionsskyddscentralen.
Genom att själv följa med arbetspensionsutdragen kan du kontrollera att din intjänade pension räknats rätt.
Om det finns fel i uppgifterna, kontakta ditt pensionsbolag eller Pensionsskyddscentralen.
Spara arbetsintyg för eventuella granskningar.
Det är också bra att spara lönekvitton.
Att beställa ett arbetspensionsutdragfinska _ svenska _ engelska _ ryska _ estniska
Du kan ansöka om folkpension om du inte har någon arbetspension eller om din arbetspension är väldigt liten. Folkpensionens belopp beror på hur länge du har bott eller arbetat i Finland.
Dina familjeförhållanden och andra kontinuerliga pensionsinkomster påverkar också folkpensionens belopp.
FPA sköter folkpensionerna och garantipensionerna.
Du kan söka folkpension och garantipension om du omfattas av Finländska socialskyddet och när du har bott i Finland minst tre år efter att du fyllde 16 år.
Också den tid som du har varit bosatt i något annat EU- eller EES-land kan delvis beaktas.
Garantipensionen tryggar ett existensminimum för pensionärer.
Garantipensionens belopp är mellanskillnaden mellan de övriga pensionerna som du får och garantipensionens fulla belopp.
Om det sammanlagda beloppet från dina övriga pensioner överskrider garantipensionens fulla belopp kan du inte få garantipension.
Mer information om garantipensionen får du vid FPA.
I vissa fall kan du få folkpension även innan du fyllt 65 år.
FPA ger mer information om förtida ålderspension och tilläggsdagar till folkpension.
linkkiPensionsskyddscentralen:
Pensionssystemet i Finlandfinska _ svenska _ engelska
Stöden för pensionärerfinska _ svenska _ engelska
Information om frågor som rör pensionfinska _ svenska _ engelska _ ryska _ estniska
Att söka pension
Alla pensioner måste sökas.
Du kan ansöka om arbets- och folkpension med samma blankett.
Du kan fylla i blanketten på nätet eller lämna in den till FPA, folkpensionsverket eller Pensionskyddscentralen.
Blanketterna finns på verksamhetsställena och på internet.
Du kan ansöka om garantipensioni FPA:s nättjänst eller på kontoret.
Du kan ansöka om FPA:s åldringspension och garantipension även per telefon.
Numret till FPA:s pensionsärenden är 020 692 202.
Pension från utlandet
Om du har bott eller arbetat i andra EU-länder än Finland eller i något land med vilket Finland har ett socialskyddsavtal, kan du ha rätt till pension från dessa länder.
Du kan ansöka om pension från dessa länder samtidigt som du ansöker om den finländska arbets- eller folkpensionen.
Bifoga till din ansökan blanketten Boende och arbete utomlands.
Du kan skriva ut blanketten på FPA:s eller Pensionsskyddscentralens webbplats.
Om du har arbetat i andra länder som Finland inte har ett socialskyddsavtal med, måste du själv ta reda på om du har rätt att få pension från dessa länder.
Om du kan få pension, måste du själv ansöka om den.
Om du ansöker om pension från utlandet, får du råd vid Pensionsskyddscentralen.
Läs mer på Pensionsskyddscentralens webbplats.
Du kan även fråga om råd hos FPA.
linkkiPensionsskyddscentralen:
Broschyren Att söka pension från utlandetfinska _ svenska _ engelska _ ryska _ estniska
Utbetalning av pension till utlandet
Arbetspension utomlands
Om du flyttar från Finland utbetalas arbetspension från Finland då du går i pension.
Pensionen kan utbetalas till vilket land som helst.
Det är viktigt att du har ett arbetsintyg från alla anställningar i Finland.
Det är också bra att spara lönekvitton.
Hur du ansöker om pension till utlandet beror på i vilket land du bor.
Du kan fråga din pensionsanstalt eller Pensionsskyddscentralen om råd.
Innan du ansöker om pension ska du begära ett arbetspensionsutdrag av din pensionsanstalt eller Pensionsskyddscentralen.
Arbetspensionsutdraget visar hur stor pension du tjänat in i Finland.
FPA:s pensioner utomlands
Du ska alltid meddela FPA om varaktig flytt utomlands eller vistelse utomlands som varar över tre månader.
Om du vistas utomlands tillfälligt, det vill säga under ett år, betalar FPA vanligtvis din pension som vanligt.
I vissa fall betalar FPA till exempel ålderspension och familjepension till vissa länder även då du flyttar till landet för över ett år.
Sådana länder är till exempel de övriga EU-länderna och EES-länderna samt en del av de länder som Finland har ett socialskyddsavtal med.
Garantipensionen betalas inte om du flyttar utomlands för över ett år.
På FPA:s webbplats finns information om i vilka fall du kan få FPA:s pensioner utomlands.
Du kan också fråga om din egen situation vid FPA:s kontor eller telefontjänst.
Partiell förtida ålderspension
Om du har fyllt 61 år kan du få partiell pension redan före din lägsta ålderspensionsålder.
Detta kallas partiell förtida ålderspension.
Du kan själv välja om du vill ta ut 25 procent eller 50 procent av beloppet på din månatliga arbetspension.
Om du vill kan du samtidigt fortsätta arbeta heltid eller komma överens om en kortare arbetstid med arbetsgivaren.
Du kan också sluta arbeta.
Du bör observera att den partiella förtida ålderspensionen permanent minskar beloppet på den slutliga ålderspensionen.
Du kan fråga mer av din pensionsanstalt.
Om du är sjuk under en längre tid får du vanligtvis först under ungefär ett års tid sjukdagpenning.
Om du inte kan återgå till arbetet på grund av sjukdom eller skada kan du ansöka om invaliditetspension (työkyvyttömyyseläke) eller rehabiliteringsstöd (kuntoutustuki).
Rehabiliteringsstöd är invaliditetspension på viss tid.
Du kan ansöka om invaliditetspension med en blankett som du får från FPA.Som bilaga till ansökan krävs B-utlåtande av läkare.
FPA och arbetspensionsanstalten bedömer din arbetsförmåga och om du har nytta av rehabilitering.
Mer information om invaliditetspension och rehabilitering får du av FPA, din pensionsanstalt eller av företagshälsovården.
Om du får invaliditetspension påverkar din lönenivå pensionen.
Du ska meddela FPA och arbetspensionsanstalten om du börjar arbeta.
Om du har en tillräckligt hög inkomst från arbetet per månad kan du låta din pension vila.
Detta innebär att du håller en paus i lyftandet av pensionen.
Pausen kan vara minst tre månader och högst två år lång.
Under denna tid förlorar du inte rätten till invaliditetspension.
Övriga förmåner för pensionärer
Utöver pension kan FPA betala ut bostadsbidrag till pensionstagare med låga inkomster.
Mer information om bostadsbidrag för pensionstagare hittar du på FPA:s webbplats.
Till långtidssjuka eller handikappade kan FPA betala ut vårdbidrag för pensionstagare.
Fråga mer på FPA.
Rabatter för pensionärer
När du har pensionerats kan du få pensionärsrabatt till exempel på tåg-, buss- och flygresor i Finland.
De som fyllt 65 år får reserabatt genom att uppvisa sitt identitetsbevis.
En pensionär som inte har fyllt 65 år kan få rabatt genom att uppvisa sitt personbevis och sitt arbetspensionskort eller folkpensionärskort.
Kontrollera villkoren för pensionärsrabatten på biljettkontoren.
Du kan även få rabatt på exempelvis olika former av motion och kultur.
Om du vill ansöka om finskt medborgarskap behöver du ett officiellt intyg över dina kunskaper i finska eller svenska.
Du kan behöva intyget också när du söker ett jobb eller en studieplats.
Du kan påvisa dina språkkunskaper:
med en allmän språkexamen (yleinen kielitutkinto)
med vitsordet i finska eller svenska på ditt avgångsbetyg (päättötodistus).
Allmän språkexamen
Allmän språkexamen, ASE, är ett språktest för vuxna.
Med en allmän språkexamen kan du påvisa dina kunskaper i finska eller svenska.
Examen är avgiftsbelagd.
När du avlagt examen får du ett intyg som anger nivån på dina språkkunskaper.
Språkexamen finns på tre olika nivåer: grundnivån, mellannivån och högsta nivån.
Varje examensnivå består av två färdighetsnivåer, vilka det alltså finns sammanlagt sex av.
Grundnivån är avsedd för personer som kan använda språket i vardagliga sammanhang.
Deras färdighetsnivå är 1–2.
Medelnivån är avsedd för personer som kan språket relativt väl. Deras färdighetsnivå är 3–4.
Den högsta nivån är avsedd för personer som kan språket mycket väl. Deras färdighetsnivå är 5–6.
Närmare beskrivningar av de olika färdighetsnivåerna finns på Utbildningsstyrelsens webbplats.
Om du vill ansöka om finskt medborgarskap (kansalaisuus) kan du påvisa att du har tillräckliga kunskaper i finska eller svenska genom att avlägga den muntliga och skriftliga delen av en allmän språkexamen minst på nivå 3.
Språkexamenstillfället pågår 3–6 timmar.
Uppgifternas ämnesområden rör det vardagliga livet såsom fritid, utbildning och vanliga situationer på arbetet.
I examen ingår olika uppgifter där följande färdigheter krävs:
textförståelse
skriftliga färdigheter
grammatik och vokabulär
talförståelse
muntliga färdigheter
Du kan avlägga examen på olika orter i Finland.
Mer information om anmälan får du på Utbildningsstyrelsens (Opetushallitus) webbplats.
Examina kategoriseras på en annan skala än kurserna.
Om du har slutfört en språkkurs som kategoriserats enligt den europeiska referensramen motsvarar kursen nivån på den allmänna språkexamen ungefär enligt följande tabell:
A1 – ASE 1
A2 – ASE 2
B1 – ASE 3
B2 – ASE 4
C1 – ASE 5
C2 – ASE 6
Innan du anmäler dig till examen ska du göra dig förtrogen med kraven på de olika examensnivåerna.
Du kan även fråga din lärare i finska.
Mer information om den allmänna språkexamen får du på Utbildningsstyrelsens webbplats.
linkkiUtbildningsstyrelsen:
Allmänna språkexaminafinska _ svenska _ engelska
linkkiUtbildningsstyrelsen:
Färdighetsnivåerna i allmänna språkexaminafinska _ svenska _ engelska
linkkiUtbildningsstyrelsen:
Att anmäla sig till en allmän språkexamen och examensavgifterfinska _ svenska _ engelska
Statsförvaltningens språkexamen om kunskaper i finska och svenska
Om du vill arbeta inom den offentliga förvaltningen behöver du vanligtvis ett intyg över dina kunskaper i finska eller svenska.
Du kan påvisa dina kunskaper i finska eller svenska med statsförvaltningens språkexamen.
Fråga din arbetsgivare hurdana språkkunskapskrav som gäller på den arbetsplats som du vill söka.
Språkexamen finns på tre olika nivåer: för nöjaktiga, goda och utmärkta språkkunskaper.
Det beror på din arbets- eller studieplats vilken examensnivå du måste avlägga.
För finskt medborgarskap behöver du ett intyg för åtminstone nöjaktiga språkkunskaper.
Du kan avlägga examen för nöjaktiga eller goda språkkunskaper olika orter i Finland.
På Utbildningsstyrelsens webbplats hittar du en förteckning över de städer där examen kan avläggas.
Examen på utmärkt nivå kan endast avläggas i Helsingfors.
Examen omfattar olika tester. I dem ska du läsa och lyssna på texter och svara på frågor.
Därtill finns det intervjuer, diskussioner och skriftliga uppgifter.
Du kan ersätta statsförvaltningens språkexamen med vissa andra studier.
Till exempel motsvarar statsförvaltningens språkexamen som gäller goda språkkunskaper ett mognadsprov (kypsyysnäyte) som du har avlagt på finska eller svenska vid universitetet.
Mer information får du på Utbildningsstyrelsens webbplats.
linkkiUtbildningsstyrelsen:
Statsförvaltningens språkexaminafinska _ svenska
linkkiUtbildningsstyrelsen:
Färdighetsnivåerna i statsförvaltningens språkexaminafinska _ svenska
linkkiUtbildningsstyrelsen:
Mottagare av statsförvaltningens språkexamina, finska språketfinska _ svenska
linkkiUtbildningsstyrelsen:
Mottagare av statsförvaltningens språkexamina, svenska språketfinska _ svenska
Intyg över språkkunskaper på basis av studier
Om du vill ansöka om finskt medborgarskap kan du påvisa dina kunskaper i finska eller svenska även med något av följande intyg:
avgångsbetyg från grundskolan med ett godkänt vitsord i finska eller svenska som modersmål eller som andra språk
avgångsbetyg från gymnasiet med ett godkänt vitsord i finska eller svenska som modersmål eller som andra språk
studentexamen på finska eller svenska med ett godkänt vitsord i finska eller svenska som modersmål eller som andra språk
intyg på yrkesinriktad grundexamen som du har avlagt på finska eller svenska
intyg på yrkesexamen som du har avlagt på finska eller svenska
intyg på studier i tjänstemannafinska eller -svenska som du har avlagt vid universitet eller högskola
intyg på mognadsprov som du har avlagt på finska eller svenska för universitetsexamen eller yrkeshögskoleexamen
Mer information får du på Migrationsverkets (Maahanmuuttovirasto) webbplats.
linkkiUtbildningsstyrelsen:
Språkkunskaper och finskt medborgarskapfinska _ svenska _ engelska
Ungefär 90 procent av finländarna har finska som modersmål.
Ungefär fem procent av finländarna har svenska som modersmål.
När du funderar på om det är finska eller svenska som du borde lära dig ska du beakta vilket språk som talas på din hemort och i din näromgivning.
Om du vill ansöka om finskt medborgarskap måste du kunna finska, svenska eller i det finska teckenspråket.
När du ansöker om medborgarskap, bifoga ett intyg över dina språkkunskaper.
Läs mer om språkkunskapskraven på InfoFinlands sida Officiellt intyg över språkkunskaper.
På de flesta arbetsplatser är det nödvändigt att kunna finska.
Om du vill studera i Finland behöver du sannolikt kunna finska.
Det kan vara bra att lära sig finska eller svenska trots att du inte tänker bo en lång tid i landet.
Även om finländarna i allmänhet behärskar engelska relativt väl har du ändå mycket nytta av att kunna finska eller svenska.
När du behärskar språket är det lättare för dig att trivas i landet och anpassa dig till livet i Finland.
Du har lättare att sköta dina ärenden med myndigheter, följa nyheter, få nya bekantskaper och vänner.
Du lär dig språket bäst om du vågar använda det.
Du behöver inte alltid förstå allting, det räcker med att du förstår det viktigaste.
Dra dig alltså inte för situationer där du har möjlighet att tala finska eller svenska.
Information om språklagenfinska _ svenska _ engelska
linkkiKommuner.net:
Svenskspråkiga och tvåspråkiga kommunerfinska _ svenska
Vem är berättigad till utkomstskydd för arbetslösa?
Du kan registrera dig som arbetssökande vid TE-byrån om
du har ett uppehållstillstånd som ger dig rätt att arbeta i Finland
ditt uppehållstillstånd inte begränsar vilken arbetsgivare du får arbeta för
eller
du är medborgare i ett EU-land, ett EES-land eller Schweiz
du är familjemedlem till en medborgare i ett EU-land, ett EES-land eller Schweiz
Då du registrerat dig som arbetssökande har du rätt till arbetslöshetsunderstöd om du
är 17–64 år gammal
är arbetslös och anmäld som arbetssökande vid TE-byrån
söker heltidsarbete
är arbetsförmögen och tillgänglig på arbetsmarknaden
uppfyller villkoren för inkomstrelaterad dagpenning, grunddagpenning eller arbetsmarknadsstöd.
För att få utkomstskydd för arbetslösa måste du aktivt söka jobb och vara beredd att ta emot ett jobb.
Du ska också ingå en sysselsättnings- och integrationsplan med TE-byrån och delta i de tjänster och åtgärder som TE-byrån erbjuder åt dig.
På full arbetslöshetsförmån ställs även andra villkor.
Du kan få full arbetslöshetsförmån om du under 65 betalningsdagar, alltså under cirka tre månaders tid, utför en viss mängd lönearbete, får inkomst som företagare eller deltar i en verksamhet eller en tjänst som främjar din sysselsättning.
Detta kallas för aktiveringsmodellen för arbetslöshetsförsäkringen (työttömyysturvan aktiivimalli).
Arbetslöshetsförmånerna är den inkomstrelaterade dagpenningen, grunddagpenningen och arbetsmarknadsstödet.
Skatt betalas på alla arbetslöshetsförmåner.
linkkiArbets- och näringsministeriet:
Om du blir arbetslösfinska _ svenska _ engelska
linkkiArbets- och näringsministeriet:
Utkomstskydd för arbetslösafinska _ svenska _ engelska
Information om utkomstskyddet för arbetslösafinska _ svenska _ engelska
linkkiArbets- och näringsministeriet:
Rådgivning om utkomstskydd för arbetslösafinska _ svenska _ engelska _ ryska
Aktiveringsmodellen för arbetslöshetsförsäkringen finska _ svenska _ engelska
Inkomstrelaterad dagpenning
Du kan få inkomstrelaterad dagpenning om du
registrerat dig som arbetslös arbetssökande vid arbets- och näringsbyrån
hör till en finländsk arbetslöshetskassa
uppfyller arbetsvillkoret, d.v.s. har arbetat tillräckligt länge före arbetslösheten
har varit medlem i arbetslöshetskassan i minst 26 veckor innan du blev arbetslös.
Den inkomstrelaterade dagpenningen beviljas och utbetalas av den arbetslöshetskassa där du är medlem.
Den inkomstrelaterade dagpenningen beräknas utgående från storleken på den lön som du hade innan du blev arbetslös.
Vanligtvis kan inkomstrelaterad dagpenning fås under 400 dagar. Undantag från detta är följande situationer:
Om du har arbetat i sammanlagt tre år eller mindre, kan du få inkomstrelaterad dagpenning i högst 300 dagar.
Om du har fyllt 58 år innan du blev arbetslös, kan du få inkomstrelaterad dagpenning i mindre än 500 dagar.
Läs mer om arbetslöshetskassan på InfoFinlands sida Fackförbund.
Information om den inkomstrelaterade dagpenningenfinska _ svenska _ engelska
Grunddagpenning
Du kan få grunddagpenning om du omfattas av den sociala tryggheten i Finland utifrån permanent boende eller arbete före arbetslösheten och
registrerat dig som arbetslös arbetssökande vid arbets- och näringsbyrån
uppfyller arbetsvillkoret, d.v.s. har arbetat tillräckligt länge före arbetslösheten
inte uppfyller villkoren för inkomstrelaterad dagpenning.
Grunddagpenningen beviljas och utbetalas av Fpa.
Vanligtvis kan du få grunddagpenning i mindre än 400 dagar. Undantag från detta är följande situationer:
Om du har arbetat i sammanlagt tre år eller mindre, kan du få grunddagpenning i högst 300 dagar.
Om du har fyllt 58 år innan du blev arbetslös, kan du få grunddagpenning i mindre än 500 dagar.
Om du får andra sociala förmåner eller arbetsinkomster under arbetslösheten, är din grunddagpenning mindre.
Grunddagpenningfinska _ svenska _ engelska
Arbetsmarknadsstöd
Du kan få arbetsmarknadsstöd om du
registrerat dig som arbetslös arbetssökande vid arbets- och näringsbyrån
bor permanent i Finland
inte uppfyller arbetsvillkoret, d.v.s. inte arbetat tillräckligt länge innan du blev arbetslös eller fått förvärvsrelaterad dagpenning eller grunddagpenning under maximitiden.
Om du har en gällande integrationsplan, kan du söka arbetsmarknadsstöd för den tid då du deltar i utbildningar och annan verksamhet som nedtecknats i planen.
Närmare uppgifter om integrationsplanen finns på InfoFinlands sida Integration i Finland.
Arbetsmarknadsstödet beviljas och utbetalas av Fpa.
Arbetsmarknadsstödet är behovsprövat.
Det betyder att till exempel sociala förmåner och lön minskar arbetsmarknadsstödets belopp.
Om du är under 25 år, kontrollera tilläggsvillkoren för arbetsmarknadsstödet för unga på TE-tjänsternas webbplats.
Arbetsmarknadsstödfinska _ svenska _ engelska
På nätet hittar du finskakurser på många olika nivåer.
På nätet kan du till exempel göra övningar, spela spel, lära dig grammatik och vokabulär och läsa texter.
De flesta webbkurser är på finska eller svenska, men det finns även andra alternativ:
Nybörjarnivån
linkkiYle:
Nybörjarkurs i finska, Easyfinnishfinska
Nybörjarkurs i finska "A Taste of Finnish"engelska
linkkiTammerfors yrkeshögskola:
Nybörjarkurs i finska, Uunofinska
Nybörjarkurs i finska, Tavataan taasengelska _ franska _ tyska _ bulgariska
Nybörjarkurs i finskafinska _ svenska _ engelska _ arabiska
linkkiWordDive:
Nybörjarkurs i finskafinska _ svenska _ engelska _ ryska _ kinesiska _ tyska
Inledningskurs i finskaengelska
Tilläggsövningar till läroboken Hyvin meneefinska
Mångsidiga övningar i finska språketfinska
Ordspel för nybörjareengelska _ franska _ japanska
Applikationen Suomipassi med flera stödspråkfinska _ engelska
Grundnivån
linkkiYle:
Övningar för allmänna språkexaminafinska
Webbkurs med många hjälpspråksvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ portugisiska
linkkiEdu.fi:
Vardagsfinska: videoinspelning med intervjuerfinska
Vokabulärövningarfinska
linkkiYle:
Läromaterial från TV-serien Supisuomeafinska
linkkiUtbildningsstyrelsen:
Finska i arbetslivetfinska
Mångsidiga övningar i finska språketfinska
Lär dig finska med hjälp av filmerfinska _ engelska _ persiska _ arabiska
Självständiga språkanvändare
linkkiYle:
Nyheter på klarspråkfinska
Information om olika ämnen på klarspråkfinska
Nyheter på lättläst finskafinska
linkkiUtbildningsstyrelsen:
linkkiUtbildningsstyrelsen:
Finska i arbetslivetfinska
Avancerade språkanvändare
Lyssna på finska dialekterfinska
linkkiWordDive:
Finskans grammatikfinska _ svenska _ engelska _ ryska _ spanska _ tyska _ japanska
Finskans grammatikengelska
Finskans grammatikengelska
Verbböjningengelska
linkkiInstitutet för de inhemska språken:
Grammatiken Iso suomen kielioppi på nätetfinska
Information om finska språketengelska
Ordböcker på nätet
Flerspråkiga ordböckerfinska
linkkiBab.la:
Flerspråkiga ordböckerfinska _ svenska _ engelska
Intern kommunikation på arbetsplatsen
Vanligen informerar man om kommande händelser och ändringar på arbetsplatsen vid möten.
Om man deltar i möten kan man påverka, föreslå ändringar och utveckla sitt eget arbete.
På varje arbetsplats finns också andra kanaler för den interna kommunikationen, såsom anslagstavlor, e-post eller de anställdas postfack.
Följ informationen på arbetsplatsen.
Pauser
I arbetsavtalet står det ofta hur långa pauser som ingår i arbetsdagen och tidpunkten för dessa.
Vanligen har man en kort kaffepaus på förmiddagen, en lunchpaus mitt på dagen och en kaffepaus till på eftermiddagen.
Längden på lunchpausen varierar mellan olika arbetsplatser.
Fråga din chef hur långa pauser du har.
Arbetsplatsbespisningen är ordnad på olika sätt på olika arbetsplatser: vissa arbetsplatser har en egen personalmatsal, på andra ställen tar de anställda med sig maten hemifrån.
På vissa arbetsplatser kan man köpa förmånliga lunchsedlar som man kan använda på matställen i närheten av arbetsplatsen.
Under lunchen arbetar man vanligtvis inte.
Att sköta egna ärenden under arbetsdagen
På arbetstid får man inte sköta sina privata angelägenheter, utan detta måste göras utanför arbetstiden.
Antalet arbetstimmar som står i arbetsavtalet är bindande och det avtalade antalet arbetstimmar ska fullgöras.
Under pauserna kan du till exempel ringa viktiga samtal.
Du kan också ansöka om oavlönad ledighet om din situation kräver att du är frånvarande en längre tid.
Om du av någon anledning inte till exempel lyckas få en läkartid utanför arbetstiden, ska du komma överens med din chef om att du är borta och hur du ersätter din frånvaro.
Företagshälsovården kan du besöka under arbetstid.
Utbildning som rör arbetet
Även om arbetstagaren har sådan utbildning som krävs för yrket redan när anställningen inleds, uppmuntrar många arbetsgivare sina anställda att skaffa sig mer utbildning.
Ofta kan du utbilda dig på arbetstid och arbetsgivaren kan betala för utbildningen.
De flesta arbetsgivare värdesätter att den anställda vill utveckla sig i sitt arbete och inhämta nya kunskaper.
Vanligen ger man inte varandra presenter på arbetsplatserna.
På viktiga bemärkelsedagar (födelsedagar, äktenskap, pensionering) uppmärksammar arbetskamraterna och arbetsgivaren festföremålet med en liten present eller en blombukett.
Arbetstid och semester
En normal arbetsdag är vanligtvis åtta timmar.
Arbetstagaren kan även komma överens om någon annan tid med arbetsgivaren.
I Finland gör arbetstagare vanligtvis inte mycket övertid.
Man arbetar de timmar som står i anställningsavtalet.
I Finland börjar semesterperioden i början av maj.
Antalet intjänade semesterdagar beror på anställningstiden i år och när anställningen har börjat.
Utöver den betalda semesterna kan du ansöka om obetald ledighet.
Jämfört med många andra länder har arbetstagare i Finland långa semestrar.
Arbetshälsa och rekreation
På många arbetsplatser vill man stödja de anställdas arbetsmotivation och -trivsel med olika rekreationsdagar och fester på arbetsplatsen. Arbetsgivaren kan också erbjuda sina anställda olika hobbymöjligheter vid sidan av arbetet.
Årliga helger
Vissa dagar är allmänna lediga dagar i Finland.
Till dem hör följande:
nyårsdagen 1.1
trettondagen 6.1
påsk: tidpunkten varierar, i mars-april
första maj 1.5
midsommarafton: i juni, alltid en fredag
självständighetsdagen 6.12
juldagen 25.12
annandag jul 26.12
Läs mer om dessa dagar på sidan Finländska helgdagar.
På vissa arbetsplatser, till exempel sjukhus, arbetar man även under helgerna.
För arbetet under helgerna betalas högre lön.
Kontrollera ersättningen i ditt kollektivavtal.
Anmäl dig som arbetslös arbetssökande
Om du blir arbetslös ska du anmäla dig hos TE-byrån senast den första dagen av din arbetslöshet.
Om du omfattas av den finländska sociala tryggheten kan du ansöka om arbetslöshetsstöd.
Du kan få arbetslöshetsstöd från och med det datum då du anmälde dig som arbetslös.
Kom ihåg att anmäla dig också direkt efter studier, arbetskraftsutbildning eller en period med sysselsättningsstöd.
Anmäl dig som arbetssökande i TE-byråns webbtjänst.
Logga in med finländska nätbankskoder eller personkort med microchip.
En anställd vid TE-byrån tar kontakt med dig om det behövs ytterligare uppgifter.
Du behöver inte ringa eller besöka TE-byrån om du inte uttryckligen ombes göra detta.
Om du saknar nätbankskoder eller personkort med microchip ska du anmäla dig som arbetssökande vid närmaste TE-byrå.
Endast medborgare i EU-länderna, Norge, Island, Liechtenstein och Schweiz kan anmäla sig som arbetssökande i webbtjänsten.
Om du är medborgare i ett annat land måste du besöka arbets- och näringsbyrån.
När du går till TE-byrån ska du ta med dig
alla dina arbetsintyg och studiebetyg
ditt pass där ditt uppehållstillstånd syns
TE-byrån undersöker uppgifterna som du lämnar.
Det finns vissa villkor för att få utkomstskydd för de arbetslösa och TE-byrån utreder om dessa villkor uppfylls i din situation.
Därefter ger TE-byrån ett utlåtande i ärendet till den instans som betalar förmånen, det vill säga till arbetslöshetskassan eller FPA.
Du kan fråga råd i ärenden som rör utkomstskyddet för arbetslösa vid din egen TE-byrå.
Du kan också ringa TE-tjänsternas rådgivning om utkomstskydd för arbetslösa:
på finska: 0295 020 701
på svenska: 0295 020 711
på engelska: 0295 030 713
på ryska: 0295 020 715
Läs också InfoFinlands sida:
Arbetslöshetsförsäkring
linkkiArbets- och näringsministeriet:
Om du blir arbetslösfinska _ svenska _ engelska
linkkiArbets- och näringsministeriet:
Att anmäla sig som arbetslös arbetssökandefinska _ svenska
linkkiArbets- och näringsministeriet:
Rådgivning om utkomstskydd för arbetslösafinska _ svenska _ engelska _ ryska
Semester, studier eller arbete under arbetslösheten
Om du börjar arbeta eller studera när du är arbetslös ska du meddela detta till TE-byrån.
Du får anvisningar om hur detta påverkar ditt utkomststöd för arbetslösa.
Om du reser i hemlandet eller utomlands ska du se till att du alltid kan nås.
Lämna till exempel ditt telefonnummer och din adress till TE-byrån och ange hur länge du ämnar vistas på resmålet.
Du kan ändå inte tacka nej till ett jobb som erbjuds till dig på grund av en utlandsresa.
Om du startar ett företag när du är arbetslös, kan du få arbetslöshetsförmån under de fyra första månaderna.
Karens
Du kan förlora din rätt till arbetslöshetsdagpenning för en viss tid om du själv har förorsakat arbetslösheten.
Du kan sättas i karens till exempel om:
du inte söker ett jobb som TE-byrån föreslår för dig
du inte tar emot ett jobb som erbjuds till dig
du säger upp dig från ditt jobb utan en godtagbar anledning
Karenstidens längd varierar från 15 dagar till 90 dagar.
Längden beror på orsaken till karensen.
I vissa fall kan du förlora rätten till utkomststöd för arbetslösa tillsvidare.
I Finland beskrivs språkkursernas nivåer på olika sätt.
Ofta använder man bedömningsskalan enligt den gemensamma europeiska referensramen (GER).
(Eurooppalainen viitekehys EVK) Denna skala omfattar följande nivåer:
nivåerna A1 och A2: grundläggande språkkunskaper (peruskielitaito)
nivåerna B1 och B2: en självständig språkanvändares språkkunskaper (itsenäisen kielenkäyttäjän kielitaito)
nivåerna C1 och C2: en avancerad språkanvändares språkkunskaper (taitavan kielenkäyttäjän kielitaito)
Dessa nivåer delas ytterligare in i undernivåer.
Till exempel omfattar nivå A1 kurserna A1.1, A1.2 och A1.3 och nivå A2 kurserna A2.1 och A2.2.
Mer information om hurdana kunskaper de olika nivåerna avser i praktiken får du på Utbildningsstyrelsens (Opetushallitus) webbplats.
Du kan också fråga direkt vid läroanstalterna.
I InfoFinland under rubriken Officiellt intyg över språkkunskaper får du information om hur du kan jämföra kursernas nivåer med nivån på den allmänna språkexamen (yleinen kielitutkinto).
linkkiUtbildningsstyrelsen:
Skala för beskrivning av språkkunskapsnivåer(pdf, 119,85 kb)finska
linkkiEuropass.eu:
Utvärdera nivån på din språkkunskapfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
I Finland värdesätts ärlighet, punktlighet och jämställdhet.
Det syns överallt i den finländska kulturen, även i arbetslivet.
På den här sidan finns mer information om den finländska arbetskulturen.
Lagar och avtal i arbetslivet
Arbetslivet i Finland styrs av många regler som arbetstagaren och arbetsgivaren måste följa.
I lagstiftningen och kollektivavtalen fastställs till exempel minimilöner, arbetstider, semester, lön under sjukskrivning och uppsägningsvillkor.
Ibland kan arbetsgivaren be arbetstagaren arbeta övertid.
Enligt lag ska arbetsgivaren betala högre lön för övertid.
Du kan även få ersättningen i form av ledighet.
Du har rätt att vägra övertidsarbete.
Information om arbetstagarnas rättigheter och skyldigheter i Finland hittar du på InfoFinlands sida Arbetstagarens rättigheter och skyldigheter.
linkkiFFC:
Arbetslivet i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ kinesiska _ arabiska
Lär dig finska eller svenska
Du kan utveckla dina språkkunskaper på kurser eller i arbetet.
Dra dig inte för att prata finska eller svenska med dina kollegor.
Läs mer om språkstudier i InfoFinlands avsnitt Finska och svenska språket.
Jämlikhet och jämställdhet i arbetslivet
Enligt finsk lag är alla slags diskriminering på arbetsplatserna förbjuden.
Arbetsgivaren ska se till att jämlikhet och jämställdhet mellan könen förverkligas på arbetsplatsen.
Läs mer på InfoFinlands sida Jämlikhet och jämställdhet i arbetslivet.
Eget initiativtagande och ansvar
På en finländsk arbetsplats övervakar chefen inte de anställdas arbete hela tiden.
Arbetstagarna tillfrågas om sina åsikter och åsikterna beaktas i planeringen av arbetet.
Man kommer överens om utförandet av arbetet på gemensamma möten och alla håller fast vid det man kommit överens om.
Chefen ger den anställda arbetsuppgifter och förväntar sig att den anställda själv fattar beslut om detaljerna i arbetets utförande.
Om den anställda inte kan eller förmår utföra arbetsuppgiften som anvisats, går han eller hon själv till andra anställda eller chefen för att be om råd.
Pålitlighet och att hålla tidtabeller
I den finländska arbetskulturen är det viktigt att hålla fast vid överenskommelser.
När man har beslutat något tillsammans förväntar sig både de anställda och arbetsgivaren att alla gör det man kommit överens om.
I Finland är det också viktigt att man håller fast vid tider.
Man kommer punktligt till arbetet på den avtalade tiden.
Klockan 8.00 betyder prick klockan 8.00, inte klockan 8.10.
Det är oartigt att komma för sent eftersom de andra då tvingas vänta på den som är försenad.
Om du vet att du kommer att bli sen till arbetet ska du tala om det för din chef.
På många arbetsplatser har man flexibel arbetstid och man kan komma till arbetet till exempel mellan klockan 7 och 9 och gå hem mellan klockan 15 och 17.
Om man har flexibel arbetstid ska den anställda själv se till att han eller hon arbetar den tid som avtalats.
Kommunikationsstil
Finländarna är ofta rakt på sak och frispråkighet upplevs inte som något oartigt.
Rättframhet är också vanligt i arbetslivet.
Om man till exempel inte har tillräckligt med tid för att göra en arbetsuppgift, är det bra att säga det uppriktigt till chefen.
På möten och vid diskussioner är det vanligt att man går rakt på sak genast efter att man hälsat på varandra.
I den finländska arbetskulturen tilltalar man varandra på ett mycket informellt sätt.
På de flesta arbetsplatserna duar alla varandra oberoende av sin ställning.
Religionens påverkan på arbetslivet
Många finländare är kristna men inte speciellt religiösa.
I den finländska kulturen följs dock fortfarande många kristna seder.
I arbetslivet syns religionens inflytande i de många lediga dagarna som anställda får.
Under de kristna helgerna, såsom på jul och påsk, har man lagstadgade lediga dagar.
Läs mer om högtidsdagarna på InfoFinlands sida Finländska helgdagar.
Religiösa seder eller ritualer hör inte hemma på den finländska arbetsplatsen.
På vissa arbetsplatser har man ordnat en plats för bön om de anställda framfört önskemål om det.
Sådan praxis är dock ovanlig på arbetsplatser.
Om en anställd till exempel vill hålla en bönestund under arbetsdagen ska detta göras under de avtalade pauserna.
Yttre religiösa symboler, såsom huvuddukar, är tillåtna i Finland, men de klädregler som gäller på arbetsplatserna måste följas.
Orsaken till detta är arbetssäkerhets- och hygienföreskrifter som anknyter till arbetsuppgifterna.
Du kan läsa mer om värderingar och seder i det finländska samhället på sidan Finländska seder.
Arbetsgivaren har rätt att:
anställa en arbetstagare
leda arbetet och ge råd och utfärda bestämmelser som ansluter till utförandet av arbetet
säga upp och häva ett arbetsavtal inom ramen för begränsningarna i lag
Arbetsgivaren har skyldighet att:
följa lagar och avtal
behandla arbetstagarna jämlikt oavsett deras härkomst, religion, kön, ålder eller politiska åsikt
sörja för arbetstagarnas säkerhet och arbetshälsa
ge arbetstagaren en skriftligt utredning om de centrala villkoren i arbetet
främja ett gott arbetsklimat, arbetstagarens arbetsprestationer och yrkesutveckling
Kollektivavtal
Arbetsgivaren måste följa kollektivavtalet.
Han eller hon kan till exempel inte betala ut en mindre lön än vad som fastställts i kollektivavtalet.
Inkomstregistret
Inkomstregistret är en databas dit arbetsgivarna anmäler lönerna som de utbetalat till sina anställda.
Anmälan ska göras senast fem dagar efter löneutbetalningen.
Uppgifterna ska skickas till inkomstregistret elektroniskt:
direkt via lönesystemet om det har en inbyggd teknisk förbindelse till Inkomstregistret eller
via Inkomstregistrets ärendehantering, till vilken man får tillträde med webbankkoder eller andra medel för elektronisk identifiering.
Löneuppgifterna kan endast i undantagsfall anmälas med ett pappersformulär.
Läs mer om Inkomstregistret och om att anmäla löner på Inkomstregistrets webbplats.
linkkiSkatteförvaltningen:
Inkomstregistretfinska _ svenska _ engelska _ ryska _ estniska _ kinesiska
Olycksfallsförsäkring
Arbetsgivaren ska teckna en olycksfallsförsäkring (tapaturmavakuutus) åt sina anställda.
Detta ska alltid göras när en anställning börjar.
Arbetstagaren kan få ersättning vid ett olycksfall.
Ersättningen kan vara en ersättning av sjukvårdskostnader och inkomstbortfall i form av dagpenning, olycksfallspension, ersättning för den skada som olyckan har orsakat, rehabilitering eller vid dödsfall familjepension till de anhöriga.
Arbetsgivaren kan utöver de lagstadgade försäkringarna även teckna olika frivilliga försäkringar åt sina anställda.
Det är bra att klarlägga med arbetsgivaren vilka försäkringar han eller hon har tecknat åt sina anställda.
Arbetsintyg
När en anställning upphör har den anställda rätt att få ett skriftligt arbetsintyg av arbetsgivaren.
Läs mer på InfoFinlands sida Arbetsintyg.
I Finland finns många möjligheter att studera finska.
Olika kurser ordnas för både barn och vuxna.
Undervisning i finska för vuxna
Du hittar information om kurser i finska till exempel hos medborgarinstitut, arbetarinstitut, universitet och sommaruniversitet.
Fråga mer vid rådgivningstjänsterna för invandrare, utbildningsväsendet i din hemkommun eller studievägledarna vid lokala läroanstalter.
På vissa orter har informationen om kurserna samlats på ett och samma ställe.
Till exempel finns det information om kurserna i finska språket i Helsingfors, Tammerfors och Åbo i tjänsten Finnishcourses.fi.
Vid läroanstalterna börjar kurserna vanligtvis i augusti eller september och i januari.
Språkkurserna är ofta fullsatta.
Därför är det viktigt att anmäla sig till kursen i god tid.
Medborgarinstitut i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Kurser i finska och svenska språketfinska _ engelska _ ryska
Språkstudier i anslutning till annan utbildning
Du kan studera finska också i arbetskraftsutbildning och i förberedande utbildning före yrkesutbildning (VALMA) eller förberedande gymnasieutbildning (LUVA).
Om du är kund vid arbets- och näringsbyrån kan du få plats på en kurs i finska via arbets- och näringsbyrån.
Hurdan språkundervisning du behöver bedöms på arbets- och näringsbyrån i samband med att du får en integrations- eller sysselsättningsplan.
Du kan studera finska som arbetskraftsutbildning.
Arbetskraftsutbildning är i huvudsak utbildning avsedd för arbetslösa arbetssökande.
Utbildningen är kostnadsfri för deltagarna.
Fråga om kurserna i finska på din egen arbets- och näringsbyrå.
linkkiArbets- och näringsministeriet:
Kontaktuppgifter till TE-byråerfinska _ svenska
linkkiArbets- och näringsministeriet:
Utbildning i finska och svenska språketfinska _ svenska _ engelska
Finska på arbetsplatsen
Vissa arbetsgivare ordnar finskundervisning för sina arbetstagare.
Fråga din arbetsgivare om du kan studera finska på din arbetsplats.
Arbetsgivaren kan ansöka om stöd för arbetstagarnas finskundervisning via arbets- och näringslivstjänsterna.
linkkiTE-tjänster:
Finska på arbetsplatsenfinska _ svenska _ engelska
Undervisning i finska för barn
Barn lär sig nya språk snabbt, även om det kan kännas svårt i början.
Finskundervisning ges på daghem, i förskola och skola.
Undervisningen kallas finska som andra språk eller S2-undervisning.
Barnet eller den unga kan även delta i förberedande undervisning.
Den är avsedd för de elever som ännu inte har särskilt bra kunskaper i finska.
Under den förberedande undervisningen studerar barnet eller den unga finska och några läroämnen.
Den förberedande undervisningen är avsedd för 7–16-åringar.
Undervisningen varar vanligtvis ett år.
Därefter flyttas eleven till en vanlig klass.
linkkiEdu.fi:
Finska som andra språk i den grundläggande undervisningenfinska
I Finland finns två pensionssystem som kompletterar varandra:
Arbetspensionen intjänas med det egna lönearbetet och företagandet.
Arbetsgivaren är skyldig att teckna pensionsförsäkring åt alla sina anställda och betala försäkringspremierna.
Privatföretagare sköter sina premier själva.
Folkpensionen och garantipensionen är avsedda för de pensionärer som inte får arbetspension eller vars pension är mycket liten.
Båda pensionssystemen omfattar ålderspension och invalidpension.
Du kan få folkpension när du har fyllt 65 år.
Ditt födelseår avgör i vilken ålder du kan få arbetspension.
Kontrollera din pensionsålder på ditt arbetspensionsutdrag eller hos din arbetspensionsanstalt.
Om man är arbetsoförmögen kan man få invalidpension före ålderspensionen.
Om man vill kan man också arbeta när man är pensionerad.
Om du är i ålderspension påverkar din arbetsinkomst inte pensionens storlek.
I Finland betalas skatt på pensionerna.
Arbetsgivarna och arbetstagarna finansierar pensionsskyddet tillsammans.
Arbetsgivaren drar av arbetstagarens andel från lönen och betalar den och sin egen andel av försäkringspremierna till pensionsanstalten.
Arbetspensionens belopp beror på hur länge du har arbetat och hur stor lön du har haft.
Arbetspensionsförsäkringsbolag, pensionskassor och -stiftelser har hand om arbetspensionsförsäkringarna.
Pensionsskyddscentralen sköter centraliserat frågor som rör pensionsskyddet.
linkkiPensionsskyddscentralen:
Arbetspensionfinska _ svenska _ engelska
Kontrollera på arbetspensionsutdraget hur stor pension du tjänat in
Din pensionsanstalt skickar regelbundet ett arbetspensionsutdrag till dig.
På arbetspensionsutdraget finns en uppskattning av din intjänade pension.
Du kan också beställa ett arbetspensionsutdrag från din pensionsanstalt eller Pensionsskyddscentralen.
Genom att själv följa med arbetspensionsutdragen kan du kontrollera att din intjänade pension räknats rätt.
Om det finns fel i uppgifterna, kontakta ditt pensionsbolag eller Pensionsskyddscentralen.
Spara arbetsintyg för eventuella granskningar.
Det är också bra att spara lönekvitton.
Att beställa ett arbetspensionsutdragfinska _ svenska _ engelska _ ryska _ estniska
Du kan ansöka om folkpension om du inte har någon arbetspension eller om din arbetspension är väldigt liten.
Folkpensionens belopp beror på hur länge du har bott eller arbetat i Finland. Dina familjeförhållanden och andra kontinuerliga pensionsinkomster påverkar också folkpensionens belopp.
FPA sköter folkpensionerna och garantipensionerna.
Du kan söka folkpension och garantipension om du omfattas av Finländska socialskyddet och när du har bott i Finland minst tre år efter att du fyllde 16 år.
Också den tid som du har varit bosatt i något annat EU- eller EES-land kan delvis beaktas.
Garantipensionen tryggar ett existensminimum för pensionärer.
Garantipensionens belopp är mellanskillnaden mellan de övriga pensionerna som du får och garantipensionens fulla belopp.
Om det sammanlagda beloppet från dina övriga pensioner överskrider garantipensionens fulla belopp kan du inte få garantipension.
Mer information om garantipensionen får du vid FPA.
I vissa fall kan du få folkpension även innan du fyllt 65 år.
FPA ger mer information om förtida ålderspension och tilläggsdagar till folkpension.
linkkiPensionsskyddscentralen:
Pensionssystemet i Finlandfinska _ svenska _ engelska
Stöden för pensionärerfinska _ svenska _ engelska
Information om frågor som rör pensionfinska _ svenska _ engelska _ ryska _ estniska
Att söka pension
Alla pensioner måste sökas.
Du kan ansöka om arbets- och folkpension med samma blankett.
Du kan fylla i blanketten på nätet eller lämna in den till FPA, folkpensionsverket eller Pensionskyddscentralen.
Blanketterna finns på verksamhetsställena och på internet.
Du kan ansöka om garantipensioni FPA:s nättjänst eller på kontoret.
Du kan ansöka om FPA:s åldringspension och garantipension även per telefon.
Numret till FPA:s pensionsärenden är 020 692 202.
Pension från utlandet
Om du har bott eller arbetat i andra EU-länder än Finland eller i något land med vilket Finland har ett socialskyddsavtal, kan du ha rätt till pension från dessa länder.
Du kan ansöka om pension från dessa länder samtidigt som du ansöker om den finländska arbets- eller folkpensionen.
Bifoga till din ansökan blanketten Boende och arbete utomlands.
Du kan skriva ut blanketten på FPA:s eller Pensionsskyddscentralens webbplats.
Om du har arbetat i andra länder som Finland inte har ett socialskyddsavtal med, måste du själv ta reda på om du har rätt att få pension från dessa länder.
Om du kan få pension, måste du själv ansöka om den.
Om du ansöker om pension från utlandet, får du råd vid Pensionsskyddscentralen.
Läs mer på Pensionsskyddscentralens webbplats.
Du kan även fråga om råd hos FPA.
linkkiPensionsskyddscentralen:
Broschyren Att söka pension från utlandetfinska _ svenska _ engelska _ ryska _ estniska
Utbetalning av pension till utlandet
Arbetspension utomlands
Om du flyttar från Finland utbetalas arbetspension från Finland då du går i pension.
Pensionen kan utbetalas till vilket land som helst.
Det är viktigt att du har ett arbetsintyg från alla anställningar i Finland.
Det är också bra att spara lönekvitton.
Hur du ansöker om pension till utlandet beror på i vilket land du bor.
Du kan fråga din pensionsanstalt eller Pensionsskyddscentralen om råd.
Innan du ansöker om pension ska du begära ett arbetspensionsutdrag av din pensionsanstalt eller Pensionsskyddscentralen.
Arbetspensionsutdraget visar hur stor pension du tjänat in i Finland.
FPA:s pensioner utomlands
Du ska alltid meddela FPA om varaktig flytt utomlands eller vistelse utomlands som varar över tre månader.
Om du vistas utomlands tillfälligt, det vill säga under ett år, betalar FPA vanligtvis din pension som vanligt.
I vissa fall betalar FPA till exempel ålderspension och familjepension till vissa länder även då du flyttar till landet för över ett år.
Sådana länder är till exempel de övriga EU-länderna och EES-länderna samt en del av de länder som Finland har ett socialskyddsavtal med.
Garantipensionen betalas inte om du flyttar utomlands för över ett år.
På FPA:s webbplats finns information om i vilka fall du kan få FPA:s pensioner utomlands.
Du kan också fråga om din egen situation vid FPA:s kontor eller telefontjänst.
Partiell förtida ålderspension
Om du har fyllt 61 år kan du få partiell pension redan före din lägsta ålderspensionsålder.
Detta kallas partiell förtida ålderspension.
Du kan själv välja om du vill ta ut 25 procent eller 50 procent av beloppet på din månatliga arbetspension.
Om du vill kan du samtidigt fortsätta arbeta heltid eller komma överens om en kortare arbetstid med arbetsgivaren.
Du kan också sluta arbeta.
Du bör observera att den partiella förtida ålderspensionen permanent minskar beloppet på den slutliga ålderspensionen.
Du kan fråga mer av din pensionsanstalt.
Om du är sjuk under en längre tid får du vanligtvis först under ungefär ett års tid sjukdagpenning.
Om du inte kan återgå till arbetet på grund av sjukdom eller skada kan du ansöka om invaliditetspension (työkyvyttömyyseläke) eller rehabiliteringsstöd (kuntoutustuki).
Rehabiliteringsstöd är invaliditetspension på viss tid.
Du kan ansöka om invaliditetspension med en blankett som du får från FPA.Som bilaga till ansökan krävs B-utlåtande av läkare.
FPA och arbetspensionsanstalten bedömer din arbetsförmåga och om du har nytta av rehabilitering.
Mer information om invaliditetspension och rehabilitering får du av FPA, din pensionsanstalt eller av företagshälsovården.
Om du får invaliditetspension påverkar din lönenivå pensionen.
Du ska meddela FPA och arbetspensionsanstalten om du börjar arbeta.
Om du har en tillräckligt hög inkomst från arbetet per månad kan du låta din pension vila.
Detta innebär att du håller en paus i lyftandet av pensionen.
Pausen kan vara minst tre månader och högst två år lång.
Under denna tid förlorar du inte rätten till invaliditetspension.
Övriga förmåner för pensionärer
Utöver pension kan FPA betala ut bostadsbidrag till pensionstagare med låga inkomster.
Mer information om bostadsbidrag för pensionstagare hittar du på FPA:s webbplats.
Till långtidssjuka eller handikappade kan FPA betala ut vårdbidrag för pensionstagare.
Fråga mer på FPA.
Rabatter för pensionärer
När du har pensionerats kan du få pensionärsrabatt till exempel på tåg-, buss- och flygresor i Finland.
De som fyllt 65 år får reserabatt genom att uppvisa sitt identitetsbevis.
En pensionär som inte har fyllt 65 år kan få rabatt genom att uppvisa sitt personbevis och sitt arbetspensionskort eller folkpensionärskort.
Kontrollera villkoren för pensionärsrabatten på biljettkontoren.
Du kan även få rabatt på exempelvis olika former av motion och kultur.
I skattedeklarationen finns uppgifter om inkomster, skatter och avdrag från föregående år.
Kontrollera uppgifterna i skattedeklarationen.
Den slutliga beskattningen fastställs utgående från uppgifterna i skattedeklarationen.
Om alla uppgifter är korrekta, och det inte saknas några uppgifter, behöver du inte göra någonting.
Om uppgifterna inte är korrekta, eller om det saknas något, komplettera och korrigera skattedeklarationen i webbtjänsten MinSkatt.
Du kan använda webbtjänsten, om du har finländska nätbankskoder eller ett mobilcertifikat.
Om du inte gör rättelserna i webbtjänsten MinSkatt, hämta pappersblanketter för rättelserna på Skatteförvaltningens webbplats eller i skattebyrån.
Skicka blanketterna per post.
Kom ihåg att kontrollera skattedeklarationen och göra de ändringar som behövs före utgången av den sista returdagen.
Beskattningsbeslut
Beskattningsbeslutet (Verotuspäätös) är en beräkning av det slutliga skattebeloppet.
På din lön eller annan inkomst har det innehållits skatt utgående från skattekortet.
Det här kallas för förskottsinnehållning (ennakonpidätys).
Förskottsinnehållningens storlek baserar sig på en uppskattning av dina inkomster.
Skattebeloppet justeras i efterskott utgående från hur stora dina inkomster och avdrag verkligen har varit.
Tillsammans med den på förhand ifyllda skattedeklarationen får du ett beskattningsbeslut.
Om du inte korrigerar skattedeklarationen, förblir det här beskattningsbeslutet i kraft.
Om du korrigerar skattedeklarationen, får du ett nytt beskattningsbeslut senare.
Kom ihåg att kontrollera också det nya beskattningsbeslutet.
Spara beskattningsbeslutet och den specifikationsdel som du fick på våren tillsammans med skattedeklarationen.
Om du beställer en ny specifikationsdel, tas det ut en avgift för den.
linkkiSkatteförvaltningen:
Skattedeklaration och beskattningsbeslutfinska _ svenska _ engelska
Avdrag
I beskattningen kan du göra avdrag (vähennykset), som minskar beskattningen.
Skatteförvaltningen gör en del avdrag automatiskt, men vissa avdrag måste du själv ansöka om.
Avdrag är till exempel:
hushållsavdrag
avdrag för resekostnader mellan bostaden och arbetsplatsen
ränteavdrag på bostadslån
Du kan avdra räntorna för bostadslånet i beskattningen då du har tagit ett lån för din stadigvarande bostad.
Du kan dra av räntorna på bostadslånet i beskattningen också då din stadigvarande bostad finns utomlands.
Om du har tagit ett lån hos en finländsk bank, får skattemyndigheten uppgifterna om lånet direkt från banken.
Om du har ett bostadslån i en utländsk bank, ska du själv ge uppgifterna om lånet till skattemyndigheten.
Du kan meddela om avdrag, när du beställer ett nytt skattekort.
Avdragen beaktas då i din skatteprocent.
Du kan också ansöka om avdrag i efterskott med skattedeklarationen.
Du får då avdragen i efterskott som en skatteåterbäring.
linkkiSkatteförvaltningen:
Avdrag vid beskattningenfinska _ svenska _ engelska
Skatteåterbäring och kvarskatt
Du ser i beskattningsbeslutet om du har betalat rätt mängd skatt.
Om du har betalat för mycket i skatt, får du skatteåterbäring (veronpalautus).
Om du har betalat för lite i skatt, blir du tvungen att betala kvarskatt (jäännösvero).
Skatteåterbäringen betalas antingen direkt på ditt bankkonto.
Meddela numret på ditt bankkonto via Skatteförvaltningens webbtjänst eller på en separat pappersblankett.
Du kan få skatteåterbäringen antingen till ett finländskt eller till ett utländsk bankkonto.
Om du blir tvungen att betala kvarskatt, får du tillsammans med beskattningsbeslutet en bankgiroblankett.
På bankgiroblanketten ser du kvarskattebeloppet, bankkontonumret, förfallodagen och referensnumret.
Du blir också tvungen att betala ränta på kvarskatten efter en viss tid.
linkkiSkatteåterbäringar:
Skatteåterbäringarfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Ange kontonummerfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Kvarskattfinska _ svenska _ engelska
Ungefär 90 procent av finländarna har finska som modersmål.
Ungefär fem procent av finländarna har svenska som modersmål.
När du funderar på om det är finska eller svenska som du borde lära dig ska du beakta vilket språk som talas på din hemort och i din näromgivning.
Om du vill ansöka om finskt medborgarskap måste du kunna finska, svenska eller i det finska teckenspråket.
När du ansöker om medborgarskap, bifoga ett intyg över dina språkkunskaper.
Läs mer om språkkunskapskraven på InfoFinlands sida Officiellt intyg över språkkunskaper.
På de flesta arbetsplatser är det nödvändigt att kunna finska.
Om du vill studera i Finland behöver du sannolikt kunna finska.
Det kan vara bra att lära sig finska eller svenska trots att du inte tänker bo en lång tid i landet.
Även om finländarna i allmänhet behärskar engelska relativt väl har du ändå mycket nytta av att kunna finska eller svenska.
När du behärskar språket är det lättare för dig att trivas i landet och anpassa dig till livet i Finland.
Du har lättare att sköta dina ärenden med myndigheter, följa nyheter, få nya bekantskaper och vänner.
Du lär dig språket bäst om du vågar använda det.
Du behöver inte alltid förstå allting, det räcker med att du förstår det viktigaste.
Dra dig alltså inte för situationer där du har möjlighet att tala finska eller svenska.
Information om språklagenfinska _ svenska _ engelska
linkkiKommuner.net:
Svenskspråkiga och tvåspråkiga kommunerfinska _ svenska
Vem är berättigad till utkomstskydd för arbetslösa?
Du kan registrera dig som arbetssökande vid TE-byrån om
du har ett uppehållstillstånd som ger dig rätt att arbeta i Finland
ditt uppehållstillstånd inte begränsar vilken arbetsgivare du får arbeta för
eller
du är medborgare i ett EU-land, ett EES-land eller Schweiz
du är familjemedlem till en medborgare i ett EU-land, ett EES-land eller Schweiz
Då du registrerat dig som arbetssökande har du rätt till arbetslöshetsunderstöd om du
är 17–64 år gammal
är arbetslös och anmäld som arbetssökande vid TE-byrån
söker heltidsarbete
är arbetsförmögen och tillgänglig på arbetsmarknaden
uppfyller villkoren för inkomstrelaterad dagpenning, grunddagpenning eller arbetsmarknadsstöd.
För att få utkomstskydd för arbetslösa måste du aktivt söka jobb och vara beredd att ta emot ett jobb.
Du ska också ingå en sysselsättnings- och integrationsplan med TE-byrån och delta i de tjänster och åtgärder som TE-byrån erbjuder åt dig.
På full arbetslöshetsförmån ställs även andra villkor.
Du kan få full arbetslöshetsförmån om du under 65 betalningsdagar, alltså under cirka tre månaders tid, utför en viss mängd lönearbete, får inkomst som företagare eller deltar i en verksamhet eller en tjänst som främjar din sysselsättning.
Detta kallas för aktiveringsmodellen för arbetslöshetsförsäkringen (työttömyysturvan aktiivimalli).
Arbetslöshetsförmånerna är den inkomstrelaterade dagpenningen, grunddagpenningen och arbetsmarknadsstödet.
Skatt betalas på alla arbetslöshetsförmåner.
linkkiArbets- och näringsministeriet:
Om du blir arbetslösfinska _ svenska _ engelska
linkkiArbets- och näringsministeriet:
Utkomstskydd för arbetslösafinska _ svenska _ engelska
Information om utkomstskyddet för arbetslösafinska _ svenska _ engelska
linkkiArbets- och näringsministeriet:
Rådgivning om utkomstskydd för arbetslösafinska _ svenska _ engelska _ ryska
Aktiveringsmodellen för arbetslöshetsförsäkringen finska _ svenska _ engelska
Inkomstrelaterad dagpenning
Du kan få inkomstrelaterad dagpenning om du
registrerat dig som arbetslös arbetssökande vid arbets- och näringsbyrån
hör till en finländsk arbetslöshetskassa
uppfyller arbetsvillkoret, d.v.s. har arbetat tillräckligt länge före arbetslösheten
har varit medlem i arbetslöshetskassan i minst 26 veckor innan du blev arbetslös.
Den inkomstrelaterade dagpenningen beviljas och utbetalas av den arbetslöshetskassa där du är medlem.
Den inkomstrelaterade dagpenningen beräknas utgående från storleken på den lön som du hade innan du blev arbetslös.
Vanligtvis kan inkomstrelaterad dagpenning fås under 400 dagar. Undantag från detta är följande situationer:
Om du har arbetat i sammanlagt tre år eller mindre, kan du få inkomstrelaterad dagpenning i högst 300 dagar.
Om du har fyllt 58 år innan du blev arbetslös, kan du få inkomstrelaterad dagpenning i mindre än 500 dagar.
Läs mer om arbetslöshetskassan på InfoFinlands sida Fackförbund.
Information om den inkomstrelaterade dagpenningenfinska _ svenska _ engelska
Grunddagpenning
Du kan få grunddagpenning om du omfattas av den sociala tryggheten i Finland utifrån permanent boende eller arbete före arbetslösheten och
registrerat dig som arbetslös arbetssökande vid arbets- och näringsbyrån
uppfyller arbetsvillkoret, d.v.s. har arbetat tillräckligt länge före arbetslösheten
inte uppfyller villkoren för inkomstrelaterad dagpenning.
Grunddagpenningen beviljas och utbetalas av Fpa.
Vanligtvis kan du få grunddagpenning i mindre än 400 dagar. Undantag från detta är följande situationer:
Om du har arbetat i sammanlagt tre år eller mindre, kan du få grunddagpenning i högst 300 dagar.
Om du har fyllt 58 år innan du blev arbetslös, kan du få grunddagpenning i mindre än 500 dagar.
Om du får andra sociala förmåner eller arbetsinkomster under arbetslösheten, är din grunddagpenning mindre.
Grunddagpenningfinska _ svenska _ engelska
Arbetsmarknadsstöd
Du kan få arbetsmarknadsstöd om du
registrerat dig som arbetslös arbetssökande vid arbets- och näringsbyrån
bor permanent i Finland
inte uppfyller arbetsvillkoret, d.v.s. inte arbetat tillräckligt länge innan du blev arbetslös eller fått förvärvsrelaterad dagpenning eller grunddagpenning under maximitiden.
Om du har en gällande integrationsplan, kan du söka arbetsmarknadsstöd för den tid då du deltar i utbildningar och annan verksamhet som nedtecknats i planen.
Närmare uppgifter om integrationsplanen finns på InfoFinlands sida Integration i Finland.
Arbetsmarknadsstödet beviljas och utbetalas av Fpa.
Arbetsmarknadsstödet är behovsprövat.
Det betyder att till exempel sociala förmåner och lön minskar arbetsmarknadsstödets belopp.
Om du är under 25 år, kontrollera tilläggsvillkoren för arbetsmarknadsstödet för unga på TE-tjänsternas webbplats.
Arbetsmarknadsstödfinska _ svenska _ engelska
Du behöver ett skattekort (verokortti), om du får lön eller har andra inkomster i Finland.
På skattekortet finns en anteckning om skatteprocenten (veroprosentti).
Av det ser arbetsgivaren, hur mycket skatt som ska betalas på lönen.
Skatteprocenten beror på hur hög din inkomst är.
Om du håller på att flytta till Finland, får du skattekortet från skattebyrån (verotoimisto).
Uppskatta för skattekortet, hur stora dina inkomster kommer att bli för hela skatteåret.
Du behöver också en finländsk personbeteckning.
Du får personbeteckningen, när du registrerar dig som invånare hos magistraten.
Du kan få en personbeteckning också från skattebyrån.
Läs mer på sidan Registrering som invånare.
När du bor i Finland stadigvarande, skickar Skatteförvaltningen ett nytt skattekort till dig varje år i januari.
Skatteförvaltningen räknar ut en lämplig skatteprocent åt dig utgående från hur mycket du förtjänade året innan.
Förete skattekortet till din arbetsgivare.
Om du inte företer skattekortet till din arbetsgivare, innehåller arbetsgivaren en skatt på 60 % på din lön.
Om dina inkomster blir mindre eller större under året, ska du beställa ett nytt skattekort.
Du får ett nytt skattekort:
från Skatteförvaltningens webbtjänst MinSkatt
på skattebyrån
Du kan även beställa skattekortet via Skatteförvaltningens telefontjänst:
finska 029 497 000
svenska 029 497 001
engelska 029 497 050
När du söker ett nytt skattekort, behöver du följande uppgifter:
en uppskattning av dina inkomster för hela året
de inkomster som du har haft från början av året
de skatter som har betalats på dina inkomster från början av året
uppgift om de avdrag som du söker i beskattningen för innevarande år
Om du betalar för mycket skatt, får du skatteåterbäring.
Om du betalar för litet i skatt, blir du tvungen att betala kvarskatt.
linkkiSkatteförvaltningen:
Nytt skattekortfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Hur beräknas skatteprocenten?finska _ svenska _ engelska
Om du har flera arbetsgivare
Om du har flera arbetsgivare ska du förete ditt skattekort till dem alla.
Du kan använda samma skattekort hos alla arbetsgivarna.
Du betalar samma skatt hos alla dina arbetsgivare.
På skattekortet anges en inkomstgräns och din skatteprocent beräknas utifrån den.
Kom ihåg att hålla ett öga på dina inkomster.
Om du får mer lön än vad du uppgett, överskrids din inkomstgräns.
Om inkomstgränsen överskrids ska du beställa ett nytt skattekort.
Skattenummer
Du behöver en skattenummer (veronumero), om du arbetar på en bygg- eller monteringsarbetsplats i Finland.
Med hjälp av skattenumret kontrolleras, att alla arbetstagare finns i Skatteförvaltningens register.
Skattenumret ska framgå av den fotoförsedda namnskylt som du får av din arbetsgivare.
Du får inte arbeta på en byggplats utan namnskylt.
Du får skattenumret från skattebyrån samtidigt som du går efter skattekortet.
Om du redan har finländsk personbeteckning och ett skattekort, hittar du skattenumret på ditt skattekort.
linkkiSkatteförvaltningen:
Skattenummerfinska _ svenska _ engelska
Intern kommunikation på arbetsplatsen
Vanligen informerar man om kommande händelser och ändringar på arbetsplatsen vid möten.
Om man deltar i möten kan man påverka, föreslå ändringar och utveckla sitt eget arbete.
På varje arbetsplats finns också andra kanaler för den interna kommunikationen, såsom anslagstavlor, e-post eller de anställdas postfack.
Följ informationen på arbetsplatsen.
Pauser
I arbetsavtalet står det ofta hur långa pauser som ingår i arbetsdagen och tidpunkten för dessa.
Vanligen har man en kort kaffepaus på förmiddagen, en lunchpaus mitt på dagen och en kaffepaus till på eftermiddagen.
Längden på lunchpausen varierar mellan olika arbetsplatser.
Fråga din chef hur långa pauser du har.
Arbetsplatsbespisningen är ordnad på olika sätt på olika arbetsplatser: vissa arbetsplatser har en egen personalmatsal, på andra ställen tar de anställda med sig maten hemifrån.
På vissa arbetsplatser kan man köpa förmånliga lunchsedlar som man kan använda på matställen i närheten av arbetsplatsen.
Under lunchen arbetar man vanligtvis inte.
Att sköta egna ärenden under arbetsdagen
På arbetstid får man inte sköta sina privata angelägenheter, utan detta måste göras utanför arbetstiden.
Antalet arbetstimmar som står i arbetsavtalet är bindande och det avtalade antalet arbetstimmar ska fullgöras.
Under pauserna kan du till exempel ringa viktiga samtal.
Du kan också ansöka om oavlönad ledighet om din situation kräver att du är frånvarande en längre tid.
Om du av någon anledning inte till exempel lyckas få en läkartid utanför arbetstiden, ska du komma överens med din chef om att du är borta och hur du ersätter din frånvaro.
Företagshälsovården kan du besöka under arbetstid.
Utbildning som rör arbetet
Även om arbetstagaren har sådan utbildning som krävs för yrket redan när anställningen inleds, uppmuntrar många arbetsgivare sina anställda att skaffa sig mer utbildning.
Ofta kan du utbilda dig på arbetstid och arbetsgivaren kan betala för utbildningen.
De flesta arbetsgivare värdesätter att den anställda vill utveckla sig i sitt arbete och inhämta nya kunskaper.
Vanligen ger man inte varandra presenter på arbetsplatserna.
På viktiga bemärkelsedagar (födelsedagar, äktenskap, pensionering) uppmärksammar arbetskamraterna och arbetsgivaren festföremålet med en liten present eller en blombukett.
Arbetstid och semester
En normal arbetsdag är vanligtvis åtta timmar.
Arbetstagaren kan även komma överens om någon annan tid med arbetsgivaren.
I Finland gör arbetstagare vanligtvis inte mycket övertid.
Man arbetar de timmar som står i anställningsavtalet.
I Finland börjar semesterperioden i början av maj.
Antalet intjänade semesterdagar beror på anställningstiden i år och när anställningen har börjat.
Utöver den betalda semesterna kan du ansöka om obetald ledighet.
Jämfört med många andra länder har arbetstagare i Finland långa semestrar.
Arbetshälsa och rekreation
På många arbetsplatser vill man stödja de anställdas arbetsmotivation och -trivsel med olika rekreationsdagar och fester på arbetsplatsen. Arbetsgivaren kan också erbjuda sina anställda olika hobbymöjligheter vid sidan av arbetet.
Årliga helger
Vissa dagar är allmänna lediga dagar i Finland.
Till dem hör följande:
nyårsdagen 1.1
trettondagen 6.1
påsk: tidpunkten varierar, i mars-april
första maj 1.5
midsommarafton: i juni, alltid en fredag
självständighetsdagen 6.12
juldagen 25.12
annandag jul 26.12
Läs mer om dessa dagar på sidan Finländska helgdagar.
På vissa arbetsplatser, till exempel sjukhus, arbetar man även under helgerna.
För arbetet under helgerna betalas högre lön.
Kontrollera ersättningen i ditt kollektivavtal.
Anmäl dig som arbetslös arbetssökande
Om du blir arbetslös ska du anmäla dig hos TE-byrån senast den första dagen av din arbetslöshet.
Om du omfattas av den finländska sociala tryggheten kan du ansöka om arbetslöshetsstöd.
Du kan få arbetslöshetsstöd från och med det datum då du anmälde dig som arbetslös.
Kom ihåg att anmäla dig också direkt efter studier, arbetskraftsutbildning eller en period med sysselsättningsstöd.
Anmäl dig som arbetssökande i TE-byråns webbtjänst.
Logga in med finländska nätbankskoder eller personkort med microchip.
En anställd vid TE-byrån tar kontakt med dig om det behövs ytterligare uppgifter.
Du behöver inte ringa eller besöka TE-byrån om du inte uttryckligen ombes göra detta.
Om du saknar nätbankskoder eller personkort med microchip ska du anmäla dig som arbetssökande vid närmaste TE-byrå.
Endast medborgare i EU-länderna, Norge, Island, Liechtenstein och Schweiz kan anmäla sig som arbetssökande i webbtjänsten.
Om du är medborgare i ett annat land måste du besöka arbets- och näringsbyrån.
När du går till TE-byrån ska du ta med dig
alla dina arbetsintyg och studiebetyg
ditt pass där ditt uppehållstillstånd syns
TE-byrån undersöker uppgifterna som du lämnar.
Det finns vissa villkor för att få utkomstskydd för de arbetslösa och TE-byrån utreder om dessa villkor uppfylls i din situation.
Därefter ger TE-byrån ett utlåtande i ärendet till den instans som betalar förmånen, det vill säga till arbetslöshetskassan eller FPA.
Du kan fråga råd i ärenden som rör utkomstskyddet för arbetslösa vid din egen TE-byrå.
Du kan också ringa TE-tjänsternas rådgivning om utkomstskydd för arbetslösa:
på finska: 0295 020 701
på svenska: 0295 020 711
på engelska: 0295 030 713
på ryska: 0295 020 715
Läs också InfoFinlands sida:
Arbetslöshetsförsäkring
linkkiArbets- och näringsministeriet:
Om du blir arbetslösfinska _ svenska _ engelska
linkkiArbets- och näringsministeriet:
Att anmäla sig som arbetslös arbetssökandefinska _ svenska
linkkiArbets- och näringsministeriet:
Rådgivning om utkomstskydd för arbetslösafinska _ svenska _ engelska _ ryska
Semester, studier eller arbete under arbetslösheten
Om du börjar arbeta eller studera när du är arbetslös ska du meddela detta till TE-byrån.
Du får anvisningar om hur detta påverkar ditt utkomststöd för arbetslösa.
Om du reser i hemlandet eller utomlands ska du se till att du alltid kan nås.
Lämna till exempel ditt telefonnummer och din adress till TE-byrån och ange hur länge du ämnar vistas på resmålet.
Du kan ändå inte tacka nej till ett jobb som erbjuds till dig på grund av en utlandsresa.
Om du startar ett företag när du är arbetslös, kan du få arbetslöshetsförmån under de fyra första månaderna.
Karens
Du kan förlora din rätt till arbetslöshetsdagpenning för en viss tid om du själv har förorsakat arbetslösheten.
Du kan sättas i karens till exempel om:
du inte söker ett jobb som TE-byrån föreslår för dig
du inte tar emot ett jobb som erbjuds till dig
du säger upp dig från ditt jobb utan en godtagbar anledning
Karenstidens längd varierar från 15 dagar till 90 dagar.
Längden beror på orsaken till karensen.
I vissa fall kan du förlora rätten till utkomststöd för arbetslösa tillsvidare.
I Finland betalar du inkomstskatt (tulovero) på lön.
Du betalar också skatt på till exempel följande inkomster:
arbetsersättning
företagsinkomst
arbetslöshetsdagpenning
föräldradagpenning
pensioner
studiestöd
För skattepengarna betalar staten och kommunerna till exempel:
hälsovård
utbildning
dagvård
försvar
I Finland är beskattningen progressiv.
Det innebär att man på en stor lön betalar en större andel skatt än på en mindre lön.
Skatteprocenten (Veroprosentti) beräknas i Finland för var och en separat.
Din makes/makas inkomster inverkar inte på din skatteprocent.
Du kan uppskatta din skatteprocent med Skatteförvaltningens skatteräknare.
Arbetsgivaren betalar skatterna direkt från din lön.
För att kunna göra det behöver arbetsgivaren ett skattekort av dig.
Skatt som betalas direkt från lönen, är förskottsskatt (ennakonpidätys).
Skatteförvaltningen räknar efter varje år om du har betalat tillräckligt med skatt på dina inkomster.
Om du har betalat för mycket i skatt, får du skatteåterbäring (veronpalautus).
Om du har betalat för lite i skatt, blir du tvungen att betala kvarskatt (jäännösvero).
Läs mer på sidan: Skattedeklaration och beskattningsbeslut.
Kontrollera i lönespecifikationen och skattedeklarationen (veroilmoitus), att arbetsgivaren har betalat skatt på din lön.
Spara lönekvittona.
Om skatten inte har betalats, blir du tvungen att betala den i efterskott.
Utöver skatt betalar arbetsgivaren försäkringspremier på din lön i händelse av arbetslöshet eller sjukdom.
linkkiSkatteförvaltningen:
Information om beskattningenfinska _ svenska _ engelska
linkkiSkattemyndigheten:
Skattekortfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Att beställa skattekort finska _ svenska _ engelska
linkkiSkatteförvaltningen:
Skatteprocenträknarefinska _ svenska _ engelska
Beskattningen när du börjar arbeta i Finland
Om du kommer till Finland för att arbeta, beror din beskattning på hur länge du vistas i Finland.
På beskattningen inverkar också huruvida din arbetsgivare är ett finländskt eller ett utländskt företag.
Om du vistas i Finland i mer än sex månader, ska du i allmänhet betala skatt på din lön till Finland.
Du ska i allmänhet också betala de obligatoriska försäkringspremierna till Finland.
Du behöver en finländsk personbeteckning och ett finländskt skattekort.
Skatteprocenten räknas på inkomsterna för hela året.
Du får skatteavdrag på samma grunder som andra som bor i Finland stadigvarande.
Om du vistas i Finland i högst sex månader och din arbetsgivare är ett utländskt företag, behöver du i allmänhet inte betala skatt till Finland.
Om din arbetsgivare är finländare eller om din utländska arbetsgivare har en arbetsplats i Finland, betalar du skatt i Finland.
Du kan söka progressiv beskattning, om du bor i ett land som hör till Europeiska ekonomiska samarbetsområdet eller i en stat, med vilken Finland har ett skatteavtal.
I annat fall betalar du en källskatt (lähdevero) på 35 % på lönen och du behöver ett källskattekort.
Källskattekort måste du ansöka med en pappersblankett.
För progressiv beskattning behöver du ett skattekort för begränsat skattskyldiga (rajoitetusti verovelvollisen verokortti).
Du får ett sådant på skattebyrån.
Du kan söka progressiv beskattning också i efterskott.
Du blir också tvungen att betala försäkringspremier, om du inte är försäkrad i det land där du bor stadigvarande.
Om du redan är försäkrad i ett annat land, behöver du ett intyg A1/E101 över försäkringen.
När du flyttar bort från Finland, kom ihåg att göra en flyttningsanmälan till magistraten.
Du får då din skattedeklaration till rätt adress.
När du håller på att flytta till Finland, får du ytterligare information i avsnittet Flytta till Finland.
linkkiSkatteförvaltningen:
Arbeta i Finlandfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Ansökan om progressiv inkomstbeskattningfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Utländsk hyrd arbetskraft och beskattningen i Finlandfinska _ svenska _ engelska
Flyttanmälanfinska _ svenska _ engelska
I Finland värdesätts ärlighet, punktlighet och jämställdhet.
Det syns överallt i den finländska kulturen, även i arbetslivet.
På den här sidan finns mer information om den finländska arbetskulturen.
Du kan läsa mer om värderingar och seder i det finländska samhället på sidan Finländska seder.
Lär dig finska eller svenska
Du kan utveckla dina språkkunskaper på kurser eller i arbetet.
Dra dig inte för att prata finska eller svenska med dina kollegor.
Läs mer om språkstudier i InfoFinlands avsnitt Finska och svenska språket.
Jämlikhet och jämställdhet i arbetslivet
Enligt finsk lag är alla slags diskriminering på arbetsplatserna förbjuden.
Arbetsgivaren ska se till att jämlikhet och jämställdhet mellan könen förverkligas på arbetsplatsen.
Läs mer på InfoFinlands sida Jämlikhet och jämställdhet i arbetslivet.
Eget initiativtagande och ansvar
På en finländsk arbetsplats övervakar chefen inte de anställdas arbete hela tiden.
Arbetstagarna tillfrågas om sina åsikter och åsikterna beaktas i planeringen av arbetet.
Man kommer överens om utförandet av arbetet på gemensamma möten och alla håller fast vid det man kommit överens om.
Chefen ger den anställda arbetsuppgifter och förväntar sig att den anställda själv fattar beslut om detaljerna i arbetets utförande.
Om den anställda inte kan eller förmår utföra arbetsuppgiften som anvisats, går han eller hon själv till andra anställda eller chefen för att be om råd.
Pålitlighet och att hålla tidtabeller
I den finländska arbetskulturen är det viktigt att hålla fast vid överenskommelser.
När man har beslutat något tillsammans förväntar sig både de anställda och arbetsgivaren att alla gör det man kommit överens om.
I Finland är det också viktigt att man håller fast vid tider.
Man kommer punktligt till arbetet på den avtalade tiden.
Klockan 8.00 betyder prick klockan 8.00, inte klockan 8.10.
Det är oartigt att komma för sent eftersom de andra då tvingas vänta på den som är försenad.
Om du vet att du kommer att bli sen till arbetet ska du tala om det för din chef.
På många arbetsplatser har man flexibel arbetstid och man kan komma till arbetet till exempel mellan klockan 7 och 9 och gå hem mellan klockan 15 och 17.
Om man har flexibel arbetstid ska den anställda själv se till att han eller hon arbetar den tid som avtalats.
Kommunikationsstil
Finländarna är ofta rakt på sak och frispråkighet upplevs inte som något oartigt.
Rättframhet är också vanligt i arbetslivet.
Om man till exempel inte har tillräckligt med tid för att göra en arbetsuppgift, är det bra att säga det uppriktigt till chefen.
På möten och vid diskussioner är det vanligt att man går rakt på sak genast efter att man hälsat på varandra.
I den finländska arbetskulturen tilltalar man varandra på ett mycket informellt sätt.
På de flesta arbetsplatserna duar alla varandra oberoende av sin ställning.
Religionens påverkan på arbetslivet
Många finländare är kristna men inte speciellt religiösa.
I den finländska kulturen följs dock fortfarande många kristna seder.
I arbetslivet syns religionens inflytande i de många lediga dagarna som anställda får.
Under de kristna helgerna, såsom på jul och påsk, har man lagstadgade lediga dagar.
Läs mer om högtidsdagarna på InfoFinlands sida Finländska helgdagar.
Religiösa seder eller ritualer hör inte hemma på den finländska arbetsplatsen.
På vissa arbetsplatser har man ordnat en plats för bön om de anställda framfört önskemål om det.
Sådan praxis är dock ovanlig på arbetsplatser.
Om en anställd till exempel vill hålla en bönestund under arbetsdagen ska detta göras under de avtalade pauserna.
Yttre religiösa symboler, såsom huvuddukar, är tillåtna i Finland, men de klädregler som gäller på arbetsplatserna måste följas.
Orsaken till detta är arbetssäkerhets- och hygienföreskrifter som anknyter till arbetsuppgifterna.
linkkiFFC:
Arbetslivet i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ kinesiska _ arabiska
Arbetsgivaren har rätt att:
anställa en arbetstagare
leda arbetet och ge råd och utfärda bestämmelser som ansluter till utförandet av arbetet
säga upp och häva ett arbetsavtal inom ramen för begränsningarna i lag
Arbetsgivaren har skyldighet att:
följa lagar och avtal
behandla arbetstagarna jämlikt oavsett deras härkomst, religion, kön, ålder eller politiska åsikt
sörja för arbetstagarnas säkerhet och arbetshälsa
ge arbetstagaren en skriftligt utredning om de centrala villkoren i arbetet
främja ett gott arbetsklimat, arbetstagarens arbetsprestationer och yrkesutveckling
Kollektivavtal
Arbetsgivaren måste följa kollektivavtalet.
Han eller hon kan till exempel inte betala ut en mindre lön än vad som fastställts i kollektivavtalet.
Inkomstregistret
Inkomstregistret är en databas dit arbetsgivarna anmäler lönerna som de utbetalat till sina anställda.
Anmälan ska göras senast fem dagar efter löneutbetalningen.
Uppgifterna ska skickas till inkomstregistret elektroniskt:
direkt via lönesystemet om det har en inbyggd teknisk förbindelse till Inkomstregistret eller
via Inkomstregistrets ärendehantering, till vilken man får tillträde med webbankkoder eller andra medel för elektronisk identifiering.
Löneuppgifterna kan endast i undantagsfall anmälas med ett pappersformulär.
Läs mer om Inkomstregistret och om att anmäla löner på Inkomstregistrets webbplats.
linkkiSkatteförvaltningen:
Inkomstregistretfinska _ svenska _ engelska _ ryska _ estniska _ kinesiska
Olycksfallsförsäkring
Arbetsgivaren ska teckna en olycksfallsförsäkring (tapaturmavakuutus) åt sina anställda.
Detta ska alltid göras när en anställning börjar.
Arbetstagaren kan få ersättning vid ett olycksfall.
Ersättningen kan vara en ersättning av sjukvårdskostnader och inkomstbortfall i form av dagpenning, olycksfallspension, ersättning för den skada som olyckan har orsakat, rehabilitering eller vid dödsfall familjepension till de anhöriga.
Arbetsgivaren kan utöver de lagstadgade försäkringarna även teckna olika frivilliga försäkringar åt sina anställda.
Det är bra att klarlägga med arbetsgivaren vilka försäkringar han eller hon har tecknat åt sina anställda.
Arbetsintyg
När en anställning upphör har den anställda rätt att få ett skriftligt arbetsintyg av arbetsgivaren.
Läs mer på InfoFinlands sida Arbetsintyg.
Intressebevakning och rådgivning för företagare
Företagarens utkomstskydd för arbetslösa
Företagarens företagshälsovård
Om en företagare blir sjuk
Intressebevakning och rådgivning för företagare
Finlands Näringsliv EK representerar alla privata branscher och företag i alla storlekar.
Branschförbunden är intressebevakningsorganisationer för företag i olika branscher.
De tillhandahåller sina medlemsföretag ofta också många slags tjänster såsom rådgivning i frågor som rör företagande och den aktuella branschen.
linkkiFinlands Näringsliv EK:
Intressebevakning för företagarefinska _ svenska _ engelska
Företagarna i Finland (Suomen Yrittäjät) är företagarnas intressebevakningsorganisation som också producerar sina medlemmar olika tjänster, som till exempel gratis telefonrådgivning i frågor som rör företagande.
linkkiFöretagarna i Finland:
Intressebevakning för företagarefinska _ svenska _ engelska
TE-byrån tillhandahåller tjänster som stöder utvecklingen av affärsverksamheten.
Via TE-byrån kan du även leta en fortsättare för din företagsverksamhet eller en partner till ditt företag.
Nyföretagarcentraler erbjuder kostnadsfri företagsrådgivning runtom i Finland.
Hos företagsrådgivningen kan du få hjälp med frågor kring företagets verksamhet eller utveckling.
linkkiNyföretagarcentralerna i Finland:
Företagsrådgivningfinska _ svenska _ engelska
Företagsfinland erbjuder en gratis telefontjänst där du får sakkunnig rådgivning om ditt företag har ekonomiska svårigheter.
Rådgivning ges på finska och svenska.
Ekonomihjälp-rådgivningen
på finska, tfn 029 502 4880
på svenska, tfn 029 502 4881
Tjänsten har öppet måndag till fredag kl. 9.00–16.00.
linkkiFöretagsFinland:
Ekonomisk rådgivning för företagarefinska _ svenska
Företagarens utkomstskydd för arbetslösa
Också företagaren har rätt till utkomstskydd för arbetslösa.
En företagare är arbetslös när han eller hon har lagt ned sin företagsverksamhet eller sålt sin andel av företaget.
Företagandet kan också upphöra om företaget säljs, avvecklas, går i konkurs, försätts i likvidation eller på grund av skilsmässa.
Företagaren betraktas som arbetslös också om man har haft ett uppehåll på minst fyra månader i företagsverksamheten.
Om du måste lägga ned din företagsverksamhet, ska du omgående anmäla dig som arbetslös arbetssökande via TE-byråns webbtjänst.
Du kan få arbetslöshetsersättning tidigast från den dag då du gjort anmälan vid TE-byrån.
Information om företagarens sociala trygghetfinska _ svenska _ engelska
Om du vill få inkomstrelaterat utkomstskydd för arbetslösa, ska du ansluta dig som medlem i företagarnas arbetslöshetskassa (yrittäjien työttömyyskassa).
Om din företagsverksamhet upphör, kan du ansöka om inkomstrelaterad dagpenning (ansiosidonnainen päiväraha) vid arbetslöshetskassan.
Du kan få inkomstrelaterad dagpenning från företagarnas arbetslöshetskassa om du har bedrivit företagsverksamhet och varit medlem i kassan tillräckligt länge innan du blev arbetslös.
Den inkomstrelaterade dagpenningen är större än grunddagpenningen eller arbetsmarknadsstödet.
Hur stor inkomstrelaterad dagpenning du får beror på hur stora förvärvsinkomster du angett som grund för arbetslöshetsförsäkringen.
linkkiFöretagarnas Arbetslöshetskassa i Finland:
Företagarnas Arbetslöshetskassa i Finlandfinska _ svenska
linkkiYrkesutövarnas och företagarnas arbetslöshetskassa:
Yrkesutövarnas och företagarnas arbetslöshetskassafinska _ svenska _ engelska _ ryska _ estniska
Grunddagpenning
Fpa kan betala grunddagpenning (peruspäiväraha) för en arbetslös företagare som inte är medlem i en arbetslöshetskassa.
Om du uppfyller arbetsvillkoret för företagare och omfattas av den sociala tryggheten i Finland kan du få grunddagpenning.
På FPA:s webbplats finns en räknare som du kan använda för att beräkna om du uppfyller arbetsvillkoret för företagare.
Arbetsmarknadsstöd
Om du inte har rätt till grunddagpenning eller inkomstrelaterad dagpenning, men omfattas av den sociala tryggheten i Finland, kan du ansöka om arbetsmarknadsstöd.
Arbetsmarknadsstödet är behovsprövat, vilket betyder att dina andra inkomster och din situation som en helhet påverkar dess belopp.
Företagarens företagshälsovård
En företagare och andra som arbetar åt sig själv kan ordna företagshälsovård för sig själv om de så önskar.
Företagare måste inte ordna företagshälsovård för sig själv, men däremot måste de ordna det för sina anställda.
Företagshälsovård kan ordnas på den lokala hälsovårdscentralen (terveyskeskus) eller till exempel en privat läkarstation.
Läs mer på InfoFinlands sida Företagshälsovård.
Information för företagare om företagshälsovårdenfinska _ svenska _ engelska
Om en företagare blir sjuk
Om du blir sjuk, kan du få sjukdagpenning (sairauspäiväraha) från Fpa. Den ersätter inkomstbortfallet på grund av arbetsoförmåga när arbetsoförmågan varar mindre än ett år.
Betalningen av dagpenning inleds efter en självrisktid (omavastuuaika).
För företagare är självrisktiden oftast dagen för insjuknandet och följande tre vardagar.
Företagarens sjukdagpenningfinska _ svenska _ engelska
I Finland finns två pensionssystem som kompletterar varandra:
Arbetspensionen intjänas med det egna lönearbetet och företagandet.
Arbetsgivaren är skyldig att teckna pensionsförsäkring åt alla sina anställda och betala försäkringspremierna.
Privatföretagare sköter sina premier själva.
Folkpensionen och garantipensionen är avsedda för de pensionärer som inte får arbetspension eller vars pension är mycket liten.
Båda pensionssystemen omfattar ålderspension och invalidpension.
Du kan få folkpension när du har fyllt 65 år.
Ditt födelseår avgör i vilken ålder du kan få arbetspension.
Kontrollera din pensionsålder på ditt arbetspensionsutdrag eller hos din arbetspensionsanstalt.
Om man är arbetsoförmögen kan man få invalidpension före ålderspensionen.
Om man vill kan man också arbeta när man är pensionerad.
Om du är i ålderspension påverkar din arbetsinkomst inte pensionens storlek.
I Finland betalas skatt på pensionerna.
Arbetsgivarna och arbetstagarna finansierar pensionsskyddet tillsammans.
Arbetsgivaren drar av arbetstagarens andel från lönen och betalar den och sin egen andel av försäkringspremierna till pensionsanstalten.
Arbetspensionens belopp beror på hur länge du har arbetat och hur stor lön du har haft.
Arbetspensionsförsäkringsbolag, pensionskassor och -stiftelser har hand om arbetspensionsförsäkringarna.
Pensionsskyddscentralen sköter centraliserat frågor som rör pensionsskyddet.
linkkiPensionsskyddscentralen:
Arbetspensionfinska _ svenska _ engelska
Kontrollera på arbetspensionsutdraget hur stor pension du tjänat in
Din pensionsanstalt skickar regelbundet ett arbetspensionsutdrag till dig.
På arbetspensionsutdraget finns en uppskattning av din intjänade pension.
Du kan också beställa ett arbetspensionsutdrag från din pensionsanstalt eller Pensionsskyddscentralen.
Genom att själv följa med arbetspensionsutdragen kan du kontrollera att din intjänade pension räknats rätt.
Om det finns fel i uppgifterna, kontakta ditt pensionsbolag eller Pensionsskyddscentralen.
Spara arbetsintyg för eventuella granskningar.
Det är också bra att spara lönekvitton.
Att beställa ett arbetspensionsutdragfinska _ svenska _ engelska _ ryska _ estniska
Du kan ansöka om folkpension om du inte har någon arbetspension eller om din arbetspension är väldigt liten. Folkpensionens belopp beror på hur länge du har bott eller arbetat i Finland.
Dina familjeförhållanden och andra kontinuerliga pensionsinkomster påverkar också folkpensionens belopp.
FPA sköter folkpensionerna och garantipensionerna.
Du kan söka folkpension och garantipension om du omfattas av Finländska socialskyddet och när du har bott i Finland minst tre år efter att du fyllde 16 år.
Också den tid som du har varit bosatt i något annat EU- eller EES-land kan delvis beaktas.
Garantipensionen tryggar ett existensminimum för pensionärer.
Garantipensionens belopp är mellanskillnaden mellan de övriga pensionerna som du får och garantipensionens fulla belopp.
Om det sammanlagda beloppet från dina övriga pensioner överskrider garantipensionens fulla belopp kan du inte få garantipension.
Mer information om garantipensionen får du vid FPA.
I vissa fall kan du få folkpension även innan du fyllt 65 år.
FPA ger mer information om förtida ålderspension och tilläggsdagar till folkpension.
linkkiPensionsskyddscentralen:
Pensionssystemet i Finlandfinska _ svenska _ engelska
Stöden för pensionärerfinska _ svenska _ engelska
Information om frågor som rör pensionfinska _ svenska _ engelska _ ryska _ estniska
Att söka pension
Alla pensioner måste sökas.
Du kan ansöka om arbets- och folkpension med samma blankett.
Du kan fylla i blanketten på nätet eller lämna in den till FPA, folkpensionsverket eller Pensionskyddscentralen.
Blanketterna finns på verksamhetsställena och på internet.
Du kan ansöka om garantipensioni FPA:s nättjänst eller på kontoret.
Du kan ansöka om FPA:s åldringspension och garantipension även per telefon.
Numret till FPA:s pensionsärenden är 020 692 202.
Pension från utlandet
Om du har bott eller arbetat i andra EU-länder än Finland eller i något land med vilket Finland har ett socialskyddsavtal, kan du ha rätt till pension från dessa länder.
Du kan ansöka om pension från dessa länder samtidigt som du ansöker om den finländska arbets- eller folkpensionen.
Bifoga till din ansökan blanketten Boende och arbete utomlands.
Du kan skriva ut blanketten på FPA:s eller Pensionsskyddscentralens webbplats.
Om du har arbetat i andra länder som Finland inte har ett socialskyddsavtal med, måste du själv ta reda på om du har rätt att få pension från dessa länder.
Om du kan få pension, måste du själv ansöka om den.
Om du ansöker om pension från utlandet, får du råd vid Pensionsskyddscentralen.
Läs mer på Pensionsskyddscentralens webbplats.
Du kan även fråga om råd hos FPA.
linkkiPensionsskyddscentralen:
Broschyren Att söka pension från utlandetfinska _ svenska _ engelska _ ryska _ estniska
Utbetalning av pension till utlandet
Arbetspension utomlands
Om du flyttar från Finland utbetalas arbetspension från Finland då du går i pension.
Pensionen kan utbetalas till vilket land som helst.
Det är viktigt att du har ett arbetsintyg från alla anställningar i Finland.
Det är också bra att spara lönekvitton.
Hur du ansöker om pension till utlandet beror på i vilket land du bor.
Du kan fråga din pensionsanstalt eller Pensionsskyddscentralen om råd.
Innan du ansöker om pension ska du begära ett arbetspensionsutdrag av din pensionsanstalt eller Pensionsskyddscentralen.
Arbetspensionsutdraget visar hur stor pension du tjänat in i Finland.
FPA:s pensioner utomlands
Du ska alltid meddela FPA om varaktig flytt utomlands eller vistelse utomlands som varar över tre månader.
Om du vistas utomlands tillfälligt, det vill säga under ett år, betalar FPA vanligtvis din pension som vanligt.
I vissa fall betalar FPA till exempel ålderspension och familjepension till vissa länder även då du flyttar till landet för över ett år.
Sådana länder är till exempel de övriga EU-länderna och EES-länderna samt en del av de länder som Finland har ett socialskyddsavtal med.
Garantipensionen betalas inte om du flyttar utomlands för över ett år.
På FPA:s webbplats finns information om i vilka fall du kan få FPA:s pensioner utomlands.
Du kan också fråga om din egen situation vid FPA:s kontor eller telefontjänst.
Partiell förtida ålderspension
Om du har fyllt 61 år kan du få partiell pension redan före din lägsta ålderspensionsålder.
Detta kallas partiell förtida ålderspension.
Du kan själv välja om du vill ta ut 25 procent eller 50 procent av beloppet på din månatliga arbetspension.
Om du vill kan du samtidigt fortsätta arbeta heltid eller komma överens om en kortare arbetstid med arbetsgivaren.
Du kan också sluta arbeta.
Du bör observera att den partiella förtida ålderspensionen permanent minskar beloppet på den slutliga ålderspensionen.
Du kan fråga mer av din pensionsanstalt.
Om du är sjuk under en längre tid får du vanligtvis först under ungefär ett års tid sjukdagpenning.
Om du inte kan återgå till arbetet på grund av sjukdom eller skada kan du ansöka om invaliditetspension (työkyvyttömyyseläke) eller rehabiliteringsstöd (kuntoutustuki).
Rehabiliteringsstöd är invaliditetspension på viss tid.
Du kan ansöka om invaliditetspension med en blankett som du får från FPA.Som bilaga till ansökan krävs B-utlåtande av läkare.
FPA och arbetspensionsanstalten bedömer din arbetsförmåga och om du har nytta av rehabilitering.
Mer information om invaliditetspension och rehabilitering får du av FPA, din pensionsanstalt eller av företagshälsovården.
Om du får invaliditetspension påverkar din lönenivå pensionen.
Du ska meddela FPA och arbetspensionsanstalten om du börjar arbeta.
Om du har en tillräckligt hög inkomst från arbetet per månad kan du låta din pension vila.
Detta innebär att du håller en paus i lyftandet av pensionen.
Pausen kan vara minst tre månader och högst två år lång.
Under denna tid förlorar du inte rätten till invaliditetspension.
Övriga förmåner för pensionärer
Utöver pension kan FPA betala ut bostadsbidrag till pensionstagare med låga inkomster.
Mer information om bostadsbidrag för pensionstagare hittar du på FPA:s webbplats.
Till långtidssjuka eller handikappade kan FPA betala ut vårdbidrag för pensionstagare.
Fråga mer på FPA.
Rabatter för pensionärer
När du har pensionerats kan du få pensionärsrabatt till exempel på tåg-, buss- och flygresor i Finland.
De som fyllt 65 år får reserabatt genom att uppvisa sitt identitetsbevis.
En pensionär som inte har fyllt 65 år kan få rabatt genom att uppvisa sitt personbevis och sitt arbetspensionskort eller folkpensionärskort.
Kontrollera villkoren för pensionärsrabatten på biljettkontoren.
Du kan även få rabatt på exempelvis olika former av motion och kultur.
I skattedeklarationen finns uppgifter om inkomster, skatter och avdrag från föregående år.
Kontrollera uppgifterna i skattedeklarationen.
Den slutliga beskattningen fastställs utgående från uppgifterna i skattedeklarationen.
Om alla uppgifter är korrekta, och det inte saknas några uppgifter, behöver du inte göra någonting.
Om uppgifterna inte är korrekta, eller om det saknas något, komplettera och korrigera skattedeklarationen i webbtjänsten MinSkatt.
Du kan använda webbtjänsten, om du har finländska nätbankskoder eller ett mobilcertifikat.
Om du inte gör rättelserna i webbtjänsten MinSkatt, hämta pappersblanketter för rättelserna på Skatteförvaltningens webbplats eller i skattebyrån.
Skicka blanketterna per post.
Kom ihåg att kontrollera skattedeklarationen och göra de ändringar som behövs före utgången av den sista returdagen.
Beskattningsbeslut
Beskattningsbeslutet (Verotuspäätös) är en beräkning av det slutliga skattebeloppet.
På din lön eller annan inkomst har det innehållits skatt utgående från skattekortet.
Det här kallas för förskottsinnehållning (ennakonpidätys).
Förskottsinnehållningens storlek baserar sig på en uppskattning av dina inkomster.
Skattebeloppet justeras i efterskott utgående från hur stora dina inkomster och avdrag verkligen har varit.
Tillsammans med den på förhand ifyllda skattedeklarationen får du ett beskattningsbeslut.
Om du inte korrigerar skattedeklarationen, förblir det här beskattningsbeslutet i kraft.
Om du korrigerar skattedeklarationen, får du ett nytt beskattningsbeslut senare.
Kom ihåg att kontrollera också det nya beskattningsbeslutet.
Spara beskattningsbeslutet och den specifikationsdel som du fick på våren tillsammans med skattedeklarationen.
Om du beställer en ny specifikationsdel, tas det ut en avgift för den.
linkkiSkatteförvaltningen:
Skattedeklaration och beskattningsbeslutfinska _ svenska _ engelska
Avdrag
I beskattningen kan du göra avdrag (vähennykset), som minskar beskattningen.
Skatteförvaltningen gör en del avdrag automatiskt, men vissa avdrag måste du själv ansöka om.
Avdrag är till exempel:
hushållsavdrag
avdrag för resekostnader mellan bostaden och arbetsplatsen
ränteavdrag på bostadslån
Du kan avdra räntorna för bostadslånet i beskattningen då du har tagit ett lån för din stadigvarande bostad.
Du kan dra av räntorna på bostadslånet i beskattningen också då din stadigvarande bostad finns utomlands.
Om du har tagit ett lån hos en finländsk bank, får skattemyndigheten uppgifterna om lånet direkt från banken.
Om du har ett bostadslån i en utländsk bank, ska du själv ge uppgifterna om lånet till skattemyndigheten.
Du kan meddela om avdrag, när du beställer ett nytt skattekort.
Avdragen beaktas då i din skatteprocent.
Du kan också ansöka om avdrag i efterskott med skattedeklarationen.
Du får då avdragen i efterskott som en skatteåterbäring.
linkkiSkatteförvaltningen:
Avdrag vid beskattningenfinska _ svenska _ engelska
Skatteåterbäring och kvarskatt
Du ser i beskattningsbeslutet om du har betalat rätt mängd skatt.
Om du har betalat för mycket i skatt, får du skatteåterbäring (veronpalautus).
Om du har betalat för lite i skatt, blir du tvungen att betala kvarskatt (jäännösvero).
Skatteåterbäringen betalas antingen direkt på ditt bankkonto.
Meddela numret på ditt bankkonto via Skatteförvaltningens webbtjänst eller på en separat pappersblankett.
Du kan få skatteåterbäringen antingen till ett finländskt eller till ett utländsk bankkonto.
Om du blir tvungen att betala kvarskatt, får du tillsammans med beskattningsbeslutet en bankgiroblankett.
På bankgiroblanketten ser du kvarskattebeloppet, bankkontonumret, förfallodagen och referensnumret.
Du blir också tvungen att betala ränta på kvarskatten efter en viss tid.
linkkiSkatteåterbäringar:
Skatteåterbäringarfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Ange kontonummerfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Kvarskattfinska _ svenska _ engelska
Tillstånd eller anmälan
Etableringsanmälan
Försäkringar
Bokföring
Beskattning
Inkomstregistret
Arbetstagarnas inskolning och säkerhet
När du inleder företagsverksamheten har du många skyldigheter.
Du ska bland annat registrera företaget, betala skatt och ordna bokföringen.
Tillstånd eller anmälan
I Finland får man driva en laglig näring som följer god sed utan ett tillstånd som beviljas av myndigheter.
I vissa fall behövs det dock ett tillstånd från myndigheter för att starta företagsverksamhet, eller också måste man anmäla verksamheten till myndigheter.
Om du till exempel har ett företag som idkar skönhetsvård eller säljer livsmedel ska företagets lokaler kontrolleras.
Ansök om tillstånd hos kommunens hälsomyndighet innan lokalerna tas i bruk.
Innan du startar företagsverksamheten, kontrollera om du behöver tillstånd för verksamheten eller om du måste anmäla verksamheten till en myndighet.
Du kan kontrollera hos regionförvaltningsverken eller på Företagsfinlands webbplats om du behöver ett tillstånd för ditt företag.
linkkiFöretagsfinland:
Tillstånd och anmälan som är anknutna till idkandet av en näringfinska _ svenska _ engelska
linkkiFinlands Näringsliv:
Företagslagstiftningfinska
Etableringsanmälan
Ny företagsverksamhet ska anmälas till handelsregistret som upprätthålls av Patent- och registerstyrelsen (Patentti- ja rekisterihallitus).
Du kan använda samma blankett när du gör etableringsanmälan för ditt företag till Patent- och registerstyrelsen och till Skatteförvaltningen.
linkkiPatent- och registerstyrelsen:
Anmälan om grundande av ett företagfinska _ svenska _ engelska
Försäkringar
Företagarpensionsförsäkringen (FöPL) (YEL-vakuutus) är obligatorisk för företagare i åldern 18–68 år, vars företagsverksamhet inbringar minst 7 799,37 euro om året som arbetsinkomst (år 2019).
Pensionsförsäkringen tryggar företagarens utkomst då företagsverksamheten upphör på grund av invaliditet eller ålder och den ger företagarens anhöriga ett familjepensionsskydd efter att företagaren har dött.
Pensionsförsäkringar fås antingen genom försäkringsbolag eller pensionskassor (eläkekassa).
Teckna en pensionsförsäkring senast när det har gått sex månader sedan du startade företagsverksamheten.
En ny företagare får en rabatt på 22 procent på pensionspremierna under de fyra första åren.
Storleken av försäkringspremierna och pensionen beror på hur stor förvärvsinkomst (työtulo) förtagaren har.
Förvärvsinkomstens storlek inverkar också på storleken av olika inkomstrelaterade förmåner (ansiosidonnanen etuus), såsom sjukdagpenningen.
linkkiPensionsskyddscentralen:
Information om företagarpensionsförsäkringenfinska _ svenska _ engelska
Du ska teckna en pensionsförsäkring (ArPL-försäkring) (eläkevakuutus (TyEL-vakuutus)) och en olycksfallsförsäkring som omfattar en grupplivförsäkring och en arbetslöshetsförsäkring för de anställda.
Arbetsgivaren betalar arbetstagarens socialskyddsavgifter till skattemyndigheten i anslutning till skatteinnehållningen.
I vissa branscher finns också andra obligatoriska försäkringar.
Du bör också överväga andra frivilliga försäkringar som till exempel företagarens olycksfallsförsäkring.
linkkiPensionsskyddscentralen:
Information om att teckna försäkringar för anställdafinska _ svenska _ engelska
linkkiFöretagsFinland:
Information om att teckna försäkringar för anställdafinska _ svenska _ engelska
Bokföring
I Finland har alla företagare bokföringsskyldighet.
Om du inte vill sköta bokföringen själv, kan du anlita en revisionsbyrå som sköter företagets bokföring åt dig.
I Finland anlitar många företag revisionsbyråer.
Beskattning
Företagsformen påverkar företagets beskattning.
Detta är det bra att beakta när du väljer företagsform.
En ny företagare kan anmäla sig till Skatteförvaltningens förskottsuppbördsregister.
Anmälan till förskottsuppbördsregistret görs med samma anmälan som görs för grundande av företaget, d.v.s. etableringsanmälan (yrityksen perustamisilmoitus).
Om ditt företag är i förskottsuppbördsregistret kan du fakturera kunder utan förskottsinnehållning.
Skatter betalas på de inkomster som företagaren eller företaget har kvar när alla kostnader för företagsverksamheten har dragits av försäljningen.
Företagets skatter betalas på basis av de beskattningsbara inkomsterna, vars belopp man uppskattar på förhand.
Uppskattningen baseras på beloppet av de beskattningsbara inkomsterna året innan.
I ett nytt företag uppskattar företagaren själv storleken av den beskattningsbara inkomsten och meddelar denna till skattmyndigheten.
linkkiSkatteförvaltningen:
Information om beskattningen av företag och företagarefinska _ svenska _ engelska
linkkiFöretagsFinland:
Information om beskattningen av företag och företagarefinska _ svenska _ engelska
Mervärdesskatt
Mervärdesskatten (arvonlisävero) är en konsumtionsskatt som i Finland betalas för nästan alla varor och tjänster.
Företagare som säljer varor och tjänster i Finland är skyldiga att betala mervärdesskatt.
Om inkomsten som man får för försäljningen av varor och tjänster är mindre än 10 000 euro per år, behöver ingen mervärdesskatt betalas på den.
Företagsformen påverkar inte mervärdesskattens belopp.
Mervärdesskattebeloppet varierar emellertid för olika produkter.
Inkomstregistret
Inkomstregistret är en databas dit arbetsgivarna anmäler lönerna som de utbetalat till sina anställda.
Anmälan ska göras senast fem dagar efter löneutbetalningen.
Uppgifterna ska skickas till inkomstregistret elektroniskt:
direkt via lönesystemet om det har en inbyggd teknisk förbindelse till Inkomstregistret eller
via Inkomstregistrets ärendehantering, till vilken man får tillträde med webbankkoder eller andra medel för elektronisk identifiering.
Löneuppgifterna kan endast i undantagsfall anmälas med ett pappersformulär.
Läs mer om Inkomstregistret och om att anmäla löner på Inkomstregistrets webbplats.
linkkiSkatteförvaltningen:
Inkomstregistretfinska _ svenska _ engelska _ ryska _ estniska _ kinesiska
Arbetstagarnas inskolning och säkerhet
Som företagare har du ansvaret för att ge arbetstagarna inskolning i arbetsuppgifterna.
Arbetsgivaren ska introducera förhållandena på arbetsplatsen och de rätta arbetsmetoderna för arbetstagaren.
Arbetsgivaren är också skyldig att sörja för arbetstagarnas säkerhet och hälsa i arbetet.
Arbetsgivaren ska utarbeta ett verksamhetsprogram för arbetarskyddet (työsuojelun toimintaohjelma) som tar upp de säkerhets- och hälsorelaterade riskerna på arbetsplatsen och hur man undgår dem.
Läs mer om att vara arbetsgivare på InfoFinlands sida Arbetsgivarens rättigheter och skyldigheter.
linkkiArbetarskyddscentralen:
Information om arbetarskyddfinska _ svenska _ engelska
Vem är berättigad till utkomstskydd för arbetslösa?
Du kan registrera dig som arbetssökande vid TE-byrån om
du har ett uppehållstillstånd som ger dig rätt att arbeta i Finland
ditt uppehållstillstånd inte begränsar vilken arbetsgivare du får arbeta för
eller
du är medborgare i ett EU-land, ett EES-land eller Schweiz
du är familjemedlem till en medborgare i ett EU-land, ett EES-land eller Schweiz
Då du registrerat dig som arbetssökande har du rätt till arbetslöshetsunderstöd om du
är 17–64 år gammal
är arbetslös och anmäld som arbetssökande vid TE-byrån
söker heltidsarbete
är arbetsförmögen och tillgänglig på arbetsmarknaden
uppfyller villkoren för inkomstrelaterad dagpenning, grunddagpenning eller arbetsmarknadsstöd.
För att få utkomstskydd för arbetslösa måste du aktivt söka jobb och vara beredd att ta emot ett jobb.
Du ska också ingå en sysselsättnings- och integrationsplan med TE-byrån och delta i de tjänster och åtgärder som TE-byrån erbjuder åt dig.
På full arbetslöshetsförmån ställs även andra villkor.
Du kan få full arbetslöshetsförmån om du under 65 betalningsdagar, alltså under cirka tre månaders tid, utför en viss mängd lönearbete, får inkomst som företagare eller deltar i en verksamhet eller en tjänst som främjar din sysselsättning.
Detta kallas för aktiveringsmodellen för arbetslöshetsförsäkringen (työttömyysturvan aktiivimalli).
Arbetslöshetsförmånerna är den inkomstrelaterade dagpenningen, grunddagpenningen och arbetsmarknadsstödet.
Skatt betalas på alla arbetslöshetsförmåner.
linkkiArbets- och näringsministeriet:
Om du blir arbetslösfinska _ svenska _ engelska
linkkiArbets- och näringsministeriet:
Utkomstskydd för arbetslösafinska _ svenska _ engelska
Information om utkomstskyddet för arbetslösafinska _ svenska _ engelska
linkkiArbets- och näringsministeriet:
Rådgivning om utkomstskydd för arbetslösafinska _ svenska _ engelska _ ryska
Aktiveringsmodellen för arbetslöshetsförsäkringen finska _ svenska _ engelska
Inkomstrelaterad dagpenning
Du kan få inkomstrelaterad dagpenning om du
registrerat dig som arbetslös arbetssökande vid arbets- och näringsbyrån
hör till en finländsk arbetslöshetskassa
uppfyller arbetsvillkoret, d.v.s. har arbetat tillräckligt länge före arbetslösheten
har varit medlem i arbetslöshetskassan i minst 26 veckor innan du blev arbetslös.
Den inkomstrelaterade dagpenningen beviljas och utbetalas av den arbetslöshetskassa där du är medlem.
Den inkomstrelaterade dagpenningen beräknas utgående från storleken på den lön som du hade innan du blev arbetslös.
Vanligtvis kan inkomstrelaterad dagpenning fås under 400 dagar. Undantag från detta är följande situationer:
Om du har arbetat i sammanlagt tre år eller mindre, kan du få inkomstrelaterad dagpenning i högst 300 dagar.
Om du har fyllt 58 år innan du blev arbetslös, kan du få inkomstrelaterad dagpenning i mindre än 500 dagar.
Läs mer om arbetslöshetskassan på InfoFinlands sida Fackförbund.
Information om den inkomstrelaterade dagpenningenfinska _ svenska _ engelska
Grunddagpenning
Du kan få grunddagpenning om du omfattas av den sociala tryggheten i Finland utifrån permanent boende eller arbete före arbetslösheten och
registrerat dig som arbetslös arbetssökande vid arbets- och näringsbyrån
uppfyller arbetsvillkoret, d.v.s. har arbetat tillräckligt länge före arbetslösheten
inte uppfyller villkoren för inkomstrelaterad dagpenning.
Grunddagpenningen beviljas och utbetalas av Fpa.
Vanligtvis kan du få grunddagpenning i mindre än 400 dagar. Undantag från detta är följande situationer:
Om du har arbetat i sammanlagt tre år eller mindre, kan du få grunddagpenning i högst 300 dagar.
Om du har fyllt 58 år innan du blev arbetslös, kan du få grunddagpenning i mindre än 500 dagar.
Om du får andra sociala förmåner eller arbetsinkomster under arbetslösheten, är din grunddagpenning mindre.
Grunddagpenningfinska _ svenska _ engelska
Arbetsmarknadsstöd
Du kan få arbetsmarknadsstöd om du
registrerat dig som arbetslös arbetssökande vid arbets- och näringsbyrån
bor permanent i Finland
inte uppfyller arbetsvillkoret, d.v.s. inte arbetat tillräckligt länge innan du blev arbetslös eller fått förvärvsrelaterad dagpenning eller grunddagpenning under maximitiden.
Om du har en gällande integrationsplan, kan du söka arbetsmarknadsstöd för den tid då du deltar i utbildningar och annan verksamhet som nedtecknats i planen.
Närmare uppgifter om integrationsplanen finns på InfoFinlands sida Integration i Finland.
Arbetsmarknadsstödet beviljas och utbetalas av Fpa.
Arbetsmarknadsstödet är behovsprövat.
Det betyder att till exempel sociala förmåner och lön minskar arbetsmarknadsstödets belopp.
Om du är under 25 år, kontrollera tilläggsvillkoren för arbetsmarknadsstödet för unga på TE-tjänsternas webbplats.
Arbetsmarknadsstödfinska _ svenska _ engelska
Du behöver ett skattekort (verokortti), om du får lön eller har andra inkomster i Finland.
På skattekortet finns en anteckning om skatteprocenten (veroprosentti).
Av det ser arbetsgivaren, hur mycket skatt som ska betalas på lönen.
Skatteprocenten beror på hur hög din inkomst är.
Om du håller på att flytta till Finland, får du skattekortet från skattebyrån (verotoimisto).
Uppskatta för skattekortet, hur stora dina inkomster kommer att bli för hela skatteåret.
Du behöver också en finländsk personbeteckning.
Du får personbeteckningen, när du registrerar dig som invånare hos magistraten.
Du kan få en personbeteckning också från skattebyrån.
Läs mer på sidan Registrering som invånare.
När du bor i Finland stadigvarande, skickar Skatteförvaltningen ett nytt skattekort till dig varje år i januari.
Skatteförvaltningen räknar ut en lämplig skatteprocent åt dig utgående från hur mycket du förtjänade året innan.
Förete skattekortet till din arbetsgivare.
Om du inte företer skattekortet till din arbetsgivare, innehåller arbetsgivaren en skatt på 60 % på din lön.
Om dina inkomster blir mindre eller större under året, ska du beställa ett nytt skattekort.
Du får ett nytt skattekort:
från Skatteförvaltningens webbtjänst MinSkatt
på skattebyrån
Du kan även beställa skattekortet via Skatteförvaltningens telefontjänst:
finska 029 497 000
svenska 029 497 001
engelska 029 497 050
När du söker ett nytt skattekort, behöver du följande uppgifter:
en uppskattning av dina inkomster för hela året
de inkomster som du har haft från början av året
de skatter som har betalats på dina inkomster från början av året
uppgift om de avdrag som du söker i beskattningen för innevarande år
Om du betalar för mycket skatt, får du skatteåterbäring.
Om du betalar för litet i skatt, blir du tvungen att betala kvarskatt.
linkkiSkatteförvaltningen:
Nytt skattekortfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Hur beräknas skatteprocenten?finska _ svenska _ engelska
Om du har flera arbetsgivare
Om du har flera arbetsgivare ska du förete ditt skattekort till dem alla.
Du kan använda samma skattekort hos alla arbetsgivarna.
Du betalar samma skatt hos alla dina arbetsgivare.
På skattekortet anges en inkomstgräns och din skatteprocent beräknas utifrån den.
Kom ihåg att hålla ett öga på dina inkomster.
Om du får mer lön än vad du uppgett, överskrids din inkomstgräns.
Om inkomstgränsen överskrids ska du beställa ett nytt skattekort.
Skattenummer
Du behöver en skattenummer (veronumero), om du arbetar på en bygg- eller monteringsarbetsplats i Finland.
Med hjälp av skattenumret kontrolleras, att alla arbetstagare finns i Skatteförvaltningens register.
Skattenumret ska framgå av den fotoförsedda namnskylt som du får av din arbetsgivare.
Du får inte arbeta på en byggplats utan namnskylt.
Du får skattenumret från skattebyrån samtidigt som du går efter skattekortet.
Om du redan har finländsk personbeteckning och ett skattekort, hittar du skattenumret på ditt skattekort.
linkkiSkatteförvaltningen:
Skattenummerfinska _ svenska _ engelska
När du grundar ett företag måste du välja företagsform och ett namn för företaget samt definiera branschen.
På valet av företagsform inverkar bland annat antalet grundare, behovet av kapital, fördelningen av ansvar och bestämmanderätt, finansieringen och beskattningen.
Olika företagsformer i Finland är enskild näringsidkare (toiminimi); öppet bolag (avoin yhtiö); kommanditbolag (kommandiittiyhtiö); aktiebolag (osakeyhtiö) och andelslag (osuuskunta).
När du funderar på vilken företagsform du ska välja, är det absolut tillrådligt att du kontaktar företagsrådgivningen.
linkkiNyföretagarcentralerna i Finland:
Företagsrådgivningfinska _ svenska _ engelska
Enskild näringsidkare (toiminimi)
Det enklaste och vanligaste sättet att starta företagsverksamhet är att som enskild näringsidkare driva en firma.
Du har bestämmanderätt över och ansvar för firmans ärenden och företaget kan anställa medarbetare precis som andra företag.
Företagsverksamhet som bisyssla lönar det sig ofta att starta som enskild näringsidkare.
Det är snabbt och enkelt att starta företagsverksamhet som enskild näringsidkare.
Aktiebolaget är den vanligaste företagsformen i Finland.
Ett aktiebolag passar för all slags affärsverksamhet.
Du kan grunda ett aktiebolag antingen själv eller tillsammans med andra delägare.
Delägarens rösträtt, avkastning och ansvar i bolaget beror på hur många aktier i bolaget hen äger.
Ett öppet bolag bildas då två eller fler personer kommer överens om att grunda ett bolag genom att teckna ett bolagsavtal.
Bolagsmännen, d.v.s. personerna som tillsammans äger bolaget, är jämställda i all verksamhet som bolaget driver och de ansvarar tillsammans och personligen för bolagets beslut, förbindelser och skulder.
Ett kommanditbolag är ett personbolag som skiljer sig från ett öppet bolag på så sätt att det i kommanditbolaget finns utöver en eller flera ansvariga bolagsmän åtminstone en tyst bolagsman, d.v.s. en person som är delägare i företaget. Vanligen är den tysta bolagsmannen en investerare.
Det behövs minst tre personer för att grunda ett andelslag.
Ett andelslag kan ha en eller fler medlemmar.
Ett andelslag är ett företag som ägs av medlemmarna.
På andelslagets stämma har varje medlem en röst. Medlemmarna ansvarar för andelslagets förpliktelser (till exempel skulder) endast med det belopp som de investerat i andelslaget.
linkkiFöretagsFinland:
Information om företagsformerfinska _ svenska _ engelska
Anmäl dig som arbetslös arbetssökande
Om du blir arbetslös ska du anmäla dig hos TE-byrån senast den första dagen av din arbetslöshet.
Om du omfattas av den finländska sociala tryggheten kan du ansöka om arbetslöshetsstöd.
Du kan få arbetslöshetsstöd från och med det datum då du anmälde dig som arbetslös.
Kom ihåg att anmäla dig också direkt efter studier, arbetskraftsutbildning eller en period med sysselsättningsstöd.
Anmäl dig som arbetssökande i TE-byråns webbtjänst.
Logga in med finländska nätbankskoder eller personkort med microchip.
En anställd vid TE-byrån tar kontakt med dig om det behövs ytterligare uppgifter.
Du behöver inte ringa eller besöka TE-byrån om du inte uttryckligen ombes göra detta.
Om du saknar nätbankskoder eller personkort med microchip ska du anmäla dig som arbetssökande vid närmaste TE-byrå.
Endast medborgare i EU-länderna, Norge, Island, Liechtenstein och Schweiz kan anmäla sig som arbetssökande i webbtjänsten.
Om du är medborgare i ett annat land måste du besöka arbets- och näringsbyrån.
När du går till TE-byrån ska du ta med dig
alla dina arbetsintyg och studiebetyg
ditt pass där ditt uppehållstillstånd syns
TE-byrån undersöker uppgifterna som du lämnar.
Det finns vissa villkor för att få utkomstskydd för de arbetslösa och TE-byrån utreder om dessa villkor uppfylls i din situation.
Därefter ger TE-byrån ett utlåtande i ärendet till den instans som betalar förmånen, det vill säga till arbetslöshetskassan eller FPA.
Du kan fråga råd i ärenden som rör utkomstskyddet för arbetslösa vid din egen TE-byrå.
Du kan också ringa TE-tjänsternas rådgivning om utkomstskydd för arbetslösa:
på finska: 0295 020 701
på svenska: 0295 020 711
på engelska: 0295 030 713
på ryska: 0295 020 715
Läs också InfoFinlands sida:
Arbetslöshetsförsäkring
linkkiArbets- och näringsministeriet:
Om du blir arbetslösfinska _ svenska _ engelska
linkkiArbets- och näringsministeriet:
Att anmäla sig som arbetslös arbetssökandefinska _ svenska
linkkiArbets- och näringsministeriet:
Rådgivning om utkomstskydd för arbetslösafinska _ svenska _ engelska _ ryska
Semester, studier eller arbete under arbetslösheten
Om du börjar arbeta eller studera när du är arbetslös ska du meddela detta till TE-byrån.
Du får anvisningar om hur detta påverkar ditt utkomststöd för arbetslösa.
Om du reser i hemlandet eller utomlands ska du se till att du alltid kan nås.
Lämna till exempel ditt telefonnummer och din adress till TE-byrån och ange hur länge du ämnar vistas på resmålet.
Du kan ändå inte tacka nej till ett jobb som erbjuds till dig på grund av en utlandsresa.
Om du startar ett företag när du är arbetslös, kan du få arbetslöshetsförmån under de fyra första månaderna.
Karens
Du kan förlora din rätt till arbetslöshetsdagpenning för en viss tid om du själv har förorsakat arbetslösheten.
Du kan sättas i karens till exempel om:
du inte söker ett jobb som TE-byrån föreslår för dig
du inte tar emot ett jobb som erbjuds till dig
du säger upp dig från ditt jobb utan en godtagbar anledning
Karenstidens längd varierar från 15 dagar till 90 dagar.
Längden beror på orsaken till karensen.
I vissa fall kan du förlora rätten till utkomststöd för arbetslösa tillsvidare.
I Finland betalar du inkomstskatt (tulovero) på lön.
Du betalar också skatt på till exempel följande inkomster:
arbetsersättning
företagsinkomst
arbetslöshetsdagpenning
föräldradagpenning
pensioner
studiestöd
För skattepengarna betalar staten och kommunerna till exempel:
hälsovård
utbildning
dagvård
försvar
I Finland är beskattningen progressiv.
Det innebär att man på en stor lön betalar en större andel skatt än på en mindre lön.
Skatteprocenten (Veroprosentti) beräknas i Finland för var och en separat.
Din makes/makas inkomster inverkar inte på din skatteprocent.
Du kan uppskatta din skatteprocent med Skatteförvaltningens skatteräknare.
Arbetsgivaren betalar skatterna direkt från din lön.
För att kunna göra det behöver arbetsgivaren ett skattekort av dig.
Skatt som betalas direkt från lönen, är förskottsskatt (ennakonpidätys).
Skatteförvaltningen räknar efter varje år om du har betalat tillräckligt med skatt på dina inkomster.
Om du har betalat för mycket i skatt, får du skatteåterbäring (veronpalautus).
Om du har betalat för lite i skatt, blir du tvungen att betala kvarskatt (jäännösvero).
Läs mer på sidan: Skattedeklaration och beskattningsbeslut.
Kontrollera i lönespecifikationen och skattedeklarationen (veroilmoitus), att arbetsgivaren har betalat skatt på din lön.
Spara lönekvittona.
Om skatten inte har betalats, blir du tvungen att betala den i efterskott.
Utöver skatt betalar arbetsgivaren försäkringspremier på din lön i händelse av arbetslöshet eller sjukdom.
linkkiSkatteförvaltningen:
Information om beskattningenfinska _ svenska _ engelska
linkkiSkattemyndigheten:
Skattekortfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Att beställa skattekort finska _ svenska _ engelska
linkkiSkatteförvaltningen:
Skatteprocenträknarefinska _ svenska _ engelska
Beskattningen när du börjar arbeta i Finland
Om du kommer till Finland för att arbeta, beror din beskattning på hur länge du vistas i Finland.
På beskattningen inverkar också huruvida din arbetsgivare är ett finländskt eller ett utländskt företag.
Om du vistas i Finland i mer än sex månader, ska du i allmänhet betala skatt på din lön till Finland.
Du ska i allmänhet också betala de obligatoriska försäkringspremierna till Finland.
Du behöver en finländsk personbeteckning och ett finländskt skattekort.
Skatteprocenten räknas på inkomsterna för hela året.
Du får skatteavdrag på samma grunder som andra som bor i Finland stadigvarande.
Om du vistas i Finland i högst sex månader och din arbetsgivare är ett utländskt företag, behöver du i allmänhet inte betala skatt till Finland.
Om din arbetsgivare är finländare eller om din utländska arbetsgivare har en arbetsplats i Finland, betalar du skatt i Finland.
Du kan söka progressiv beskattning, om du bor i ett land som hör till Europeiska ekonomiska samarbetsområdet eller i en stat, med vilken Finland har ett skatteavtal.
I annat fall betalar du en källskatt (lähdevero) på 35 % på lönen och du behöver ett källskattekort.
Källskattekort måste du ansöka med en pappersblankett.
För progressiv beskattning behöver du ett skattekort för begränsat skattskyldiga (rajoitetusti verovelvollisen verokortti).
Du får ett sådant på skattebyrån.
Du kan söka progressiv beskattning också i efterskott.
Du blir också tvungen att betala försäkringspremier, om du inte är försäkrad i det land där du bor stadigvarande.
Om du redan är försäkrad i ett annat land, behöver du ett intyg A1/E101 över försäkringen.
När du flyttar bort från Finland, kom ihåg att göra en flyttningsanmälan till magistraten.
Du får då din skattedeklaration till rätt adress.
När du håller på att flytta till Finland, får du ytterligare information i avsnittet Flytta till Finland.
linkkiSkatteförvaltningen:
Arbeta i Finlandfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Ansökan om progressiv inkomstbeskattningfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Utländsk hyrd arbetskraft och beskattningen i Finlandfinska _ svenska _ engelska
Flyttanmälanfinska _ svenska _ engelska
Uppehållstillstånd eller registrering av uppehållsrätt?
Kom på en affärsidé
Gör en affärsverksamhetsplan
Fråga om råd på företagsrådgivningen
Ordna finansiering
Välj företagsform
Du kan grunda ett företag i Finland oavsett ditt medborgarskap.
Det viktiga är att du har uppehållsrätt i Finland, de yrkeskunskaper som krävs och tillräckliga kunskaper i finska.
Uppehållstillstånd eller registrering av uppehållsrätt?
Om du är medborgare i ett nordiskt land och flyttar till Finland ska du registrera dig vid magistraten.
Du behöver inget uppehållstillstånd i Finland.
Läs mer på InfoFinlands sida Nordisk medborgare.
Om du är medborgare i något EU-land, Liechtenstein eller Schweiz och flyttar till Finland permanent, ska du registrera dig vid Migrationsverket och magistraten.
Läs mer på InfoFinlands sida EU-medborgare.
Om du är medborgare i något land som inte tillhör EU och flyttar till Finland som företagare, behöver du antingen ett uppehållstillstånd för företagare, ett uppehållstillstånd för arbetstagare eller ett uppehållstillstånd för uppstartsföretagare.
Läs mer på InfoFinlands sida Till Finland som företagare.
Som företagare till Finland:
Vilka tillstånd behöver du?(pdf, 384 kt)finska _ engelska
Tillstånd och anmälningar för utländska företagarefinska _ svenska _ engelska
Kom på en affärsidé
Processen för att grunda ett företag är likadant som för finska medborgare.
När du vill grunda ett företag ska du noga fundera på om du har en bra affärsidé.
Fundera också på om du har tillräckliga yrkeskunskaper och erfarenhet.
Det är viktigt att du känner väl till din bransch och de lagar som styr företagande.
Det är också viktigt att känna till sina kunder och försäljningsmetoder.
Kom ihåg att företagande även medför risker.
Tillräcklig finansiering och noggrann planering är nödvändiga.
linkkiFöretagsfinland:
Att grunda ett företagfinska _ svenska _ engelska
Gör en affärsverksamhetsplan
I affärsverksamhetsplanen funderar du på styrkorna och svagheterna i ditt kunnande och egenskaperna hos den produkt, vara eller tjänst som du erbjuder.
Fundera på vilka som är dina kunder och vilka önskemål de har.
Fundera också på vilka som är dina konkurrenter och hurdana produkter och verksamhetssätt de har.
Den viktigaste delen i affärsverksamhetsplanen är verksamhetsplanen för ditt eget företag.
Fundera noga hur företaget drivs och var och hurdana lokaler företaget har.
Fundera på vilka produktionsmedel eller vilken arbetskraft du behöver.
Vilka reklammedel ska du använda för att främja försäljningen?
Ta också reda på om försäkringar täcker de risker som förknippas med verksamheten.
Fundera också på hur du ordnar bokföringen och planerar ekonomin.
Hur avser du följa upp hur dina planer förverkligas?
Anteckna allt detta i din affärsverksamhetsplan.
Hjälp med att upprätta en affärsverksamhetsplan
Du får närmare anvisningar om hur du upprättar en affärsverksamhetsplan vid företagsrådgivningscentra.
På deras webbplatser kan du även ladda ned företagarguider åtminstone på finska och engelska.
Där får du även en mall för affärsverksamhetsplanen och andra dokumentmallar.
Guide om att grunda ett företagfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ turkiska _ kinesiska _ arabiska
Fråga om råd på företagsrådgivningen
I Finland har alla möjlighet att få kostnadsfri företagsrådgivning.
Rådgivning erbjuds vid till exempel:
Nyföretagarcentraler
Närings-, trafik- och miljöcentralerna (NTM-centralerna)
Arbets- och näringsbyråer (TE-byråer)
FöretagsFinland (via webbplatsen och per telefon)
När du får en bra affärsidé, kontakta närmaste företagsservicecenter.
Där hjälper experterna dig att utveckla affärsidén, göra en marknadsundersökning, beräkna lönsamheten och kartlägga finansieringen.
Du får även stöd när du funderar på om du ska starta ett företag.
Företagsrådgivning fås på finska och svenska och åtminstone i de större städerna även på engelska.
Ibland kan det finnas möjlighet att få rådgivning även på något annat språk.
linkkiFöretagsFinland:
Företagsrådgivningfinska _ svenska _ engelska
Företagarkurser
Olika instanser ordnar företagarkurser och informationsmöten som är mycket nyttiga för dig som ska grunda ett företag.
På kurserna behandlas till exempel upprättande av affärsverksamhetsplan, start av företagsverksamheten, bokföring, företagsbeskattning, juridiska frågor, marknadsföring, försäljning och kundtjänst.
Ordna finansiering
Planera företagets finansiering noga innan du grundar företaget.
Det är viktigt att du har tillräckligt stort kapital i början.
En del av företagets finansiering kan bestå av en gåva eller ett lån.
När du ansöker om finansiering måste du ha en ordentlig affärsverksamhetsplan färdig.
Lån
Banker och Finnvera beviljar lån till företagare som startar ett företag.
Finnvera är ett finansieringsbolag som ägs av finska staten.
Det ger lån till nya företag och redan aktiva företag.
Om ditt företag har förutsättningarna för en lönsam verksamhet men du inte har tillräckligt mycket pengar eller säkerheter för att få ett banklån, ska du fråga om du kan få ett lån eller borgen hos Finnvera.
linkkiFöretagsFinland:
Finansiering för ett företagfinska _ svenska _ engelska
linkkiFinnvera:
Finansiering för ett företagfinska _ svenska _ engelska
Startpenning
När du blir företagare, kan du få startpenning för att trygga försörjningen när företagsverksamheten precis har börjat.
Du ansöker om startpenning vid den arbets- och näringsbyrå där du är kund.
Du kan få startpenning för högst tolv månader.
När du ansöker om startpenning utreder arbets- och näringsbyrån om företagande är ett lämpligt alternativ för dig.
Du kan få startpenning om
du är arbetslös arbetssökande
du inte är arbetslös, men går från till exempel lönearbete, studier eller hemmaarbete till företagare
du har företagande som bisyssla och utvidgar företagsverksamheten till din huvudsyssla.
Förutsättningar för att få startpenning är till exempel:
företagande som huvudsyssla
tillräckliga kunskaper, färdigheter och resurser för den företagsverksamhet som du planerar
arbets- och näringsbyrån uppskattar att företagsverksamheten kan vara lönsam
du behöver startpenningen för din försörjning
Företagsverksamheten startas först när stödet har beviljats.
Om du avser ansöka om startpenning ska du kontakta arbets- och näringsbyrån i ett så tidigt skede som möjligt.
Det finns även andra stödformer för nya företagare.
FöretagsFinland ger dig information om olika finansieringsalternativ.
linkkiArbets- och näringsministeriet:
Information om startpengenfinska _ svenska _ engelska
Välj företagsform
När du ska grunda ett företag, måste du välja företagsform och ett namn för företaget samt ange bransch.
När du väljer företagsformen ska du beakta bland annat antalet grundare, behovet av kapital, fördelningen av ansvar och beslutsmakt samt finansiering och beskattning.
Olika företagsformer i Finland är firma, öppet bolag, kommanditbolag, aktiebolag och andelslag.
När du funderar på vilken företagsform du ska välja, är det absolut tillrådligt att du kontaktar företagsrådgivningen.
Läs mer på InfoFinlands sida Företagsformer.
Arbetsgivaren har rätt att:
anställa en arbetstagare
leda arbetet och ge råd och utfärda bestämmelser som ansluter till utförandet av arbetet
säga upp och häva ett arbetsavtal inom ramen för begränsningarna i lag
Arbetsgivaren har skyldighet att:
följa lagar och avtal
behandla arbetstagarna jämlikt oavsett deras härkomst, religion, kön, ålder eller politiska åsikt
sörja för arbetstagarnas säkerhet och arbetshälsa
ge arbetstagaren en skriftligt utredning om de centrala villkoren i arbetet
främja ett gott arbetsklimat, arbetstagarens arbetsprestationer och yrkesutveckling
Kollektivavtal
Arbetsgivaren måste följa kollektivavtalet.
Han eller hon kan till exempel inte betala ut en mindre lön än vad som fastställts i kollektivavtalet.
Inkomstregistret
Inkomstregistret är en databas dit arbetsgivarna anmäler lönerna som de utbetalat till sina anställda.
Anmälan ska göras senast fem dagar efter löneutbetalningen.
Uppgifterna ska skickas till inkomstregistret elektroniskt:
direkt via lönesystemet om det har en inbyggd teknisk förbindelse till Inkomstregistret eller
via Inkomstregistrets ärendehantering, till vilken man får tillträde med webbankkoder eller andra medel för elektronisk identifiering.
Löneuppgifterna kan endast i undantagsfall anmälas med ett pappersformulär.
Läs mer om Inkomstregistret och om att anmäla löner på Inkomstregistrets webbplats.
linkkiSkatteförvaltningen:
Inkomstregistretfinska _ svenska _ engelska _ ryska _ estniska _ kinesiska
Olycksfallsförsäkring
Arbetsgivaren ska teckna en olycksfallsförsäkring (tapaturmavakuutus) åt sina anställda.
Detta ska alltid göras när en anställning börjar.
Arbetstagaren kan få ersättning vid ett olycksfall.
Ersättningen kan vara en ersättning av sjukvårdskostnader och inkomstbortfall i form av dagpenning, olycksfallspension, ersättning för den skada som olyckan har orsakat, rehabilitering eller vid dödsfall familjepension till de anhöriga.
Arbetsgivaren kan utöver de lagstadgade försäkringarna även teckna olika frivilliga försäkringar åt sina anställda.
Det är bra att klarlägga med arbetsgivaren vilka försäkringar han eller hon har tecknat åt sina anställda.
Arbetsintyg
När en anställning upphör har den anställda rätt att få ett skriftligt arbetsintyg av arbetsgivaren.
Läs mer på InfoFinlands sida Arbetsintyg.
Intressebevakning och rådgivning för företagare
Företagarens utkomstskydd för arbetslösa
Företagarens företagshälsovård
Om en företagare blir sjuk
Intressebevakning och rådgivning för företagare
Finlands Näringsliv EK representerar alla privata branscher och företag i alla storlekar.
Branschförbunden är intressebevakningsorganisationer för företag i olika branscher.
De tillhandahåller sina medlemsföretag ofta också många slags tjänster såsom rådgivning i frågor som rör företagande och den aktuella branschen.
linkkiFinlands Näringsliv EK:
Intressebevakning för företagarefinska _ svenska _ engelska
Företagarna i Finland (Suomen Yrittäjät) är företagarnas intressebevakningsorganisation som också producerar sina medlemmar olika tjänster, som till exempel gratis telefonrådgivning i frågor som rör företagande.
linkkiFöretagarna i Finland:
Intressebevakning för företagarefinska _ svenska _ engelska
TE-byrån tillhandahåller tjänster som stöder utvecklingen av affärsverksamheten.
Via TE-byrån kan du även leta en fortsättare för din företagsverksamhet eller en partner till ditt företag.
Nyföretagarcentraler erbjuder kostnadsfri företagsrådgivning runtom i Finland.
Hos företagsrådgivningen kan du få hjälp med frågor kring företagets verksamhet eller utveckling.
linkkiNyföretagarcentralerna i Finland:
Företagsrådgivningfinska _ svenska _ engelska
Företagsfinland erbjuder en gratis telefontjänst där du får sakkunnig rådgivning om ditt företag har ekonomiska svårigheter.
Rådgivning ges på finska och svenska.
Ekonomihjälp-rådgivningen
på finska, tfn 029 502 4880
på svenska, tfn 029 502 4881
Tjänsten har öppet måndag till fredag kl. 9.00–16.00.
linkkiFöretagsFinland:
Ekonomisk rådgivning för företagarefinska _ svenska
Företagarens utkomstskydd för arbetslösa
Också företagaren har rätt till utkomstskydd för arbetslösa.
En företagare är arbetslös när han eller hon har lagt ned sin företagsverksamhet eller sålt sin andel av företaget.
Företagandet kan också upphöra om företaget säljs, avvecklas, går i konkurs, försätts i likvidation eller på grund av skilsmässa.
Företagaren betraktas som arbetslös också om man har haft ett uppehåll på minst fyra månader i företagsverksamheten.
Om du måste lägga ned din företagsverksamhet, ska du omgående anmäla dig som arbetslös arbetssökande via TE-byråns webbtjänst.
Du kan få arbetslöshetsersättning tidigast från den dag då du gjort anmälan vid TE-byrån.
Information om företagarens sociala trygghetfinska _ svenska _ engelska
Om du vill få inkomstrelaterat utkomstskydd för arbetslösa, ska du ansluta dig som medlem i företagarnas arbetslöshetskassa (yrittäjien työttömyyskassa).
Om din företagsverksamhet upphör, kan du ansöka om inkomstrelaterad dagpenning (ansiosidonnainen päiväraha) vid arbetslöshetskassan.
Du kan få inkomstrelaterad dagpenning från företagarnas arbetslöshetskassa om du har bedrivit företagsverksamhet och varit medlem i kassan tillräckligt länge innan du blev arbetslös.
Den inkomstrelaterade dagpenningen är större än grunddagpenningen eller arbetsmarknadsstödet.
Hur stor inkomstrelaterad dagpenning du får beror på hur stora förvärvsinkomster du angett som grund för arbetslöshetsförsäkringen.
linkkiFöretagarnas Arbetslöshetskassa i Finland:
Företagarnas Arbetslöshetskassa i Finlandfinska _ svenska
linkkiYrkesutövarnas och företagarnas arbetslöshetskassa:
Yrkesutövarnas och företagarnas arbetslöshetskassafinska _ svenska _ engelska _ ryska _ estniska
Grunddagpenning
Fpa kan betala grunddagpenning (peruspäiväraha) för en arbetslös företagare som inte är medlem i en arbetslöshetskassa.
Om du uppfyller arbetsvillkoret för företagare och omfattas av den sociala tryggheten i Finland kan du få grunddagpenning.
På FPA:s webbplats finns en räknare som du kan använda för att beräkna om du uppfyller arbetsvillkoret för företagare.
Arbetsmarknadsstöd
Om du inte har rätt till grunddagpenning eller inkomstrelaterad dagpenning, men omfattas av den sociala tryggheten i Finland, kan du ansöka om arbetsmarknadsstöd.
Arbetsmarknadsstödet är behovsprövat, vilket betyder att dina andra inkomster och din situation som en helhet påverkar dess belopp.
Företagarens företagshälsovård
En företagare och andra som arbetar åt sig själv kan ordna företagshälsovård för sig själv om de så önskar.
Företagare måste inte ordna företagshälsovård för sig själv, men däremot måste de ordna det för sina anställda.
Företagshälsovård kan ordnas på den lokala hälsovårdscentralen (terveyskeskus) eller till exempel en privat läkarstation.
Läs mer på InfoFinlands sida Företagshälsovård.
Information för företagare om företagshälsovårdenfinska _ svenska _ engelska
Om en företagare blir sjuk
Om du blir sjuk, kan du få sjukdagpenning (sairauspäiväraha) från Fpa. Den ersätter inkomstbortfallet på grund av arbetsoförmåga när arbetsoförmågan varar mindre än ett år.
Betalningen av dagpenning inleds efter en självrisktid (omavastuuaika).
För företagare är självrisktiden oftast dagen för insjuknandet och följande tre vardagar.
Företagarens sjukdagpenningfinska _ svenska _ engelska
Var får jag hjälp med problem i arbetslivet?
Prata först med din chef.
Om det inte hjälper, kontakta arbetsplatsens förtroendeman.
Om det inte finns en förtroendeman på arbetsplatsen och du är medlem i facket, kontakta ditt fackförbund.
Finlands Fackförbunds Centralorganisation FFC erbjuder gratis anställningsrådgivning.
Du kan få rådgivning även om du inte är medlem i ett fackförbund.
Juristerna svarar på dina frågor på finska och engelska.
Rådgivning ges både per telefon och via e-post:
Tfn 0800 414 004, tis. och ons. kl. 9–11 och 12–15
Du kan även ringa arbetarskyddsmyndigheternas riksomfattande rådgivningstelefon:
Tfn 0295 016 620
Mån.–fre. kl. 9–15
linkkiArbetarskyddsförvaltning:
Kontaktuppgifter till arbetarskyddsmyndigheternafinska _ svenska _ engelska
Min anställning upphör inom kort.
Hur påverkar det mitt uppehållstillstånd?
Detta beror på vilket slags uppehållstillstånd du har.
Om ditt uppehållstillstånd är kopplat till endast en arbetsgivare, ska du ansöka om ett nytt uppehållstillstånd för arbetstagare.
För att kunna ansöka om ett nytt uppehållstillstånd för arbetstagare måste du ha ett nytt jobb.
Du kan även ansöka om uppehållstillstånd på någon annan grund.
Läs mer om grunderna för uppehållstillstånd i InfoFinlands avsnitt Icke EU-medborgare.
Om din anställning upphör innan ditt uppehållstillstånd går ut, ska du meddela detta skriftligt till Migrationsverket.
Också din arbetsgivare kan göra anmälan.
Om ditt uppehållstillstånd är beviljat för en viss bransch, kan du byta jobb inom samma bransch.
Information om uppehållstillstånd för arbetstagare och företagare hittar du på sidorna Arbeta i Finland och Till Finland som företagare.
Läs mer om att söka jobb i Finland på sidan Var hittar jag jobb?
Mer information om att söka arbetslöshetsersättning hittar du på sidan Arbetslöshetsförsäkring.
Information om uppehållstillståndfinska _ svenska _ engelska
Jag har fått för lite lön utbetalad.
Vad ska jag göra?
Kontrollera alltid i lönespecifikationen att du har fått rätt belopp.
Om du har fått för lite lön, ska du be din arbetsgivare att rätta till löneutbetalningen.
Om arbetsgivaren inte betalar ut rätt lön, ska du fråga om råd hos regionförvaltningsverkets arbetarskydd eller ditt fackförbund.
Om du inte kan komma överens om löneutbetalningen med din arbetsgivare måste ärendet avgöras i domstol.
Detta är dock det sista alternativet.
linkkiArbetarskyddsförvaltning:
Information om löneutbetalningfinska _ svenska _ engelska
Min arbetsgivare vill endast betala ut lönen i kontanter.
Får man göra så?
Din arbetsgivare borde betala ut lönen till ditt bankkonto.
Lönen får endast betalas ut i kontanter om inga andra alternativ finns.
Så gör man till exempel om du inte har ett bankkonto.
Om du får lönen utbetalad i kontanter, ska du ge din arbetsgivare ett skriftligt intyg om löneutbetalningen.
På så sätt kan man bevisa att lönen verkligen har betalats till dig.
Min tillsvidareanställning upphörde, men min sista lön betalades inte ut.
Vad bör jag göra?
Fråga arbetsgivaren varför lönen blivit försenad.
Kräv att arbetsgivaren betalar ut lönen.
Framför kravet skriftligt.
Om du är medlem i ett fackförbund kan du be förbundet om hjälp.
Om du inte är medlem i ett fackförbund, kontakta till exempel arbetarskyddsmyndigheterna.
Jag avslutade mitt jobb hos min förra arbetsgivare, men jag har inte fått ett arbetsintyg.
Hur får jag arbetsintyget?
Arbetsgivare behöver inte ge dig ett arbetsintyg på eget bevåg.
Om du vill ha ett arbetsintyg ska du be om det.
Intyget ska lämnas till dig så snart som möjligt.
Om du har bett om ett arbetsintyg men inte fått det, ska du kontakta arbetarskyddsmyndigheterna.
Läs mer på InfoFinlands sida Arbetsintyg.
Jag upplever att jag blir osakligt bemött på min arbetsplats.
Vad kan jag göra?
Alla arbetstagare ska behandlas jämlikt och lika.
Enligt lag får ingen diskrimineras till exempel av följande orsaker:
anställningsform
ålder
kön
etnisk bakgrund
hälsotillstånd
religion
sexuell läggning.
Läs mer på InfoFinlands sida Diskriminering och rasism.
Förutom diskriminering kan det även förekomma andra typer av osakligt bemötande på arbetsplatser, till exempel mobbning eller sexuella trakasserier.
Om hen inte kan hjälpa dig, ska du kontakta arbetsplatsens arbetarskyddsfullmäktige eller förtroendeman.
Om ärendet inte kan lösas på arbetsplatsen, kontakta arbetarskyddsmyndigheterna eller ditt fackförbund.
Om din chef behandlar dig osakligt, anmäl detta till arbetarskyddsmyndigheterna.
Du kan göra anmälan med ditt eget namn eller anonymt.
Jag tvingas att utföra ett jobb utan att få betalt.
Min arbetsgivare hotar mig dessutom med våld.
Var kan jag få hjälp?
Du har rätt till hjälp och skydd.
Enligt lagen i Finland måste arbetstagarna behandlas väl och de ska betalas lön.
Människohandel är ett brott i Finland.
Läs mer på InfoFinlands sida Människohandel och tvångsarbete.
Du hittar information om arbetstagarens rättigheter och skyldigheter i Finland på InfoFinlands sida Arbetstagarens rättigheter och skyldigheter.
Hjälp till offer för människohandelfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska _ polska _ rumänska _ bulgariska
I skattedeklarationen finns uppgifter om inkomster, skatter och avdrag från föregående år.
Kontrollera uppgifterna i skattedeklarationen.
Den slutliga beskattningen fastställs utgående från uppgifterna i skattedeklarationen.
Om alla uppgifter är korrekta, och det inte saknas några uppgifter, behöver du inte göra någonting.
Om uppgifterna inte är korrekta, eller om det saknas något, komplettera och korrigera skattedeklarationen i webbtjänsten MinSkatt.
Du kan använda webbtjänsten, om du har finländska nätbankskoder eller ett mobilcertifikat.
Om du inte gör rättelserna i webbtjänsten MinSkatt, hämta pappersblanketter för rättelserna på Skatteförvaltningens webbplats eller i skattebyrån.
Skicka blanketterna per post.
Kom ihåg att kontrollera skattedeklarationen och göra de ändringar som behövs före utgången av den sista returdagen.
Beskattningsbeslut
Beskattningsbeslutet (Verotuspäätös) är en beräkning av det slutliga skattebeloppet.
På din lön eller annan inkomst har det innehållits skatt utgående från skattekortet.
Det här kallas för förskottsinnehållning (ennakonpidätys).
Förskottsinnehållningens storlek baserar sig på en uppskattning av dina inkomster.
Skattebeloppet justeras i efterskott utgående från hur stora dina inkomster och avdrag verkligen har varit.
Tillsammans med den på förhand ifyllda skattedeklarationen får du ett beskattningsbeslut.
Om du inte korrigerar skattedeklarationen, förblir det här beskattningsbeslutet i kraft.
Om du korrigerar skattedeklarationen, får du ett nytt beskattningsbeslut senare.
Kom ihåg att kontrollera också det nya beskattningsbeslutet.
Spara beskattningsbeslutet och den specifikationsdel som du fick på våren tillsammans med skattedeklarationen.
Om du beställer en ny specifikationsdel, tas det ut en avgift för den.
linkkiSkatteförvaltningen:
Skattedeklaration och beskattningsbeslutfinska _ svenska _ engelska
Avdrag
I beskattningen kan du göra avdrag (vähennykset), som minskar beskattningen.
Skatteförvaltningen gör en del avdrag automatiskt, men vissa avdrag måste du själv ansöka om.
Avdrag är till exempel:
hushållsavdrag
avdrag för resekostnader mellan bostaden och arbetsplatsen
ränteavdrag på bostadslån
Du kan avdra räntorna för bostadslånet i beskattningen då du har tagit ett lån för din stadigvarande bostad.
Du kan dra av räntorna på bostadslånet i beskattningen också då din stadigvarande bostad finns utomlands.
Om du har tagit ett lån hos en finländsk bank, får skattemyndigheten uppgifterna om lånet direkt från banken.
Om du har ett bostadslån i en utländsk bank, ska du själv ge uppgifterna om lånet till skattemyndigheten.
Du kan meddela om avdrag, när du beställer ett nytt skattekort.
Avdragen beaktas då i din skatteprocent.
Du kan också ansöka om avdrag i efterskott med skattedeklarationen.
Du får då avdragen i efterskott som en skatteåterbäring.
linkkiSkatteförvaltningen:
Avdrag vid beskattningenfinska _ svenska _ engelska
Skatteåterbäring och kvarskatt
Du ser i beskattningsbeslutet om du har betalat rätt mängd skatt.
Om du har betalat för mycket i skatt, får du skatteåterbäring (veronpalautus).
Om du har betalat för lite i skatt, blir du tvungen att betala kvarskatt (jäännösvero).
Skatteåterbäringen betalas antingen direkt på ditt bankkonto.
Meddela numret på ditt bankkonto via Skatteförvaltningens webbtjänst eller på en separat pappersblankett.
Du kan få skatteåterbäringen antingen till ett finländskt eller till ett utländsk bankkonto.
Om du blir tvungen att betala kvarskatt, får du tillsammans med beskattningsbeslutet en bankgiroblankett.
På bankgiroblanketten ser du kvarskattebeloppet, bankkontonumret, förfallodagen och referensnumret.
Du blir också tvungen att betala ränta på kvarskatten efter en viss tid.
linkkiSkatteåterbäringar:
Skatteåterbäringarfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Ange kontonummerfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Kvarskattfinska _ svenska _ engelska
Tillstånd eller anmälan
Etableringsanmälan
Försäkringar
Bokföring
Beskattning
Inkomstregistret
Arbetstagarnas inskolning och säkerhet
När du inleder företagsverksamheten har du många skyldigheter.
Du ska bland annat registrera företaget, betala skatt och ordna bokföringen.
Tillstånd eller anmälan
I Finland får man driva en laglig näring som följer god sed utan ett tillstånd som beviljas av myndigheter.
I vissa fall behövs det dock ett tillstånd från myndigheter för att starta företagsverksamhet, eller också måste man anmäla verksamheten till myndigheter.
Om du till exempel har ett företag som idkar skönhetsvård eller säljer livsmedel ska företagets lokaler kontrolleras.
Ansök om tillstånd hos kommunens hälsomyndighet innan lokalerna tas i bruk.
Innan du startar företagsverksamheten, kontrollera om du behöver tillstånd för verksamheten eller om du måste anmäla verksamheten till en myndighet.
Du kan kontrollera hos regionförvaltningsverken eller på Företagsfinlands webbplats om du behöver ett tillstånd för ditt företag.
linkkiFöretagsfinland:
Tillstånd och anmälan som är anknutna till idkandet av en näringfinska _ svenska _ engelska
linkkiFinlands Näringsliv:
Företagslagstiftningfinska
Etableringsanmälan
Ny företagsverksamhet ska anmälas till handelsregistret som upprätthålls av Patent- och registerstyrelsen (Patentti- ja rekisterihallitus).
Du kan använda samma blankett när du gör etableringsanmälan för ditt företag till Patent- och registerstyrelsen och till Skatteförvaltningen.
linkkiPatent- och registerstyrelsen:
Anmälan om grundande av ett företagfinska _ svenska _ engelska
Försäkringar
Företagarpensionsförsäkringen (FöPL) (YEL-vakuutus) är obligatorisk för företagare i åldern 18–68 år, vars företagsverksamhet inbringar minst 7 799,37 euro om året som arbetsinkomst (år 2019).
Pensionsförsäkringen tryggar företagarens utkomst då företagsverksamheten upphör på grund av invaliditet eller ålder och den ger företagarens anhöriga ett familjepensionsskydd efter att företagaren har dött.
Pensionsförsäkringar fås antingen genom försäkringsbolag eller pensionskassor (eläkekassa).
Teckna en pensionsförsäkring senast när det har gått sex månader sedan du startade företagsverksamheten.
En ny företagare får en rabatt på 22 procent på pensionspremierna under de fyra första åren.
Storleken av försäkringspremierna och pensionen beror på hur stor förvärvsinkomst (työtulo) förtagaren har.
Förvärvsinkomstens storlek inverkar också på storleken av olika inkomstrelaterade förmåner (ansiosidonnanen etuus), såsom sjukdagpenningen.
linkkiPensionsskyddscentralen:
Information om företagarpensionsförsäkringenfinska _ svenska _ engelska
Du ska teckna en pensionsförsäkring (ArPL-försäkring) (eläkevakuutus (TyEL-vakuutus)) och en olycksfallsförsäkring som omfattar en grupplivförsäkring och en arbetslöshetsförsäkring för de anställda.
Arbetsgivaren betalar arbetstagarens socialskyddsavgifter till skattemyndigheten i anslutning till skatteinnehållningen.
I vissa branscher finns också andra obligatoriska försäkringar.
Du bör också överväga andra frivilliga försäkringar som till exempel företagarens olycksfallsförsäkring.
linkkiPensionsskyddscentralen:
Information om att teckna försäkringar för anställdafinska _ svenska _ engelska
linkkiFöretagsFinland:
Information om att teckna försäkringar för anställdafinska _ svenska _ engelska
Bokföring
I Finland har alla företagare bokföringsskyldighet.
Om du inte vill sköta bokföringen själv, kan du anlita en revisionsbyrå som sköter företagets bokföring åt dig.
I Finland anlitar många företag revisionsbyråer.
Beskattning
Företagsformen påverkar företagets beskattning.
Detta är det bra att beakta när du väljer företagsform.
En ny företagare kan anmäla sig till Skatteförvaltningens förskottsuppbördsregister.
Anmälan till förskottsuppbördsregistret görs med samma anmälan som görs för grundande av företaget, d.v.s. etableringsanmälan (yrityksen perustamisilmoitus).
Om ditt företag är i förskottsuppbördsregistret kan du fakturera kunder utan förskottsinnehållning.
Skatter betalas på de inkomster som företagaren eller företaget har kvar när alla kostnader för företagsverksamheten har dragits av försäljningen.
Företagets skatter betalas på basis av de beskattningsbara inkomsterna, vars belopp man uppskattar på förhand.
Uppskattningen baseras på beloppet av de beskattningsbara inkomsterna året innan.
I ett nytt företag uppskattar företagaren själv storleken av den beskattningsbara inkomsten och meddelar denna till skattmyndigheten.
linkkiSkatteförvaltningen:
Information om beskattningen av företag och företagarefinska _ svenska _ engelska
linkkiFöretagsFinland:
Information om beskattningen av företag och företagarefinska _ svenska _ engelska
Mervärdesskatt
Mervärdesskatten (arvonlisävero) är en konsumtionsskatt som i Finland betalas för nästan alla varor och tjänster.
Företagare som säljer varor och tjänster i Finland är skyldiga att betala mervärdesskatt.
Om inkomsten som man får för försäljningen av varor och tjänster är mindre än 10 000 euro per år, behöver ingen mervärdesskatt betalas på den.
Företagsformen påverkar inte mervärdesskattens belopp.
Mervärdesskattebeloppet varierar emellertid för olika produkter.
Inkomstregistret
Inkomstregistret är en databas dit arbetsgivarna anmäler lönerna som de utbetalat till sina anställda.
Anmälan ska göras senast fem dagar efter löneutbetalningen.
Uppgifterna ska skickas till inkomstregistret elektroniskt:
direkt via lönesystemet om det har en inbyggd teknisk förbindelse till Inkomstregistret eller
via Inkomstregistrets ärendehantering, till vilken man får tillträde med webbankkoder eller andra medel för elektronisk identifiering.
Löneuppgifterna kan endast i undantagsfall anmälas med ett pappersformulär.
Läs mer om Inkomstregistret och om att anmäla löner på Inkomstregistrets webbplats.
linkkiSkatteförvaltningen:
Inkomstregistretfinska _ svenska _ engelska _ ryska _ estniska _ kinesiska
Arbetstagarnas inskolning och säkerhet
Som företagare har du ansvaret för att ge arbetstagarna inskolning i arbetsuppgifterna.
Arbetsgivaren ska introducera förhållandena på arbetsplatsen och de rätta arbetsmetoderna för arbetstagaren.
Arbetsgivaren är också skyldig att sörja för arbetstagarnas säkerhet och hälsa i arbetet.
Arbetsgivaren ska utarbeta ett verksamhetsprogram för arbetarskyddet (työsuojelun toimintaohjelma) som tar upp de säkerhets- och hälsorelaterade riskerna på arbetsplatsen och hur man undgår dem.
Läs mer om att vara arbetsgivare på InfoFinlands sida Arbetsgivarens rättigheter och skyldigheter.
linkkiArbetarskyddscentralen:
Information om arbetarskyddfinska _ svenska _ engelska
Arbetstagaren har rätt att på begäran få ett arbetsintyg av arbetsgivaren när anställningen upphör.
Arbetsintyget är ett viktigt dokument där anställningens längd och arbetsuppgifterna nämns.
Arbetstagaren kan också be att orsaken till att anställningen upphört och en bedömning av arbetstagarens färdigheter och uppförande antecknas i intyget.
Arbetsgivaren är skyldig att utfärda ett arbetsintyg ännu tio år efter att anställningen har upphört och efter detta endast om detta inte medför en orimlig olägenhet för arbetsgivaren.
Om arbetstagaren vill att en bedömning av färdigheterna och uppförandet antecknas i arbetsintyget måste arbetsgivaren utfärda ett sådant intyg ännu fem år efter att anställningen har upphört till arbetstagaren på hans eller hennes begäran.
Arbetsgivare måste också ge arbetstagaren ett nytt arbetsintyg om arbetstagarens arbetsintyg kommer bort eller förstörs.
En arbetsgivare som avsiktligt eller av vårdslöshet inte utfärdar ett arbetsintyg bryter mot arbetsavtalslagen.
Arbetsavtalslagenfinska _ svenska _ engelska
linkkiArbetarskyddsförvaltningen:
Information om rätten till arbetsintygfinska _ svenska _ engelska
Du behöver ett skattekort (verokortti), om du får lön eller har andra inkomster i Finland.
På skattekortet finns en anteckning om skatteprocenten (veroprosentti).
Av det ser arbetsgivaren, hur mycket skatt som ska betalas på lönen.
Skatteprocenten beror på hur hög din inkomst är.
Om du håller på att flytta till Finland, får du skattekortet från skattebyrån (verotoimisto).
Uppskatta för skattekortet, hur stora dina inkomster kommer att bli för hela skatteåret.
Du behöver också en finländsk personbeteckning.
Du får personbeteckningen, när du registrerar dig som invånare hos magistraten.
Du kan få en personbeteckning också från skattebyrån.
Läs mer på sidan Registrering som invånare.
När du bor i Finland stadigvarande, skickar Skatteförvaltningen ett nytt skattekort till dig varje år i januari.
Skatteförvaltningen räknar ut en lämplig skatteprocent åt dig utgående från hur mycket du förtjänade året innan.
Förete skattekortet till din arbetsgivare.
Om du inte företer skattekortet till din arbetsgivare, innehåller arbetsgivaren en skatt på 60 % på din lön.
Om dina inkomster blir mindre eller större under året, ska du beställa ett nytt skattekort.
Du får ett nytt skattekort:
från Skatteförvaltningens webbtjänst MinSkatt
när du ringer numret 029 497 000 (betjäningsspråk: finska, svenska, engelska)
på skattebyrån
När du söker ett nytt skattekort, behöver du följande uppgifter:
en uppskattning av dina inkomster för hela året
de inkomster som du har haft från början av året
de skatter som har betalats på dina inkomster från början av året
uppgift om de avdrag som du söker i beskattningen för innevarande år
Om du betalar för mycket skatt, får du skatteåterbäring.
Om du betalar för litet i skatt, blir du tvungen att betala kvarskatt.
linkkiSkatteförvaltningen:
Nytt skattekortfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Hur beräknas skatteprocenten?finska _ svenska
Om du har flera arbetsgivare
Om du har flera arbetsgivare ska du förete ditt skattekort till dem alla.
Du kan använda samma skattekort hos alla arbetsgivarna.
Du betalar samma skatt hos alla dina arbetsgivare.
På skattekortet anges en inkomstgräns och din skatteprocent beräknas utifrån den.
Kom ihåg att hålla ett öga på dina inkomster.
Om du får mer lön än vad du uppgett, överskrids din inkomstgräns.
Om inkomstgränsen överskrids ska du beställa ett nytt skattekort.
Skattenummer
Du behöver en skattenummer (veronumero), om du arbetar på en bygg- eller monteringsarbetsplats i Finland.
Med hjälp av skattenumret kontrolleras, att alla arbetstagare finns i Skatteförvaltningens register.
Skattenumret ska framgå av den fotoförsedda namnskylt som du får av din arbetsgivare.
Du får inte arbeta på en byggplats utan namnskylt.
Du får skattenumret från skattebyrån samtidigt som du går efter skattekortet.
Om du redan har finländsk personbeteckning och ett skattekort, hittar du skattenumret på ditt skattekort.
linkkiSkatteförvaltningen:
Skattenummerfinska _ svenska _ engelska
När du grundar ett företag måste du välja företagsform och ett namn för företaget samt definiera branschen.
På valet av företagsform inverkar bland annat antalet grundare, behovet av kapital, fördelningen av ansvar och bestämmanderätt, finansieringen och beskattningen.
Olika företagsformer i Finland är enskild näringsidkare (toiminimi); öppet bolag (avoin yhtiö); kommanditbolag (kommandiittiyhtiö); aktiebolag (osakeyhtiö) och andelslag (osuuskunta).
När du funderar på vilken företagsform du ska välja, är det absolut tillrådligt att du kontaktar företagsrådgivningen.
linkkiNyföretagarcentralerna i Finland:
Företagsrådgivningfinska _ svenska _ engelska
Enskild näringsidkare (toiminimi)
Det enklaste och vanligaste sättet att starta företagsverksamhet är att som enskild näringsidkare driva en firma.
Du har bestämmanderätt över och ansvar för firmans ärenden och företaget kan anställa medarbetare precis som andra företag.
Företagsverksamhet som bisyssla lönar det sig ofta att starta som enskild näringsidkare.
Det är snabbt och enkelt att starta företagsverksamhet som enskild näringsidkare.
Aktiebolaget är den vanligaste företagsformen i Finland.
Ett aktiebolag passar för all slags affärsverksamhet.
Du kan grunda ett aktiebolag antingen själv eller tillsammans med andra delägare.
Delägarens rösträtt, avkastning och ansvar i bolaget beror på hur många aktier i bolaget hen äger.
Ett öppet bolag bildas då två eller fler personer kommer överens om att grunda ett bolag genom att teckna ett bolagsavtal.
Bolagsmännen, d.v.s. personerna som tillsammans äger bolaget, är jämställda i all verksamhet som bolaget driver och de ansvarar tillsammans och personligen för bolagets beslut, förbindelser och skulder.
Ett kommanditbolag är ett personbolag som skiljer sig från ett öppet bolag på så sätt att det i kommanditbolaget finns utöver en eller flera ansvariga bolagsmän åtminstone en tyst bolagsman, d.v.s. en person som är delägare i företaget. Vanligen är den tysta bolagsmannen en investerare.
Det behövs minst tre personer för att grunda ett andelslag.
Ett andelslag är ett företag som ägs av medlemmarna.
På andelslagets stämma har varje medlem en röst.
Medlemmarna ansvarar för andelslagets förpliktelser (till exempel skulder) endast med det belopp som de investerat i andelslaget.
linkkiFöretagsFinland:
Information om företagsformerfinska _ svenska _ engelska
När ett barn föds till familjen har föräldrarna rätt att ta familjeledighet, det vill säga stanna hemma för att ta hand om barnet.
Med familjeledighet avses
moderskapsledighet
faderskapsledighet
föräldraledighet
vårdledighet
Meddela din arbetsgivare om familjeledigheten senast två månader innan den börjar.
Familjeledigheterna är vanligen oavlönad ledighet.
Huruvida du får lön under familjeledigheten beror på ditt kollektivavtal.
Kontrollera detta med din arbetsgivare.
FPA betalar ut familjeförmåner för familjeledigheten: föräldrapenning och stöd för hemvård av barn.
Läs om villkoren för familjeförmånerna på InfoFinlands sida Stöd efter barnets födelse och Stöd för vård av barn i hemmet.
När familjeledigheterna upphör har arbetstagaren rätt att återvända till sitt eget arbete eller motsvarande arbete på den gamla arbetsplatsen.
Arbetsavtalet för en gravid kvinna får inte hävas och hon får inte diskrimineras på grund av sin graviditet.
I Finland känner arbetsgivarna och arbetstagarna till familjeledigheterna och de används allmänt.
linkkiArbets- och näringsministeriet:
Familjeledigheterfinska _ svenska _ engelska
Information om stöd till barnfamiljerfinska _ svenska _ engelska
Moderskapsledighet
Moderskapsledigheten är 105 vardagar.
Arbete under moderskapsledigheten är tillåtet om det kan utföras utan att moderns, fostrets eller barnets säkerhet äventyras.
Under moderskapsledigheten får man dock inte arbeta under de två veckor som föregår det beräknade födelsedatumet och under två veckor efter förlossningen.
Faderskapsledighet
Faderskapsledigheten är den del av föräldraledigheten som är avsedd att tas ut av fadern.
Faderskapsledigheten är allt som allt 54 vardagar.
Dessa dagar kan inte överföras till modern.
Du kan ta ut högst 18 dagar av din faderskapsledighet samtidigt som barnets mor är moderskaps- eller föräldraledig.
Dessa dagar kan du dela upp på högst fyra perioder.
De återstående 36 dagarna kan du dela upp på högst två perioder.
Under dessa dagar kan modern inte vara moderskapsledig samtidigt.
Avsikten är att fadern tar hand om barnet.
Du kan också ta ut alla 54 dagar av din faderskapsledighet vid olika tider med modern.
Du kan själv bestämma om du tar ut hela faderskapsledigheten eller bara en del av dagarna.
Faderskapsledigheten får endast tas ut före barnet har fyllt två år.
När barnet fyller två år kan du inte längre ta ut faderskapsledighet trots att du har dagar kvar.
Föräldraledighet
Efter moderskapsledigheten kan antingen modern eller fadern stanna hemma för att ta hand om barnet. Föräldraledigheten varar 158 vardagar.
Båda föräldrarna kan inte vara föräldralediga samtidigt.
Däremot kan man dela upp föräldraledigheten så att modern eller fadern stannar hemma växelvis för att ta hand om barnet.
Vårdledighet
Efter föräldraledigheten kan antingen modern eller fadern ta ut en oavlönad vårdledighet för att ta hand om barnet tills barnet fyller tre år.
Det förutsätter att modern eller fadern varit anställd hos samma arbetsgivare minst sex månader under det senaste året.
Under vårdledigheten betalar FPA stöd för hemvård av barn.
Se villkoren för stödet för hemvård av barn på InfoFinlands sida Stöd för vård av barn i hemmet.
Partiell vårdledighet
Du kan också vara vårdledig på deltid.
Då arbetar du kortare dagar och får på motsvarande sätt mindre lön.
Makarna kan vara partiellt vårdlediga samtidigt så att den ena förkortar sin arbetstid från morgonen och den andra från eftermiddagen.
Du kan vara partiellt vårdledig tills barnet har gått ut årskurs två.
Om du har hemkommun i Finland kan du ansöka om partiell vårdpenning hos FPA för hemvård av barn under tre år eller skolbarn i årskurserna 1 eller 2.
Partiell vårdpenning betalas inte för vård av ett barn som fyllt tre men ännu inte går i skolan.
Läs mer om partiell vårdpenning på InfoFinlands sida Stöd för vård av barn i hemmet.
I Finland betalar du inkomstskatt (tulovero) på lön.
Du betalar också skatt på till exempel följande inkomster:
arbetslöshetsdagpenning
föräldradagpenning
pensioner
studiestöd
För skattepengarna betalar staten och kommunerna till exempel:
hälsovård
utbildning
dagvård
försvar
I Finland är beskattningen progressiv.
Det innebär att man på en stor lön betalar en större andel skatt än på en mindre lön.
Skatteprocenten (Veroprosentti) beräknas i Finland för var och en separat.
Din makes/makas inkomster inverkar inte på din skatteprocent.
Du kan uppskatta din skatteprocent med Skatteförvaltningens skatteräknare.
Arbetsgivaren betalar skatterna direkt från din lön.
För att kunna göra det behöver arbetsgivaren ett skattekort av dig.
Skatt som betalas direkt från lönen, är förskottsskatt (ennakonpidätys).
Skatteförvaltningen räknar efter varje år om du har betalat tillräckligt med skatt på dina inkomster.
Om du har betalat för mycket i skatt, får du skatteåterbäring (veronpalautus).
Om du har betalat för lite i skatt, blir du tvungen att betala kvarskatt (jäännösvero).
Läs mer på sidan: Skattedeklaration och beskattningsbeslut.
Kontrollera i lönespecifikationen och skattedeklarationen (veroilmoitus), att arbetsgivaren har betalat skatt på din lön.
Spara lönekvittona.
Om skatten inte har betalats, blir du tvungen att betala den i efterskott.
Utöver skatt betalar arbetsgivaren försäkringspremier på din lön i händelse av arbetslöshet eller sjukdom.
linkkiSkatteförvaltningen:
Information om beskattningenfinska _ svenska _ engelska
linkkiSkattemyndigheten:
Skattekortfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Skatteprocenträknarefinska _ svenska _ engelska
Beskattningen när du börjar arbeta i Finland
Om du kommer till Finland för att arbeta, beror din beskattning på hur länge du vistas i Finland.
På beskattningen inverkar också huruvida din arbetsgivare är ett finländskt eller ett utländskt företag.
Om du vistas i Finland i mer än sex månader, ska du i allmänhet betala skatt på din lön till Finland.
Du ska i allmänhet också betala de obligatoriska försäkringspremierna till Finland.
Du behöver en finländsk personbeteckning och ett finländskt skattekort.
Skatteprocenten räknas på inkomsterna för hela året.
Du får skatteavdrag på samma grunder som andra som bor i Finland stadigvarande.
Om du vistas i Finland i högst sex månader och din arbetsgivare är ett utländskt företag, behöver du i allmänhet inte betala skatt till Finland.
Om din arbetsgivare är finländare eller om din utländska arbetsgivare har en arbetsplats i Finland, betalar du skatt i Finland.
Du kan söka progressiv beskattning, om du bor i ett land som hör till Europeiska ekonomiska samarbetsområdet eller i en stat, med vilken Finland har ett skatteavtal.
I annat fall betalar du en källskatt (lähdevero) på 35 % på lönen och du behöver ett källskattekort.
Källskattekort måste du ansöka med en pappersblankett.
För progressiv beskattning behöver du ett skattekort för begränsat skattskyldiga (rajoitetusti verovelvollisen verokortti).
Du får ett sådant på skattebyrån.
Du kan söka progressiv beskattning också i efterskott.
Du blir också tvungen att betala försäkringspremier, om du inte är försäkrad i det land där du bor stadigvarande.
Om du redan är försäkrad i ett annat land, behöver du ett intyg A1/E101 över försäkringen.
När du flyttar bort från Finland, kom ihåg att göra en flyttningsanmälan till magistraten.
Du får då din skattedeklaration till rätt adress.
När du håller på att flytta till Finland, får du ytterligare information i avsnittet Flytta till Finland.
linkkiSkatteförvaltningen:
Arbeta i Finlandfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Ansökan om progressiv inkomstbeskattningfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Utländsk hyrd arbetskraft och beskattningen i Finlandfinska _ svenska _ engelska
Flyttanmälanfinska _ svenska _ engelska
Uppehållstillstånd eller registrering av uppehållsrätt?
Kom på en affärsidé
Gör en affärsverksamhetsplan
Fråga om råd på företagsrådgivningen
Ordna finansiering
Välj företagsform
Du kan grunda ett företag i Finland oavsett ditt medborgarskap.
Det viktiga är att du har uppehållsrätt i Finland, de yrkeskunskaper som krävs och tillräckliga kunskaper i finska.
Uppehållstillstånd eller registrering av uppehållsrätt?
Om du är medborgare i ett nordiskt land och flyttar till Finland ska du registrera dig vid magistraten.
Du behöver inget uppehållstillstånd i Finland.
Läs mer på InfoFinlands sida Nordisk medborgare.
Om du är medborgare i något EU-land, Liechtenstein eller Schweiz och flyttar till Finland permanent, ska du registrera dig vid Migrationsverket och magistraten.
Läs mer på InfoFinlands sida EU-medborgare.
Om du är medborgare i något land som inte tillhör EU och flyttar till Finland som företagare, behöver du antingen ett uppehållstillstånd för företagare, ett uppehållstillstånd för arbetstagare eller ett uppehållstillstånd för uppstartsföretagare.
Läs mer på InfoFinlands sida Till Finland som företagare.
Som företagare till Finland:
Vilka tillstånd behöver du?(pdf, 384 kt)finska _ engelska
Tillstånd och anmälningar för utländska företagarefinska _ svenska _ engelska
Kom på en affärsidé
Processen för att grunda ett företag är likadant som för finska medborgare.
När du vill grunda ett företag ska du noga fundera på om du har en bra affärsidé.
Fundera också på om du har tillräckliga yrkeskunskaper och erfarenhet.
Det är viktigt att du känner väl till din bransch och de lagar som styr företagande.
Det är också viktigt att känna till sina kunder och försäljningsmetoder.
Kom ihåg att företagande även medför risker.
Tillräcklig finansiering och noggrann planering är nödvändiga.
linkkiFöretagsfinland:
Att grunda ett företagfinska _ svenska _ engelska
Gör en affärsverksamhetsplan
I affärsverksamhetsplanen funderar du på styrkorna och svagheterna i ditt kunnande och egenskaperna hos den produkt, vara eller tjänst som du erbjuder.
Fundera på vilka som är dina kunder och vilka önskemål de har.
Fundera också på vilka som är dina konkurrenter och hurdana produkter och verksamhetssätt de har.
Den viktigaste delen i affärsverksamhetsplanen är verksamhetsplanen för ditt eget företag.
Fundera noga hur företaget drivs och var och hurdana lokaler företaget har.
Fundera på vilka produktionsmedel eller vilken arbetskraft du behöver.
Vilka reklammedel ska du använda för att främja försäljningen?
Ta också reda på om försäkringar täcker de risker som förknippas med verksamheten.
Fundera också på hur du ordnar bokföringen och planerar ekonomin.
Hur avser du följa upp hur dina planer förverkligas?
Anteckna allt detta i din affärsverksamhetsplan.
Hjälp med att upprätta en affärsverksamhetsplan
Du får närmare anvisningar om hur du upprättar en affärsverksamhetsplan vid företagsrådgivningscentra.
På deras webbplatser kan du även ladda ned företagarguider åtminstone på finska och engelska.
Där får du även en mall för affärsverksamhetsplanen och andra dokumentmallar.
Guide om att grunda ett företagfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ turkiska _ kinesiska _ arabiska
Fråga om råd på företagsrådgivningen
I Finland har alla möjlighet att få kostnadsfri företagsrådgivning.
Rådgivning erbjuds vid till exempel:
Nyföretagarcentraler
Närings-, trafik- och miljöcentralerna (NTM-centralerna)
Arbets- och näringsbyråer (TE-byråer)
FöretagsFinland (via webbplatsen och per telefon)
När du får en bra affärsidé, kontakta närmaste företagsservicecenter.
Där hjälper experterna dig att utveckla affärsidén, göra en marknadsundersökning, beräkna lönsamheten och kartlägga finansieringen.
Du får även stöd när du funderar på om du ska starta ett företag.
Företagsrådgivning fås på finska och svenska och åtminstone i de större städerna även på engelska.
Ibland kan det finnas möjlighet att få rådgivning även på något annat språk.
linkkiFöretagsFinland:
Företagsrådgivningfinska _ svenska _ engelska
Företagarkurser
Olika instanser ordnar företagarkurser och informationsmöten som är mycket nyttiga för dig som ska grunda ett företag.
På kurserna behandlas till exempel upprättande av affärsverksamhetsplan, start av företagsverksamheten, bokföring, företagsbeskattning, juridiska frågor, marknadsföring, försäljning och kundtjänst.
Ordna finansiering
Planera företagets finansiering noga innan du grundar företaget.
Det är viktigt att du har tillräckligt stort kapital i början.
En del av företagets finansiering kan bestå av en gåva eller ett lån.
När du ansöker om finansiering måste du ha en ordentlig affärsverksamhetsplan färdig.
Lån
Banker och Finnvera beviljar lån till företagare som startar ett företag.
Finnvera är ett finansieringsbolag som ägs av finska staten.
Det ger lån till nya företag och redan aktiva företag.
Om ditt företag har förutsättningarna för en lönsam verksamhet men du inte har tillräckligt mycket pengar eller säkerheter för att få ett banklån, ska du fråga om du kan få ett lån eller borgen hos Finnvera.
linkkiFöretagsFinland:
Finansiering för ett företagfinska _ svenska _ engelska
linkkiFinnvera:
Finansiering för ett företagfinska _ svenska _ engelska
Startpenning
När du blir företagare, kan du få startpenning för att trygga försörjningen när företagsverksamheten precis har börjat.
Du ansöker om startpenning vid den arbets- och näringsbyrå där du är kund.
Du kan få startpenning för högst tolv månader.
När du ansöker om startpenning utreder arbets- och näringsbyrån om företagande är ett lämpligt alternativ för dig.
Du kan få startpenning om
du är arbetslös arbetssökande
du inte är arbetslös, men går från till exempel lönearbete, studier eller hemmaarbete till företagare
du har företagande som bisyssla och utvidgar företagsverksamheten till din huvudsyssla.
Förutsättningar för att få startpenning är till exempel:
företagande som huvudsyssla
tillräckliga kunskaper, färdigheter och resurser för den företagsverksamhet som du planerar
arbets- och näringsbyrån uppskattar att företagsverksamheten kan vara lönsam
du behöver startpenningen för din försörjning
Företagsverksamheten startas först när stödet har beviljats.
Om du avser ansöka om startpenning ska du kontakta arbets- och näringsbyrån i ett så tidigt skede som möjligt.
Det finns även andra stödformer för nya företagare.
FöretagsFinland ger dig information om olika finansieringsalternativ.
linkkiArbets- och näringsministeriet:
Information om startpengenfinska _ svenska _ engelska
Välj företagsform
När du ska grunda ett företag, måste du välja företagsform och ett namn för företaget samt ange bransch.
När du väljer företagsformen ska du beakta bland annat antalet grundare, behovet av kapital, fördelningen av ansvar och beslutsmakt samt finansiering och beskattning.
Olika företagsformer i Finland är firma, öppet bolag, kommanditbolag, aktiebolag och andelslag.
När du funderar på vilken företagsform du ska välja, är det absolut tillrådligt att du kontaktar företagsrådgivningen.
Läs mer på InfoFinlands sida Företagsformer.
Om du blir sjuk eller råkar ut för en olycka har du rätt att stanna hemma från arbetet.
Arbetsgivaren är skyldig att betala lön för sjukledigheten.
Om din anställning varat över en månad före insjuknandet får du lönen till fullt belopp för minst den dag då du insjuknade och nio därefter följande dagar.
Om du fortfarande inte kan återvända till arbetet kan du söka sjukdagpenning (sairauspäiväraha) hos FPA om du omfattas av den finländska sjukförsäkringen.
Läs mer på InfoFinlands sida Den sociala tryggheten i Finland.
Det kan hända att man i kollektivavtalet har kommit överens om andra villkor och du får lön för en längre tid.
Arbetsgivaren har rätt att kräva ett läkarintyg för den tid då du är sjuk.
Om du blir sjuk och inte kan arbeta ska du utan dröjsmål meddela detta till din chef.
Din chef berättar för dig om du behöver ett läkarintyg om sjukdomen direkt eller först från och med den fjärde sjukledighetsdagen.
Sjukledighet är ingen semester utan den beviljas för att du ska återhämta dig från din sjukdom.
Därför får du under dessa dagar inte göra något som kan äventyra ditt tillfrisknande.
Sjukdagpenningfinska _ svenska _ engelska
Att ansöka om sjukdagpenningfinska _ svenska _ engelska
Du kan rådfråga om sådant som rör företagets verksamhet eller utveckling av företaget hos företagsrådgivningen.
Läs mer på InfoFinlands sida Företagsrådgivning.
Intressebevakning (edunvalvonta) och andra tjänster för företagare
Finlands Näringsliv EK representerar alla privata branscher och företag i alla storlekar.
Branschförbunden är intressebevakningsorganisationer för företag i olika branscher.
De tillhandahåller sina medlemsföretag ofta också många slags tjänster såsom rådgivning i frågor som rör företagande och den aktuella branschen.
Företagarna i Finland (Suomen Yrittäjät) är företagarnas intressebevakningsorganisation som också producerar sina medlemmar olika tjänster, som till exempel gratis telefonrådgivning i frågor som rör företagande.
Företagarnas stödnät (Yrittäjän tukiverkko) är en gratis webbtjänst som Företagarna i Finland upprätthåller. Tjänsten innehåller mycket nyttig information för företagare.
Tjänsten finns på finska och svenska.
TE-byrån tillhandahåller tjänster som stöder utvecklingen av affärsverksamheten.
Via TE-byrån kan du även leta en fortsättare för din företagsverksamhet eller en partner till ditt företag.
linkkiFinlands Näringsliv EK:
Intressebevakning för företagarefinska _ svenska _ engelska
linkkiFöretagarna i Finland:
Intressebevakning för företagarefinska _ svenska _ engelska
linkkiArbets- och näringsministeriet:
Tjänster för företagarefinska _ svenska _ engelska
Företagsfinland erbjuder en gratis telefontjänst där du får sakkunnig rådgivning om ditt företag har ekonomiska svårigheter.
Rådgivning ges på finska och svenska.
Ekonomihjälp-rådgivningen
på finska, tfn 029 502 4880
på svenska, tfn 029 502 4881
Tjänsten har öppet måndag till fredag kl. 9.00–16.00.
linkkiFöretagsFinland:
Ekonomisk rådgivning för företagarefinska _ svenska
Företagarens utkomstskydd för arbetslösa
Också företagaren har rätt till utkomstskydd för arbetslösa.
En företagare är arbetslös när han eller hon har lagt ned sin företagsverksamhet eller sålt sin andel av företaget.
Företagandet kan också upphöra om företaget säljs, avvecklas, går i konkurs, försätts i likvidation eller på grund av skilsmässa.
Företagaren betraktas som arbetslös också om man har haft ett uppehåll på minst fyra månader i företagsverksamheten.
Om du måste lägga ned din företagsverksamhet, ska du omgående anmäla dig som arbetslös arbetssökande via TE-byråns webbtjänst.
Du kan få arbetslöshetsersättning tidigast från den dag då du gjort anmälan vid TE-byrån.
Information om företagarens sociala trygghetfinska _ svenska _ engelska
Information om arbetsgivarens socialskyddsavgifterfinska _ svenska
linkkiFöretagsFinland:
Information om utkomstskyddet för arbetslösafinska _ svenska _ engelska
Information om utkomstskyddet för arbetslösafinska _ svenska _ engelska
Om du vill få inkomstrelaterat utkomstskydd för arbetslösa, ska du ansluta dig som medlem i företagarnas arbetslöshetskassa (yrittäjien työttömyyskassa).
Om din företagsverksamhet upphör, kan du ansöka om inkomstrelaterad dagpenning (ansiosidonnainen päiväraha) vid arbetslöshetskassan.
Du kan få inkomstrelaterad dagpenning från företagarnas arbetslöshetskassa om du har bedrivit företagsverksamhet och varit medlem i kassan tillräckligt länge innan du blev arbetslös.
Den inkomstrelaterade dagpenningen är större än grunddagpenningen eller arbetsmarknadsstödet.
Hur stor inkomstrelaterad dagpenning du får beror på hur stora förvärvsinkomster du angett som grund för arbetslöshetsförsäkringen.
linkkiFöretagarnas Arbetslöshetskassa i Finland:
Företagarnas Arbetslöshetskassa i Finlandfinska _ svenska
linkkiYrkesutövarnas och företagarnas arbetslöshetskassa:
Yrkesutövarnas och företagarnas arbetslöshetskassafinska _ svenska _ engelska _ ryska _ estniska
Grunddagpenning
Fpa kan betala grunddagpenning (peruspäiväraha) för en arbetslös företagare som inte är medlem i en arbetslöshetskassa.
Om du uppfyller arbetsvillkoret för företagare och omfattas av den sociala tryggheten i Finland kan du få grunddagpenning.
På FPA:s webbplats finns en räknare som du kan använda för att beräkna om du uppfyller arbetsvillkoret för företagare.
Arbetsmarknadsstöd
Om du inte har rätt till grunddagpenning eller inkomstrelaterad dagpenning, men omfattas av den sociala tryggheten i Finland, kan du ansöka om arbetsmarknadsstöd.
Arbetsmarknadsstödet är behovsprövat, vilket betyder att dina andra inkomster och din situation som en helhet påverkar dess belopp.
Företagarens företagshälsovård (työterveyshuolto)
En företagare och andra som arbetar åt sig själv kan ordna företagshälsovård för sig själv om de så önskar.
Företagare måste inte ordna företagshälsovård för sig själv, men däremot måste de ordna det för sina anställda.
Företagshälsovård kan ordnas på den lokala hälsovårdscentralen (terveyskeskus) eller till exempel en privat läkarstation.
Läs mer på InfoFinlands sida Företagshälsovård.
Information för företagare om företagshälsovårdenfinska _ svenska _ engelska
Om en företagare blir sjuk
Om du blir sjuk, kan du få sjukdagpenning (sairauspäiväraha) från Fpa. Den ersätter inkomstbortfallet på grund av arbetsoförmåga när arbetsoförmågan varar mindre än ett år.
Betalningen av dagpenning inleds efter en självrisktid (omavastuuaika).
För företagare är självrisktiden oftast dagen för insjuknandet och följande tre vardagar.
Företagarens sjukdagpenningfinska _ svenska _ engelska
Var får jag hjälp med problem i arbetslivet?
Prata först med din chef.
Om det inte hjälper, kontakta arbetsplatsens förtroendeman.
Om det inte finns en förtroendeman på arbetsplatsen och du är medlem i facket, kontakta ditt fackförbund.
Finlands Fackförbunds Centralorganisation FFC erbjuder gratis anställningsrådgivning.
Du kan få rådgivning även om du inte är medlem i ett fackförbund.
Juristerna svarar på dina frågor på finska och engelska.
Rådgivning ges både per telefon och via e-post:
Tfn 0800 414 004, tis. och ons. kl. 9–11 och 12–15
Du kan även ringa arbetarskyddsmyndigheternas riksomfattande rådgivningstelefon:
Tfn 0295 016 620
Mån.–fre. kl. 9–15
linkkiArbetarskyddsförvaltning:
Kontaktuppgifter till arbetarskyddsmyndigheternafinska _ svenska _ engelska
Min anställning upphör inom kort.
Hur påverkar det mitt uppehållstillstånd?
Detta beror på vilket slags uppehållstillstånd du har.
Om ditt uppehållstillstånd är kopplat till endast en arbetsgivare, ska du ansöka om ett nytt uppehållstillstånd för arbetstagare.
För att kunna ansöka om ett nytt uppehållstillstånd för arbetstagare måste du ha ett nytt jobb.
Du kan även ansöka om uppehållstillstånd på någon annan grund.
Läs mer om grunderna för uppehållstillstånd i InfoFinlands avsnitt Icke EU-medborgare.
Om din anställning upphör innan ditt uppehållstillstånd går ut, ska du meddela detta skriftligt till Migrationsverket.
Också din arbetsgivare kan göra anmälan.
Om ditt uppehållstillstånd är beviljat för en viss bransch, kan du byta jobb inom samma bransch.
Information om uppehållstillstånd för arbetstagare och företagare hittar du på sidorna Arbeta i Finland och Till Finland som företagare.
Läs mer om att söka jobb i Finland på sidan Var hittar jag jobb?
Mer information om att söka arbetslöshetsersättning hittar du på sidan Arbetslöshetsförsäkring.
Information om uppehållstillståndfinska _ svenska _ engelska
Jag har fått för lite lön utbetalad.
Vad ska jag göra?
Kontrollera alltid i lönespecifikationen att du har fått rätt belopp.
Om du har fått för lite lön, ska du be din arbetsgivare att rätta till löneutbetalningen.
Om arbetsgivaren inte betalar ut rätt lön, ska du fråga om råd hos regionförvaltningsverkets arbetarskydd eller ditt fackförbund.
Om du inte kan komma överens om löneutbetalningen med din arbetsgivare måste ärendet avgöras i domstol.
Detta är dock det sista alternativet.
linkkiArbetarskyddsförvaltning:
Information om löneutbetalningfinska _ svenska _ engelska
Min arbetsgivare vill endast betala ut lönen i kontanter.
Får man göra så?
Din arbetsgivare borde betala ut lönen till ditt bankkonto.
Lönen får endast betalas ut i kontanter om inga andra alternativ finns.
Så gör man till exempel om du inte har ett bankkonto.
Om du får lönen utbetalad i kontanter, ska du ge din arbetsgivare ett skriftligt intyg om löneutbetalningen.
På så sätt kan man bevisa att lönen verkligen har betalats till dig.
Min tillsvidareanställning upphörde, men min sista lön betalades inte ut.
Vad bör jag göra?
Fråga arbetsgivaren varför lönen blivit försenad.
Kräv att arbetsgivaren betalar ut lönen.
Framför kravet skriftligt.
Om du är medlem i ett fackförbund kan du be förbundet om hjälp.
Om du inte är medlem i ett fackförbund, kontakta till exempel arbetarskyddsmyndigheterna.
Jag avslutade mitt jobb hos min förra arbetsgivare, men jag har inte fått ett arbetsintyg.
Hur får jag arbetsintyget?
Arbetsgivare behöver inte ge dig ett arbetsintyg på eget bevåg.
Om du vill ha ett arbetsintyg ska du be om det.
Intyget ska lämnas till dig så snart som möjligt.
Om du har bett om ett arbetsintyg men inte fått det, ska du kontakta arbetarskyddsmyndigheterna.
Läs mer på InfoFinlands sida Arbetsintyg.
Jag upplever att jag blir osakligt bemött på min arbetsplats.
Vad kan jag göra?
Alla arbetstagare ska behandlas jämlikt och lika.
Enligt lag får ingen diskrimineras till exempel av följande orsaker:
anställningsform
ålder
kön
etnisk bakgrund
hälsotillstånd
religion
sexuell läggning.
Läs mer på InfoFinlands sida Diskriminering och rasism.
Förutom diskriminering kan det även förekomma andra typer av osakligt bemötande på arbetsplatser, till exempel mobbning eller sexuella trakasserier.
Om hen inte kan hjälpa dig, ska du kontakta arbetsplatsens arbetarskyddsfullmäktige eller förtroendeman.
Om ärendet inte kan lösas på arbetsplatsen, kontakta arbetarskyddsmyndigheterna eller ditt fackförbund.
Om din chef behandlar dig osakligt, anmäl detta till arbetarskyddsmyndigheterna.
Du kan göra anmälan med ditt eget namn eller anonymt.
Jag tvingas att utföra ett jobb utan att få betalt.
Min arbetsgivare hotar mig dessutom med våld.
Var kan jag få hjälp?
Du har rätt till hjälp och skydd.
Enligt lagen i Finland måste arbetstagarna behandlas väl och de ska betalas lön.
Människohandel är ett brott i Finland.
Läs mer på InfoFinlands sida Människohandel och tvångsarbete.
Du hittar information om arbetstagarens rättigheter och skyldigheter i Finland på InfoFinlands sida Arbetstagarens rättigheter och skyldigheter.
Hjälp till offer för människohandelfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska _ polska _ rumänska _ bulgariska
Alla har rätt till företagshälsovård
I Finland är arbetsgivare skyldiga att ordna förebyggande företagshälsovård för sina anställda.
Arbetsgivaren kan också ordna sjukvårdstjänster för sina anställda.
Inom företagshälsovården har arbetstagaren tillgång till hälsovårdarens, företagsläkarens och företagspsykologens tjänster.
Ofta finns det i företagshälsovården också fysioterapeuter.
Specialisternas tjänster ingår vanligen inte i företagshälsovården.
Fråga din arbetsgivare vad företagshälsovården på din arbetsplats omfattar.
Rätten till företagshälsovårdens tjänster omfattar inte den anställdas familj.
Avsikten med företagshälsovården är att främja hälsan och arbetsförmågan och samarbetet på arbetsplatserna.
Anställda inom företagshälsovården har sekretessplikt.
De lämnar inte ut information om din situation till din arbetsgivare, om inte du själv har gett tillstånd till det.
Företagshälsovården kan dock ge din arbetsgivare en bedömning av huruvida ditt hälsotillstånd tillåter att du fortsätter att arbeta.
Fpa ersätter arbetsgivaren och företagaren en del av kostnaderna för företagshälsovården, om dessa är nödvändiga och rimliga.
linkkiArbetarskyddsförvaltningen:
Information om företagshälsovårdenfinska _ svenska _ engelska
linkkiArbetshälsoinstitutet:
Information om företagshälsovårdenfinska _ svenska
linkkiSocial- och hälsovårdsministeriet:
Företagshälsovårdfinska _ svenska _ engelska
Lagen om företagshälsovårdfinska _ svenska _ engelska
Sjukdagpenningfinska _ svenska _ engelska
Tillstånd eller anmälan
Etableringsanmälan
Försäkringar
Bokföring
Beskattning
Inkomstregistret
Ansvar för arbetstagarnas inskolning och säkerhet
När du inleder företagsverksamheten har du många skyldigheter, bland annat ska du registrera företaget och ordna beskattning och bokföring.
Tillstånd eller anmälan
I Finland får man driva en laglig näring som följer god sed utan ett tillstånd som beviljas av myndigheter.
I vissa fall behövs det dock ett tillstånd från myndigheter för att starta företagsverksamhet, eller också måste man anmäla verksamheten till myndigheter.
Till exempel ska lokaler där man säljer livsmedel eller idkar skönhetsvård kontrolleras och tillstånd sökas hos kommunens hälsomyndighet innan lokalerna tas i bruk.
Innan du startar företagsverksamheten, kontrollera om du behöver tillstånd för verksamheten eller om du måste anmäla verksamheten till en myndighet.
Du kan kontrollera hos regionförvaltningsverken eller på Företagsfinlands webbplats om du behöver ett tillstånd för ditt företag.
linkkiFöretagsfinland:
Tillstånd och anmälan som är anknutna till idkandet av en näringfinska _ svenska _ engelska
Etableringsanmälan
Ny företagsverksamhet ska anmälas till handelsregistret som upprätthålls av Patent- och registerstyrelsen (Patentti- ja rekisterihallitus).
Du kan använda samma blankett när du gör etableringsanmälan för ditt företag till Patent- och registerstyrelsen och till Skatteförvaltningen.
linkkiPatent- och registerstyrelsen:
Anmälan om grundande av ett företagfinska _ svenska _ engelska
Försäkringar
Företagarpensionsförsäkringen (FöPL) (YEL-vakuutus) är obligatorisk för företagare i åldern 18–68 år, vars företagsverksamhet inbringar minst 7 645,25 euro om året som arbetsinkomst (år 2018).
Pensionsförsäkringen tryggar företagarens utkomst då företagsverksamheten upphör på grund av invaliditet eller ålder och den ger företagarens anhöriga ett familjepensionsskydd efter att företagaren har dött.
Pensionsförsäkringar fås antingen genom försäkringsbolag eller pensionskassor (eläkekassa).
Teckna en pensionsförsäkring senast när det har gått sex månader sedan du startade företagsverksamheten.
En ny företagare får en rabatt på 22 procent på pensionspremierna under de fyra första åren.
Storleken av försäkringspremierna och pensionen beror på hur stor förvärvsinkomst (työtulo) förtagaren har.
Den som ger försäkringen och företagaren kommer överens om förvärvsinkomstens storlek när företagaren tecknar företagarpensionsförsäkringen.
Förvärvsinkomsten ska vara ungefär lika stor som företagarens genomsnittliga lön skulle vara om han eller hon skulle utföra liknande arbete som anställd.
Förvärvsinkomstens storlek inverkar också på storleken av olika inkomstrelaterade förmåner (ansiosidonnanen etuus), såsom sjukdagpenningen.
Du ska teckna en pensionsförsäkring (ArPL-försäkring) (eläkevakuutus (TyEL-vakuutus)) och en olycksfallsförsäkring som omfattar en grupplivförsäkring och en arbetslöshetsförsäkring för de anställda.
Arbetsgivaren betalar arbetstagarens socialskyddsavgifter till skattemyndigheten i anslutning till skatteinnehållningen.
I vissa branscher finns också andra obligatoriska försäkringar.
Du bör också överväga andra frivilliga försäkringar som till exempel företagarens olycksfallsförsäkring.
linkkiPensionsskyddscentralen:
Information om företagarpensionsförsäkringenfinska _ svenska _ engelska
linkkiPensionsskyddscentralen:
Information om att teckna försäkringar för anställdafinska _ svenska _ engelska
linkkiFöretagsFinland:
Information om att teckna försäkringar för anställdafinska _ svenska _ engelska
Bokföring
I Finland har alla företagare bokföringsskyldighet.
Om du inte vill sköta bokföringen själv, kan du anlita en revisionsbyrå som sköter företagets bokföring åt dig.
I Finland anlitar många företag revisionsbyråer.
Beskattning
Företagsformen påverkar företagets beskattning.
Detta är det bra att beakta när du väljer företagsform.
En ny företagare kan anmäla sig till Skatteförvaltningens förskottsuppbördsregister.
Anmälan till förskottsuppbördsregistret görs med samma anmälan som görs för grundande av företaget, d.v.s. etableringsanmälan (yrityksen perustamisilmoitus).
Om ditt företag är i förskottsuppbördsregistret kan du fakturera kunder utan förskottsinnehållning.
Skatter betalas på de inkomster som företagaren eller företaget har kvar när alla kostnader för företagsverksamheten har dragits av försäljningen.
Företagets skatter betalas på basis av de beskattningsbara inkomsterna, vars belopp man uppskattar på förhand.
Uppskattningen baseras på beloppet av de beskattningsbara inkomsterna året innan.
I ett nytt företag uppskattar företagaren själv storleken av den beskattningsbara inkomsten och meddelar denna till skattmyndigheten.
linkkiSkatteförvaltningen:
Information om beskattningen av företag och företagarefinska _ svenska _ engelska
linkkiFöretagsFinland:
Information om beskattningen av företag och företagarefinska _ svenska _ engelska
Mervärdesskatt
Mervärdesskatten (arvonlisävero) är en konsumtionsskatt som i Finland betalas för nästan alla varor och tjänster.
Företagare som säljer varor och tjänster i Finland är skyldiga att betala mervärdesskatt.
Om inkomsten som man får för försäljningen av varor och tjänster är mindre än 10 000 euro per år, behöver ingen mervärdesskatt betalas på den.
Företagsformen påverkar inte mervärdesskattens belopp.
Mervärdesskattebeloppet varierar emellertid för olika produkter.
Beskattning av en enskild näringsidkare
Den vanligaste företagsformen är en enskild näringsidkare, vilket betyder att man driver företagsverksamhet utan ett skilt grundat företag.
Den som är en enskild näringsidkare beskattas på så sätt att alla inkomster som återstår efter att man har dragit av kostnaderna för företagsverksamheten är beskattningsbara inkomster.
Företagaren betalar alltså inte skilt ut en lön åt sig.
Inkomsten beskattas utifrån företagets förmögenhet antingen som kapitalinkomst (pääomatulo) eller som förvärvsinkomst (ansiotulo).
Skatteprocenten på kapitalinkomsten är alltid densamma.
Förvärvsinkomsten beskattas progressivt, d.v.s. ju större inkomster man har, desto mer skatt betalar man.
Inkomstregistret
Inkomstregistret är en databas dit arbetsgivarna anmäler lönerna som de utbetalat till sina anställda.
Anmälan ska göras senast fem dagar efter löneutbetalningen.
Uppgifterna ska skickas till inkomstregistret elektroniskt:
direkt via lönesystemet om det har en inbyggd teknisk förbindelse till Inkomstregistret eller
via Inkomstregistrets ärendehantering, till vilken man får tillträde med webbankkoder eller andra medel för elektronisk identifiering.
Löneuppgifterna kan endast i undantagsfall anmälas med ett pappersformulär.
Läs mer om Inkomstregistret och om att anmäla löner på Inkomstregistrets webbplats.
linkkiSkatteförvaltningen:
Inkomstregistretfinska _ svenska _ engelska _ ryska _ estniska _ kinesiska
Ansvar för arbetstagarnas inskolning och säkerhet
Som företagare har du ansvaret för att ge arbetstagarna inskolning i arbetsuppgifterna.
Arbetsgivaren ska introducera förhållandena på arbetsplatsen och de rätta arbetsmetoderna för arbetstagaren.
Arbetsgivaren är också skyldig att sörja för arbetstagarnas säkerhet och hälsa i arbetet.
Arbetsgivaren ska utarbeta ett verksamhetsprogram för arbetarskyddet (työsuojelun toimintaohjelma) som tar upp de säkerhets- och hälsorelaterade riskerna på arbetsplatsen och hur man undgår dem.
linkkiArbetarskyddscentralen:
Information om arbetarskyddfinska _ svenska _ engelska
Arbetstagaren har rätt att på begäran få ett arbetsintyg av arbetsgivaren när anställningen upphör.
Arbetsintyget är ett viktigt dokument där anställningens längd och arbetsuppgifterna nämns.
Arbetstagaren kan också be att orsaken till att anställningen upphört och en bedömning av arbetstagarens färdigheter och uppförande antecknas i intyget.
Arbetsgivaren är skyldig att utfärda ett arbetsintyg ännu tio år efter att anställningen har upphört och efter detta endast om detta inte medför en orimlig olägenhet för arbetsgivaren.
Om arbetstagaren vill att en bedömning av färdigheterna och uppförandet antecknas i arbetsintyget måste arbetsgivaren utfärda ett sådant intyg ännu fem år efter att anställningen har upphört till arbetstagaren på hans eller hennes begäran.
Arbetsgivare måste också ge arbetstagaren ett nytt arbetsintyg om arbetstagarens arbetsintyg kommer bort eller förstörs.
En arbetsgivare som avsiktligt eller av vårdslöshet inte utfärdar ett arbetsintyg bryter mot arbetsavtalslagen.
Arbetsavtalslagenfinska _ svenska _ engelska
linkkiArbetarskyddsförvaltningen:
Information om rätten till arbetsintygfinska _ svenska _ engelska
Arbetarskyddsverksamhet på arbetsplatsen
I Finland fästs stor uppmärksamhet vid arbetssäkerhet.
Arbetsgivaren ansvarar för att alla kan arbeta tryggt.
Arbetsgivaren ska ordna arbetsplatsintroduktion för nya anställda.
Arbetsgivaren är också skyldig att göra de anställda förtrogna med arbetsplatsens säkerhetsanvisningar och lära dem korrekta arbetssätt.
De anställda ska också själva sörja för arbetssäkerheten.
Arbetet ska utföras enligt anvisningarna.
Om arbetet är uppenbart farligt kan den anställda vägra att utföra det.
På arbetsplatserna ska det finnas tillräckligt många personer med kunskaper i första hjälpen, första hjälpen-utrustning samt instruktioner för olycksfall.
Arbetsgivarna ordnar utbildning i första hjälpen på arbetsplatsen.
Om det finns minst tio anställda på en arbetsplats väljer dessa ut en arbetarskyddsfullmäktig som representerar dem.
Arbetarskyddsfullmäktige gör sig insatt i arbetarskyddsfrågor som gäller arbetsplatsen, deltar i arbetsplatsens arbetarskyddsinspektioner och informerar de anställda om ärenden som rör arbetets säkerhet och hälsa.
Arbetsgivaren utser för varje arbetsplats en arbetarskyddschef, som bistår arbetsgivaren i samarbetet med anställda och arbetarskyddsmyndigheter.
Arbetarskyddsmyndigheter
I Finland finns det fem ansvarsområden för arbetarskydd som lyder under Regionförvaltningsverket (RFV).
Ansvarsområdena övervakar att de lagenliga arbetarskyddsföreskrifterna följs på arbetsplatserna.
Ansvarsområdena för arbetarskydd ger både arbetstagare och arbetsgivare råd i frågor som gäller arbetets säkerhet och hälsa samt i frågor som rör anställningsvillkor.
Arbetarskyddsinspektörerna utför kontroller på arbetsplatser.
De kontrollerar bland annat om säkerhetsföreskrifterna följs på arbetsplatsen, om man har gett tillräcklig introduktion i arbetet och huruvida utländska arbetstagares arbetsförhållanden och anställningsvillkor följer finländska lagar och avtal.
Arbetarskyddsinspektören har rätt att få tillträde till varje arbetsplats och tillgång till de dokument som är väsentliga för övervakningen av arbetarskyddet.
Arbetarskyddsmyndigheten kan förplikta arbetsgivaren att rätta till brister i arbetssäkerheten som förekommer på arbetsplatsen
linkkiArbetarskyddsförvaltningen:
Information om arbetarskydd och råd vid problemfinska _ svenska _ engelska
linkkiEuropeiska arbetsmiljöbyrån:
Information om arbetarskyddfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Företagarens skyldigheter
Behöver jag ett tillstånd för företaget?
Vilka försäkringar måste jag ha?
Läs mer om dessa och andra viktiga frågor som en företagare bör veta på InfoFinlands sida Företagarens skyldigheter.
Stöd till företagare
Vem sköter företagarnas intressebevakning i Finland?
Hurdant utkomstskydd för arbetslösa får företagare i Finland?
Läs mer på InfoFinlands sida Stöd till företagare.
Den finländska företagskulturen
Om du vill driva ett framgångsrikt företag i Finland, är det viktigt att du känner till den finländska företagskulturen.
När du känner igen grundläggande drag i den finländska företagskulturen kan du bättre betjäna dina kunder. Du har också bättre insikt i vad folk förväntar av dig.
Läs mer på InfoFinlands sida Den finländska arbetskulturen.
När ett barn föds till familjen har föräldrarna rätt att ta familjeledighet, det vill säga stanna hemma för att ta hand om barnet.
Med familjeledighet avses
moderskapsledighet
faderskapsledighet
föräldraledighet
vårdledighet
Meddela din arbetsgivare om familjeledigheten senast två månader innan den börjar.
Familjeledigheterna är vanligen oavlönad ledighet.
Huruvida du får lön under familjeledigheten beror på ditt kollektivavtal.
Kontrollera detta med din arbetsgivare.
FPA betalar ut familjeförmåner för familjeledigheten: föräldrapenning och stöd för hemvård av barn.
Läs om villkoren för familjeförmånerna på InfoFinlands sida Stöd efter barnets födelse och Stöd för vård av barn i hemmet.
När familjeledigheterna upphör har arbetstagaren rätt att återvända till sitt eget arbete eller motsvarande arbete på den gamla arbetsplatsen.
Arbetsavtalet för en gravid kvinna får inte hävas och hon får inte diskrimineras på grund av sin graviditet.
I Finland känner arbetsgivarna och arbetstagarna till familjeledigheterna och de används allmänt.
linkkiArbets- och näringsministeriet:
Familjeledigheterfinska _ svenska _ engelska
Information om stöd till barnfamiljerfinska _ svenska _ engelska
Moderskapsledighet
Moderskapsledigheten är 105 vardagar.
Arbete under moderskapsledigheten är tillåtet om det kan utföras utan att moderns, fostrets eller barnets säkerhet äventyras.
Under moderskapsledigheten får man dock inte arbeta under de två veckor som föregår det beräknade födelsedatumet och under två veckor efter förlossningen.
Faderskapsledighet
Faderskapsledigheten är den del av föräldraledigheten som är avsedd att tas ut av fadern.
Faderskapsledigheten är allt som allt 54 vardagar.
Dessa dagar kan inte överföras till modern.
Du kan ta ut högst 18 dagar av din faderskapsledighet samtidigt som barnets mor är moderskaps- eller föräldraledig.
Dessa dagar kan du dela upp på högst fyra perioder.
De återstående 36 dagarna kan du dela upp på högst två perioder.
Under dessa dagar kan modern inte vara moderskapsledig samtidigt.
Avsikten är att fadern tar hand om barnet.
Du kan också ta ut alla 54 dagar av din faderskapsledighet vid olika tider med modern.
Du kan själv bestämma om du tar ut hela faderskapsledigheten eller bara en del av dagarna.
Faderskapsledigheten får endast tas ut före barnet har fyllt två år.
När barnet fyller två år kan du inte längre ta ut faderskapsledighet trots att du har dagar kvar.
Föräldraledighet
Efter moderskapsledigheten kan antingen modern eller fadern stanna hemma för att ta hand om barnet. Föräldraledigheten varar 158 vardagar.
Båda föräldrarna kan inte vara föräldralediga samtidigt.
Däremot kan man dela upp föräldraledigheten så att modern eller fadern stannar hemma växelvis för att ta hand om barnet.
Vårdledighet
Efter föräldraledigheten kan antingen modern eller fadern ta ut en oavlönad vårdledighet för att ta hand om barnet tills barnet fyller tre år.
Det förutsätter att modern eller fadern varit anställd hos samma arbetsgivare minst sex månader under det senaste året.
Under vårdledigheten betalar FPA stöd för hemvård av barn.
Se villkoren för stödet för hemvård av barn på InfoFinlands sida Stöd för vård av barn i hemmet.
Partiell vårdledighet
Du kan också vara vårdledig på deltid.
Då arbetar du kortare dagar och får på motsvarande sätt mindre lön.
Makarna kan vara partiellt vårdlediga samtidigt så att den ena förkortar sin arbetstid från morgonen och den andra från eftermiddagen.
Du kan vara partiellt vårdledig tills barnet har gått ut årskurs två.
Om du har hemkommun i Finland kan du ansöka om partiell vårdpenning hos FPA för hemvård av barn under tre år eller skolbarn i årskurserna 1 eller 2.
Partiell vårdpenning betalas inte för vård av ett barn som fyllt tre men ännu inte går i skolan.
Läs mer om partiell vårdpenning på InfoFinlands sida Stöd för vård av barn i hemmet.
Allmänt om fackförbund
I Finland tryggar lagen arbetstagarnas rätt att höra till ett fackförbund (ammattiliitto).
Denna rätt kan inte begränsas med avtal.
Diskriminering av arbetstagare på grund av deras medlemskap i fackförbund är straffbart.
De flesta finländare är med i något fackförbund.
Fackförbunden strävar efter att trygga sina medlemmars intressen och rättigheter, försöker förbättra lönerna och anställningsskyddet samt förbättra arbetslivets kvalitet.
Arbetstagarförbunden är organiserade under tre centralförbund för löntagare.
Dessa är Finlands Fackförbunds Centralorganisation FFC, Tjänstemannacentralorganisationen STTK och Centralorganisationen för högutbildade i Finland Akava.
linkkiFCC, STTK och AKAVA:
Fackets ABC-bokfinska _ engelska _ ryska _ estniska
linkkiCentralorganisationen för högutbildade i Finland Akava:
Information om fackförbundsverksamhetfinska _ svenska _ engelska
Information om fackförbundsverksamhetfinska _ svenska _ engelska
linkkiTjänstemannacentralorganisationen STTK:
Information om fackförbundsverksamhetfinska _ svenska _ engelska
Att ansluta sig till ett fackförbund och medlemsavgiften
Om du vill kan du ansluta dig till fackförbundet i din egen bransch.
Du kan ansluta dig till ett fackförbund genom att ta kontakt med förtroendemannen på din egen arbetsplats eller genom att kontakta fackförbundet direkt.
Till de flesta fackförbund kan man också ansluta sig genom att fylla i en anslutningsblankett på fackets webbplats.
Fackförbundets medlemmar betalar förbundet en medlemsavgift som vanligen är cirka 1–2 procent av lönen.
Medlemsavgiften får dras av i beskattningen.
Fackförbundets medlemmar kan delta i utbildning och fritidsaktiviteter som förbundet ordnar.
De får också stöd av förbundets förtroendeman vid konflikter på arbetsplatsen.
Vid behov får man också råd eller förhandlingsstöd från fackförbundet.
Arbetslöshetskassa
I Finland finns ett frivilligt system med arbetslöshetskassor.
En arbetstagare som är medlem i en arbetslöshetskassa betalar en medlemsavgift till arbetslöshetskassan när han eller hon förvärvsarbetar.
Om arbetet upphör och arbetstagaren blir arbetslös kan han eller hon ansöka om inkomstrelaterad arbetslöshetsdagpenning från kassan.
Det lönar sig att ansluta sig till en arbetslöshetskassa, eftersom den inkomstrelaterade dagpenningen är större än det vanliga utkomstskyddet för arbetslösa.
När du ansluter dig till ett fackförbund kan du samtidigt ansluta dig till förbundets arbetslöshetskassa.
Fackförbundet och arbetslöshetskassan är dock två separata system.
Det finns också arbetslöshetskassor som man kan ansluta sig till utan att vara medlem i något fackförbund.
För att få inkomstrelaterad dagpenning finns några villkor som måste uppfyllas innan det är möjligt att få dagpenning.
Till exempel ska man ha varit med i arbetslöshetskassan en viss tid före man blir arbetslös.
Ta reda på dessa villkor genast när du ansluter dig till arbetslöshetskassan.
Läs mer på InfoFinlands sida Utkomstskydd för arbetslösa.
linkkiArbetslöshetskassornas samorganisation:
information om arbetslöshetskassorfinska _ svenska _ engelska
Fackförbundets representant på arbetsplatsen
På arbetsplatsen representeras fackförbundet och de anställda som är medlemmar i det av förtroendemannen.
Förtroendemannen väljs av de anställda.
Förtroendemannen agerar som förhandlare, medlare och informationsförmedlare mellan arbetsgivaren och anställda.
Man kan också vända sig till förtroendemannen till exempel med frågor om kollektivavtalet.
När du grundar ett företag måste du välja företagsform och ett namn för företaget samt definiera branschen.
På valet av företagsform inverkar bland annat antalet grundare, behovet av kapital, fördelningen av ansvar och bestämmanderätt, finansieringen och beskattningen.
Olika företagsformer i Finland är enskild näringsidkare (toiminimi); öppet bolag (avoin yhtiö); kommanditbolag (kommandiittiyhtiö); aktiebolag (osakeyhtiö) och andelslag (osuuskunta).
När du funderar på vilken företagsform du ska välja, är det absolut tillrådligt att du kontaktar företagsrådgivningen.
Enskild näringsidkare (toiminimi)
Det enklaste och vanligaste sättet att starta företagsverksamhet är att som enskild näringsidkare driva en firma.
Du har bestämmanderätt över och ansvar för firmans ärenden och företaget kan anställa medarbetare precis som andra företag.
Företagsverksamhet som bisyssla lönar det sig ofta att starta som enskild näringsidkare.
Det är snabbt och enkelt att starta företagsverksamhet som enskild näringsidkare.
För att grunda ett aktiebolag behövs minst en person eller ett samfund med ett minsta aktiekapital på 2 500 euro, med andra ord ska det sammanlagda värdet av aktierna uppgå till minst 2 500 euro.
Aktieägarens rösträtt, vinster och ansvar i företaget beror på hur många av bolagets aktier han eller hon äger.
Ett öppet bolag bildas då två eller fler personer kommer överens om att grunda ett bolag genom att teckna ett bolagsavtal.
Bolagsmännen, d.v.s. personerna som tillsammans äger bolaget, är jämställda i all verksamhet som bolaget driver och de ansvarar tillsammans och personligen för bolagets beslut, förbindelser och skulder.
Ett kommanditbolag är ett personbolag som skiljer sig från ett öppet bolag på så sätt att det i kommanditbolaget finns utöver en eller flera ansvariga bolagsmän åtminstone en tyst bolagsman, d.v.s. en person som är delägare i företaget. Vanligen är den tysta bolagsmannen en investerare.
Det behövs minst tre personer för att grunda ett andelslag.
Ett andelslag kan ha en eller fler medlemmar.
På andelslagets stämma har varje medlem en röst.
Medlemmarna ansvarar för andelslagets förpliktelser (till exempel skulder) endast med det belopp som de investerat i andelslaget.
linkkiFöretagsFinland:
Information om företagsformerfinska _ svenska _ engelska
Om du blir sjuk eller råkar ut för en olycka har du rätt att stanna hemma från arbetet.
Arbetsgivaren är skyldig att betala lön för sjukledigheten.
Om din anställning varat över en månad före insjuknandet får du lönen till fullt belopp för minst den dag då du insjuknade och nio därefter följande dagar.
Om du fortfarande inte kan återvända till arbetet kan du söka sjukdagpenning (sairauspäiväraha) hos FPA om du omfattas av den finländska sjukförsäkringen.
Läs mer på InfoFinlands sida Den sociala tryggheten i Finland.
Det kan hända att man i kollektivavtalet har kommit överens om andra villkor och du får lön för en längre tid.
Arbetsgivaren har rätt att kräva ett läkarintyg för den tid då du är sjuk.
Om du blir sjuk och inte kan arbeta ska du utan dröjsmål meddela detta till din chef.
Din chef berättar för dig om du behöver ett läkarintyg om sjukdomen direkt eller först från och med den fjärde sjukledighetsdagen.
Sjukledighet är ingen semester utan den beviljas för att du ska återhämta dig från din sjukdom.
Därför får du under dessa dagar inte göra något som kan äventyra ditt tillfrisknande.
Sjukdagpenningfinska _ svenska _ engelska
Att ansöka om sjukdagpenningfinska _ svenska _ engelska
Arbetsavtalet upprättas i två exemplar, ett till den anställda och ett till arbetsgivaren.
Arbetsavtalet innehåller vanligen åtminstone följande punkter:
Parterna som ingår arbetsavtalet
Både arbetsgivaren och den anställda undertecknar arbetsavtalet.
Tidpunkten då arbetet inletts
Om avtalet är tillsvidare gällande eller tidsbundet
Huvudregeln är att arbetsavtalet gäller tillsvidare.
Detta innebär att arbetet pågår tills den anställda säger upp sig eller tills arbetsgivaren säger upp den anställda.
Arbetsgivaren ska ha en välgrundad orsak för att säga upp en anställd.
Godtagbara orsaker för uppsägning definieras i arbetsavtalslagen.
När arbetsavtalet gäller tillsvidare har arbetstagaren en fast eller permanent anställning.
Ett tidsbundet avtal innebär att man har avtalat om tidpunkten då arbetet inleds och avslutas.
Arbetsavtalet kan vara tidsbundet om det finns en välgrundad orsak till detta.
Lagar och kollektivavtal reglerar exakt när tidsbundna anställningar får tillämpas.
En anställning kan vara tidsbunden om orsaken är till exempel
vikariat
praktik
projekt
efterfrågan eller säsongtopp
Om arbetsavtalet är tidsbundet binder det båda parterna en bestämd tid, om man inte har kommit överens om möjligheten till uppsägning.
Ett tidsbundet avtal kan hävas endast av mycket vägande skäl.
Prövotid och längden på den
Man kan komma överens om en prövotid i anställningens början.
Prövotiden kan vara högst sex månader.
Vid en tidsbunden anställning kan prövotiden vara högst hälften av den tid anställningen pågår.
Under prövotiden kan arbetstagaren bedöma om arbetet lämpar sig för honom eller henne och arbetsgivaren kan bedöma om arbetstagaren är lämplig för arbetet.
Under prövotiden kan arbetstagaren och arbetsgivaren häva arbetsavtalet utan uppsägningstid.
Grunderna för hävande av ett arbetsavtal under prövotiden får inte vara diskriminerande.
Arbetstagaren får normal lön under prövotiden.
Platsen för utförandet av arbetet
Arbetsuppgifterna
Lönen och utbetalning av lönen
Lönen bestäms enligt kollektivavtalet.
Om branschen inte har ett kollektivavtal har arbetstagaren rätt till en skälig lön.
Arbetsgivaren får inte betala en lön som är mindre än vad som fastställs i kollektivavtalet.
Lönen kan innehålla olika förmåner.
Typiska lönetillägg i Finland är erfarenhetstillägg, övertidstillägg och skiftarbetstillägg.
Avlöningsdagen är vanligen en eller två gånger i månaden.
Arbetsgivaren betalar in lönen på bankkontot.
Arbetstagaren har rätt att få en lönespecifikation där det står vad lönen består av.
När man talar om lön avser man oftast bruttolönen (bruttopalkka) från vilken skatter och personalbikostnader dras av.
Den lön som betalas till arbetstagaren är nettolönen (nettopalkka).
Arbetstid
I avtalet ska den regelbundna arbetstiden nedtecknas.
Arbetstiden ska följa arbetslagstiftningen och kollektivavtalet.
Semester och semesterpenning
Arbetstagaren har rätt att få samma lön under semestern som under arbetet.
Dessutom betalas en semesterpenning.
Utbetalningen av semesterpenning baserar sig på kollektivavtalet.
När anställningen upphör har arbetstagaren rätt att få semesterersättning för de dagar som han eller hon inte har fått semester eller semesterersättning för vid tidpunkten för anställningens upphörande.
Uppsägningstid
Ett tillsvidare gällande arbetsavtal upphör antingen när arbetstagarens eller arbetsgivarens uppsägningstid har gått ut.
Uppsägningstiden är den tid som arbetstagaren är skyldig att arbeta innan arbetet upphör.
Under uppsägningstiden har arbetstagaren samma rättigheter och skyldigheter och han eller hon får normal lön.
Om arbetsgivaren säger upp en arbetstagare måste arbetsgivaren ange orsaken till detta.
Arbetsavtalslagen beskriver vilka orsaker som är godtagbara för uppsägning.
Omnämnande om viket kollektivavtal arbetsavtalet följer
linkkiArbets- och näringsministeriet:
Arbetsavtal och anställningfinska _ svenska _ engelska
Planera noga
Planera finansieringen för ditt företag noga innan du grundar företaget.
Det är viktigt att du har tillräckligt med kapital i startskedet.
Företagets finansiering kan också delvis bestå av pengar man fått eller lånat. För att ansöka om finansiering ska man ha en ordentlig affärsverksamhetsplan.
Lån
Lån som beviljas av banker eller Finnvera är vanliga finansieringskällor för många nya företagare.
Finnvera är ett specialfinansieringsbolag som ägs av finska staten.
Bolaget beviljar lån och borgen åt nya företag eller företag som redan är verksamma.
Företag som har förutsättningar för lönsam verksamhet, men inte den egenfinansieringsandel eller de garantier som bankerna kräver, kan få ett lån eller borgen för ett lån vid Finnvera.
Vid Företagsfinland får du information om olika finansieringsalternativ.
Fråga även vid arbets- och näringsbyrån om du kan få startstöd för ditt företag.
linkkiFöretagsFinland:
Finansiering för ett företagfinska _ svenska _ engelska
linkkiFinnvera:
Finansiering för ett företagfinska _ svenska _ engelska
Startpeng (starttiraha)
När du startar ett eget företag kan du beviljas en startpeng som tryggar din utkomst under den tid då du inleder din företagsverksamhet.
Startpengen beviljas av den TE-byrå där du är kund.
Den kan beviljas för högst 12 månader.
När du ansöker om startpeng undersöker TE-byrån om företagandet är ett lämpligt alternativ för dig.
Du kan få startpeng om
du är arbetslös arbetssökande
du inte är arbetslös, men du ska gå över till företagande på heltid till exempel från lönearbete, studier eller arbete i hemmet.
Förutsättningar för att få startpeng är bland annat att:
företagsverksamheten är din huvudsyssla
du har tillräckliga kunskaper, färdigheter och resurser för den företagsverksamhet som du planerar
TE-byrån bedömer att företagsverksamheten kan vara lönsam
du behöver startpengen för ditt uppehälle
du startar företagsverksamheten först när stödet har beviljats.
Ta kontakt med TE-byrån så tidigt som möjligt om du ämnar ansöka om startpeng.
Även andra stödformer för nya företagare finns tillgängliga.
Företagsfinland ger upplysningar om olika finansieringsalternativ.
linkkiArbets- och näringsministeriet:
Information om startpengenfinska _ svenska _ engelska
Alla har rätt till företagshälsovård
I Finland är arbetsgivare skyldiga att ordna förebyggande företagshälsovård för sina anställda.
Arbetsgivaren kan också ordna sjukvårdstjänster för sina anställda.
Inom företagshälsovården har arbetstagaren tillgång till hälsovårdarens, företagsläkarens och företagspsykologens tjänster.
Ofta finns det i företagshälsovården också fysioterapeuter.
Specialisternas tjänster ingår vanligen inte i företagshälsovården.
Fråga din arbetsgivare vad företagshälsovården på din arbetsplats omfattar.
Rätten till företagshälsovårdens tjänster omfattar inte den anställdas familj.
Avsikten med företagshälsovården är att främja hälsan och arbetsförmågan och samarbetet på arbetsplatserna.
Anställda inom företagshälsovården har sekretessplikt.
De lämnar inte ut information om din situation till din arbetsgivare, om inte du själv har gett tillstånd till det.
Företagshälsovården kan dock ge din arbetsgivare en bedömning av huruvida ditt hälsotillstånd tillåter att du fortsätter att arbeta.
Fpa ersätter arbetsgivaren och företagaren en del av kostnaderna för företagshälsovården, om dessa är nödvändiga och rimliga.
linkkiArbetarskyddsförvaltningen:
Information om företagshälsovårdenfinska _ svenska _ engelska
linkkiArbetshälsoinstitutet:
Information om företagshälsovårdenfinska _ svenska
linkkiSocial- och hälsovårdsministeriet:
Företagshälsovårdfinska _ svenska _ engelska
Lagen om företagshälsovårdfinska _ svenska _ engelska
Sjukdagpenningfinska _ svenska _ engelska
I Finland bestäms arbetstagarnas rättigheter enligt arbetslagstiftningen och kollektivavtalen (työehtosopimukset).
I dessa fastställs till exempel minimilöner, arbetstider, semestrar, lön för sjukdomstid och uppsägningsvillkor.
Arbetsgivarförbundet och arbetstagarförbundet kommer gemensamt överens om anställningsvillkoren i en viss bransch.
På detta sätt uppstår ett kollektivavtal för branschen.
I den offentliga sektorn (arbetsgivaren är en kommun eller staten) ingås tjänstekollektivavtal eller allmänt kommunalt tjänste- och arbetskollektivavtal.
Förmånerna som man har avtalat om med ett kollektivavtal är alltid minimiförmåner.
Dessa kan inte underskridas i arbetsavtalet.
Lönen kan till exempel inte vara lägre än vad som avtalats med kollektivavtalet.
Arbetsgivaren och arbetstagaren kan ändå i arbetsavtalet komma överens om villkor som är bättre än villkoren i kollektivavtalet.
Kollektivavtalen uppgörs för en viss tid, vanligen för ett eller två år eller också för en längre tid.
Kollektiv- och tjänstekollektivavtalet är bindande för de löntagar- och arbetsgivarförbund som slutit dem och för deras medlemmar.
Ett kollektivavtal kan också vara allmänt bindande.
Då måste även de arbetsgivare som inte hör till arbetsgivarförbundet följa avtalet med sina anställda.
I platsannonser och arbetsavtal kan det stå: ”palkkaus TES:in mukainen” (”avlöning enligt kollektivavtalet”).
Det är bra att ta reda på hur stora lönerna är i den egna branschen i Finland.
Det är viktigt att känna till kollektivavtalet, eftersom det i Finland inte finns till exempel en lag om minimilöner, utan minimilönerna fastställs alltid enligt kollektivavtalet.
linkkiArbets- och näringsministeriet:
Arbetslagstiftningfinska _ svenska _ engelska
Arbetsavtal
Arbetsgivaren ingår vanligen ett skriftligt arbetsavtal med en ny anställd.
I arbetsavtalet fastställs arbetsuppgifterna och lönen samt andra förmåner och villkor.
Avtalet kan också vara muntligt.
Om man inte har uppgjort ett skriftligt arbetsavtal ska arbetsgivaren utan särskild begäran ge en skriftlig redogörelse för de centrala villkoren i arbetet.
Det är rekommendabelt att arbetsavtalet är skriftligt.
När allt finns på papper kan både den anställda och arbetsgivaren kontrollera i avtalet vad man gemensamt har avtalat.
Detta hjälper om det uppstår konflikter i arbetet.
Läs mer om upprättandet av arbetsavtalet på InfoFinlands sida Innehållet i arbetsavtalet.
linkkiArbetarskyddsförvaltningen:
Att uppgöra ett arbetsavtalfinska _ svenska _ engelska
Ett skriftligt avtal om de centrala villkoren i arbetet
Arbetsgivaren ska ge den anställda en skriftlig redogörelse för de centrala villkoren i arbetet vid tillsvidare gällande anställningar samt anställningar som varar över en månad.
Av redogörelsen ska det åtminstone framgå
arbetsgivarens och arbetstagarens hemort eller driftställe
tidpunkten då arbetet inletts
längden på ett tidsbundet arbetsavtal och orsaken till att avtalet är tidsbundet
prövotidens längd
stället där arbetet utförs
den anställdas arbetsuppgifter
kollektivavtalet som tillämpas på arbetet
de grunder enligt vilka lön eller andra vederlag bestäms samt löneperioden
den regelbundna arbetstiden
hur semestern bestäms
uppsägningstiden eller grunden för bestämmande av den
Om arbetsgivaren inte ger en redogörelse för de centrala villkoren i arbetet till den anställda kan han eller hon dömas till böter.
Det viktigaste i affärsverksamhetsplanen är verksamhetsplanen för ditt eget företag. Fundera noga på hurudan verksamhet ditt företag bedriver samt var ditt företag har lokaler och hurudana lokaler det har.
Tänk också på vilka produktionsmedel eller hurudan arbetskraft du behöver.
Anteckna i affärsverksamhetsplanen också hur du tänker ordna bokföringen och ekonomiplaneringen och hur du följer upp realiseringen av dina planer.
Hjälp med att utarbeta affärsverksamhetsplanen
På deras webbplatser kan du också ladda ned företagarhandböcker åtminstone på finska och på engelska.
Där kan du även hämta en mall för affärsverksamhetsplanen och andra dokumentmallar.
Arbetarskyddsverksamhet på arbetsplatsen
I Finland fästs stor uppmärksamhet vid arbetssäkerhet.
Arbetsgivaren ansvarar för att alla kan arbeta tryggt.
Arbetsgivaren ska ordna arbetsplatsintroduktion för nya anställda.
Arbetsgivaren är också skyldig att göra de anställda förtrogna med arbetsplatsens säkerhetsanvisningar och lära dem korrekta arbetssätt.
De anställda ska också själva sörja för arbetssäkerheten.
Arbetet ska utföras enligt anvisningarna.
Om arbetet är uppenbart farligt kan den anställda vägra att utföra det.
På arbetsplatserna ska det finnas tillräckligt många personer med kunskaper i första hjälpen, första hjälpen-utrustning samt instruktioner för olycksfall.
Arbetsgivarna ordnar utbildning i första hjälpen på arbetsplatsen.
Om det finns minst tio anställda på en arbetsplats väljer dessa ut en arbetarskyddsfullmäktig som representerar dem.
Arbetarskyddsfullmäktige gör sig insatt i arbetarskyddsfrågor som gäller arbetsplatsen, deltar i arbetsplatsens arbetarskyddsinspektioner och informerar de anställda om ärenden som rör arbetets säkerhet och hälsa.
Arbetsgivaren utser för varje arbetsplats en arbetarskyddschef, som bistår arbetsgivaren i samarbetet med anställda och arbetarskyddsmyndigheter.
Arbetarskyddsmyndigheter
I Finland finns det fem ansvarsområden för arbetarskydd som lyder under Regionförvaltningsverket (RFV).
Ansvarsområdena övervakar att de lagenliga arbetarskyddsföreskrifterna följs på arbetsplatserna.
Ansvarsområdena för arbetarskydd ger både arbetstagare och arbetsgivare råd i frågor som gäller arbetets säkerhet och hälsa samt i frågor som rör anställningsvillkor.
Arbetarskyddsinspektörerna utför kontroller på arbetsplatser.
De kontrollerar bland annat om säkerhetsföreskrifterna följs på arbetsplatsen, om man har gett tillräcklig introduktion i arbetet och huruvida utländska arbetstagares arbetsförhållanden och anställningsvillkor följer finländska lagar och avtal.
Arbetarskyddsinspektören har rätt att få tillträde till varje arbetsplats och tillgång till de dokument som är väsentliga för övervakningen av arbetarskyddet.
Arbetarskyddsmyndigheten kan förplikta arbetsgivaren att rätta till brister i arbetssäkerheten som förekommer på arbetsplatsen
linkkiArbetarskyddsförvaltningen:
Information om arbetarskydd och råd vid problemfinska _ svenska _ engelska
linkkiEuropeiska arbetsmiljöbyrån:
Information om arbetarskyddfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Jämlikheten är nedtecknad i lagar
Finlands grundlag garanterar jämlikt bemötande för alla.
Jämlikhet (yhdenvertaisuus) betyder att alla människor är likvärdiga oberoende av kön, ålder, etnisk eller nationell härkomst, nationalitet, språk, religion och övertygelse, åsikt, handikapp, hälsotillstånd, sexuell läggning eller någon annan orsak som gäller hans eller hennes person.
Om jämlikhet i arbetslivet föreskrivs i lagen om likabehandling och i arbetsavtalslagen.
Enligt dessa ska anställda behandlas lika när det gäller anställning, arbetsförhållanden, anställningsvillkor, utbildning för personalen och avancemang i karriären.
Finlands grundlagfinska _ svenska _ engelska _ ryska _ franska _ spanska _ tyska
Lag om likabehandlingfinska _ svenska _ engelska
Jämlikhet i rekryteringen
Lagen om likabehandling (yhdenvertaisuuslaki) förutsätter att alla arbetssökande behandlas lika.
Arbetsgivaren ska välja den sökande som har de bästa meriterna för uppgiften.
Arbetsgivaren ska också kunna bevisa att det finns godtagbara grunder för valet som anknyter till arbetets karaktär och att valet inte har varit diskriminerande.
Man får inte kräva sådana egenskaper av arbetssökanden som inte är nödvändiga i utförandet av arbetet.
Jämlikhet på arbetsplatsen
Arbetsgivaren får inte diskriminera de anställda när han eller hon fattar beslut om fördelning av arbetsuppgifter, erbjudande av möjligheter till avancemang eller upphävande av anställningen.
Arbetsdiskriminering är ett brott.
Om du misstänker att du har fallit offer för arbetsdiskriminering kan du ta kontakt med arbetarskyddsmyndigheterna eller ditt eget fackförbund.
Vid problem kan du fråga råd hos arbetarskyddsfullmäktige eller förtroendemannen.
linkkiArbetarskyddsförvaltningen:
Arbetarskyddfinska _ svenska _ engelska
linkkiRegionförvaltningsverket:
Arbetarskyddfinska _ svenska _ engelska
linkkiArbets- och näringsministeriet:
Likabehandling och förebyggande av diskriminering på arbetsplatserfinska _ svenska _ engelska
Jämställdhet (tasa-arvo) mellan könen
Enligt Finlands lag är män och kvinnor jämställda.
Män och kvinnor ska behandlas lika vid anställning och beträffande arbetsförhållanden och lönesättning.
En anställd får inte särbehandlas i arbetslivet på grund av graviditet eller föräldraskap.
I Finland finns en lag om likabehandling, som föreskriver att arbetsgivaren ska övervaka att jämställdheten på arbetsplatsen realiseras och att ingen diskrimineras på arbetsplatsen.
Jämställdhetsombudsmannen övervakar att lagen om likabehandling av män och kvinnor följs.
Om du misstänker att din arbetsgivare har diskriminerat dig på grund av ditt kön kan du be jämställdhetsombudsmannen om råd och anvisningar samt hjälp med att reda ut saken.
linkkiJämställdhetsombudsmannens byrå:
Information om jämställdhet i arbetslivetfinska _ svenska _ engelska _ ryska _ samiska
Jämställdhetslagenfinska _ svenska
I Finland har alla möjlighet att få avgiftsfri företagsrådgivning.
Rådgivning tillhandahålls till exempel av:
Företagsfinland (Yritys-Suomi) (webbplats och telefontjänst)
Dessa aktörer handleder alla som är intresserade av företagande i hela Finland.
När du får en bra affärsidé, ta kontakt med det närmaste företagsservicecentret.
Experterna där hjälper dig att utveckla affärsidén. Du får hjälp med att utarbeta preliminära marknadsundersökningar, lönsamhetskalkyler och en kartläggning om tillgången till finansiering.
Du får också råd om utarbetandet av en affärsverksamhetsplan och stöd för ditt beslut att starta ett företag.
Företagsrådgivning kan fås på finska och svenska och åtminstone i större städer också på engelska och andra språk.
Företagsfinland ger företagsrådgivning telefonledes på finska och svenska.
Företagsfinlands telefonrådgivningsnummer är:
på finska 0295 020 500
på svenska 0295 020 501
Om du vill ha rådgivning på engelska, ska du skicka in din fråga via Företagsfinlands engelskspråkiga webbplats.
Telefontjänsten har öppet måndag till fredag kl. 9.00–16.15.
linkkiFöretagsFinland:
Företagsrådgivningfinska _ svenska _ engelska
Företagarkurser
Olika instanser anordnar företagarkurser och informationsmöten som man har mycket nytta av om man vill starta ett företag.
Ämnen som behandlas på kurserna är till exempel utarbetande av en affärsverksamhetsplan, startande av företagsverksamhet, bokföring, företagsbeskattning, juridiska frågor, marknadsföring, försäljning och kundtjänst.
Guide om att grunda ett företagfinska _ engelska _ kinesiska
linkkiFöretagsfinland:
Att grunda ett företagfinska _ svenska _ engelska
linkkiArbets- och näringsministeriet:
Tjänster för företagarefinska _ svenska _ engelska
linkkiEuropeiska unionen:
Information om att arbeta och driva ett företag i den europeiska unionenfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
Kurssökningfinska _ svenska _ engelska
Allmänt om fackförbund
I Finland tryggar lagen arbetstagarnas rätt att höra till ett fackförbund (ammattiliitto).
Denna rätt kan inte begränsas med avtal.
Diskriminering av arbetstagare på grund av deras medlemskap i fackförbund är straffbart.
De flesta finländare är med i något fackförbund.
Fackförbunden strävar efter att trygga sina medlemmars intressen och rättigheter, försöker förbättra lönerna och anställningsskyddet samt förbättra arbetslivets kvalitet.
Arbetstagarförbunden är organiserade under tre centralförbund för löntagare.
Dessa är Finlands Fackförbunds Centralorganisation FFC, Tjänstemannacentralorganisationen STTK och Centralorganisationen för högutbildade i Finland Akava.
linkkiFCC, STTK och AKAVA:
Fackets ABC-bokfinska _ engelska _ ryska _ estniska
linkkiCentralorganisationen för högutbildade i Finland Akava:
Information om fackförbundsverksamhetfinska _ svenska _ engelska _ ryska _ estniska _ franska
Information om fackförbundsverksamhetfinska _ svenska _ engelska
linkkiTjänstemannacentralorganisationen STTK:
Information om fackförbundsverksamhetfinska _ svenska _ engelska
Att ansluta sig till ett fackförbund och medlemsavgiften
Om du vill kan du ansluta dig till fackförbundet i din egen bransch.
Du kan ansluta dig till ett fackförbund genom att ta kontakt med förtroendemannen på din egen arbetsplats eller genom att kontakta fackförbundet direkt.
Till de flesta fackförbund kan man också ansluta sig genom att fylla i en anslutningsblankett på fackets webbplats.
Fackförbundets medlemmar betalar förbundet en medlemsavgift som vanligen är cirka 1–2 procent av lönen.
Medlemsavgiften får dras av i beskattningen.
Fackförbundets medlemmar kan delta i utbildning och fritidsaktiviteter som förbundet ordnar.
De får också stöd av förbundets förtroendeman vid konflikter på arbetsplatsen.
Vid behov får man också råd eller förhandlingsstöd från fackförbundet.
Arbetslöshetskassa
I Finland finns ett frivilligt system med arbetslöshetskassor.
En arbetstagare som är medlem i en arbetslöshetskassa betalar en medlemsavgift till arbetslöshetskassan när han eller hon förvärvsarbetar.
Om arbetet upphör och arbetstagaren blir arbetslös kan han eller hon ansöka om inkomstrelaterad arbetslöshetsdagpenning från kassan.
Det lönar sig att ansluta sig till en arbetslöshetskassa, eftersom den inkomstrelaterade dagpenningen är större än det vanliga utkomstskyddet för arbetslösa.
När du ansluter dig till ett fackförbund kan du samtidigt ansluta dig till förbundets arbetslöshetskassa.
Fackförbundet och arbetslöshetskassan är dock två separata system.
Det finns också arbetslöshetskassor som man kan ansluta sig till utan att vara medlem i något fackförbund.
För att få inkomstrelaterad dagpenning finns några villkor som måste uppfyllas innan det är möjligt att få dagpenning.
Till exempel ska man ha varit med i arbetslöshetskassan en viss tid före man blir arbetslös.
Ta reda på dessa villkor genast när du ansluter dig till arbetslöshetskassan.
Läs mer på InfoFinlands sida Utkomstskydd för arbetslösa.
linkkiArbetslöshetskassornas samorganisation:
information om arbetslöshetskassorfinska _ svenska _ engelska
Fackförbundets representant på arbetsplatsen
På arbetsplatsen representeras fackförbundet och de anställda som är medlemmar i det av förtroendemannen.
Förtroendemannen väljs av de anställda.
Förtroendemannen agerar som förhandlare, medlare och informationsförmedlare mellan arbetsgivaren och anställda.
Man kan också vända sig till förtroendemannen till exempel med frågor om kollektivavtalet.
I Finland har en arbetstagare rätt:
till lön och övriga minimivillkor enligt kollektivavtalet
till skydd utgående från lagar och avtal
att organisera sig
till en sund och trygg arbetsmiljö.
En arbetstagare är skyldig att
utföra arbetet omsorgsfullt
följa de överenskomna arbetstiderna
följa arbetsledningens anvisningar
vägra att delta i verksamhet som konkurrerar med arbetsgivaren
hålla affärs- och yrkeshemligheter
ta hänsyn till arbetsgivarens intresse.
Anställningsrådgivning för invandrare
Om du har frågor om eller problem med din anställning, kan du kontakta anställningsrådgivningen för invandrare.
Rådgivningen ges av Finlands Fackförbunds Centralorganisation FFC.
Du kan få rådgivning även om du inte är medlem i fackförbundet.
En jurist svarar på dina frågor till exempel om arbetsavtal, lön eller arbetstider.
Den kostnadsfria rådgivningen ges på finska och engelska.
Anställningsrådgivningen har öppet på tisdagar och onsdagar klockan 9–11 och 12–15.
Telefon: 0800 414 004
Du kan även ringa arbetarskyddsmyndigheternas riksomfattande rådgivningstelefon:
Tfn 0295 016 620
Mån.–fre. kl. 9–15
linkkiFFC:
Anställningsrådgivning för invandrarefinska _ svenska _ engelska
linkkiFFC:
Arbetslivet i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ kinesiska _ arabiska
linkkiArbetshälsoinstitutet:
Handboken Jobba i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ kurdiska _ tyska _ thai _ vietnamesiska
linkkiBrottsofferjouren:
Video om arbetstagarens rättigheter i Finlandengelska _ kinesiska _ arabiska _ thai _ hindi
Arbetstagarnas rättigheter tryggas med lagar och avtal
Arbetslagstiftningen och kollektivavtalen föreskriver vilka rättigheter och skyldigheter arbetstagare har.
Arbetstagar- och arbetsgivarförbunden förhandlar gemensamt fram branschspecifika kollektivavtal.
I lagstiftningen och kollektivavtalet fastställs till exempel minimilöner, arbetstider, semestrar, lön för sjukdomstid och uppsägningsvillkor.
Läs mer på InfoFinlands sidor Att komma överens om anställningsvillkoren och Innehållet i arbetsavtalet.
linkkiArbets- och näringsministeriet:
Broschyrer om arbetslagstiftningenfinska _ svenska _ engelska
Jämlikhet
Varje anställd har rätt till ett jämlikt och icke-diskriminerande bemötande när de söker jobb och på arbetsplatsen.
Läs mer på InfoFinlands sida Jämlikhet och jämställdhet i arbetslivet.
Arbetsavtal
Ett arbetsavtal uppstår när arbetstagaren och arbetsgivaren kommer överens om utförandet av ett arbete och lönen som betalas för det samt övriga förmåner och villkor.
Anställningsvillkoren bestäms enligt arbetslagstiftningen och kollektivavtalet.
Arbetsavtalet är bindande för båda parterna.
Läs mer om arbetsavtalet på InfoFinlands sidor Att komma överens om anställningsvillkoren och Innehållet i arbetsavtalet.
Fackförbund
I Finland är facklig organisering vanligt och aktiva fackförbundsmedlemmar trakasseras inte.
Du kan ansluta dig till fackförbundet i din egen bransch.
Förbundet strävar efter att trygga sina medlemmars intressen i arbetslivet.
Läs mer på InfoFinlands sida Fackförbund.
Arbetarskydd
Arbetsgivaren är skyldig att trygga de anställdas säkerhet.
Arbetarskyddsförvaltningen övervakar att de i lagen stadgade arbetarskyddsföreskrifterna följs på arbetsplatserna.
Läs mer på InfoFinlands sida Arbetarskydd.
Utkomstskydd för arbetslösa
När en person som är fast bosatt i Finland blir arbetslös, har han eller hon rätt att få utkomstskydd för arbetslösa.
Läs mer på InfoFinlands sida Utkomstskydd för arbetslösa.
En invandrare som har bott tillräckligt länge i Finland kan få pension på grund av sin ålder eller arbetsoförmögenhet.
Läs mer på InfoFinlands sida Pension.
Beskattning
När du arbetar i Finland måste du betala skatter.
Läs mer på InfoFinlands sida Beskattning.
Företagshälsovård
Varje arbetsgivare är skyldig att ordna förebyggande företagshälsovård för sina anställda.
Läs mer på InfoFinlands sida Företagshälsovård.
Familjeledigheter
När ett barn föds till familjen kan modern eller fadern enligt lag stanna hemma för att ta hand om barnet.
Läs mer på InfoFinlands sida Familjeledigheter.
Arbetsintyg
När en anställning upphör har den anställda rätt att få ett skriftligt arbetsintyg av arbetsgivaren.
Läs mer på InfoFinlands sida Arbetsintyg.
Hur grundar jag ett företag?
Du hittar grundläggande information om att starta ett företag i Finland på dessa sidor i InfoFinland.
De centrala stegen när man startar ett företag:
Kom på en bra affärsidé
Gör en affärsverksamhetsplan
Ordna finansiering
Välj företagsform
Ta reda på vilka tillstånd du behöver
Gör anmälan till handelsregistret och skattemyndigheten
Teckna försäkringar
Ordna bokföringen
Förbered dig på företagande
Företagande kräver yrkeskunnighet och utbildning. Det är viktigt att du är väl insatt i din bransch och lagarna som gäller företagande.
Också kännedom om de egna kunderna och försäljningsmetoderna är viktig.
Tillräcklig finansiering och noggrann planering är oumbärliga.
Förbered dig på företagande genom att skaffa så goda kunskaper och färdigheter som möjligt, eftersom det är riskabelt att starta ett företag utan tillräckligt kunnande och tillräckliga språkkunskaper.
När du vill starta ett företag ska du fundera noga på om du har en bra affärsidé.
Fundera också om du har tillräcklig yrkeskunnighet och erfarenhet och planera hur du ska ordna finansiering.
Du kan be om hjälp i frågor som rör startandet av ett företag hos nyföretagarcentralerna.
Läs mer på InfoFinlands sida Företagsrådgivning.
Kom även ihåg att en underskrift är ett bindande avtal. Läs noga igenom alla dokument innan du undertecknar något.
Guide om att grunda ett företagfinska _ engelska _ kinesiska
Som företagare till Finland:
Vilka tillstånd behöver du?(pdf, 384 kt)finska _ engelska
linkkiFöretagsfinland:
Att grunda ett företagfinska _ svenska _ engelska
ABC för restaurangbranschen:
Anvisningar för dig som ska grunda ett café eller en restaurang finska _ engelska
Arbetsavtalet upprättas i två exemplar, ett till den anställda och ett till arbetsgivaren.
Arbetsavtalet innehåller vanligen åtminstone följande punkter:
Parterna som ingår arbetsavtalet
Både arbetsgivaren och den anställda undertecknar arbetsavtalet.
Tidpunkten då arbetet inletts
Om avtalet är tillsvidare gällande eller tidsbundet
Huvudregeln är att arbetsavtalet gäller tillsvidare.
Detta innebär att arbetet pågår tills den anställda säger upp sig eller tills arbetsgivaren säger upp den anställda.
Arbetsgivaren ska ha en välgrundad orsak för att säga upp en anställd.
Godtagbara orsaker för uppsägning definieras i arbetsavtalslagen.
När arbetsavtalet gäller tillsvidare har arbetstagaren en fast eller permanent anställning.
Ett tidsbundet avtal innebär att man har avtalat om tidpunkten då arbetet inleds och avslutas.
Arbetsavtalet kan vara tidsbundet om det finns en välgrundad orsak till detta.
Lagar och kollektivavtal reglerar exakt när tidsbundna anställningar får tillämpas.
En anställning kan vara tidsbunden om orsaken är till exempel
vikariat
praktik
projekt
efterfrågan eller säsongtopp
Om arbetsavtalet är tidsbundet binder det båda parterna en bestämd tid, om man inte har kommit överens om möjligheten till uppsägning.
Ett tidsbundet avtal kan hävas endast av mycket vägande skäl.
Prövotid och längden på den
Man kan komma överens om en prövotid i anställningens början.
Prövotiden kan vara högst sex månader.
Vid en tidsbunden anställning kan prövotiden vara högst hälften av den tid anställningen pågår.
Under prövotiden kan arbetstagaren bedöma om arbetet lämpar sig för honom eller henne och arbetsgivaren kan bedöma om arbetstagaren är lämplig för arbetet.
Under prövotiden kan arbetstagaren och arbetsgivaren häva arbetsavtalet utan uppsägningstid.
Grunderna för hävande av ett arbetsavtal under prövotiden får inte vara diskriminerande.
Arbetstagaren får normal lön under prövotiden.
Platsen för utförandet av arbetet
Arbetsuppgifterna
Lönen och utbetalning av lönen
Lönen bestäms enligt kollektivavtalet.
Om branschen inte har ett kollektivavtal har arbetstagaren rätt till en skälig lön.
Arbetsgivaren får inte betala en lön som är mindre än vad som fastställs i kollektivavtalet.
Lönen kan innehålla olika förmåner.
Typiska lönetillägg i Finland är erfarenhetstillägg, övertidstillägg och skiftarbetstillägg.
Avlöningsdagen är vanligen en eller två gånger i månaden.
Arbetsgivaren betalar in lönen på bankkontot.
Arbetstagaren har rätt att få en lönespecifikation där det står vad lönen består av.
När man talar om lön avser man oftast bruttolönen (bruttopalkka) från vilken skatter och personalbikostnader dras av.
Den lön som betalas till arbetstagaren är nettolönen (nettopalkka).
Arbetstid
I avtalet ska den regelbundna arbetstiden nedtecknas.
Arbetstiden ska följa arbetslagstiftningen och kollektivavtalet.
Semester och semesterpenning
Arbetstagaren har rätt att få samma lön under semestern som under arbetet.
Dessutom betalas en semesterpenning.
Utbetalningen av semesterpenning baserar sig på kollektivavtalet.
När anställningen upphör har arbetstagaren rätt att få semesterersättning för de dagar som han eller hon inte har fått semester eller semesterersättning för vid tidpunkten för anställningens upphörande.
Uppsägningstid
Ett tillsvidare gällande arbetsavtal upphör antingen när arbetstagarens eller arbetsgivarens uppsägningstid har gått ut.
Uppsägningstiden är den tid som arbetstagaren är skyldig att arbeta innan arbetet upphör.
Under uppsägningstiden har arbetstagaren samma rättigheter och skyldigheter och han eller hon får normal lön.
Om arbetsgivaren säger upp en arbetstagare måste arbetsgivaren ange orsaken till detta.
Arbetsavtalslagen beskriver vilka orsaker som är godtagbara för uppsägning.
Omnämnande om viket kollektivavtal arbetsavtalet följer
linkkiArbets- och näringsministeriet:
Arbetsavtal och anställningfinska _ svenska _ engelska
Om du har avlagt examen i något annat land kan du behöva beslut om erkännande av examen för att kunna arbeta eller studera i Finland.
I de flesta situationerna bedömer arbetsgivaren, läroanstalten eller högskolan vilken behörighet och kompetens din utländska examen ger.
Du behöver Utbildningsstyrelsens eller någon annan myndighets beslut om erkännande av examen om du vill arbeta inom ett reglerat yrke eller en uppgift som kräver högskoleexamen på viss nivå.
linkkiUtbildningsstyrelsen:
Erkännande av en examenfinska _ svenska _ engelska
linkkiUtbildningsstyrelsen :
Broschyr om erkännande av examen(pdf, 102,14 kt)finska _ svenska _ engelska _ ryska _ estniska _ franska _ spanska _ kinesiska _ persiska _ arabiska _ portugisiska
linkkiUtbildningsstyrelsen :
Diagram över erkännande av examen(pdf, 410,87 kt)finska _ svenska _ engelska
linkkiUtbildningsstyrelsen:
Servicepriserfinska _ svenska _ engelska
Om du vill fortsätta dina studier i Finland
Högskolor och läroanstalter beslutar om antagning av studerande.
De beslutar också huruvida dina utländska studier och din övriga kompetens kan godkännas som en del av den examen du avlägger i Finland.
Om du har avlagt högskolestudier utomlands och vill fortsätta dina studier i Finland kan du få information och handledning vid högskolornas tjänster för studerande och SIMHE-tjänsterna.
Högskolor som erbjuder SIMHE-tjänsterfinska _ svenska _ engelska
Uppgifter som inte kräver en viss utbildning
Enligt Finlands lag kräver inte alla uppgifter en viss utbildning eller examen på en viss nivå.
Till exempel bedömer arbetsgivare i privatsektorn oftast själv huruvida en utländsk examen ger tillräckliga kvalifikationer för uppgiften.
Jämställande av nivån på en högskolexamen
För uppgifter inom den offentliga sektorn (kommun eller stat) krävs ofta examen på en viss nivå, till exempel en högre högskoleexamen.
Om du har avlagt en högskoleexamen utomlands kan du ansöka om beslut om jämställande av nivån på en högskolexamen vid Utbildningsstyrelsen.
Beslutet är avgiftsbelagt.
När din examensnivå har jämställts med en finländsk högskoleexamen, kan du söka till uppgifter som kräver den nivå på högskoleexamen som du har.
linkkiUtbildningsstyrelsen:
Jämställande av nivån på en högskolexamenfinska _ svenska _ engelska
Reglerade yrken
I Finland är vissa yrken reglerade.
Det betyder att det stadgas i lag vilken utbildning som krävs för dessa yrken.
Sådana uppgifter är till exempel fysioterapeut, läkare, tandläkare, provisor, sjukskötare, advokat, revisor, klasslärare och sotare.
Branschspecifika myndigheter beslutar om rätten att utöva ett reglerat yrke eller använda en yrkesbeteckning.
Till exempel inom social- och hälsovårdsbranschen fattas beslutet av Valvira, och inom undervisningssektorn av Utbildningsstyrelsen.
Beslutet är avgiftsbelagt.
På Utbildningsstyrelsens webbplats hittar du en förteckning över reglerade yrken och de myndigheter som fattar beslut.
linkkiUtbildningsstyrelsen:
Reglerade yrken och ansvariga myndigheterfinska _ svenska _ engelska
Information om erkännande av examen för yrken inom hälsovårdenfinska _ svenska _ engelska
Reglerade yrken och examen från ett annat EU-land
Om
du är medborgare i ett EU-land, EES-land eller Schweiz och du har
förvärvat kvalifikationer för ett yrke som är reglerat i Finland i ett EU-land, EES-land eller Schweiz,
kan du ansöka om erkännande av yrkeskvalifikationer för detta yrke hos den branschspecifika myndigheten.
Om din utbildning skiljer sig mycket från den utbildning som krävs i Finland måste du eventuellt avlägga en anpassningsperiod eller ett lämplighetsprov.
linkkiUtbildningsstyrelsen:
Erkännande av yrkeskvalifikationer som förvärvats i ett EU-landfinska _ svenska _ engelska
linkkiEuropeiska kommissionen:
Information om reglerade yrken i EU-ländernaengelska
Utländsk yrkesexamen
Om du har avlagt en yrkesexamen utomlands kan du ansöka om ett utlåtande om det hos Utbildningsstyrelsen.
I utlåtandet beskrivs examensnivån och innehåll samt för vilka uppgifter examen ger kvalifikationer i det land där du har avlagt examen.
Utlåtandet ger dig dock inte kvalifikationer att utöva ett reglerat yrke i Finland.
linkkiUtbildningsstyrelsen:
Utlåtanden om utländska yrkesexamenfinska _ svenska _ engelska
Översättning av handlingar
Om originalspråket för ditt betyg inte är finska, svenska eller engelska behöver du vanligtvis en officiell översättning av handlingarna som görs av en auktoriserad översättare.
Vissa myndigheter godkänner även handlingar på andra europeiska språk.
Läs noga anvisningarna om ansökning från den branschspecifika myndigheten.
Var får jag hjälp med problem i arbetslivet?
Prata först med din chef.
Om det inte hjälper, kontakta arbetsplatsens förtroendeman.
Om det inte finns en förtroendeman på arbetsplatsen och du är medlem i facket, kontakta ditt fackförbund.
Finlands Fackförbunds Centralorganisation FFC erbjuder gratis anställningsrådgivning.
Du kan få rådgivning även om du inte är medlem i ett fackförbund.
Juristerna svarar på dina frågor på finska och engelska.
Rådgivning ges både per telefon och via e-post:
Tfn 0800 414 004, tis. och ons. kl. 9–11 och 12–15
Du kan även ringa arbetarskyddsmyndigheternas riksomfattande rådgivningstelefon:
Tfn 0295 016 620
Mån.–fre. kl. 9–15
linkkiArbetarskyddsförvaltning:
Kontaktuppgifter till arbetarskyddsmyndigheternafinska _ svenska _ engelska
Min anställning upphör inom kort.
Hur påverkar det mitt uppehållstillstånd?
Detta beror på vilket slags uppehållstillstånd du har.
Om ditt uppehållstillstånd är kopplat till endast en arbetsgivare, ska du ansöka om ett nytt uppehållstillstånd för arbetstagare.
För att kunna ansöka om ett nytt uppehållstillstånd för arbetstagare måste du ha ett nytt jobb.
Du kan även ansöka om uppehållstillstånd på någon annan grund.
Läs mer om grunderna för uppehållstillstånd i InfoFinlands avsnitt Icke EU-medborgare.
Om din anställning upphör innan ditt uppehållstillstånd går ut, ska du meddela detta skriftligt till Migrationsverket.
Också din arbetsgivare kan göra anmälan.
Om ditt uppehållstillstånd är beviljat för en viss bransch, kan du byta jobb inom samma bransch.
Information om uppehållstillstånd för arbetstagare och företagare hittar du på sidorna Arbeta i Finland och Till Finland som företagare.
Läs mer om att söka jobb i Finland på sidan Var hittar jag jobb?
Mer information om att söka arbetslöshetsersättning hittar du på sidan Arbetslöshetsförsäkring.
Information om uppehållstillståndfinska _ svenska _ engelska
Jag har fått för lite lön utbetalad.
Vad ska jag göra?
Kontrollera alltid i lönespecifikationen att du har fått rätt belopp.
Om du har fått för lite lön, ska du be din arbetsgivare att rätta till löneutbetalningen.
Om arbetsgivaren inte betalar ut rätt lön, ska du fråga om råd hos regionförvaltningsverkets arbetarskydd eller ditt fackförbund.
Om du inte kan komma överens om löneutbetalningen med din arbetsgivare måste ärendet avgöras i domstol.
Detta är dock det sista alternativet.
linkkiArbetarskyddsförvaltning:
Information om löneutbetalningfinska _ svenska _ engelska
Min arbetsgivare vill endast betala ut lönen i kontanter.
Får man göra så?
Din arbetsgivare borde betala ut lönen till ditt bankkonto.
Lönen får endast betalas ut i kontanter om inga andra alternativ finns.
Så gör man till exempel om du inte har ett bankkonto.
Om du får lönen utbetalad i kontanter, ska du ge din arbetsgivare ett skriftligt intyg om löneutbetalningen.
På så sätt kan man bevisa att lönen verkligen har betalats till dig.
Min tillsvidareanställning upphörde, men min sista lön betalades inte ut.
Vad bör jag göra?
Fråga arbetsgivaren varför lönen blivit försenad.
Kräv att arbetsgivaren betalar ut lönen.
Framför kravet skriftligt.
Om du är medlem i ett fackförbund kan du be förbundet om hjälp.
Om du inte är medlem i ett fackförbund, kontakta till exempel arbetarskyddsmyndigheterna.
Jag avslutade mitt jobb hos min förra arbetsgivare, men jag har inte fått ett arbetsintyg.
Hur får jag arbetsintyget?
Arbetsgivare behöver inte ge dig ett arbetsintyg på eget bevåg.
Om du vill ha ett arbetsintyg ska du be om det.
Intyget ska lämnas till dig så snart som möjligt.
Om du har bett om ett arbetsintyg men inte fått det, ska du kontakta arbetarskyddsmyndigheterna.
Läs mer på InfoFinlands sida Arbetsintyg.
Jag upplever att jag blir osakligt bemött på min arbetsplats.
Vad kan jag göra?
Alla arbetstagare ska behandlas jämlikt och lika.
Enligt lag får ingen diskrimineras till exempel av följande orsaker:
anställningsform
ålder
kön
etnisk bakgrund
hälsotillstånd
religion
sexuell läggning.
Läs mer på InfoFinlands sida Diskriminering och rasism.
Förutom diskriminering kan det även förekomma andra typer av osakligt bemötande på arbetsplatser, till exempel mobbning eller sexuella trakasserier.
Om hen inte kan hjälpa dig, ska du kontakta arbetsplatsens arbetarskyddsfullmäktige eller förtroendeman.
Om ärendet inte kan lösas på arbetsplatsen, kontakta arbetarskyddsmyndigheterna eller ditt fackförbund.
Om din chef behandlar dig osakligt, anmäl detta till arbetarskyddsmyndigheterna.
Du kan göra anmälan med ditt eget namn eller anonymt.
Jag tvingas att utföra ett jobb utan att få betalt.
Min arbetsgivare hotar mig dessutom med våld.
Var kan jag få hjälp?
Du har rätt till hjälp och skydd.
Enligt lagen i Finland måste arbetstagarna behandlas väl och de ska betalas lön.
Människohandel är ett brott i Finland.
Läs mer på InfoFinlands sida Människohandel och tvångsarbete.
Du hittar information om arbetstagarens rättigheter och skyldigheter i Finland på InfoFinlands sida Arbetstagarens rättigheter och skyldigheter.
Hjälp till offer för människohandelfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska _ polska _ rumänska _ bulgariska
I Finland bestäms arbetstagarnas rättigheter enligt arbetslagstiftningen och kollektivavtalen (työehtosopimukset).
I dessa fastställs till exempel minimilöner, arbetstider, semestrar, lön för sjukdomstid och uppsägningsvillkor.
Arbetsgivarförbundet och arbetstagarförbundet kommer gemensamt överens om anställningsvillkoren i en viss bransch.
På detta sätt uppstår ett kollektivavtal för branschen.
I den offentliga sektorn (arbetsgivaren är en kommun eller staten) ingås tjänstekollektivavtal eller allmänt kommunalt tjänste- och arbetskollektivavtal.
Förmånerna som man har avtalat om med ett kollektivavtal är alltid minimiförmåner.
Dessa kan inte underskridas i arbetsavtalet.
Lönen kan till exempel inte vara lägre än vad som avtalats med kollektivavtalet.
Arbetsgivaren och arbetstagaren kan ändå i arbetsavtalet komma överens om villkor som är bättre än villkoren i kollektivavtalet.
Kollektivavtalen uppgörs för en viss tid, vanligen för ett eller två år eller också för en längre tid.
Kollektiv- och tjänstekollektivavtalet är bindande för de löntagar- och arbetsgivarförbund som slutit dem och för deras medlemmar.
Ett kollektivavtal kan också vara allmänt bindande.
Då måste även de arbetsgivare som inte hör till arbetsgivarförbundet följa avtalet med sina anställda.
I platsannonser och arbetsavtal kan det stå: ”palkkaus TES:in mukainen” (”avlöning enligt kollektivavtalet”).
Det är bra att ta reda på hur stora lönerna är i den egna branschen i Finland.
Det är viktigt att känna till kollektivavtalet, eftersom det i Finland inte finns till exempel en lag om minimilöner, utan minimilönerna fastställs alltid enligt kollektivavtalet.
linkkiArbets- och näringsministeriet:
Arbetslagstiftningfinska _ svenska _ engelska
Arbetsavtal
Arbetsgivaren ingår vanligen ett skriftligt arbetsavtal med en ny anställd.
I arbetsavtalet fastställs arbetsuppgifterna och lönen samt andra förmåner och villkor.
Avtalet kan också vara muntligt.
Om man inte har uppgjort ett skriftligt arbetsavtal ska arbetsgivaren utan särskild begäran ge en skriftlig redogörelse för de centrala villkoren i arbetet.
Det är rekommendabelt att arbetsavtalet är skriftligt.
När allt finns på papper kan både den anställda och arbetsgivaren kontrollera i avtalet vad man gemensamt har avtalat.
Detta hjälper om det uppstår konflikter i arbetet.
Läs mer om upprättandet av arbetsavtalet på InfoFinlands sida Innehållet i arbetsavtalet.
linkkiArbetarskyddsförvaltningen:
Att uppgöra ett arbetsavtalfinska _ svenska _ engelska
Ett skriftligt avtal om de centrala villkoren i arbetet
Arbetsgivaren ska ge den anställda en skriftlig redogörelse för de centrala villkoren i arbetet vid tillsvidare gällande anställningar samt anställningar som varar över en månad.
Av redogörelsen ska det åtminstone framgå
arbetsgivarens och arbetstagarens hemort eller driftställe
tidpunkten då arbetet inletts
längden på ett tidsbundet arbetsavtal och orsaken till att avtalet är tidsbundet
prövotidens längd
stället där arbetet utförs
den anställdas arbetsuppgifter
kollektivavtalet som tillämpas på arbetet
de grunder enligt vilka lön eller andra vederlag bestäms samt löneperioden
den regelbundna arbetstiden
hur semestern bestäms
uppsägningstiden eller grunden för bestämmande av den
Om arbetsgivaren inte ger en redogörelse för de centrala villkoren i arbetet till den anställda kan han eller hon dömas till böter.
Läs jobbannonsen noga
Innan du skriver din jobbansökan, läs jobbannonsen noga och fundera på vilka färdigheter och vilket kunnande arbetsgivaren är ute efter.
Fundera på hur ditt kunnande motsvarar arbetsgivarens önskemål och krav.
Du kan också kontakta arbetsgivaren och begära mer information, om du undrar över något som inte framgår av jobbannonsen.
Ring arbetsgivaren bara om du har en konkret fråga om arbetsplatsen.
Jobbansökan
Vanligtvis när du söker ett jobb, skickar du en jobbansökan och ditt CV, alltså din meritförteckning, till arbetsgivaren.
Ibland kan jobbansökningen vara en video, en portfölj eller till exempel en webbsida.
Skriv ansökan och CV på samma språk som används i annonsen.
Skriv en ny ansökan och uppdatera ditt CV varje gång när du ansöker om ett nytt jobb.
Du kan skriva ansökningstexten direkt i e-postmeddelandet eller bifoga den till e-postmeddelandet tillsammans med ditt CV.
Lägg till bilagorna alltid i PDF-format.
Ofta kan du skicka in ansökan och CV via arbetsgivarens webbplats.
Syftet med din jobbansökan är att väcka arbetsgivarens intresse så att du blir kallad till anställningsintervju.
Ansökningen är ett svar på jobbannonsen.
Du ska svara på de önskemål och krav som nämns i jobbannonsen.
Lyft fram sådant som är viktigt i arbetsuppgiften.
Ge konkreta exempel på ditt kunnande.
Intyga arbetsgivaren om att du är lämplig för uppgiften.
En jobbansökan är oftast en knapp sida.
Be någon att läsa igenom och granska din ansökan.
Löneanspråk
Ofta ska man ange sitt löneanspråk i ansökningen.
Det är ofta svårt att uppskatta rätt belopp.
Löneanspråket får inte vara för stort, men inte heller för litet.
Från fackförbund får du mer information om lönenivån i olika branscher.
Lönejämförelse finska _ engelska
Gå igenom dina utbildningar och din arbetserfarenhet och fundera på vilka färdigheter du lärt dig i dem.
Vilka är dina styrkor?
Fundera också på vilket kunnande du har fått från dina fritidsintressen eller andra erfarenheter.
Tidsenliga intyg
Spara intygen från dina tidigare jobb och studier.
Kom ihåg att alltid begära ett intyg när du haft ett jobb, avlagt en praktik eller studerat.
Arbetsgivaren har skyldighet att utfärda ett intyg ännu tio år efter att anställningen upphört.
Du behöver vanligtvis inte skicka in dina arbetsintyg i förväg till arbetsgivaren, men det är bra att ta med dem till anställningsintervjun för det fall att arbetsgivaren vill se dem.
Det skulle vara bra att ha översättningar till finska eller svenska av alla intyg som du fått utomlands.
Mer information om detta finns på InfoFinlands sida Arbetsintyg.
Erkännande av examen
Det är lättare att söka jobb om du vet hur en examen som du avlagt utomlands motsvarar en finländsk examen.
Du kan ansöka om erkännande av utländsk examen vid Utbildningsstyrelsen.
Erkännande av examen är avgiftsbelagt.
Mer information om detta finns på InfoFinlands sida Utländsk examen i Finland.
linkkiUtbildningsstyrelsen:
Erkännande av en examenfinska _ svenska _ engelska
Öppen ansökan
Du kan ta direkt kontakt med en arbetsplats som du är intresserad av.
Du kan skicka in en öppen ansökan eller ringa arbetsgivaren, trots att de inte har några lediga jobb just nu.
I den öppna ansökan ska du berätta vad du kan och hurdana uppgifter du skulle kunna utföra.
Bifoga din meritförteckning, alltså CV, till ansökan.
Meritförteckning eller CV
En meritförteckning, eller ett CV, är en kortfattad och tydlig sammanfattning av ditt kunnande, din arbetserfarenhet och din utbildning.
Det finns olika CV-mallar.
I ett kompetensbaserat CV kan du gruppera dina färdigheter i olika kompetensområden.
CV:t kan även vara en video, en portfölj eller en webbsida.
Bekanta dig med olika CV-mallar och forma ditt eget CV såsom det passar dig.
Ett CV är vanligtvis 1–2 sidor långt.
Kom ihåg att uppdatera ditt CV för varje ny ansökan.
Vad innehåller ett CV?
Namn och kontaktuppgifter – Adress, e-postadress, telefonnummer
Arbetserfarenhet – Lista dina tidigare anställningar, den senaste först.
Ange också anställningens längd.
Beskriv dina arbetsuppgifter och de färdigheter som du lärt dig i arbetet.
Utbildning – Lista dina examina i kronologisk ordning, den senaste först.
Lägg till namnet på examen, utbildningsprogrammet och läroanstalten och när du tog examen.
Kurser – Lista kurserna i finska och andra kurser som du avlagt under en egen rubrik.
Övrigt kunnande – Språkkunskaper, IT-kunskaper, avlagda tillståndskort, till exempel hygienpass.
Publikationer eller andra arbetsprov
– Om du vill kan du även lista dina publikationer eller arbetsprov.
Fritidsintressen, förtroendeuppdrag
– Du kan även lyfta fram dina intressen.
Referenser – Du kan lägga till namnen på personer som har lovat att rekommendera dig för arbetsuppgiften.
Lägg till kontaktuppgifterna till dem.
Kom ihåg att be personen om tillstånd för detta.
I början av CV:t kan du tillfoga en sammanfattning eller profil där du beskriver din bakgrund och din kärnkompetens med några ord.
Du kan berätta vilka målsättningar du har med jobbsökningen eller vilken specialkompetens du besitter.
Du kan också lägga till ett fotografi.
linkkiArbets- och näringsministeriet:
Så här skriver du en jobbansökan och ett CVfinska _ svenska _ engelska
Kompetensbaserat CV
Ett kompetensbaserat CV lyfter fram ditt kunnande, dina färdigheter och dina erfarenheter.
Välj några kompetensområden och beskriv under rubrikerna dina erfarenheter, färdigheter och prestationer inom dem.
Du kan också lägga till sådant kunnande som du har införskaffat till exempel i frivilligarbete, fritidsintressen eller studier.
Dessutom kan du lista din arbetserfarenhet och utbildning i kronologisk ordning.
I början av CV:t kan du tillfoga en sammanfattning eller profil där du beskriver din bakgrund och din kärnkompetens med några ord.
Du kan berätta vilka målsättningar du har med jobbsökningen eller vilken specialkompetens du besitter.
Skriv ett eget CV för varje arbetsplats.
Lyft fram sådana färdigheter som behövs i uppgiften.
Fundera på vad arbetsgivaren bör veta om dina färdigheter och ditt kunnande.
Europass-CV
Europass är ett allmäneuropeiskt CV, alltså en allmäneuropeisk meritförteckning.
Det består av fem dokument som har till syfte att hjälpa arbetstagare och studerande att presentera sitt kunnande i Europa.
Dokumenten används i alla EU/EES-länderna.
Du kan använda Europass när du söker jobb eller studieplats.
Europass är särskilt nyttigt om du ansöker om ett jobb eller en utbildningsplats i Finland från ett annat EU-land.
linkkiEuropass.eu:
Information om CVfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Förbered dig på anställningsintervjun
Bekanta dig med arbetsgivaren i förväg till exempel med hjälp av webbplatsen.
Fundera på hur du ska lyfta fram ditt kunnande och din lämplighet för uppgiften.
Öva på att beskriva din bakgrund och din yrkeskunnighet med några meningar.
Fundera i förväg på vilka frågor arbetsgivaren kan ställa till dig.
Öva på att besvara allmänna frågor som ingår i en anställningsintervju.
Arbetsgivaren får inte fråga om din familj, vilken religion du har eller om du är politiskt aktiv.
Visa att du har bekantat dig med arbetsgivarens organisation och arbetsuppgiften i förväg och att du har ett äkta intresse för jobbet.
Fundera också på vilka frågor du vill ställa till arbetsgivaren.
linkkiArbets- och näringsministeriet:
Anvisningar för jobbintervjunfinska _ svenska _ engelska
Att börja på ett nytt jobb
Skriv alltid ett skriftligt anställningsavtal innan du börjar på ett nytt jobb.
Kom överens om anställningsavtalets innehåll med arbetsgivaren.
Läs avtalet noga innan du undertecknar det.
Läs mer på InfoFinlands sida Att komma överens om anställningsvillkoren.
När du börjar på ett nytt jobb ska du lämna ditt skattekort till arbetsgivaren.
Läs mer på InfoFinlands sida Skattekort.
Arbetstagaren har rätt att på begäran få ett arbetsintyg av arbetsgivaren när anställningen upphör.
Arbetsintyget är ett viktigt dokument där anställningens längd och arbetsuppgifterna nämns.
Arbetstagaren kan också be att orsaken till att anställningen upphört och en bedömning av arbetstagarens färdigheter och uppförande antecknas i intyget.
Arbetsgivaren är skyldig att utfärda ett arbetsintyg ännu tio år efter att anställningen har upphört och efter detta endast om detta inte medför en orimlig olägenhet för arbetsgivaren.
Om arbetstagaren vill att en bedömning av färdigheterna och uppförandet antecknas i arbetsintyget måste arbetsgivaren utfärda ett sådant intyg ännu fem år efter att anställningen har upphört till arbetstagaren på hans eller hennes begäran.
Arbetsgivare måste också ge arbetstagaren ett nytt arbetsintyg om arbetstagarens arbetsintyg kommer bort eller förstörs.
En arbetsgivare som avsiktligt eller av vårdslöshet inte utfärdar ett arbetsintyg bryter mot arbetsavtalslagen.
Arbetsavtalslagenfinska _ svenska _ engelska
linkkiArbetarskyddsförvaltningen:
Information om rätten till arbetsintygfinska _ svenska _ engelska
Jämlikheten är nedtecknad i lagar
Finlands grundlag garanterar jämlikt bemötande för alla.
Jämlikhet (yhdenvertaisuus) betyder att alla människor är likvärdiga oberoende av kön, ålder, etnisk eller nationell härkomst, nationalitet, språk, religion och övertygelse, åsikt, handikapp, hälsotillstånd, sexuell läggning eller någon annan orsak som gäller hans eller hennes person.
Om jämlikhet i arbetslivet föreskrivs i lagen om likabehandling och i arbetsavtalslagen.
Enligt dessa ska anställda behandlas lika när det gäller anställning, arbetsförhållanden, anställningsvillkor, utbildning för personalen och avancemang i karriären.
Finlands grundlagfinska _ svenska _ engelska _ ryska _ franska _ spanska _ tyska
Lag om likabehandlingfinska _ svenska _ engelska
Jämlikhet i rekryteringen
Lagen om likabehandling (yhdenvertaisuuslaki) förutsätter att alla arbetssökande behandlas lika.
Arbetsgivaren ska välja den sökande som har de bästa meriterna för uppgiften.
Arbetsgivaren ska också kunna bevisa att det finns godtagbara grunder för valet som anknyter till arbetets karaktär och att valet inte har varit diskriminerande.
Man får inte kräva sådana egenskaper av arbetssökanden som inte är nödvändiga i utförandet av arbetet.
Jämlikhet på arbetsplatsen
Arbetsgivaren får inte diskriminera de anställda när han eller hon fattar beslut om fördelning av arbetsuppgifter, erbjudande av möjligheter till avancemang eller upphävande av anställningen.
Arbetsdiskriminering är ett brott.
Om du misstänker att du har fallit offer för arbetsdiskriminering kan du ta kontakt med arbetarskyddsmyndigheterna eller ditt eget fackförbund.
Vid problem kan du fråga råd hos arbetarskyddsfullmäktige eller förtroendemannen.
linkkiArbetarskyddsförvaltningen:
Arbetarskyddfinska _ svenska _ engelska
linkkiRegionförvaltningsverket:
Arbetarskyddfinska _ svenska _ engelska
linkkiArbets- och näringsministeriet:
Likabehandling och förebyggande av diskriminering på arbetsplatserfinska _ svenska _ engelska
Jämställdhet (tasa-arvo) mellan könen
Enligt Finlands lag är män och kvinnor jämställda.
Män och kvinnor ska behandlas lika vid anställning och beträffande arbetsförhållanden och lönesättning.
En anställd får inte särbehandlas i arbetslivet på grund av graviditet eller föräldraskap.
I Finland finns en lag om likabehandling, som föreskriver att arbetsgivaren ska övervaka att jämställdheten på arbetsplatsen realiseras och att ingen diskrimineras på arbetsplatsen.
Jämställdhetsombudsmannen övervakar att lagen om likabehandling av män och kvinnor följs.
Om du misstänker att din arbetsgivare har diskriminerat dig på grund av ditt kön kan du be jämställdhetsombudsmannen om råd och anvisningar samt hjälp med att reda ut saken.
linkkiJämställdhetsombudsmannens byrå:
Information om jämställdhet i arbetslivetfinska _ svenska _ engelska _ ryska _ samiska
Jämställdhetslagenfinska _ svenska
Lediga jobb
Sök lediga jobb på jobbförmedlingssidor på internet, i tidningar eller på sociala medier (till exempel Facebook och LinkedIn).
Du hittar jobbförmedlingssidor när du skriver "avoimet työpaikat" (lediga jobb) i sökmotorns sökfält.
linkkiArbets- och näringsministeriet:
Lediga jobbfinska _ svenska
linkkiArbets- och näringsförvaltningen:
Länkar till jobbsajterfinska _ svenska _ engelska
linkkiArbets- och näringsministeriet:
Sysselsättningsutsikter för olika yrken i Finlandfinska _ svenska _ engelska
linkkiEures-portalen:
information om arbetsplatser i Europafinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiArbets- och näringsministeriet:
Tips för jobbsökningenfinska _ svenska _ engelska
Skapa nätverk och upprätthåll ditt kunnande
Du har nytta av nätverk när du söker jobb.
Identifiera och dra nytta av dina nätverk.
Lärare, studiekamrater, bekanta, tidigare kollegor och chefer kan också ingå i ditt nätverk.
Be om tips till jobbsökningen och hjälp med att skriva ansökningar av andra.
Fundera också på om du har någon i ditt nätverk som kan berätta om jobbtillfällen eller rekommendera dig.
Var aktiv.
Upprätthåll ditt kunnande, följ aktuella händelser och nyheter i din bransch, delta i kompletteringsutbildning och utveckla tidigare kunskaper.
Upprätthåll och utvidga ditt nätverk.
Även korta anställningar eller en praktik kan hjälpa dig att bygga ut ditt nätverk.
Besök fackevenemang i din bransch, gör frivilligarbete eller sök till ett mentorprogram.
Tänk på att frivilligarbete kan påverka din arbetslöshetsförsäkring.
Läs mer om frivilligarbete på InfoFinlands sida Frivilligarbete.
Lär dig finska eller svenska
När du kan språket är det lättare för dig att hitta jobb och sköta dina ärenden i det finländska samhället.
Du kan studera finska och svenska på olika kurser eller på egen hand via internet.
Läs mer om språkstudier i InfoFinlands avsnitt Finska och svenska språket.
Utnyttja sociala medier i jobbsökningen
Sociala nätverk på internet, såsom Facebook och LinkedIn, är bra verktyg för jobbsökningen.
Många arbetsgivare använder även Twitter som kommunikationskanal.
I tjänsterna kan du söka information om lediga jobb och bygga upp fackliga nätverk.
Du kan få viktig information om olika organisationers verksamhet och aktuella händelser i olika branscher eller delta i diskussioner.
Kontakta arbetsgivarna direkt
Du kan kontakta intressanta organisationer direkt och fråga om de har lediga jobb.
De flesta jobben är dolda jobb.
De annonseras inte ut öppet, utan arbetsgivarna söker arbetstagare via sina egna nätverk.
Du kan ringa en arbetsgivare direkt eller skicka en öppen ansökan via e-post.
Ofta kan du även skicka in en öppen ansökan via företagets webbplats.
Arbetsförmedlingstjänster
Du kan även söka jobb via företag som erbjuder arbetsförmedlingstjänster.
Arbetet kan vara kortvarigt, men det kan ge dig värdefull erfarenhet och du kan utvidga dina nätverk.
Du ingår ett avtal med företaget och företaget skickar dig till arbete för en annan arbetsgivare.
Via dessa företag kan du även få en fast anställning.
linkkiArbets- och näringsministeriet:
Hyrarbetsguidefinska _ svenska _ engelska
linkkiFörbundet för personaltjänsteföretag:
Personalbranschens regler om rekrytering av utlänningarfinska _ engelska
Sysselsätt dig som freelancer eller företagare
Arbete som freelancer innebär att du arbetar för flera uppdragsgivare utan fast anställning.
En freelancer måste själv sköta beskattningen och pensionsbetalningar.
Du kan fakturera vi en faktureringstjänst utan att starta ett eget företag.
Det kallas för lättföretagande.
Du kan även starta ett eget företag.
Tänk på att arbete som freelancer eller företagare kan påverka din arbetslöshetsförsäkring.
linkkiFreelanceri.info:
Länkar för frilansarefinska
Arbets- och näringsbyrån stöttar dig i jobbsökningen
Arbets- och näringsbyrån eller TE-byrån (TE-toimisto) ger dig handledning i jobbsökningen och information om lediga jobb och tillgängliga utbildningar.
Om du inte har ett jobb eller om du blir arbetslös, anmäl dig på arbets- och näringsbyrån senast på din första dag som arbetslös.
Läs mer på InfoFinlands sida Om du blir arbetslös.
Att anmäla sig som kund
Du kan anmäla dig som kund vid TE-byrån antingen vid den lokala TE-byrån eller på TE-byråns webbplats.
Om du är arbetslös arbetssökande, upprättar ni en integrationsplan eller en sysselsättningsplan.
Om du arbetar deltid eller bara lite, bedömer TE-byrån om du kan få en arbetslöshetsförmån samtidigt.
TE-byrån ordnar
yrkesutbildning
integrationsutbildning
utbildningsförsök
arbetsförsök
arbete med lönebidrag
arbetsträning
yrkesvägledning och karriärvägledning
linkkiArbets- och näringsministeriet:
Anmälan till arbets- och näringsbyrån finska _ svenska
linkkiTE-tjänster:
Videoklipp och broschyrer för invandrarefinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska
Integrationsutbildning
Om du har flyttat till Finland nyligen och behöver stöd med integrationen, kan du få plats i en integrationsutbildning via TE-byrån.
Integrationsutbildningen kan omfatta studier i finska, andra studier eller arbetsförsök.
Du kan även ansöka till utbildningen själv.
Du måste avtala om utbildningen med TE-byrån innan du inleder utbildningen.
Läs mer på InfoFinlands sida Integration i Finland.
linkkiArbets- och näringsministeriet:
Integrationstjänster för invandrarefinska _ svenska _ engelska
Stöd med jobbsökningen för under 30-åringar vid Navigatorn
Om du är under 30 år kan du få information om arbete, studier och annat som hör vardagslivet till vid Navigatorn.
Ohjaamofinska _ svenska _ engelska
Utbildnings- och arbetslivsguide för unga(pdf, 26 MB)finska _ svenska _ engelska _ ryska _ estniska _ somaliska
Välkommen till arbetslivet finska
Arbetslivets ABC finska
linkkiFFC:
Arbetslivet i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ kinesiska _ arabiska
linkkiArbets- och näringsministeriet:
Hitta jobb med hjälp av sysselsättningsprogrammet Kotouttamisen SIB finska _ engelska
När ett barn föds till familjen har föräldrarna rätt att ta familjeledighet, det vill säga stanna hemma för att ta hand om barnet.
Med familjeledighet avses
moderskapsledighet
faderskapsledighet
föräldraledighet
vårdledighet
Meddela din arbetsgivare om familjeledigheten senast två månader innan den börjar.
Familjeledigheterna är vanligen oavlönad ledighet.
Huruvida du får lön under familjeledigheten beror på ditt kollektivavtal.
Kontrollera detta med din arbetsgivare.
FPA betalar ut familjeförmåner för familjeledigheten: föräldrapenning och stöd för hemvård av barn.
Läs om villkoren för familjeförmånerna på InfoFinlands sida Stöd efter barnets födelse och Stöd för vård av barn i hemmet.
När familjeledigheterna upphör har arbetstagaren rätt att återvända till sitt eget arbete eller motsvarande arbete på den gamla arbetsplatsen.
Arbetsavtalet för en gravid kvinna får inte hävas och hon får inte diskrimineras på grund av sin graviditet.
I Finland känner arbetsgivarna och arbetstagarna till familjeledigheterna och de används allmänt.
linkkiArbets- och näringsministeriet:
Familjeledigheterfinska _ svenska _ engelska
Information om stöd till barnfamiljerfinska _ svenska _ engelska
Moderskapsledighet
Moderskapsledigheten är 105 vardagar.
Arbete under moderskapsledigheten är tillåtet om det kan utföras utan att moderns, fostrets eller barnets säkerhet äventyras.
Under moderskapsledigheten får man dock inte arbeta under de två veckor som föregår det beräknade födelsedatumet och under två veckor efter förlossningen.
Faderskapsledighet
Faderskapsledigheten är den del av föräldraledigheten som är avsedd att tas ut av fadern.
Faderskapsledigheten är allt som allt 54 vardagar.
Dessa dagar kan inte överföras till modern.
Du kan ta ut högst 18 dagar av din faderskapsledighet samtidigt som barnets mor är moderskaps- eller föräldraledig.
Dessa dagar kan du dela upp på högst fyra perioder.
De återstående 36 dagarna kan du dela upp på högst två perioder.
Under dessa dagar kan modern inte vara moderskapsledig samtidigt.
Avsikten är att fadern tar hand om barnet.
Du kan också ta ut alla 54 dagar av din faderskapsledighet vid olika tider med modern.
Du kan själv bestämma om du tar ut hela faderskapsledigheten eller bara en del av dagarna.
Faderskapsledigheten får endast tas ut före barnet har fyllt två år.
När barnet fyller två år kan du inte längre ta ut faderskapsledighet trots att du har dagar kvar.
Föräldraledighet
Efter moderskapsledigheten kan antingen modern eller fadern stanna hemma för att ta hand om barnet. Föräldraledigheten varar 158 vardagar.
Båda föräldrarna kan inte vara föräldralediga samtidigt.
Däremot kan man dela upp föräldraledigheten så att modern eller fadern stannar hemma växelvis för att ta hand om barnet.
Vårdledighet
Efter föräldraledigheten kan antingen modern eller fadern ta ut en oavlönad vårdledighet för att ta hand om barnet tills barnet fyller tre år.
Det förutsätter att modern eller fadern varit anställd hos samma arbetsgivare minst sex månader under det senaste året.
Under vårdledigheten betalar FPA stöd för hemvård av barn.
Se villkoren för stödet för hemvård av barn på InfoFinlands sida Stöd för vård av barn i hemmet.
Partiell vårdledighet
Du kan också vara vårdledig på deltid.
Då arbetar du kortare dagar och får på motsvarande sätt mindre lön.
Makarna kan vara partiellt vårdlediga samtidigt så att den ena förkortar sin arbetstid från morgonen och den andra från eftermiddagen.
Du kan vara partiellt vårdledig tills barnet har gått ut årskurs två.
Om du har hemkommun i Finland kan du ansöka om partiell vårdpenning hos FPA för hemvård av barn under tre år eller skolbarn i årskurserna 1 eller 2.
Partiell vårdpenning betalas inte för vård av ett barn som fyllt tre men ännu inte går i skolan.
Läs mer om partiell vårdpenning på InfoFinlands sida Stöd för vård av barn i hemmet.
I Finland har en arbetstagare rätt:
till lön och övriga minimivillkor enligt kollektivavtalet
till skydd utgående från lagar och avtal
att organisera sig
till en sund och trygg arbetsmiljö.
En arbetstagare är skyldig att
utföra arbetet omsorgsfullt
följa de överenskomna arbetstiderna
följa arbetsledningens anvisningar
vägra att delta i verksamhet som konkurrerar med arbetsgivaren
hålla affärs- och yrkeshemligheter
ta hänsyn till arbetsgivarens intresse.
Anställningsrådgivning för invandrare
Om du har frågor om eller problem med din anställning, kan du kontakta anställningsrådgivningen för invandrare.
Rådgivningen ges av Finlands Fackförbunds Centralorganisation FFC.
Du kan få rådgivning även om du inte är medlem i fackförbundet.
En jurist svarar på dina frågor till exempel om arbetsavtal, lön eller arbetstider.
Den kostnadsfria rådgivningen ges på finska och engelska.
Anställningsrådgivningen har öppet på tisdagar och onsdagar klockan 9–11 och 12–15.
Telefon: 0800 414 004
Du kan även ringa arbetarskyddsmyndigheternas riksomfattande rådgivningstelefon:
Tfn 0295 016 620
Mån.–fre. kl. 9–15
linkkiFFC:
Anställningsrådgivning för invandrarefinska _ svenska _ engelska
linkkiFFC:
Arbetslivet i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ kinesiska _ arabiska
linkkiArbetshälsoinstitutet:
Handboken Jobba i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ kurdiska _ tyska _ thai _ vietnamesiska
linkkiBrottsofferjouren:
Video om arbetstagarens rättigheter i Finlandengelska _ kinesiska _ arabiska _ thai _ hindi
Arbetstagarnas rättigheter tryggas med lagar och avtal
Arbetslagstiftningen och kollektivavtalen föreskriver vilka rättigheter och skyldigheter arbetstagare har.
Arbetstagar- och arbetsgivarförbunden förhandlar gemensamt fram branschspecifika kollektivavtal.
I lagstiftningen och kollektivavtalet fastställs till exempel minimilöner, arbetstider, semestrar, lön för sjukdomstid och uppsägningsvillkor.
Läs mer på InfoFinlands sidor Att komma överens om anställningsvillkoren och Innehållet i arbetsavtalet.
linkkiArbets- och näringsministeriet:
Broschyrer om arbetslagstiftningenfinska _ svenska _ engelska
Jämlikhet
Varje anställd har rätt till ett jämlikt och icke-diskriminerande bemötande när de söker jobb och på arbetsplatsen.
Läs mer på InfoFinlands sida Jämlikhet och jämställdhet i arbetslivet.
Arbetsavtal
Ett arbetsavtal uppstår när arbetstagaren och arbetsgivaren kommer överens om utförandet av ett arbete och lönen som betalas för det samt övriga förmåner och villkor.
Anställningsvillkoren bestäms enligt arbetslagstiftningen och kollektivavtalet.
Arbetsavtalet är bindande för båda parterna.
Läs mer om arbetsavtalet på InfoFinlands sidor Att komma överens om anställningsvillkoren och Innehållet i arbetsavtalet.
Fackförbund
I Finland är facklig organisering vanligt och aktiva fackförbundsmedlemmar trakasseras inte.
Du kan ansluta dig till fackförbundet i din egen bransch.
Förbundet strävar efter att trygga sina medlemmars intressen i arbetslivet.
Läs mer på InfoFinlands sida Fackförbund.
Arbetarskydd
Arbetsgivaren är skyldig att trygga de anställdas säkerhet.
Arbetarskyddsförvaltningen övervakar att de i lagen stadgade arbetarskyddsföreskrifterna följs på arbetsplatserna.
Läs mer på InfoFinlands sida Arbetarskydd.
Utkomstskydd för arbetslösa
När en person som är fast bosatt i Finland blir arbetslös, har han eller hon rätt att få utkomstskydd för arbetslösa.
Läs mer på InfoFinlands sida Utkomstskydd för arbetslösa.
En invandrare som har bott tillräckligt länge i Finland kan få pension på grund av sin ålder eller arbetsoförmögenhet.
Läs mer på InfoFinlands sida Pension.
Beskattning
När du arbetar i Finland måste du betala skatter.
Läs mer på InfoFinlands sida Beskattning.
Företagshälsovård
Varje arbetsgivare är skyldig att ordna förebyggande företagshälsovård för sina anställda.
Läs mer på InfoFinlands sida Företagshälsovård.
Familjeledigheter
När ett barn föds till familjen kan modern eller fadern enligt lag stanna hemma för att ta hand om barnet.
Läs mer på InfoFinlands sida Familjeledigheter.
Arbetsintyg
När en anställning upphör har den anställda rätt att få ett skriftligt arbetsintyg av arbetsgivaren.
Läs mer på InfoFinlands sida Arbetsintyg.
Anmäl flyttningen till myndigheterna
När du flyttar utomlands från Finland ska du göra en flyttanmälan till magistraten (maistraatti)
Du kan göra flyttanmälan på internet eller med en blankett som du får i magistraten eller på posten.
Om du flyttar permanent från Finland eller vistas utomlands två år utan avbrott återkallas ditt uppehållstillstånd.
Du kan ställa Migrationsverket (Maahanmuuttovirasto) en ansökan om att inte återkalla ditt uppehållstillstånd.
Ansökan ska göras innan du har vistats utomlands över två år.
Mer information om detta hittar du på InfoFinlands sida Kan jag förlora mitt uppehållstillstånd?.
Flytt utomlands och den sociala tryggheten
När du flyttar utomlands måste du meddela detta till FPA, om du får FPA:s förmåner eller om du har det europeiska sjukvårdskortet.
Om du får FPA:s förmåner har du vanligtvis rätt till dem även i fortsättningen om din utlandsvistelse varar sex månader eller mindre.
Då anses din utlandsvistelse vara tillfällig och du behöver inte nödvändigtvis anmäla den till FPA.
En utlandsvistelse som varar 3–6 månader bör du anmäla den till FPA, om
du får det allmänna bostadsbidraget
du får stöd för hemvård av barn eller
om du måste köpa receptbelagda läkemedel på apoteket för över tre månaders tid.
Om du ska arbeta i ett EU-/EES-land omfattas du av den sociala tryggheten i arbetslandet under den tid då du arbetar i landet, även om arbetet pågår mindre än sex månader.
Då har du inte rätt till FPA:s förmåner.
Om du flyttar utomlands för över sex månader anses din flytt vara permanent.
Din rätt till FPA:s förmåner upphör då samma dag som du flyttar.
I vissa situationer kan du behålla din rätt till FPA:s förmåner även om du vistas utomlands längre än sex månader.
När du är utomlands och har rätt till FPA:s förmåner ska du alltid anmäla ändringar i dina förhållanden till FPA.
Till exempel ändrade familjeförhållanden eller att du börjar arbeta kan påverka din rätt till FPA:s förmåner.
Du hittar mer information om den sociala tryggheten i Finland på FPA:s webbplats och på InfoFinlands sida Den sociala tryggheten i Finland.
Frivillig återflyttning av flyktingar, asylsökande och emigranter
Om du vill återvända till ditt hemland kan du i vissa fall få stöd för frivilligt återvändande.
Stödet består antingen av pengar eller tjänster.
Penningsummans storlek beror på vilket land du återvänder till.
Tjänsten kan till exempel vara att du får hjälp med att leta efter en bostad eller arbetsplats i det land dit du återvänder.
Du kan få stöd om:
du är asylsökande och handläggningen av din ansökan är oavslutad
du har fått ett negativt beslut på din asylansökan
du är ett offer för människohandel och du inte har en hemkommun i Finland
du har ett tillfälligt uppehållstillstånd på grund av hinder för avlägsnande ur landet
du har fått tillfälligt skydd
din flyktingstatus i Finland har upphört eller återkallats eller det har fattats beslut om att avvisa dig.
Om du är kund hos en mottagningscentral kan du ansöka om stöd för frivilligt återvändande vid din egen mottagningscentral.
Om du inte är kund hos en mottagningscentral kan du ansöka om stöd hos Migrationsverket.
Flyttanmälanfinska _ svenska _ engelska
Återkallelse av uppehållstillståndfinska _ svenska _ engelska
Flytt utomlands och social trygghetfinska _ svenska _ engelska
Frivillig återflyttningfinska _ svenska _ engelska
Om du blir sjuk eller råkar ut för en olycka har du rätt att stanna hemma från arbetet.
Arbetsgivaren är skyldig att betala lön för sjukledigheten.
Om din anställning varat över en månad före insjuknandet får du lönen till fullt belopp för minst den dag då du insjuknade och nio därefter följande dagar.
Om du fortfarande inte kan återvända till arbetet kan du söka sjukdagpenning (sairauspäiväraha) hos FPA om du omfattas av den finländska sjukförsäkringen.
Läs mer på InfoFinlands sida Den sociala tryggheten i Finland.
Det kan hända att man i kollektivavtalet har kommit överens om andra villkor och du får lön för en längre tid.
Arbetsgivaren har rätt att kräva ett läkarintyg för den tid då du är sjuk.
Om du blir sjuk och inte kan arbeta ska du utan dröjsmål meddela detta till din chef.
Din chef berättar för dig om du behöver ett läkarintyg om sjukdomen direkt eller först från och med den fjärde sjukledighetsdagen.
Sjukledighet är ingen semester utan den beviljas för att du ska återhämta dig från din sjukdom.
Därför får du under dessa dagar inte göra något som kan äventyra ditt tillfrisknande.
Sjukdagpenningfinska _ svenska _ engelska
Att ansöka om sjukdagpenningfinska _ svenska _ engelska
Om du har avlagt examen i något annat land kan du behöva beslut om erkännande av examen för att kunna arbeta eller studera i Finland.
I de flesta situationerna bedömer arbetsgivaren, läroanstalten eller högskolan vilken behörighet och kompetens din utländska examen ger.
Du behöver Utbildningsstyrelsens eller någon annan myndighets beslut om erkännande av examen om du vill arbeta inom ett reglerat yrke eller en uppgift som kräver högskoleexamen på viss nivå.
linkkiUtbildningsstyrelsen:
Erkännande av en examenfinska _ svenska _ engelska
linkkiUtbildningsstyrelsen :
Broschyr om erkännande av examen(pdf, 102,14 kt)finska _ svenska _ engelska _ ryska _ estniska _ franska _ spanska _ kinesiska _ persiska _ arabiska
linkkiUtbildningsstyrelsen :
Diagram över erkännande av examen(pdf, 410,87 kt)finska _ svenska _ engelska _ ryska
linkkiUtbildningsstyrelsen:
Servicepriserfinska _ svenska _ engelska
Om du vill fortsätta dina studier i Finland
Högskolor och läroanstalter beslutar om antagning av studerande.
De beslutar också huruvida dina utländska studier och din övriga kompetens kan godkännas som en del av den examen du avlägger i Finland.
Om du har avlagt högskolestudier utomlands och vill fortsätta dina studier i Finland kan du få information och handledning vid högskolornas tjänster för studerande och SIMHE-tjänsterna.
linkkiUtbildningsstyrelsen:
Högskolor som erbjuder SIMHE-tjänsterfinska _ svenska _ engelska
Uppgifter som inte kräver en viss utbildning
Enligt Finlands lag kräver inte alla uppgifter en viss utbildning eller examen på en viss nivå.
Till exempel bedömer arbetsgivare i privatsektorn oftast själv huruvida en utländsk examen ger tillräckliga kvalifikationer för uppgiften.
Jämställande av nivån på en högskolexamen
För uppgifter inom den offentliga sektorn (kommun eller stat) krävs ofta examen på en viss nivå, till exempel en högre högskoleexamen.
Om du har avlagt en högskoleexamen utomlands kan du ansöka om beslut om jämställande av nivån på en högskolexamen vid Utbildningsstyrelsen.
Beslutet är avgiftsbelagt.
När din examensnivå har jämställts med en finländsk högskoleexamen, kan du söka till uppgifter som kräver den nivå på högskoleexamen som du har.
linkkiUtbildningsstyrelsen:
Jämställande av nivån på en högskolexamenfinska _ svenska _ engelska
Reglerade yrken
I Finland är vissa yrken reglerade.
Det betyder att det stadgas i lag vilken utbildning som krävs för dessa yrken.
Sådana uppgifter är till exempel fysioterapeut, läkare, tandläkare, provisor, sjukskötare, advokat, revisor, klasslärare och sotare.
Branschspecifika myndigheter beslutar om rätten att utöva ett reglerat yrke eller använda en yrkesbeteckning.
Till exempel inom social- och hälsovårdsbranschen fattas beslutet av Valvira, och inom undervisningssektorn av Utbildningsstyrelsen.
Beslutet är avgiftsbelagt.
På Utbildningsstyrelsens webbplats hittar du en förteckning över reglerade yrken och de myndigheter som fattar beslut.
linkkiUtbildningsstyrelsen:
Reglerade yrken och ansvariga myndigheterfinska _ svenska _ engelska
Information om erkännande av examen för yrken inom hälsovårdenfinska _ svenska _ engelska
Reglerade yrken och examen från ett annat EU-land
Om
du är medborgare i ett EU-land, EES-land eller Schweiz och du har
förvärvat kvalifikationer för ett yrke som är reglerat i Finland i ett EU-land, EES-land eller Schweiz,
kan du ansöka om erkännande av yrkeskvalifikationer för detta yrke hos den branschspecifika myndigheten.
Om din utbildning skiljer sig mycket från den utbildning som krävs i Finland måste du eventuellt avlägga en anpassningsperiod eller ett lämplighetsprov.
linkkiUtbildningsstyrelsen:
Erkännande av yrkeskvalifikationer som förvärvats i ett EU-landfinska _ svenska _ engelska
linkkiEuropeiska kommissionen:
Information om reglerade yrken i EU-ländernaengelska
Utländsk yrkesexamen
Om du har avlagt en yrkesexamen utomlands kan du ansöka om ett utlåtande om det hos Utbildningsstyrelsen.
I utlåtandet beskrivs examensnivån och innehåll samt för vilka uppgifter examen ger kvalifikationer i det land där du har avlagt examen.
Utlåtandet ger dig dock inte kvalifikationer att utöva ett reglerat yrke i Finland.
linkkiUtbildningsstyrelsen:
Utlåtanden om utländska yrkesexamenfinska _ svenska _ engelska
Översättning av handlingar
Om originalspråket för ditt betyg inte är finska, svenska eller engelska behöver du vanligtvis en officiell översättning av handlingarna som görs av en auktoriserad översättare.
Vissa myndigheter godkänner även handlingar på andra europeiska språk.
Läs noga anvisningarna om ansökning från den branschspecifika myndigheten.
Många länder har en beskickning i Finland.
Beskickningen kan antingen vara en ambassad eller ett konsulat.
Ambassaderna finns i Helsingfors.
Vissa länder har också konsulat i andra städer.
Om du behöver sköta ett ärende med myndigheterna i ditt hemland ska du ta kontakt med ditt lands beskickning.
Via beskickningen kan du ofta uträtta till exempel följande ärenden:
Få en födelseattest
Ansöka om medborgarskap i ditt hemland om du har förlorat det eller avstått från det
Anmäla födelsen av ditt barn till myndigheterna i ditt hemland om barnet föds i Finland
Ansöka om medborgarskap i ditt hemland för ditt barn om barnet har fötts i Finland
Registrera ett äktenskap i ditt hemland om du har gift dig i Finland
Rösta i val i ditt hemland
Observera att alla beskickningar inte erbjuder samma tjänster.
Det är inte nödvändigtvis möjligt att sköta alla ovannämnda ärenden i alla beskickningar.
Vilka tjänster ditt lands beskickning tillhandahåller beror på lagen i ditt hemland.
Mer information får du från ditt hemlands beskickning.
Alla länder har inte en beskickning i Finland.
I detta fall betjänas du ofta av ditt hemlands beskickning i något av Finlands grannländer.
På det finska utrikesministeriets webbplats finns en förteckning över andra länders beskickningar i Finland.
Där hittar du även kontaktuppgifterna till beskickningarna.
Andra länders beskickningar i Finlandfinska _ svenska _ engelska
Alla har rätt till företagshälsovård
I Finland är arbetsgivare skyldiga att ordna förebyggande företagshälsovård för sina anställda.
Arbetsgivaren kan också ordna sjukvårdstjänster för sina anställda.
Inom företagshälsovården har arbetstagaren tillgång till hälsovårdarens, företagsläkarens och företagspsykologens tjänster.
Ofta finns det i företagshälsovården också fysioterapeuter.
Specialisternas tjänster ingår vanligen inte i företagshälsovården.
Fråga din arbetsgivare vad företagshälsovården på din arbetsplats omfattar.
Rätten till företagshälsovårdens tjänster omfattar inte den anställdas familj.
Avsikten med företagshälsovården är att främja hälsan och arbetsförmågan och samarbetet på arbetsplatserna.
Anställda inom företagshälsovården har sekretessplikt.
De lämnar inte ut information om din situation till din arbetsgivare, om inte du själv har gett tillstånd till det.
Företagshälsovården kan dock ge din arbetsgivare en bedömning av huruvida ditt hälsotillstånd tillåter att du fortsätter att arbeta.
Fpa ersätter arbetsgivaren och företagaren en del av kostnaderna för företagshälsovården, om dessa är nödvändiga och rimliga.
linkkiArbetarskyddsförvaltningen:
Information om företagshälsovårdenfinska _ svenska _ engelska
linkkiArbetshälsoinstitutet:
Information om företagshälsovårdenfinska _ svenska
linkkiSocial- och hälsovårdsministeriet:
Företagshälsovårdfinska _ svenska _ engelska
Lagen om företagshälsovårdfinska _ svenska _ engelska
Sjukdagpenningfinska _ svenska _ engelska
Läs jobbannonsen noga
Innan du skriver din jobbansökan, läs jobbannonsen noga och fundera på vilka färdigheter och vilket kunnande arbetsgivaren är ute efter.
Fundera på hur ditt kunnande motsvarar arbetsgivarens önskemål och krav.
Du kan också kontakta arbetsgivaren och begära mer information, om du undrar över något som inte framgår av jobbannonsen.
Ring arbetsgivaren bara om du har en konkret fråga om arbetsplatsen.
Jobbansökan
Vanligtvis när du söker ett jobb, skickar du en jobbansökan och ditt CV, alltså din meritförteckning, till arbetsgivaren.
Ibland kan jobbansökningen vara en video, en portfölj eller till exempel en webbsida.
Skriv ansökan och CV på samma språk som används i annonsen.
Skriv en ny ansökan och uppdatera ditt CV varje gång när du ansöker om ett nytt jobb.
Du kan skriva ansökningstexten direkt i e-postmeddelandet eller bifoga den till e-postmeddelandet tillsammans med ditt CV.
Lägg till bilagorna alltid i PDF-format.
Ofta kan du skicka in ansökan och CV via arbetsgivarens webbplats.
Syftet med din jobbansökan är att väcka arbetsgivarens intresse så att du blir kallad till anställningsintervju.
Ansökningen är ett svar på jobbannonsen.
Du ska svara på de önskemål och krav som nämns i jobbannonsen.
Lyft fram sådant som är viktigt i arbetsuppgiften.
Ge konkreta exempel på ditt kunnande.
Intyga arbetsgivaren om att du är lämplig för uppgiften.
En jobbansökan är oftast en knapp sida.
Be någon att läsa igenom och granska din ansökan.
Löneanspråk
Ofta ska man ange sitt löneanspråk i ansökningen.
Det är ofta svårt att uppskatta rätt belopp.
Löneanspråket får inte vara för stort, men inte heller för litet.
Från fackförbund får du mer information om lönenivån i olika branscher.
Lönejämförelse finska _ engelska
Gå igenom dina utbildningar och din arbetserfarenhet och fundera på vilka färdigheter du lärt dig i dem.
Vilka är dina styrkor?
Fundera också på vilket kunnande du har fått från dina fritidsintressen eller andra erfarenheter.
Tidsenliga intyg
Spara intygen från dina tidigare jobb och studier.
Kom ihåg att alltid begära ett intyg när du haft ett jobb, avlagt en praktik eller studerat.
Arbetsgivaren har skyldighet att utfärda ett intyg ännu tio år efter att anställningen upphört.
Du behöver vanligtvis inte skicka in dina arbetsintyg i förväg till arbetsgivaren, men det är bra att ta med dem till anställningsintervjun för det fall att arbetsgivaren vill se dem.
Det skulle vara bra att ha översättningar till finska eller svenska av alla intyg som du fått utomlands.
Mer information om detta finns på InfoFinlands sida Arbetsintyg.
Erkännande av examen
Det är lättare att söka jobb om du vet hur en examen som du avlagt utomlands motsvarar en finländsk examen.
Du kan ansöka om erkännande av utländsk examen vid Utbildningsstyrelsen.
Erkännande av examen är avgiftsbelagt.
Mer information om detta finns på InfoFinlands sida Utländsk examen i Finland.
linkkiUtbildningsstyrelsen:
Erkännande av en examenfinska _ svenska _ engelska
Öppen ansökan
Du kan ta direkt kontakt med en arbetsplats som du är intresserad av.
Du kan skicka in en öppen ansökan eller ringa arbetsgivaren, trots att de inte har några lediga jobb just nu.
I den öppna ansökan ska du berätta vad du kan och hurdana uppgifter du skulle kunna utföra.
Bifoga din meritförteckning, alltså CV, till ansökan.
Meritförteckning eller CV
En meritförteckning, eller ett CV, är en kortfattad och tydlig sammanfattning av ditt kunnande, din arbetserfarenhet och din utbildning.
Det finns olika CV-mallar.
I ett kompetensbaserat CV kan du gruppera dina färdigheter i olika kompetensområden.
CV:t kan även vara en video, en portfölj eller en webbsida.
Bekanta dig med olika CV-mallar och forma ditt eget CV såsom det passar dig.
Ett CV är vanligtvis 1–2 sidor långt.
Kom ihåg att uppdatera ditt CV för varje ny ansökan.
Vad innehåller ett CV?
Namn och kontaktuppgifter – Adress, e-postadress, telefonnummer
Arbetserfarenhet – Lista dina tidigare anställningar, den senaste först.
Ange också anställningens längd.
Beskriv dina arbetsuppgifter och de färdigheter som du lärt dig i arbetet.
Utbildning – Lista dina examina i kronologisk ordning, den senaste först.
Lägg till namnet på examen, utbildningsprogrammet och läroanstalten och när du tog examen.
Kurser – Lista kurserna i finska och andra kurser som du avlagt under en egen rubrik.
Övrigt kunnande – Språkkunskaper, IT-kunskaper, avlagda tillståndskort, till exempel hygienpass.
Publikationer eller andra arbetsprov
– Om du vill kan du även lista dina publikationer eller arbetsprov.
Fritidsintressen, förtroendeuppdrag
– Du kan även lyfta fram dina intressen.
Referenser – Du kan lägga till namnen på personer som har lovat att rekommendera dig för arbetsuppgiften.
Lägg till kontaktuppgifterna till dem.
Kom ihåg att be personen om tillstånd för detta.
I början av CV:t kan du tillfoga en sammanfattning eller profil där du beskriver din bakgrund och din kärnkompetens med några ord.
Du kan berätta vilka målsättningar du har med jobbsökningen eller vilken specialkompetens du besitter.
Du kan också lägga till ett fotografi.
linkkiArbets- och näringsministeriet:
Så här skriver du en jobbansökan och ett CVfinska _ svenska _ engelska
Kompetensbaserat CV
Ett kompetensbaserat CV lyfter fram ditt kunnande, dina färdigheter och dina erfarenheter.
Välj några kompetensområden och beskriv under rubrikerna dina erfarenheter, färdigheter och prestationer inom dem.
Du kan också lägga till sådant kunnande som du har införskaffat till exempel i frivilligarbete, fritidsintressen eller studier.
Dessutom kan du lista din arbetserfarenhet och utbildning i kronologisk ordning.
I början av CV:t kan du tillfoga en sammanfattning eller profil där du beskriver din bakgrund och din kärnkompetens med några ord.
Du kan berätta vilka målsättningar du har med jobbsökningen eller vilken specialkompetens du besitter.
Skriv ett eget CV för varje arbetsplats.
Lyft fram sådana färdigheter som behövs i uppgiften.
Fundera på vad arbetsgivaren bör veta om dina färdigheter och ditt kunnande.
Europass-CV
Europass är ett allmäneuropeiskt CV, alltså en allmäneuropeisk meritförteckning.
Det består av fem dokument som har till syfte att hjälpa arbetstagare och studerande att presentera sitt kunnande i Europa.
Dokumenten används i alla EU/EES-länderna.
Du kan använda Europass när du söker jobb eller studieplats.
Europass är särskilt nyttigt om du ansöker om ett jobb eller en utbildningsplats i Finland från ett annat EU-land.
linkkiEuropass.eu:
Information om CVfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Förbered dig på anställningsintervjun
Bekanta dig med arbetsgivaren i förväg till exempel med hjälp av webbplatsen.
Fundera på hur du ska lyfta fram ditt kunnande och din lämplighet för uppgiften.
Öva på att beskriva din bakgrund och din yrkeskunnighet med några meningar.
Fundera i förväg på vilka frågor arbetsgivaren kan ställa till dig.
Öva på att besvara allmänna frågor som ingår i en anställningsintervju.
Arbetsgivaren får inte fråga om din familj, vilken religion du har eller om du är politiskt aktiv.
Visa att du har bekantat dig med arbetsgivarens organisation och arbetsuppgiften i förväg och att du har ett äkta intresse för jobbet.
Fundera också på vilka frågor du vill ställa till arbetsgivaren.
linkkiArbets- och näringsministeriet:
Anvisningar för jobbintervjunfinska _ svenska _ engelska
Att börja på ett nytt jobb
Skriv alltid ett skriftligt anställningsavtal innan du börjar på ett nytt jobb.
Kom överens om anställningsavtalets innehåll med arbetsgivaren.
Läs avtalet noga innan du undertecknar det.
Läs mer på InfoFinlands sida Att komma överens om anställningsvillkoren.
När du börjar på ett nytt jobb ska du lämna ditt skattekort till arbetsgivaren.
Läs mer på InfoFinlands sida Skattekort.
Finska medborgare har vissa rättigheter och skyldigheter som utlänningar bosatta i Finland inte nödvändigtvis har.
Rättigheter
rätt att få finskt pass
rätt att resa till Finland och vägra att bli utlämnad till ett annat land
rätt att rösta i presidentval, riksdagsval och folkomröstningar då man fyllt 18 år.
rätt att ställa upp som kandidat i riksdagsval då man fyllt 18 år.
möjlighet att bli utnämnd till sådana statliga ämbeten för vilka det krävs finskt medborgarskap
EU-medborgarnas rättigheter som rätten att fritt röra sig och arbeta inom EU:s område och rätten att rösta och ställa upp som kandidat i EU-val
Skyldigheter
Skyldighet att delta i landets försvar eller bistå i det.
Män som har fyllt 18 år har värnplikt (asevelvollisuus).
Skyldighet att följa Finlands lagar även annanstans än i Finland.
Finska medborgare kan i Finland dömas för brott som begåtts utomlands.
Observera att dessa är rättigheter och skyldigheter som ingår i det finska medborgarskapet.
Information om rättigheter och skyldigheter som gäller alla som är bosatta i Finland finns på InfoFinlands sida Dina rättigheter och skyldigheter i Finland.
Finska medborgares rättigheter och skyldigheterfinska _ svenska _ engelska
linkkiFörsvarsmakten:
Värnpliktfinska _ svenska _ engelska
Att ansöka om finskt passfinska _ svenska _ engelska
Att ansöka om finskt pass utomlandsfinska _ svenska _ engelska
Arbetarskyddsverksamhet på arbetsplatsen
I Finland fästs stor uppmärksamhet vid arbetssäkerhet.
Arbetsgivaren ansvarar för att alla kan arbeta tryggt.
Arbetsgivaren ska ordna arbetsplatsintroduktion för nya anställda.
Arbetsgivaren är också skyldig att göra de anställda förtrogna med arbetsplatsens säkerhetsanvisningar och lära dem korrekta arbetssätt.
De anställda ska också själva sörja för arbetssäkerheten.
Arbetet ska utföras enligt anvisningarna.
Om arbetet är uppenbart farligt kan den anställda vägra att utföra det.
På arbetsplatserna ska det finnas tillräckligt många personer med kunskaper i första hjälpen, första hjälpen-utrustning samt instruktioner för olycksfall.
Arbetsgivarna ordnar utbildning i första hjälpen på arbetsplatsen.
Om det finns minst tio anställda på en arbetsplats väljer dessa ut en arbetarskyddsfullmäktig som representerar dem.
Arbetarskyddsfullmäktige gör sig insatt i arbetarskyddsfrågor som gäller arbetsplatsen, deltar i arbetsplatsens arbetarskyddsinspektioner och informerar de anställda om ärenden som rör arbetets säkerhet och hälsa.
Arbetsgivaren utser för varje arbetsplats en arbetarskyddschef, som bistår arbetsgivaren i samarbetet med anställda och arbetarskyddsmyndigheter.
Arbetarskyddsmyndigheter
I Finland finns det fem ansvarsområden för arbetarskydd som lyder under Regionförvaltningsverket (RFV).
Ansvarsområdena övervakar att de lagenliga arbetarskyddsföreskrifterna följs på arbetsplatserna.
Ansvarsområdena för arbetarskydd ger både arbetstagare och arbetsgivare råd i frågor som gäller arbetets säkerhet och hälsa samt i frågor som rör anställningsvillkor.
Arbetarskyddsinspektörerna utför kontroller på arbetsplatser.
De kontrollerar bland annat om säkerhetsföreskrifterna följs på arbetsplatsen, om man har gett tillräcklig introduktion i arbetet och huruvida utländska arbetstagares arbetsförhållanden och anställningsvillkor följer finländska lagar och avtal.
Arbetarskyddsinspektören har rätt att få tillträde till varje arbetsplats och tillgång till de dokument som är väsentliga för övervakningen av arbetarskyddet.
Arbetarskyddsmyndigheten kan förplikta arbetsgivaren att rätta till brister i arbetssäkerheten som förekommer på arbetsplatsen
linkkiArbetarskyddsförvaltningen:
Information om arbetarskydd och råd vid problemfinska _ svenska _ engelska
linkkiEuropeiska arbetsmiljöbyrån:
Information om arbetarskyddfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Lediga jobb
Sök lediga jobb på jobbförmedlingssidor på internet, i tidningar eller på sociala medier (till exempel Facebook och LinkedIn).
Du hittar jobbförmedlingssidor när du skriver "avoimet työpaikat" (lediga jobb) i sökmotorns sökfält.
linkkiArbets- och näringsministeriet:
Lediga jobbfinska _ svenska
linkkiArbets- och näringsförvaltningen:
Länkar till jobbsajterfinska _ svenska _ engelska
linkkiArbets- och näringsministeriet:
Yrkesbarometern finska _ svenska _ engelska
linkkiEures-portalen:
information om arbetsplatser i Europafinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiArbets- och näringsministeriet:
Tips för jobbsökningenfinska _ svenska _ engelska
Skapa nätverk och upprätthåll ditt kunnande
Du har nytta av nätverk när du söker jobb.
Identifiera och dra nytta av dina nätverk.
Lärare, studiekamrater, bekanta, tidigare kollegor och chefer kan också ingå i ditt nätverk.
Be om tips till jobbsökningen och hjälp med att skriva ansökningar av andra.
Fundera också på om du har någon i ditt nätverk som kan berätta om jobbtillfällen eller rekommendera dig.
Var aktiv.
Upprätthåll ditt kunnande, följ aktuella händelser och nyheter i din bransch, delta i kompletteringsutbildning och utveckla tidigare kunskaper.
Upprätthåll och utvidga ditt nätverk.
Även korta anställningar eller en praktik kan hjälpa dig att bygga ut ditt nätverk.
Besök fackevenemang i din bransch, gör frivilligarbete eller sök till ett mentorprogram.
Tänk på att frivilligarbete kan påverka din arbetslöshetsförsäkring.
Läs mer om frivilligarbete på InfoFinlands sida Frivilligarbete.
Lär dig finska eller svenska
När du kan språket är det lättare för dig att hitta jobb och sköta dina ärenden i det finländska samhället.
Du kan studera finska och svenska på olika kurser eller på egen hand via internet.
Läs mer om språkstudier i InfoFinlands avsnitt Finska och svenska språket.
Utnyttja sociala medier i jobbsökningen
Sociala nätverk på internet, såsom Facebook och LinkedIn, är bra verktyg för jobbsökningen.
Många arbetsgivare använder även Twitter som kommunikationskanal.
I tjänsterna kan du söka information om lediga jobb och bygga upp fackliga nätverk.
Du kan få viktig information om olika organisationers verksamhet och aktuella händelser i olika branscher eller delta i diskussioner.
Kontakta arbetsgivarna direkt
Du kan kontakta intressanta organisationer direkt och fråga om de har lediga jobb.
De flesta jobben är dolda jobb.
De annonseras inte ut öppet, utan arbetsgivarna söker arbetstagare via sina egna nätverk.
Du kan ringa en arbetsgivare direkt eller skicka en öppen ansökan via e-post.
Ofta kan du även skicka in en öppen ansökan via företagets webbplats.
Arbetsförmedlingstjänster
Du kan även söka jobb via företag som erbjuder arbetsförmedlingstjänster.
Arbetet kan vara kortvarigt, men det kan ge dig värdefull erfarenhet och du kan utvidga dina nätverk.
Du ingår ett avtal med företaget och företaget skickar dig till arbete för en annan arbetsgivare.
Via dessa företag kan du även få en fast anställning.
linkkiArbets- och näringsministeriet:
Hyrarbetsguidefinska _ svenska _ engelska
linkkiFörbundet för personaltjänsteföretag:
Personalbranschens regler om rekrytering av utlänningarfinska _ engelska
Sysselsätt dig som freelancer eller företagare
Arbete som freelancer innebär att du arbetar för flera uppdragsgivare utan fast anställning.
En freelancer måste själv sköta beskattningen och pensionsbetalningar.
Du kan fakturera vi en faktureringstjänst utan att starta ett eget företag.
Det kallas för lättföretagande.
Du kan även starta ett eget företag.
Tänk på att arbete som freelancer eller företagare kan påverka din arbetslöshetsförsäkring.
linkkiFreelanceri.info:
Länkar för frilansarefinska
Arbets- och näringsbyrån stöttar dig i jobbsökningen
Arbets- och näringsbyrån eller TE-byrån (TE-toimisto) ger dig handledning i jobbsökningen och information om lediga jobb och tillgängliga utbildningar.
Om du inte har ett jobb eller om du blir arbetslös, anmäl dig på arbets- och näringsbyrån senast på din första dag som arbetslös.
Läs mer på InfoFinlands sida Om du blir arbetslös.
Att anmäla sig som kund
Du kan anmäla dig som kund vid TE-byrån antingen vid den lokala TE-byrån eller på TE-byråns webbplats.
Om du är arbetslös arbetssökande, upprättar ni en integrationsplan eller en sysselsättningsplan.
Om du arbetar deltid eller bara lite, bedömer TE-byrån om du kan få en arbetslöshetsförmån samtidigt.
TE-byrån ordnar
yrkesutbildning
integrationsutbildning
utbildningsförsök
arbetsförsök
arbete med lönebidrag
arbetsträning
yrkesvägledning och karriärvägledning
linkkiArbets- och näringsministeriet:
Anmälan till arbets- och näringsbyrån finska _ svenska
linkkiTE-tjänster:
Videoklipp och broschyrer för invandrarefinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska
Integrationsutbildning
Om du har flyttat till Finland nyligen och behöver stöd med integrationen, kan du få plats i en integrationsutbildning via TE-byrån.
Integrationsutbildningen kan omfatta studier i finska, andra studier eller arbetsförsök.
Du kan även ansöka till utbildningen själv.
Du måste avtala om utbildningen med TE-byrån innan du inleder utbildningen.
Läs mer på InfoFinlands sida Integration i Finland.
linkkiArbets- och näringsministeriet:
Integrationstjänster för invandrarefinska _ svenska _ engelska
Stöd med jobbsökningen för under 30-åringar vid Navigatorn
Om du är under 30 år kan du få information om arbete, studier och annat som hör vardagslivet till vid Navigatorn.
Ohjaamofinska _ svenska _ engelska
Utbildnings- och arbetslivsguide för unga(pdf, 26 MB)finska _ svenska _ engelska _ ryska _ estniska _ somaliska
Välkommen till arbetslivet finska
Arbetslivets ABC finska
linkkiFFC:
Arbetslivet i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ kinesiska _ arabiska
linkkiArbets- och näringsministeriet:
Hitta jobb med hjälp av sysselsättningsprogrammet Kotouttamisen SIB finska _ engelska
För att få finskt medborgarskap genom en medborgarskapsansökan krävs något av följande:
Du kan tillförlitligt intyga din identitet.
Du är minst 18 år gammal eller gift.
Du har bott i Finland tillräckligt länge.
Hur lång boendetid som krävs beror på din situation, vanligtvis ska du ha bott här minst 4–7 år.
Du har inte begått brott.
Du har inte lämnat till exempel skatter, böter, underhållsbidrag eller sjukhusavgifter obetalda.
Du kan redogöra för hur du försörjer dig i Finland.
Du kan finska, svenska eller det finska eller finlandssvenska teckenspråket åtminstone nöjaktigt.
Läs mer om att bevisa dina språkkunskaper på InfoFinlands sida Officiellt intyg över språkkunskaper.
Läs mer om att studera finska och svenska på InfoFinlands sida Finska och svenska språket.
Du kan ansöka om medborgarskap elektroniskt i tjänsten Enter Finland.
Fyll i en ansökan och lägg till bilagorna.
För en ansökan behöver du åtminstone följande dokument:
Ett giltigt identitetsbevis
En utredning om dina språkkunskaper
En utredning om ditt uppehälle.
Betala samtidigt också ansökningens handläggningsavgift.
När du fyllt i ansökningen i tjänsten har du tre månader på dig att styrka din identitet.
Boka en tid vid Migrationsverkets tjänsteställe på Migrationsverkets webbplats.
När du besöker tjänstestället för att styrka din identitet ska du ta med dig ditt identitetsbevis och ansökningsbilagorna i original.
Om du även ansöker om medborgarskap för ditt barn ska barnet följa med till tjänstestället för att styrka sin identitet.
När du fyllt i ansökningen, kom ihåg att följa ditt konto i Enter Finland-tjänsten.
Om Migrationsverket behöver ytterligare utredningar av dig, meddelas detta i Enter Finland-tjänsten.
Ansökningen kan avslås om du inte lämnar in begärda utredningar i tid.
När ett beslut har fattats får du ett meddelande.
Om du inte kan ansöka om medborgarskap elektroniskt eller inte vet hur man gör det kan du även ansöka om medborgarskap med en pappersblankett.
Skriv ut blanketten på Migrationsverkets webbplats och fyll i den färdigt.
Lämna den ifyllda ansökningen och ansökningsbilagorna personligen till Migrationsverkets tjänsteställe.
Mer information om medborgarskapsansökan och om annat som rör medborgarskap får du på Migrationsverkets webbplats.
Finskt medborgarskap är inte samma sak som uppehållstillstånd.
Om du först planerar att flytta till Finland, läs mer på InfoFinlands sida Flytta till Finland.
Att ansöka om finskt medborgarskapfinska _ svenska _ engelska
Barnets medborgarskapfinska _ svenska _ engelska
Medborgarskapsansökanfinska _ svenska _ engelska
Elektroniska tjänsterfinska _ svenska _ engelska
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Allmänt om fackförbund
I Finland tryggar lagen arbetstagarnas rätt att höra till ett fackförbund (ammattiliitto).
Denna rätt kan inte begränsas med avtal.
Diskriminering av arbetstagare på grund av deras medlemskap i fackförbund är straffbart.
De flesta finländare är med i något fackförbund.
Fackförbunden strävar efter att trygga sina medlemmars intressen och rättigheter, försöker förbättra lönerna och anställningsskyddet samt förbättra arbetslivets kvalitet.
Arbetstagarförbunden är organiserade under tre centralförbund för löntagare.
Dessa är Finlands Fackförbunds Centralorganisation FFC, Tjänstemannacentralorganisationen STTK och Centralorganisationen för högutbildade i Finland Akava.
linkkiFCC, STTK och AKAVA:
Fackets ABC-bokfinska _ engelska _ ryska _ estniska
linkkiCentralorganisationen för högutbildade i Finland Akava:
Information om fackförbundsverksamhetfinska _ svenska _ engelska _ ryska _ estniska _ franska
Information om fackförbundsverksamhetfinska _ svenska _ engelska
linkkiTjänstemannacentralorganisationen STTK:
Information om fackförbundsverksamhetfinska _ svenska _ engelska
Att ansluta sig till ett fackförbund och medlemsavgiften
Om du vill kan du ansluta dig till fackförbundet i din egen bransch.
Du kan ansluta dig till ett fackförbund genom att ta kontakt med förtroendemannen på din egen arbetsplats eller genom att kontakta fackförbundet direkt.
Till de flesta fackförbund kan man också ansluta sig genom att fylla i en anslutningsblankett på fackets webbplats.
Fackförbundets medlemmar betalar förbundet en medlemsavgift som vanligen är cirka 1–2 procent av lönen.
Medlemsavgiften får dras av i beskattningen.
Fackförbundets medlemmar kan delta i utbildning och fritidsaktiviteter som förbundet ordnar.
De får också stöd av förbundets förtroendeman vid konflikter på arbetsplatsen.
Vid behov får man också råd eller förhandlingsstöd från fackförbundet.
Arbetslöshetskassa
I Finland finns ett frivilligt system med arbetslöshetskassor.
En arbetstagare som är medlem i en arbetslöshetskassa betalar en medlemsavgift till arbetslöshetskassan när han eller hon förvärvsarbetar.
Om arbetet upphör och arbetstagaren blir arbetslös kan han eller hon ansöka om inkomstrelaterad arbetslöshetsdagpenning från kassan.
Det lönar sig att ansluta sig till en arbetslöshetskassa, eftersom den inkomstrelaterade dagpenningen är större än det vanliga utkomstskyddet för arbetslösa.
När du ansluter dig till ett fackförbund kan du samtidigt ansluta dig till förbundets arbetslöshetskassa.
Fackförbundet och arbetslöshetskassan är dock två separata system.
Det finns också arbetslöshetskassor som man kan ansluta sig till utan att vara medlem i något fackförbund.
För att få inkomstrelaterad dagpenning finns några villkor som måste uppfyllas innan det är möjligt att få dagpenning.
Till exempel ska man ha varit med i arbetslöshetskassan en viss tid före man blir arbetslös.
Ta reda på dessa villkor genast när du ansluter dig till arbetslöshetskassan.
Läs mer på InfoFinlands sida Utkomstskydd för arbetslösa.
linkkiArbetslöshetskassornas samorganisation:
information om arbetslöshetskassorfinska _ svenska _ engelska
Fackförbundets representant på arbetsplatsen
På arbetsplatsen representeras fackförbundet och de anställda som är medlemmar i det av förtroendemannen.
Förtroendemannen väljs av de anställda.
Förtroendemannen agerar som förhandlare, medlare och informationsförmedlare mellan arbetsgivaren och anställda.
Man kan också vända sig till förtroendemannen till exempel med frågor om kollektivavtalet.
Anmäl flyttningen till myndigheterna
När du flyttar utomlands från Finland ska du göra en flyttanmälan till magistraten (maistraatti)
Du kan göra flyttanmälan på internet eller med en blankett som du får i magistraten eller på posten.
Om du flyttar permanent från Finland eller vistas utomlands två år utan avbrott återkallas ditt uppehållstillstånd.
Du kan ställa Migrationsverket (Maahanmuuttovirasto) en ansökan om att inte återkalla ditt uppehållstillstånd.
Ansökan ska göras innan du har vistats utomlands över två år.
Mer information om detta hittar du på InfoFinlands sida Kan jag förlora mitt uppehållstillstånd?.
Flytt utomlands och den sociala tryggheten
När du flyttar utomlands måste du meddela detta till FPA, om du får FPA:s förmåner eller om du har det europeiska sjukvårdskortet.
Om du får FPA:s förmåner har du vanligtvis rätt till dem även i fortsättningen om din utlandsvistelse varar sex månader eller mindre.
Då anses din utlandsvistelse vara tillfällig och du behöver inte nödvändigtvis anmäla den till FPA.
En utlandsvistelse som varar 3–6 månader bör du anmäla den till FPA, om
du får det allmänna bostadsbidraget
du får stöd för hemvård av barn eller
om du måste köpa receptbelagda läkemedel på apoteket för över tre månaders tid.
Om du ska arbeta i ett EU-/EES-land omfattas du av den sociala tryggheten i arbetslandet under den tid då du arbetar i landet, även om arbetet pågår mindre än sex månader.
Då har du inte rätt till FPA:s förmåner.
Om du flyttar utomlands för över sex månader anses din flytt vara permanent.
Din rätt till FPA:s förmåner upphör då samma dag som du flyttar.
I vissa situationer kan du behålla din rätt till FPA:s förmåner även om du vistas utomlands längre än sex månader.
När du är utomlands och har rätt till FPA:s förmåner ska du alltid anmäla ändringar i dina förhållanden till FPA.
Till exempel ändrade familjeförhållanden eller att du börjar arbeta kan påverka din rätt till FPA:s förmåner.
Du hittar mer information om den sociala tryggheten i Finland på FPA:s webbplats och på InfoFinlands sida Den sociala tryggheten i Finland.
Frivillig återflyttning av flyktingar, asylsökande och emigranter
Om du vill återvända till ditt hemland kan du i vissa fall få stöd för frivilligt återvändande.
Stödet består antingen av pengar eller tjänster.
Penningsummans storlek beror på vilket land du återvänder till.
Tjänsten kan till exempel vara att du får hjälp med att leta efter en bostad eller arbetsplats i det land dit du återvänder.
Du kan få stöd om:
du är asylsökande och handläggningen av din ansökan är oavslutad
du har fått ett negativt beslut på din asylansökan
du är ett offer för människohandel och du inte har en hemkommun i Finland
du har ett tillfälligt uppehållstillstånd på grund av hinder för avlägsnande ur landet
du har fått tillfälligt skydd
din flyktingstatus i Finland har upphört eller återkallats eller det har fattats beslut om att avvisa dig.
Om du är kund hos en mottagningscentral kan du ansöka om stöd för frivilligt återvändande vid din egen mottagningscentral.
Om du inte är kund hos en mottagningscentral kan du ansöka om stöd hos Migrationsverket.
Flyttanmälanfinska _ svenska _ engelska
Återkallelse av uppehållstillståndfinska _ svenska _ engelska
Flytt utomlands och social trygghetfinska _ svenska _ engelska
Frivillig återflyttningfinska _ svenska _ engelska
Du kan få finskt medborgarskap
om du har en förälder som är finsk medborgare,
genom ansökan eller anmälan om medborgarskap.
I vissa undantagsfall kan man dessutom få medborgarskap på grundval av att man är född i Finland.
Ansöka om medborgarskap
Du kan ansöka om finskt medborgarskap när du har fyllt 18 år, har bott permanent i Finland i tillräckligt många år, har nöjaktiga muntliga och skriftliga kunskaper i finska eller svenska eller motsvarande kunskaper i finskt eller finlandssvenskt teckenspråk och din identitet är tillförlitligt utredd.
Det finns också andra villkor; till exempel måste du kunna visa hur du försörjer dig.
Du kan samtidigt ansöka om medborgarskap för ett minderårigt barn som du har vårdnaden om.
Om du har begått ett brott eller till exempel inte har betalat dina skatter, kan detta utgöra ett hinder för att få finskt medborgarskap.
Läs mer på InfoFinlands sida Hur kan man ansöka om finskt medborgarskap?
Finskt medborgarskap är inte samma sak som uppehållstillstånd.
Om du först planerar att flytta till Finland, läs mer på InfoFinlands sida Flytta till Finland.
Finskt medborgarskapfinska _ svenska _ engelska
Barnets medborgarskap
Samtidigt som du ansöker om medborgarskap för dig själv, kan du ansöka om det för ett minderårigt barn som du har vårdnaden om.
Läs mer på InfoFinlands sida Hur kan man ansöka om finskt medborgarskap?
Ett ofött barns medborgarskap
Barnet får automatiskt finskt medborgarskap vid födseln i följande fall:
Barnets mor är finsk medborgare.
Barnets far är finsk medborgare, men modern är inte det och föräldrarna är gifta med varandra.
Om föräldrarna inte är gifta, får barnet finskt medborgarskap av sin far enligt följande:
Vid födseln, då barnet föds i Finland och faderskapet bekräftas.
Genom medborgarskapsanmälan, då barnet föds i något annat land och faderskapet har bekräftats.
Också ett barn till utländska föräldrar som föds i Finland kan få finskt medborgarskap, om hen inte får medborgarskap i något annat land av sina föräldrar.
På InfoFinlands sida När ett barn föds i Finland finns mer information för föräldrar vars barn föds i Finland.
Barnets medborgarskapfinska _ svenska _ engelska
Finskt medborgarskap genom anmälan
Du kan få finskt medborgarskap genom medborgarskapsanmälan (kansalaisuusilmoitus) om du är
en före detta finska medborgare
utlänning och din far är finsk medborgare,
18–22 år och har bott i Finland i flera år
12–17 år och adoptivbarn till en finsk medborgare
medborgare i ett nordiskt land och har varit bosatt i Finland de senaste fem åren
Du kan göra en anmälan om medborgarskap på internet.
Fyll i blanketten i Enter Finland-tjänsten.
Lägg till bilagorna till ansökningen.
Betala samtidigt också ansökningens handläggningsavgift.
När du fyllt i anmälan, kom ihåg att följa ditt konto i tjänsten Enter Finland.
Du har tre månader på dig att styrka din identitet efter att du fyllt i blanketten i Enter Finland-tjänsten.
Du kan styrka din identitet vid Migrationsverkets tjänsteställe eller utomlands vid Finlands beskickning.
Fråga utrikesministeriet vilken beskickning du kan besöka för att styrka din identitet.
Boka en tid i förväg.
Ta med dig ett identitetsbevis och ansökningsbilagorna i original.
Om du inte kan göra din ansökan elektroniskt eller inte vet hur man gör det kan du också lämna in anmälan på en pappersblankett.
Mer information om hur du gör medborgarskapsanmälan hittar du på Migrationsverkets webbplats.
Medborgarskapsanmälanfinska _ svenska _ engelska
Flerfaldigt medborgarskap
Finland godkänner flerfaldigt medborgarskap, d.v.s. att du utöver ditt finska medborgarskap även har medborgarskap i ett annat land.
Alla stater godkänner dock inte flerfaldigt medborgarskap.
Innan du ansöker om finskt medborgarskap är det bra att ta reda på om flerfaldigt medborgarskap också är tillåtet i det land där du är medborgare.
Om denna stat inte tillåter flerfaldigt medborgarskap kan du förlora ditt nuvarande medborgarskap när du får finskt medborgarskap.
Flerfaldigt medborgarskap kan vara en fördel, men också en nackdel.
Det lönar sig att till exempel ta reda på om man tvingas göra värnplikten i flera medborgarskapsstater eller om det räcker med ett intyg över fullgjord värnplikt i ett land.
Flerfaldigt medborgarskap kan vara en fördel när man till exempel flyttar från ett land till ett annat.
Migrationsverket ger råd i frågor som rör medborgarskap:
Telefon 0295 419 626 tisdag, onsdag och fredag kl. 10.00–11.00
Barnets flerfaldiga medborgarskap
Barnet kan ha finskt medborgarskap och medborgarskap i något annat land.
Detta beror på huruvida det andra landet godkänner flerfaldigt medborgarskap för barnet.
Fråga mer om detta vid beskickningen för ditt eget land.
Kan man förlora sitt finska medborgarskap?
Man kan förlora sitt finska medborgarskap om man
är 22 år gammal, har medborgarskap också i en annan stat och saknar tillräcklig anknytning till Finland
har angett felaktiga uppgifter i medborgarskapsansökan eller medborgarskapsanmälan
har förvärvat sitt medborgarskap på grund av faderns finska medborgarskap och faderskapet upphävs.
Att förlora sitt finska medborgarskapfinska _ svenska _ engelska
Arbetsavtalet upprättas i två exemplar, ett till den anställda och ett till arbetsgivaren.
Arbetsavtalet innehåller vanligen åtminstone följande punkter:
Parterna som ingår arbetsavtalet
Både arbetsgivaren och den anställda undertecknar arbetsavtalet.
Tidpunkten då arbetet inletts
Om avtalet är tillsvidare gällande eller tidsbundet
Huvudregeln är att arbetsavtalet gäller tillsvidare.
Detta innebär att arbetet pågår tills den anställda säger upp sig eller tills arbetsgivaren säger upp den anställda.
Arbetsgivaren ska ha en välgrundad orsak för att säga upp en anställd.
Godtagbara orsaker för uppsägning definieras i arbetsavtalslagen.
När arbetsavtalet gäller tillsvidare har arbetstagaren en fast eller permanent anställning.
Ett tidsbundet avtal innebär att man har avtalat om tidpunkten då arbetet inleds och avslutas.
Arbetsavtalet kan vara tidsbundet om det finns en välgrundad orsak till detta.
Lagar och kollektivavtal reglerar exakt när tidsbundna anställningar får tillämpas.
En anställning kan vara tidsbunden om orsaken är till exempel
vikariat
praktik projekt
efterfrågan eller säsongtopp
Om arbetsavtalet är tidsbundet binder det båda parterna en bestämd tid, om man inte har kommit överens om möjligheten till uppsägning.
Ett tidsbundet avtal kan hävas endast av mycket vägande skäl.
Prövotid och längden på den
Man kan komma överens om en prövotid i anställningens början.
Prövotiden kan vara högst sex månader.
Vid en tidsbunden anställning kan prövotiden vara högst hälften av den tid anställningen pågår.
Under prövotiden kan arbetstagaren bedöma om arbetet lämpar sig för honom eller henne och arbetsgivaren kan bedöma om arbetstagaren är lämplig för arbetet.
Under prövotiden kan arbetstagaren och arbetsgivaren häva arbetsavtalet utan uppsägningstid.
Grunderna för hävande av ett arbetsavtal under prövotiden får inte vara diskriminerande.
Arbetstagaren får normal lön under prövotiden.
Platsen för utförandet av arbetet
Arbetsuppgifterna
Lönen och utbetalning av lönen
Lönen bestäms enligt kollektivavtalet.
Om branschen inte har ett kollektivavtal har arbetstagaren rätt till en skälig lön.
Arbetsgivaren får inte betala en lön som är mindre än vad som fastställs i kollektivavtalet.
Lönen kan innehålla olika förmåner.
Typiska lönetillägg i Finland är erfarenhetstillägg, övertidstillägg och skiftarbetstillägg.
Avlöningsdagen är vanligen en eller två gånger i månaden.
Arbetsgivaren betalar in lönen på bankkontot.
Arbetstagaren har rätt att få en lönespecifikation där det står vad lönen består av.
När man talar om lön avser man oftast bruttolönen (bruttopalkka) från vilken skatter och personalbikostnader dras av.
Den lön som betalas till arbetstagaren är nettolönen (nettopalkka).
Arbetstid
I avtalet ska den regelbundna arbetstiden nedtecknas.
Arbetstiden ska följa arbetslagstiftningen och kollektivavtalet.
Semester och semesterpenning
Arbetstagaren har rätt att få samma lön under semestern som under arbetet.
Dessutom betalas en semesterpenning.
Utbetalningen av semesterpenning baserar sig på kollektivavtalet.
När anställningen upphör har arbetstagaren rätt att få semesterersättning för de dagar som han eller hon inte har fått semester eller semesterersättning för vid tidpunkten för anställningens upphörande.
Uppsägningstid
Ett tillsvidare gällande arbetsavtal upphör antingen när arbetstagarens eller arbetsgivarens uppsägningstid har gått ut.
Uppsägningstiden är den tid som arbetstagaren är skyldig att arbeta innan arbetet upphör.
Under uppsägningstiden har arbetstagaren samma rättigheter och skyldigheter och han eller hon får normal lön.
Om arbetsgivaren säger upp en arbetstagare måste arbetsgivaren ange orsaken till detta.
Arbetsavtalslagen beskriver vilka orsaker som är godtagbara för uppsägning.
Omnämnande om viket kollektivavtal arbetsavtalet följer
linkkiArbets- och näringsministeriet:
Arbetsavtal och anställningfinska _ svenska _ engelska
Många länder har en beskickning i Finland.
Beskickningen kan antingen vara en ambassad eller ett konsulat.
Ambassaderna finns i Helsingfors.
Vissa länder har också konsulat i andra städer.
Om du behöver sköta ett ärende med myndigheterna i ditt hemland ska du ta kontakt med ditt lands beskickning.
Via beskickningen kan du ofta uträtta till exempel följande ärenden:
Få en födelseattest
Ansöka om medborgarskap i ditt hemland om du har förlorat det eller avstått från det
Anmäla födelsen av ditt barn till myndigheterna i ditt hemland om barnet föds i Finland
Ansöka om medborgarskap i ditt hemland för ditt barn om barnet har fötts i Finland
Registrera ett äktenskap i ditt hemland om du har gift dig i Finland
Rösta i val i ditt hemland
Observera att alla beskickningar inte erbjuder samma tjänster.
Det är inte nödvändigtvis möjligt att sköta alla ovannämnda ärenden i alla beskickningar.
Vilka tjänster ditt lands beskickning tillhandahåller beror på lagen i ditt hemland.
Mer information får du från ditt hemlands beskickning.
Alla länder har inte en beskickning i Finland.
I detta fall betjänas du ofta av ditt hemlands beskickning i något av Finlands grannländer.
På det finska utrikesministeriets webbplats finns en förteckning över andra länders beskickningar i Finland.
Där hittar du även kontaktuppgifterna till beskickningarna.
Andra länders beskickningar i Finlandfinska _ svenska _ engelska
På den här sidan finns information om den bosättningsbaserade sociala tryggheten som hör till FPA:s ansvarsområde.
På sidan finns information om de situationer då du betraktas ha rätt till den sociala trygghet som grundar sig på boende.
På InfoFinlands sida Utkomstskydd för arbetslösa får du mer information om vem som har rätt till utkomstskydd för arbetslösa.
FPA har bland annat hand om folkpensionen, barnbidrag, det grundläggande utkomstskyddet för arbetslösa, sjuk- och föräldradagpenningar, utkomststöd och rehabilitering.
FPA sköter även de sjukvårdsersättningar som betalas för privat sjukvård.
Om du är sjukförsäkrad i Finland, får du ett FPA-kort.
Grunderna för FPA:s bidrag definieras i lagen.
När du ansöker om en förmån, utreder FPA om du har rätt till FPA:s förmåner.
På detta inverkar ditt stadigvarande boende och arbete i Finland.
Varje sökandes livssituation behandlas individuellt när FPA fattar beslut om bidrag.
Sökandens livssituation och behov av understöd är ofta mycket olika.
Därför varierar även bidragens belopp och grunder.
Du ska alltid utreda din egen situation individuellt.
Offentliga hälso- och sjukvårdstjänster samt socialtjänster är kommunernas ansvar i Finland.
Läs mer på InfoFinlands sida Hälsovårdstjänster i Finland.
Mer information om rätten till hemkommun finns på InfoFinlands sida Hemkommun i Finland.
Information om social trygghetfinska _ svenska _ engelska
Social trygghet för dig som flyttar till Finland(pdf, 560 kb)finska _ svenska _ engelska _ ryska _ estniska
Information om sjukförsäkringfinska _ svenska _ engelska
linkkiSocial- och hälsovårdsministeriet:
Information om den sociala tryggheten i Finlandfinska _ svenska _ engelska
Rätten till FPA:s förmåner
Huvudregeln är att om du bor stadigvarande i Finland, kan du få FPA:s förmåner.
Vad stadigvarande boende betyder definieras i lagen.
Du kan också få rätt till FPA:s förmåner genom att arbeta i Finland.
Har du rätt till förmåner?
På detta inverkar om du flyttar till Finland från
ett land inom Europeiska unionen (EU), ett land inom det Europeiska ekonomiska samarbetsområdet (EES) eller Schweiz eller
från något annat land.
EES-länderna är Europeiska unionens medlemsländer samt Norge, Island och Liechtenstein.
Huruvida du får förmåner påverkas dessutom av om du flyttar till Finland till exempel som
arbetstagare eller företagare
studerande
familjemedlem
utsänd arbetstagare.
Finland har ingått avtal om den sociala tryggheten med ett antal länder.
Dessa länder är de nordiska länderna, USA, Kanada och Quebec, Chile, Israel, Indien, Kina, Sydkorea och Australien.
Avtalen rör främst pensioner.
En del avtal gäller även sjukvård.
Om du kommer från ett av dessa länder ska du kontrollera hos FPA om avtalen påverkar din sociala trygghet.
Lag om hemkommunfinska _ svenska
Information om internationella socialskyddsavtalfinska _ svenska _ engelska
Information om den sociala tryggheten i Finland för EU-medborgarefinska _ svenska _ engelska
Stadigvarande flytt till Finland och stadigvarande boende i Finland
När du flyttar till Finland bedömer FPA alltid först om din flytt till Finland är stadigvarande boende i den mening som avses i lagstiftningen om social trygghet.
Om din flytt till Finland inte anses vara stadigvarande, kan du ändå ha rätt till FPA:s förmåner på grund av att du arbetar.
Din flytt till Finland kan betraktas som stadigvarande i följande situationer:
du är återflyttare, det vill säga återvänder till Finland från utlandet
du har en fast anställning eller motsvarande avtal för ett arbete som du utför i Finland
du är gift eller annars i ett nära familjeförhållande till en person som redan bor stadigvarande i Finland.
Dessutom krävs det i allmänhet att ditt uppehållstillstånd är giltigt, om du är skyldig att ha ett uppehållstillstånd.
Din situation bedöms i sin helhet.
På basis av bedömningen beslutas om boendet är stadigvarande eller inte.
Om du flyttar till Finland tillfälligt har du vanligtvis inte rätt till FPA:s förmåner.
Från och med den 1 april 2019 kan studerande från länder utanför EU och EES ha rätt till vissa förmåner, till exempel förmåner som ingår i sjukförsäkringen.
När det finns ett avgörande om att ditt boende i Finland är stadigvarande, anses du bo stadigvarande i Finland så länge som
du har din egentliga bostad och ditt hem här och så länge du huvudsakligen vistas här
eller
du har en annan grund för den stadigvarande vistelsen, till exempel ett familjeband eller arbete.
Om du emellertid börjar arbeta i ett annat land eller reser utomlands för över sex månader, kan din rätt till FPA:s förmåner upphöra.
Mer information om sådana situationer får du vid FPA.
Det finns även bidrag som du inte kan få om du inte bor stadigvarande i Finland eller har gjort det tidigare.
Till exempel kan föräldrar få föräldradagpenning endast om de har bott i Finland minst 180 dagar före barnets beräknade förlossningsdatum.
Om du kommer från ett annat EU-land kan du i vissa fall utnyttja de försäkringsperioder som du har ackumulerat i andra EU-länder.
Fråga mer hos FPA:s center för internationella ärenden.
tfn 020 634 0200
kl. 9–16
Social trygghet för dig som flyttar till Finlandfinska _ svenska _ engelska
Flytt utomlands och social trygghetfinska _ svenska _ engelska
Kontaktuppgifter till FPAfinska _ svenska _ engelska
Arbete ger dig åtminstone delvis rätt till den sociala tryggheten i Finland
EU-länderna, EES-länderna och Schweiz
Om du flyttar till Finland för att arbeta får du vanligtvis rätt till FPA:s förmåner under din anställning, även när din anställning är kortvarig.
Om din lön uppgår till minst 696,60 € i månaden är du berättigad till de flesta av FPA:s förmåner.
Hur många timmar per vecka du arbetar eller hur lång din anställning är spelar ingen roll.
Arbetstagaren och den sociala tryggheten i Finlandfinska _ svenska _ engelska
Asylsökande
Asylsökande har inte rätt till finskt socialskydd.
Detta innebär att de inte har rätt till FPA:s förmåner.
Mottagningscentralen betalar mottagningspenning till asylsökande.
Den utbetalas så länge som asylansökan behandlas.
Mottagningspenningen är ett litet belopp som är avsett för ofrånkomliga utgifter.
Om den asylsökande beviljas uppehållstillstånd och är fast bosatt i Finland har han eller hon rätt till finskt socialskydd.
Man kan ansöka om att omfattas av det finska socialskyddet av FPA då uppehållstillstånd har beviljats.
I Finland bestäms arbetstagarnas rättigheter enligt arbetslagstiftningen och kollektivavtalen (työehtosopimukset).
I dessa fastställs till exempel minimilöner, arbetstider, semestrar, lön för sjukdomstid och uppsägningsvillkor.
Arbetsgivarförbundet och arbetstagarförbundet kommer gemensamt överens om anställningsvillkoren i en viss bransch.
På detta sätt uppstår ett kollektivavtal för branschen.
I den offentliga sektorn (arbetsgivaren är en kommun eller staten) ingås tjänstekollektivavtal eller allmänt kommunalt tjänste- och arbetskollektivavtal.
Förmånerna som man har avtalat om med ett kollektivavtal är alltid minimiförmåner.
Dessa kan inte underskridas i arbetsavtalet.
Lönen kan till exempel inte vara lägre än vad som avtalats med kollektivavtalet.
Arbetsgivaren och arbetstagaren kan ändå i arbetsavtalet komma överens om villkor som är bättre än villkoren i kollektivavtalet.
Kollektivavtalen uppgörs för en viss tid, vanligen för ett eller två år eller också för en längre tid.
Kollektiv- och tjänstekollektivavtalet är bindande för de löntagar- och arbetsgivarförbund som slutit dem och för deras medlemmar.
Ett kollektivavtal kan också vara allmänt bindande.
Då måste även de arbetsgivare som inte hör till arbetsgivarförbundet följa avtalet med sina anställda.
I platsannonser och arbetsavtal kan det stå: ”palkkaus TES:in mukainen” (”avlöning enligt kollektivavtalet”).
Det är bra att ta reda på hur stora lönerna är i den egna branschen i Finland.
Det är viktigt att känna till kollektivavtalet, eftersom det i Finland inte finns till exempel en lag om minimilöner, utan minimilönerna fastställs alltid enligt kollektivavtalet.
linkkiArbets- och näringsministeriet:
Arbetslagstiftningfinska _ svenska _ engelska
Arbetsavtal
Arbetsgivaren ingår vanligen ett skriftligt arbetsavtal med en ny anställd.
I arbetsavtalet fastställs arbetsuppgifterna och lönen samt andra förmåner och villkor.
Avtalet kan också vara muntligt.
Om man inte har uppgjort ett skriftligt arbetsavtal ska arbetsgivaren utan särskild begäran ge en skriftlig redogörelse för de centrala villkoren i arbetet.
Det är rekommendabelt att arbetsavtalet är skriftligt.
När allt finns på papper kan både den anställda och arbetsgivaren kontrollera i avtalet vad man gemensamt har avtalat.
Detta hjälper om det uppstår konflikter i arbetet.
Läs mer om upprättandet av arbetsavtalet på InfoFinlands sida Innehållet i arbetsavtalet.
linkkiArbetarskyddsförvaltningen:
Att uppgöra ett arbetsavtalfinska _ svenska _ engelska
Ett skriftligt avtal om de centrala villkoren i arbetet
Arbetsgivaren ska ge den anställda en skriftlig redogörelse för de centrala villkoren i arbetet vid tillsvidare gällande anställningar samt anställningar som varar över en månad.
Av redogörelsen ska det åtminstone framgå
arbetsgivarens och arbetstagarens hemort eller driftställe
tidpunkten då arbetet inletts
längden på ett tidsbundet arbetsavtal och orsaken till att avtalet är tidsbundet
prövotidens längd
stället där arbetet utförs
den anställdas arbetsuppgifter
kollektivavtalet som tillämpas på arbetet
de grunder enligt vilka lön eller andra vederlag bestäms samt löneperioden
den regelbundna arbetstiden
hur semestern bestäms
uppsägningstiden eller grunden för bestämmande av den
Om arbetsgivaren inte ger en redogörelse för de centrala villkoren i arbetet till den anställda kan han eller hon dömas till böter.
Finska medborgare har vissa rättigheter och skyldigheter som utlänningar bosatta i Finland inte nödvändigtvis har.
Rättigheter
rätt att få finskt pass
rätt att resa till Finland och vägra att bli utlämnad till ett annat land
rätt att rösta i presidentval, riksdagsval och folkomröstningar då man fyllt 18 år.
rätt att ställa upp som kandidat i riksdagsval då man fyllt 18 år.
möjlighet att bli utnämnd till sådana statliga ämbeten för vilka det krävs finskt medborgarskap
EU-medborgarnas rättigheter som rätten att fritt röra sig och arbeta inom EU:s område och rätten att rösta och ställa upp som kandidat i EU-val
Skyldigheter
Skyldighet att delta i landets försvar eller bistå i det.
Män som har fyllt 18 år har värnplikt (asevelvollisuus).
Skyldighet att följa Finlands lagar även annanstans än i Finland.
Finska medborgare kan i Finland dömas för brott som begåtts utomlands.
Observera att dessa är rättigheter och skyldigheter som ingår i det finska medborgarskapet.
Information om rättigheter och skyldigheter som gäller alla som är bosatta i Finland finns på InfoFinlands sida Dina rättigheter och skyldigheter i Finland.
Finska medborgares rättigheter och skyldigheterfinska _ svenska _ engelska
linkkiFörsvarsmakten:
Värnpliktfinska _ svenska _ engelska
Att ansöka om finskt passfinska _ svenska _ engelska
Att ansöka om finskt pass utomlandsfinska _ svenska _ engelska
Utlänningar som bor i Finland har nästan samma rättigheter och skyldigheter som finländarna.
Följande rättigheter och skyldigheter gäller även utlänningar som bor i Finland.
Rättigheter
Alla har rätt till likabehandling.
Ingen får särbehandlas till exempel på grund av kön, ålder, religion eller handikapp.
Var och en får fritt yttra sina åsikter i tal och skrift.
Människor får ordna möten och demonstrationer och delta i dem.
Demonstrationer ska anmälas till polisen på förhand.
Ingen får dömas till döden eller torteras.
Alla får själva välja sin bostadsort och röra sig fritt i Finland.
Alla har rätt till integritetsskydd.
Ett brev som tillhör en annan person får inte läsas och en annan persons telefonsamtal får inte avlyssnas.
Var och en får själv välja sin egen religion.
Om man inte vill behöver man inte välja någon religion alls.
Utlänningar som bor stadigvarande i Finland och som har fyllt 18 år har rätt att rösta i kommunalval.
Utlänningar som har rösträtt i kommunalval har även rätt att ställa upp som kandidat i kommunalval.
EU-medborgare som har hemort i Finland kan rösta i Europaparlamentsvalet om de har anmält sig till rösträttsregistret (äänioikeusrekisteri).
EU-medborgare som är i det finska rösträttsregistret kan också ställa upp som kandidat i Finlands Europaparlamentsval.
Läs mer om utlänningars rösträtt i Finland på InfoFinlands sida Val i Finland.
Skyldigheter
Alla som bor eller vistas i Finland måste följa Finlands lagar.
7–17-åringar har läroplikt (oppivelvollisuus), d.v.s. skyldighet att avlägga grundskolans (peruskoulu) lärokurs.
Ofta måste de som arbetar i Finland betalar skatt på sin lön i Finland.
Alla har skyldighet att vittna inför domstol om de blir kallade.
Föräldrar är skyldiga att ta hand om sina barn.
Alla har skyldighet att hjälpa vid en olycka.
Läs mer om beskattningen på InfoFinlands sida Beskattning.
Finska medborgares rättigheter och skyldigheter
Finska medborgare har utöver de ovannämnda också några ytterligare rättigheter och skyldigheter som utlänningar bosatta i Finland inte har.
Läs mer om finska medborgarnas rättigheter och skyldigheter på InfoFinlands sida Finskt medborgarskap.
Finlands grundlagfinska _ svenska _ engelska
Information om demokratin i Finlandfinska _ svenska _ engelska
Val i Finlandfinska _ svenska _ engelska
Jämlikheten är nedtecknad i lagar
Finlands grundlag garanterar jämlikt bemötande för alla.
Jämlikhet (yhdenvertaisuus) betyder att alla människor är likvärdiga oberoende av kön, ålder, etnisk eller nationell härkomst, nationalitet, språk, religion och övertygelse, åsikt, handikapp, hälsotillstånd, sexuell läggning eller någon annan orsak som gäller hans eller hennes person.
Om jämlikhet i arbetslivet föreskrivs i lagen om likabehandling och i arbetsavtalslagen.
Enligt dessa ska anställda behandlas lika när det gäller anställning, arbetsförhållanden, anställningsvillkor, utbildning för personalen och avancemang i karriären.
Finlands grundlagfinska _ svenska _ engelska _ ryska _ franska _ spanska _ tyska
Lag om likabehandlingfinska _ svenska _ engelska
Jämlikhet i rekryteringen
Lagen om likabehandling (yhdenvertaisuuslaki) förutsätter att alla arbetssökande behandlas lika.
Arbetsgivaren ska välja den sökande som har de bästa meriterna för uppgiften.
Arbetsgivaren ska också kunna bevisa att det finns godtagbara grunder för valet som anknyter till arbetets karaktär och att valet inte har varit diskriminerande.
Man får inte kräva sådana egenskaper av arbetssökanden som inte är nödvändiga i utförandet av arbetet.
Jämlikhet på arbetsplatsen
Arbetsgivaren får inte diskriminera de anställda när han eller hon fattar beslut om fördelning av arbetsuppgifter, erbjudande av möjligheter till avancemang eller upphävande av anställningen.
Arbetsdiskriminering är ett brott.
Om du misstänker att du har fallit offer för arbetsdiskriminering kan du ta kontakt med arbetarskyddsmyndigheterna eller ditt eget fackförbund.
Vid problem kan du fråga råd hos arbetarskyddsfullmäktige eller förtroendemannen.
linkkiArbetarskyddsförvaltningen:
Arbetarskyddfinska _ svenska _ engelska
linkkiRegionförvaltningsverket:
Arbetarskyddfinska _ svenska _ engelska
linkkiArbets- och näringsministeriet:
Likabehandling och förebyggande av diskriminering på arbetsplatserfinska _ svenska _ engelska
Jämställdhet (tasa-arvo) mellan könen
Enligt Finlands lag är män och kvinnor jämställda.
Män och kvinnor ska behandlas lika vid anställning och beträffande arbetsförhållanden och lönesättning.
En anställd får inte särbehandlas i arbetslivet på grund av graviditet eller föräldraskap.
I Finland finns en lag om likabehandling, som föreskriver att arbetsgivaren ska övervaka att jämställdheten på arbetsplatsen realiseras och att ingen diskrimineras på arbetsplatsen.
Jämställdhetsombudsmannen övervakar att lagen om likabehandling av män och kvinnor följs.
Om du misstänker att din arbetsgivare har diskriminerat dig på grund av ditt kön kan du be jämställdhetsombudsmannen om råd och anvisningar samt hjälp med att reda ut saken.
linkkiJämställdhetsombudsmannens byrå:
Information om jämställdhet i arbetslivetfinska _ svenska _ engelska _ ryska _ samiska
Jämställdhetslagenfinska _ svenska
För att få finskt medborgarskap genom en medborgarskapsansökan krävs något av följande:
Du kan tillförlitligt intyga din identitet.
Du är minst 18 år gammal eller gift.
Du har bott i Finland tillräckligt länge.
Hur lång boendetid som krävs beror på din situation, vanligtvis ska du ha bott här minst 4–7 år.
Du har inte begått brott.
Du har inte lämnat till exempel skatter, böter, underhållsbidrag eller sjukhusavgifter obetalda.
Du kan redogöra för hur du försörjer dig i Finland.
Du kan finska, svenska eller det finska eller finlandssvenska teckenspråket åtminstone nöjaktigt.
Läs mer om att bevisa dina språkkunskaper på InfoFinlands sida Officiellt intyg över språkkunskaper.
Läs mer om att studera finska och svenska på InfoFinlands sida Finska och svenska språket.
Du kan ansöka om medborgarskap elektroniskt i tjänsten Enter Finland.
Fyll i en ansökan och lägg till bilagorna.
För en ansökan behöver du åtminstone följande dokument:
Ett giltigt identitetsbevis
En utredning om dina språkkunskaper
En utredning om ditt uppehälle.
Betala samtidigt också ansökningens handläggningsavgift.
När du fyllt i ansökningen i tjänsten har du tre månader på dig att styrka din identitet.
Boka en tid vid Migrationsverkets tjänsteställe på Migrationsverkets webbplats.
När du besöker tjänstestället för att styrka din identitet ska du ta med dig ditt identitetsbevis och ansökningsbilagorna i original.
Om du även ansöker om medborgarskap för ditt barn ska barnet följa med till tjänstestället för att styrka sin identitet.
När du fyllt i ansökningen, kom ihåg att följa ditt konto i Enter Finland-tjänsten.
Om Migrationsverket behöver ytterligare utredningar av dig, meddelas detta i Enter Finland-tjänsten.
Ansökningen kan avslås om du inte lämnar in begärda utredningar i tid.
När ett beslut har fattats får du ett meddelande.
Om du inte kan ansöka om medborgarskap elektroniskt eller inte vet hur man gör det kan du även ansöka om medborgarskap med en pappersblankett.
Skriv ut blanketten på Migrationsverkets webbplats och fyll i den färdigt.
Lämna den ifyllda ansökningen och ansökningsbilagorna personligen till Migrationsverkets tjänsteställe.
Mer information om medborgarskapsansökan och om annat som rör medborgarskap får du på Migrationsverkets webbplats.
Finskt medborgarskap är inte samma sak som uppehållstillstånd.
Om du först planerar att flytta till Finland, läs mer på InfoFinlands sida Flytta till Finland.
Att ansöka om finskt medborgarskapfinska _ svenska _ engelska
Barnets medborgarskapfinska _ svenska _ engelska
Medborgarskapsansökanfinska _ svenska _ engelska
Elektroniska tjänsterfinska _ svenska _ engelska
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Om du måste sköta ärenden med finländska myndigheter, men inte kan finska eller svenska och det inte heller finns något annat språk som både du och myndigheten talar, kan du i vissa fall ha rätt till tolkning.
Då beställer myndigheten tolken och betalar för tolkningen.
Myndigheten kan ordna och betala tolkningen när det gäller skötsel av ärenden som behandlas på myndighetens initiativ.
Detta är dock inte alltid möjligt.
Om du behöver en tolk för den inledande kartläggningen och integrationsplanen, måste myndigheten beställa en tolk.
Du kan på förhand fråga myndigheten om detta.
Om du söker asyl i Finland har du rätt till tolkning i ärenden som rör behandlingen av din asylansökan.
Du har rätt att få information om ett beslut gällande dig på ditt modersmål eller ett annat språk som du förstår.
Information om beslutet ges genom tolkning eller översättning.
Om du själv bokar tolken och betalar tolkningen, kan du anlita en tolk när som helst.
Tolktjänsterfinska _ svenska _ engelska
Vad gör tolken?
Tolken är med på möten mellan dig och myndigheten.
Han eller hon tolkar det som du och myndigheten säger.
Tolken är antingen på plats eller också kan tolkningen ordnas via telefon eller video.
Tolken har som uppgift att tolka det som du och myndigheten säger.
Tolken sköter inga andra uppgifter utöver tolkningen.
Han eller hon kan således inte hjälpa dig med annat.
Tolken är en neutral, utomstående person som varken är på din eller på myndighetens sida.
Tolken har sekretessplikt och får inte berätta inte om dina angelägenheter för andra.
Var kan man beställa en tolk?
I Finland finns åtta kommunala tolkcentraler (tulkkikeskus).
Tolkcentralernas tjänster är främst avsedda för myndigheter som arbetar med invandrare.
Också många företag erbjuder tolktjänster.
linkkiFinlands översättar- och tolkförbund:
Sök tolk eller översättarefinska _ svenska _ engelska
Kommunala tolkcentraler
Tolkningfinska
linkkiMellersta Finlands tolkcentral:
Tolkningfinska _ svenska _ engelska
Tolkningfinska
Tolkningfinska _ engelska
linkkiÖsterbottens tolkcentral:
Tolkningfinska
linkkiNorra Finlands tolktjänst:
Tolkningfinska
linkkiÅboregionens tolkcentral:
Tolkningfinska _ svenska
Tolkningfinska
I Finland har en arbetstagare rätt:
till lön och övriga minimivillkor enligt kollektivavtalet
till skydd utgående från lagar och avtal
att organisera sig
till en sund och trygg arbetsmiljö.
En arbetstagare är skyldig att
utföra arbetet omsorgsfullt
följa de överenskomna arbetstiderna
följa arbetsledningens anvisningar
vägra att delta i verksamhet som konkurrerar med arbetsgivaren
hålla affärs- och yrkeshemligheter
ta hänsyn till arbetsgivarens intresse.
Anställningsrådgivning för invandrare
Om du har frågor om eller problem med din anställning, kan du kontakta anställningsrådgivningen för invandrare.
Rådgivningen ges av Finlands Fackförbunds Centralorganisation FFC.
Du kan få rådgivning även om du inte är medlem i fackförbundet.
En jurist svarar på dina frågor till exempel om arbetsavtal, lön eller arbetstider.
Den kostnadsfria rådgivningen ges på finska och engelska.
Anställningsrådgivningen har öppet på tisdagar och onsdagar klockan 9–11 och 12–15.
Telefon: 0800 414 004
Du kan även ringa arbetarskyddsmyndigheternas riksomfattande rådgivningstelefon:
Tfn 0295 016 620
Mån.–fre. kl. 9–15
linkkiFFC:
Anställningsrådgivning för invandrarefinska _ svenska _ engelska
linkkiFFC:
Arbetslivet i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ kinesiska _ arabiska
linkkiArbetshälsoinstitutet:
Handboken Jobba i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ kurdiska _ tyska _ thai _ vietnamesiska
linkkiBrottsofferjouren:
Video om arbetstagarens rättigheter i Finlandengelska _ kinesiska _ arabiska _ thai _ hindi
Arbetstagarnas rättigheter tryggas med lagar och avtal
Arbetslagstiftningen och kollektivavtalen föreskriver vilka rättigheter och skyldigheter arbetstagare har.
Arbetstagar- och arbetsgivarförbunden förhandlar gemensamt fram branschspecifika kollektivavtal.
I lagstiftningen och kollektivavtalet fastställs till exempel minimilöner, arbetstider, semestrar, lön för sjukdomstid och uppsägningsvillkor.
Läs mer på InfoFinlands sidor Att komma överens om anställningsvillkoren och Innehållet i arbetsavtalet.
linkkiArbets- och näringsministeriet:
Broschyrer om arbetslagstiftningenfinska _ svenska _ engelska
Jämlikhet
Varje anställd har rätt till ett jämlikt och icke-diskriminerande bemötande när de söker jobb och på arbetsplatsen.
Läs mer på InfoFinlands sida Jämlikhet och jämställdhet i arbetslivet.
Arbetsavtal
Ett arbetsavtal uppstår när arbetstagaren och arbetsgivaren kommer överens om utförandet av ett arbete och lönen som betalas för det samt övriga förmåner och villkor.
Anställningsvillkoren bestäms enligt arbetslagstiftningen och kollektivavtalet.
Arbetsavtalet är bindande för båda parterna.
Läs mer om arbetsavtalet på InfoFinlands sidor Att komma överens om anställningsvillkoren och Innehållet i arbetsavtalet.
Fackförbund
I Finland är facklig organisering vanligt och aktiva fackförbundsmedlemmar trakasseras inte.
Du kan ansluta dig till fackförbundet i din egen bransch.
Förbundet strävar efter att trygga sina medlemmars intressen i arbetslivet.
Läs mer på InfoFinlands sida Fackförbund.
Arbetarskydd
Arbetsgivaren är skyldig att trygga de anställdas säkerhet.
Arbetarskyddsförvaltningen övervakar att de i lagen stadgade arbetarskyddsföreskrifterna följs på arbetsplatserna.
Läs mer på InfoFinlands sida Arbetarskydd.
Utkomstskydd för arbetslösa
När en person som är fast bosatt i Finland blir arbetslös, har han eller hon rätt att få utkomstskydd för arbetslösa.
Läs mer på InfoFinlands sida Utkomstskydd för arbetslösa.
En invandrare som har bott tillräckligt länge i Finland kan få pension på grund av sin ålder eller arbetsoförmögenhet.
Läs mer på InfoFinlands sida Pension.
Beskattning
När du arbetar i Finland måste du betala skatter.
Läs mer på InfoFinlands sida Beskattning.
Företagshälsovård
Varje arbetsgivare är skyldig att ordna förebyggande företagshälsovård för sina anställda.
Läs mer på InfoFinlands sida Företagshälsovård.
Familjeledigheter
När ett barn föds till familjen kan modern eller fadern enligt lag stanna hemma för att ta hand om barnet.
Läs mer på InfoFinlands sida Familjeledigheter.
Arbetsintyg
När en anställning upphör har den anställda rätt att få ett skriftligt arbetsintyg av arbetsgivaren.
Läs mer på InfoFinlands sida Arbetsintyg.
Du kan få finskt medborgarskap
om du har en förälder som är finsk medborgare,
genom ansökan eller anmälan om medborgarskap.
I vissa undantagsfall kan man dessutom få medborgarskap på grundval av att man är född i Finland.
Ansöka om medborgarskap
Du kan ansöka om finskt medborgarskap när du har fyllt 18 år, har bott permanent i Finland i tillräckligt många år, har nöjaktiga muntliga och skriftliga kunskaper i finska eller svenska eller motsvarande kunskaper i finskt eller finlandssvenskt teckenspråk och din identitet är tillförlitligt utredd.
Det finns också andra villkor; till exempel måste du kunna visa hur du försörjer dig.
Du kan samtidigt ansöka om medborgarskap för ett minderårigt barn som du har vårdnaden om.
Om du har begått ett brott eller till exempel inte har betalat dina skatter, kan detta utgöra ett hinder för att få finskt medborgarskap.
Läs mer på InfoFinlands sida Hur kan man ansöka om finskt medborgarskap?
Finskt medborgarskap är inte samma sak som uppehållstillstånd.
Om du först planerar att flytta till Finland, läs mer på InfoFinlands sida Flytta till Finland.
Finskt medborgarskapfinska _ svenska _ engelska
Barnets medborgarskap
Samtidigt som du ansöker om medborgarskap för dig själv, kan du ansöka om det för ett minderårigt barn som du har vårdnaden om.
Läs mer på InfoFinlands sida Hur kan man ansöka om finskt medborgarskap?
Ett ofött barns medborgarskap
Barnet får automatiskt finskt medborgarskap vid födseln i följande fall:
Barnets mor är finsk medborgare.
Barnets far är finsk medborgare, men modern är inte det och föräldrarna är gifta med varandra.
Om föräldrarna inte är gifta, får barnet finskt medborgarskap av sin far enligt följande:
Vid födseln, då barnet föds i Finland och faderskapet bekräftas.
Genom medborgarskapsanmälan, då barnet föds i något annat land och faderskapet har bekräftats.
Också ett barn till utländska föräldrar som föds i Finland kan få finskt medborgarskap, om hen inte får medborgarskap i något annat land av sina föräldrar.
På InfoFinlands sida När ett barn föds i Finland finns mer information för föräldrar vars barn föds i Finland.
Barnets medborgarskapfinska _ svenska _ engelska
Finskt medborgarskap genom anmälan
Du kan få finskt medborgarskap genom medborgarskapsanmälan (kansalaisuusilmoitus) om du är
en före detta finska medborgare
utlänning och din far är finsk medborgare,
18–22 år och har bott i Finland i flera år
12–17 år och adoptivbarn till en finsk medborgare
medborgare i ett nordiskt land och har varit bosatt i Finland de senaste fem åren
Du kan göra en anmälan om medborgarskap på internet.
Fyll i blanketten i Enter Finland-tjänsten.
Lägg till bilagorna till ansökningen.
Betala samtidigt också ansökningens handläggningsavgift.
När du fyllt i anmälan, kom ihåg att följa ditt konto i tjänsten Enter Finland.
Du har tre månader på dig att styrka din identitet efter att du fyllt i blanketten i Enter Finland-tjänsten.
Du kan styrka din identitet vid Migrationsverkets tjänsteställe eller utomlands vid Finlands beskickning.
Fråga utrikesministeriet vilken beskickning du kan besöka för att styrka din identitet.
Boka en tid i förväg.
Ta med dig ett identitetsbevis och ansökningsbilagorna i original.
Om du inte kan göra din ansökan elektroniskt eller inte vet hur man gör det kan du också lämna in anmälan på en pappersblankett.
Mer information om hur du gör medborgarskapsanmälan hittar du på Migrationsverkets webbplats.
Medborgarskapsanmälanfinska _ svenska _ engelska
Flerfaldigt medborgarskap
Finland godkänner flerfaldigt medborgarskap, d.v.s. att du utöver ditt finska medborgarskap även har medborgarskap i ett annat land.
Alla stater godkänner dock inte flerfaldigt medborgarskap.
Innan du ansöker om finskt medborgarskap är det bra att ta reda på om flerfaldigt medborgarskap också är tillåtet i det land där du är medborgare.
Om denna stat inte tillåter flerfaldigt medborgarskap kan du förlora ditt nuvarande medborgarskap när du får finskt medborgarskap.
Flerfaldigt medborgarskap kan vara en fördel, men också en nackdel.
Det lönar sig att till exempel ta reda på om man tvingas göra värnplikten i flera medborgarskapsstater eller om det räcker med ett intyg över fullgjord värnplikt i ett land.
Flerfaldigt medborgarskap kan vara en fördel när man till exempel flyttar från ett land till ett annat.
Migrationsverket ger råd i frågor som rör medborgarskap:
Telefon 0295 419 626 tisdag, onsdag och fredag kl. 10.00–11.00
Barnets flerfaldiga medborgarskap
Barnet kan ha finskt medborgarskap och medborgarskap i något annat land.
Detta beror på huruvida det andra landet godkänner flerfaldigt medborgarskap för barnet.
Fråga mer om detta vid beskickningen för ditt eget land.
Kan man förlora sitt finska medborgarskap?
Man kan förlora sitt finska medborgarskap om man
är 22 år gammal, har medborgarskap också i en annan stat och saknar tillräcklig anknytning till Finland
har angett felaktiga uppgifter i medborgarskapsansökan eller medborgarskapsanmälan
har förvärvat sitt medborgarskap på grund av faderns finska medborgarskap och faderskapet upphävs.
Att förlora sitt finska medborgarskapfinska _ svenska _ engelska
Bankkonto
Du behöver ett bankkonto för att sköta din dagliga ekonomi.
Det lönar sig att jämföra tjänsterna och priserna som olika banker tillhandahåller så att du hittar det alternativ som är förmånligast för dig.
När du öppnar ett bankkonto behöver du ett pass, ett identitetskort för utlänningar eller någon annan officiell identitetshandling.
Om du saknar pass eller ett identitetskort för utlänningar kan du ta reda på vilken typ av identitetshandling banken kan godta.
Vissa banker godtar främlingspass, som de finska myndigheterna har utfärdat, resedokument för flykting eller någon annan identitetshandling som kan godtas som resedokument.
I vissa fall kan banken även kräva andra utredningar av identiteten, om du har en notering i din handling som anger att din identitet inte har kunnat fastställas.
Du kan inte identifiera dig med ett körkort.
När du öppnar ett bankkonto har banken en lagstadgad skyldighet att fråga vad ditt konto ska användas till.
Banken har även rätt att kontrollera om du har betalningsanmärkningar.
Banken behöver följande uppgifter från dig:
personnummer
adress i Finland eller i ett annat land
om du betalar skatt i ett annat land än Finland, din adress i det landet
samma uppgifter för de personer som har rätt att använda kontot.
När du öppnar ett bankkonto lönar det sig att även skaffa webbankkoder.
Med hjälp av webbankkoderna kan du till exempel uträtta många myndighetsärenden på nätet.
För dessa koder gäller dock hårdare krav än för öppning av ett bankkonto.
I vissa fall kan du alltså inte få webbankkoder även om du har ett bankkonto.
Vill du ha råd i bankfrågor kan du ringa till Försäkrings- och finansrådgivningen (Fine).
Tjänsten är kostnadsfri för kunderna, dvs. du betalar endast din egen samtalskostnad.
Tjänsten tillhandahålls på finska, svenska och engelska.
Försäkrings- och finansrådgivningen
tfn. 09 6850 120
linkkiFinansbranschens Centralförbund:
Utländska medborgares bankärendenfinska _ engelska
Identitetskort för utlänningar
Polisen kan utfärda dig ett identitetskort för utlänningar om du har identifierats och din identitet har verifierats på ett tillförlitligt sätt.
Din identitet kan verifieras från en handling som styrker identiteten.
Om du inte har en sådan handling, kan dina fingeravtryck jämföras med de fingeravtryck som lagrats i uppehållstillståndskortet eller uppehållskortet.
Dessutom krävs att:
du har ett giltigt uppehållstillstånd eller uppehållskort eller att din uppehållsrätt är registrerad,
du har hemkommun i Finland och
uppgifter om dig har registrerats i befolkningsdatasystemet.
Med ett identitetskort för utlänningar kan du styrka din identitet i Finland.
Du kan använda det till exempel när du ska öppna ett bankkonto i Finland.
Du kan emellertid inte använda det som resedokument på utlandsresor.
ID-kortfinska _ svenska _ engelska
Försäkringar
När du har en bostad är det bra att ta en hemförsäkring.
Hemförsäkringen ersätter till exempel skador på möbler och andra ägodelar.
Hemförsäkringar säljs av försäkringsbolag.
Om du använder en egen bil ska du enligt lagen ha en trafikförsäkring.
Om du vill ta en personförsäkring i ett finländskt försäkringsbolag ska du vanligtvis ha ett finländskt FPA-kort.
Personförsäkringar kan vara till exempel olycksfallsförsäkring, vårdkostnadsförsäkring och livförsäkring.
Försäkringsbolag i Finlandfinska
Telefon
När du tecknar ett telefonabonnemang i Finland får du ett finskt telefonnummer.
Många företag erbjuder telefonabonnemang.
För att teckna ett abonnemang behöver du ett finländskt identitetsnummer och du måste ha en adress i Finland.
Du ska vanligtvis även kunna visa ditt betalningsbeteende, dvs. uppgifter som visar att du har betalat dina räkningar och inte har några betalningsanmärkningar.
I annat fall måste du betala abonnemanget i förskott.
Du kan också köpa ett prepaid-abonnemang.
Då behöver du inte ha en finländsk identitetshandling eller adress i Finland.
Prepaid-kortet är i förväg laddat med en summa som man sedan kan ringa för.
Prepaid-abonnemang kan köpas till exempel i R-kiosker, en del snabbköp och på Internet.
När du ringer till utlandet med telefon lönar det sig att kontrollera vilket utlandsprefix du ringer förmånligast med.
Många företag erbjuder förmånliga utlandsprefix.
Observera att samtalspriset ändå alltid beror på vilket land du ringer till.
Kontrollera vilket alternativ som är förmånligast för dig.
Telefonoperatörer i Finlandfinska
Förmånliga utlandssamtalfinska _ engelska
linkkiSkype:
Förmånliga utlandssamtalfinska _ svenska _ engelska _ ryska _ estniska _ franska _ spanska _ turkiska _ kinesiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ japanska _ italienska
_ danska
_ bulgariska
_ grekiska
_ tjeckiska
Internet
I Finland kan du sköta många ärenden via Internet.
Man kan ofta uträtta ärenden hos myndigheter eller företag via deras webbsidor.
Det är bra att skaffa sig en Internetanslutning så fort som möjligt efter att du har flyttat till Finland.
Du får en Internetanslutning hem till dig genom att teckna ett avtal med en Internettjänsteleverantör.
Det lönar sig att jämföra olika tjänsteleverantörers priser innan man ingår ett avtal.
I Finland finns många företag som erbjuder olika typer av Internetanslutningar.
Dessa företag hittar till exempel genom sökning på nätet när du skriver ”internetliittymä” i sökmaskinens sökfält.
Anslutningarnas priser varierar mycket.
Om du har ett bibliotekskort kan du också använda internet gratis på biblioteken.
Ett bibliotekskort får du gratis på biblioteket.
Läs mer på InfoFinlands sida Bibliotek.
Det finns också caféer där kunderna har möjlighet att använda Internet.
linkkiKommunikationsverket:
Internet- och telefonabonnemangfinska _ svenska _ engelska
Prisnivån i Finland
Prisnivån är hög i Finland.
Till exempel mat och många typer av tjänster kostar i genomsnitt mer i Finland än i övriga Europa.
Boendekostnaderna varierar mycket.
I storstäderna kostar boendet mycket mer än på mindre orter.
Konsumentpriser i de Europeiska ländernafinska _ svenska
Priser på icke subventionerade hyresbostäderengelska
Priser på hyresbostäder med statliga stödengelska
Information om priser på sålda bostäderfinska _ svenska
Köp och konsumentens rättigheter
Alla som köper varor och tjänster är konsumenter.
Konsumentskyddslagen tryggar konsumentens rättigheter i Finland.
Du har rätt till gottgörelse till exempel då varan som du köpt har fel som inte du har orsakat.
Du kan till exempel ersättas med en felfri vara eller få dina pengar tillbaka.
Om en vara som du köpt har brister ska du först kontakt säljaren.
Om du inte kan komma överens om saken med säljaren, ta då kontakt med konsumentrådgivningen.
linkkiKonkurrens- och konsumentverket:
Konsumentrådgivningfinska _ svenska _ engelska
Information om konsumenträttigheterfinska _ svenska _ engelska
Kollektivtrafik
Kollektivtrafiken fungerar väl i Finland.
Man kan resa nästan över allt i Finland med tåg eller buss.
Man kan också flyga till många städer.
I stora städer och deras näromgivning finns en välfungerande lokaltrafik.
Lokaltrafiken trafikeras vanligtvis med bussar.
Läs mer på InfoFinlands sida Trafiken i Finland.
Körkort
Du kan ta körkort i Finland när du har fyllt 18 år.
Om du har ett körkort som beviljats i ett annat land, beror det på situationen hur du ska gå tillväga.
Läs mer på InfoFinlands sida Trafiken i Finland.
Klimat och kläder
Klimatet i Finland är kallare än i många andra länder.
I Finland ligger medeltemperaturen på vintern under noll Celsiusgrader och på sommaren över +10 Celsiusgrader.
På våren och hösten ligger temperaturerna här emellan.
På vintern ska man klä sig varmt i Finland.
Läs mer om klimatet i Finland på InfoFinlands sida Klimatet i Finland.
Medier
I Finland utkommer nästan 200 tidningar.
Läs mer på InfoFinlands sida Medier i Finland.
Kulturen i Finland
Du hittar information om den finländska kulturen på InfoFinlands sidor Finländska seder och Den finländska arbetskulturen.
Om du har avlagt en examen utomlands kan du ha nytta av jämställande av examen, erkännande av yrkeskompetens eller av att skaffa dig rätt till yrkesutövning eller en fristående examen.
Erkännande och motsvarighet av examen
Erkännande av examen betyder ett avgörande om vilken behörighet en utländsk examen ger när man söker jobb eller studieplats i Finland.
Erkännande av examen är avgiftsbelagt och söks hos Utbildningsstyrelsen.
När du söker en studieplats krävs inte nödvändigtvis erkännande av examen.
Professionellt erkännande och rätt till yrkesutövning
Personer som söker till uppgifter inom den offentliga sektorn (staten och kommunerna) måste ofta uppfylla vissa behörighetsvillkor beträffande utbildningen.
När någon som studerat utomlands söker till dessa uppgifter behöver han eller hon oftast Utbildningsstyrelsens avgörande om den tjänstebehörighet som hans eller hennes examen ger.
Ett reglerat yrke avser en uppgift som endast kan sökas av personer som har avlagt en viss lagstadgad examen eller vissa studier.
Till reglerade yrken hör både uppdrag inom den offentliga sektorn och yrken för vilka det krävs rätt till yrkesutövning.
Rätt till yrkesutövning krävs till exempel i yrken inom hälsovården och sjöfarten.
Om du har en utländsk examen i något yrke som är reglerat i Finland behöver du ett beslut från någon behörig myndighet innan du kan utöva yrket Finland.
På Utbildningsstyrelsens webbplats finns en förteckning över de reglerade yrkena och de ansvariga myndigheterna.
I den privata sektorn kan arbetsgivaren själv bedöma huruvida den anställdas utländska examen godtas.
I den privata sektorn krävs inget beslut om erkännande, men beslutet kan vara nyttigt då man söker jobb.
Utbildningsstyrelsen ger också expertutlåtanden om utländska yrkesexamina.
Ett sådant utlåtande ger inte tjänstebehörighet i Finland, men det kan ändå vara till hjälp när man ansöker om ett arbete eller en studieplats, eftersom det beskriver innehållet i och nivån på utbildningen som man har avlagt utomlands.
Akademiskt erkännande
Om du vill fortsätta dina studier i Finland kan de studier som du avlagt utomlands tillgodoräknas med hjälp av akademiskt erkännande.
Akademiskt erkännande av examina betyder
att man söker sig till en utbildning på basis av sin utländska utbildning
att de utländska studierna tillgodoräknas som en del av en finländsk examen.
Läroanstalterna beslutar själva om antagningen av studerande och om de tillgodoräknar utländska studier som en del av en examen som avläggs i Finland.
Fråga mer vid den läroanstalt där du vill studera.
linkkiUtbildningsstyrelsen:
Erkännande av en examenfinska _ svenska _ engelska
linkkiUtbildningsstyrelsen :
Broschyr om erkännande av examen(pdf, 102,14 kt)finska _ svenska _ engelska _ ryska _ estniska _ franska _ spanska _ kinesiska _ persiska _ arabiska
linkkiUtbildningsstyrelsen :
Diagram över erkännande av examen(pdf, 410,87 kt)finska _ svenska _ engelska _ ryska
linkkiArbets- och näringsministeriet:
Erkännande av examenfinska _ svenska _ engelska
linkkiUtbildningsstyrelsen:
Reglerade yrkenfinska _ svenska _ engelska
linkkiUtbildningsstyrelsen:
Utlåtanden om utländska yrkesexamenfinska _ svenska _ engelska
På den här sidan finns information om den bosättningsbaserade sociala tryggheten som hör till FPA:s ansvarsområde.
På sidan finns information om de situationer då du betraktas ha rätt till den sociala trygghet som grundar sig på boende.
På InfoFinlands sida Utkomstskydd för arbetslösa får du mer information om vem som har rätt till utkomstskydd för arbetslösa.
FPA har bland annat hand om folkpensionen, barnbidrag, det grundläggande utkomstskyddet för arbetslösa, sjuk- och föräldradagpenningar, utkomststöd och rehabilitering.
FPA sköter även de sjukvårdsersättningar som betalas för privat sjukvård.
Om du är sjukförsäkrad i Finland, får du ett FPA-kort.
Grunderna för FPA:s bidrag definieras i lagen.
När du ansöker om en förmån, utreder FPA om du har rätt till FPA:s förmåner.
På detta inverkar ditt stadigvarande boende och arbete i Finland.
Varje sökandes livssituation behandlas individuellt när FPA fattar beslut om bidrag.
Sökandens livssituation och behov av understöd är ofta mycket olika.
Därför varierar även bidragens belopp och grunder.
Du ska alltid utreda din egen situation individuellt.
Offentliga hälso- och sjukvårdstjänster samt socialtjänster är kommunernas ansvar i Finland.
Läs mer på InfoFinlands sida Hälsovårdstjänster i Finland.
Mer information om rätten till hemkommun finns på InfoFinlands sida Hemkommun i Finland.
Information om social trygghetfinska _ svenska _ engelska
Social trygghet för dig som flyttar till Finland(pdf, 560 kb)finska _ svenska _ engelska _ ryska _ estniska
Information om sjukförsäkringfinska _ svenska _ engelska
linkkiSocial- och hälsovårdsministeriet:
Information om den sociala tryggheten i Finlandengelska
Rätten till FPA:s förmåner
Huvudregeln är att om du bor stadigvarande i Finland, kan du få FPA:s förmåner.
Vad stadigvarande boende betyder definieras i lagen.
Du kan också få rätt till FPA:s förmåner genom att arbeta i Finland.
Har du rätt till förmåner?
På detta inverkar om du flyttar till Finland från
ett land inom Europeiska unionen (EU), ett land inom det Europeiska ekonomiska samarbetsområdet (EES) eller Schweiz eller
från något annat land.
EES-länderna är Europeiska unionens medlemsländer samt Norge, Island och Liechtenstein.
Huruvida du får förmåner påverkas dessutom av om du flyttar till Finland till exempel som
arbetstagare eller företagare
studerande
familjemedlem
utsänd arbetstagare.
Finland har ingått avtal om den sociala tryggheten med ett antal länder.
Dessa länder är de nordiska länderna, USA, Kanada och Quebec, Chile, Israel, Indien, Kina, Sydkorea och Australien.
Avtalen rör främst pensioner.
En del avtal gäller även sjukvård.
Om du kommer från ett av dessa länder ska du kontrollera hos FPA om avtalen påverkar din sociala trygghet.
Lag om hemkommunfinska _ svenska
Information om internationella socialskyddsavtalfinska _ svenska _ engelska
Information om den sociala tryggheten i Finland för EU-medborgarefinska _ svenska _ engelska
Stadigvarande flytt till Finland och stadigvarande boende i Finland
När du flyttar till Finland bedömer FPA alltid först om din flytt till Finland är stadigvarande boende i den mening som avses i lagstiftningen om social trygghet.
Om din flytt till Finland inte anses vara stadigvarande, kan du ändå ha rätt till FPA:s förmåner på grund av att du arbetar.
Din flytt till Finland kan betraktas som stadigvarande i följande situationer:
du är återflyttare, det vill säga återvänder till Finland från utlandet
du har en fast anställning eller motsvarande avtal för ett arbete som du utför i Finland
du är gift eller annars i ett nära familjeförhållande till en person som redan bor stadigvarande i Finland.
Dessutom krävs det i allmänhet att ditt uppehållstillstånd är giltigt, om du är skyldig att ha ett uppehållstillstånd.
Din situation bedöms i sin helhet.
På basis av bedömningen beslutas om boendet är stadigvarande eller inte.
Om du flyttar till Finland tillfälligt har du vanligtvis inte rätt till FPA:s förmåner.
Från och med den 1 april 2019 kan studerande från länder utanför EU och EES ha rätt till vissa förmåner, till exempel förmåner som ingår i sjukförsäkringen.
När det finns ett avgörande om att ditt boende i Finland är stadigvarande, anses du bo stadigvarande i Finland så länge som
du har din egentliga bostad och ditt hem här och så länge du huvudsakligen vistas här
eller
du har en annan grund för den stadigvarande vistelsen, till exempel ett familjeband eller arbete.
Om du emellertid börjar arbeta i ett annat land eller reser utomlands för över sex månader, kan din rätt till FPA:s förmåner upphöra.
Mer information om sådana situationer får du vid FPA.
Det finns även bidrag som du inte kan få om du inte bor stadigvarande i Finland eller har gjort det tidigare.
Till exempel kan föräldrar få föräldradagpenning endast om de har bott i Finland minst 180 dagar före barnets beräknade förlossningsdatum.
Om du kommer från ett annat EU-land kan du i vissa fall utnyttja de försäkringsperioder som du har ackumulerat i andra EU-länder.
Fråga mer hos FPA:s center för internationella ärenden.
tfn 020 634 0200
kl. 9–16
Social trygghet för dig som flyttar till Finlandfinska _ svenska _ engelska
Flytt utomlands och social trygghetfinska _ svenska _ engelska
Kontaktuppgifter till FPAfinska _ svenska _ engelska
Arbete ger dig åtminstone delvis rätt till den sociala tryggheten i Finland
EU-länderna, EES-länderna och Schweiz
Om du flyttar till Finland för att arbeta får du vanligtvis rätt till FPA:s förmåner under din anställning, även när din anställning är kortvarig.
Om din lön uppgår till minst 696,60 € i månaden är du berättigad till de flesta av FPA:s förmåner.
Hur många timmar per vecka du arbetar eller hur lång din anställning är spelar ingen roll.
Arbetstagaren och den sociala tryggheten i Finlandfinska _ svenska _ engelska
Asylsökande
Asylsökande har inte rätt till finskt socialskydd.
Detta innebär att de inte har rätt till FPA:s förmåner.
Mottagningscentralen betalar mottagningspenning till asylsökande.
Den utbetalas så länge som asylansökan behandlas.
Mottagningspenningen är ett litet belopp som är avsett för ofrånkomliga utgifter.
Om den asylsökande beviljas uppehållstillstånd och är fast bosatt i Finland har han eller hon rätt till finskt socialskydd.
Man kan ansöka om att omfattas av det finska socialskyddet av FPA då uppehållstillstånd har beviljats.
Med integration (kotoutuminen) avses att du bosätter dig i Finland och skaffar kunskaper och färdigheter som du behöver i det finländska samhället.
Integrationen underlättas t.ex. av att
du lär dig språket,
hittar en arbetsplats eller studieplats,
får kontakter till det finländska samhället.
I Finland finns det olika tjänster som främjar din integration, hjälper dig att hitta sysselsättning och lära dig språket.
Också dina familjemedlemmar kan ha rätt till dessa tjänster om de flyttar till Finland tillsammans med dig.
Det är viktigt att du även själv aktivt främjar din integration.
Integrationsfrämjande tjänster
Grundläggande information om Finland
Alla invandrare har rätt att få grundläggande information om Finland.
När du får uppehållstillstånd eller registrerar din uppehållsrätt, får du samtidigt skriftlig information om
det finländska samhället och arbetslivet,
dina rättigheter och skyldigheter
tjänster som främjar din integration.
Invandrarrådgivning
Arbets- och näringsbyråerna och kommunerna tillhandahåller invandrarrådgivning.
De hjälper dig att integrera dig i Finland.
integration och integrationsfrämjande tjänster
arbetslivet
utbildning och studier.
Inledande kartläggning
Vid den inledande kartläggningen görs en utvärdering av det tjänster som kan främja din integration.
Vid den inledande kartläggningen utreds t.ex. din utbildning, din arbetserfarenhet och dina språkkunskaper.
Den inledande kartläggningen görs vid arbets- och näringsbyrån eller vid kommunen.
Den kan också göras på ett annat ställe, t.ex. vid en läroinrättning.
Detta beror på vilken kommun du bor i.
Du kan framföra en begäran om en inledande kartläggning av din situation t.ex. till arbets- och näringsbyrån eller socialbyrån i din kommun.
Invandrarrådgivningen ger dig närmare information om den inledande kartläggningen och hur den ordnas i din hemkommun.
Om du behöver stöd för din integration, utarbetas en integrationsplan för dig efter den inledande kartläggningen.
En integrationsplan utarbetas för dig åtminstone om
du är arbetslös arbetssökande eller
får utkomststöd eller
du inte fyllt 18 år och inte har en vårdnadshavare i Finland.
I integrationsplanen antecknas åtgärder som främjar din integration.
Planen kan omfatta t.ex. studier i finska, andra studier eller arbetspraktik.
Du kan utarbeta en integrationsplan t.ex. med en arbetskraftsrådgivare vid arbets- och näringsbyrån, alltså TE-byrån (TE-toimisto), eller med en socialarbetare på socialbyrån.
Integrationsplanen ska utarbetas senast tre år efter att du fått ditt första uppehållstillstånd eller din uppehållsrätt registrerades.
Integrationsplanens längd beror på hur lång tid du behöver stöd för din integration.
Integrationsplanen gäller vanligen i högst tre år.
I vissa specialfall kan den gälla i fem år.
När en integrationsplan har utarbetats för dig, är det viktigt att du följer planen.
TE-byrån eller kommunen anvisar dig vid behov till integrationsutbildning.
I utbildningen ingår studier i finska eller svenska och introduktion i det finländska samhället och arbetslivet samt den finländska kulturen.
I utbildningen kan även andra studier och praktik ingå.
TE-byrån, FPA eller kommunen utreder din rätt till arbetslöshetstförmån eller utkomststöd under integrationsplanen.
Om du har en arbetsplats kan din arbetsgivare eventuellt stöda din integration.
Arbetsgivaren kan t.ex. betala avgifter för en kurs i finska för din räkning.
Ibland kan arbetsgivaren också hjälpa dig med praktiska ärenden, t.ex. leta efter en bostad åt dig.
Fråga mer om detta av din arbetsgivare.
linkkiArbets- och näringsministeriet:
Inledande kartläggning och integrationsplanfinska _ svenska _ engelska
Stöd till arbetslösa invandrarefinska _ svenska _ engelska
Integrationsutbildning
När en integrationsplan utarbetats kan du få integrationsutbildning.
Integrationsutbildning ordnas av kommuner, arbets- och näringsbyråer och många läroanstalter.
Arbets- och näringsbyrån eller kommunen hänvisar dig till integrationsutbildningen.
Integrationsutbildningen omfattar vanligen studier i finska eller svenska. I utbildningen bekantar du dig med det finländska samhället och arbetslivet och den finländska kulturen.
Studier i finska och svenska
På InfoFinlands sida Finska och svenska språket hittar du information om möjligheterna att studera finska eller svenska.
Din kultur i Finland
Din kultur, ditt språk och din religion kan fortfarande utgöra en viktig del av ditt liv också i Finland.
En invandrarförening kan hjälpa dig att bevara och utveckla din kultur.
I Finland finns många föreningar för invandrare.
Du hitar mer information om föreningar på InfoFinlands sida Föreningar.
Barn med invandrarbakgrund kan få undervisning i det egna modersmålet.
Du hitar mer information på InfoFinlands sida Grundläggande utbildning.
I Finland råder religionsfrihet (uskonnonvapaus).
Var och en har alltså rätt att bekänna och utöva sin religion.
Var och en får själv välja sin religion.
Om du vill, kan du låta att bli att välja en religion.
Du hittar mer information om religionsutövning i Finland på InfoFinlands sida Kulturer och religioner i Finland.
linkkiArbets- och näringsministeriet:
Guiden Välkommen till Finland(pdf, 3,40 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
linkkiArbets- och näringsbyrån:
Information om integrationfinska _ svenska _ engelska
linkkiArbets- och näringsbyrån:
Broschyren Jobba i Finland(pdf, 5,51 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ polska
Läs jobbannonsen noga
Innan du skriver din jobbansökan, läs jobbannonsen noga och fundera på vilka färdigheter och vilket kunnande arbetsgivaren är ute efter.
Fundera på hur ditt kunnande motsvarar arbetsgivarens önskemål och krav.
Du kan också kontakta arbetsgivaren och begära mer information, om du undrar över något som inte framgår av jobbannonsen.
Ring arbetsgivaren bara om du har en konkret fråga om arbetsplatsen.
Jobbansökan
Vanligtvis när du söker ett jobb, skickar du en jobbansökan och ditt CV, alltså din meritförteckning, till arbetsgivaren.
Ibland kan jobbansökningen vara en video, en portfölj eller till exempel en webbsida.
Skriv ansökan och CV på samma språk som används i annonsen.
Skriv en ny ansökan och uppdatera ditt CV varje gång när du ansöker om ett nytt jobb.
Du kan skriva ansökningstexten direkt i e-postmeddelandet eller bifoga den till e-postmeddelandet tillsammans med ditt CV.
Lägg till bilagorna alltid i PDF-format.
Ofta kan du skicka in ansökan och CV via arbetsgivarens webbplats.
Syftet med din jobbansökan är att väcka arbetsgivarens intresse så att du blir kallad till anställningsintervju.
Ansökningen är ett svar på jobbannonsen.
Du ska svara på de önskemål och krav som nämns i jobbannonsen.
Lyft fram sådant som är viktigt i arbetsuppgiften.
Ge konkreta exempel på ditt kunnande.
Intyga arbetsgivaren om att du är lämplig för uppgiften.
En jobbansökan är oftast en knapp sida.
Be någon att läsa igenom och granska din ansökan.
Löneanspråk
Ofta ska man ange sitt löneanspråk i ansökningen.
Det är ofta svårt att uppskatta rätt belopp.
Löneanspråket får inte vara för stort, men inte heller för litet.
Från fackförbund får du mer information om lönenivån i olika branscher.
Lönejämförelse finska _ engelska
Gå igenom dina utbildningar och din arbetserfarenhet och fundera på vilka färdigheter du lärt dig i dem.
Vilka är dina styrkor?
Fundera också på vilket kunnande du har fått från dina fritidsintressen eller andra erfarenheter.
Tidsenliga intyg
Spara intygen från dina tidigare jobb och studier.
Kom ihåg att alltid begära ett intyg när du haft ett jobb, avlagt en praktik eller studerat.
Arbetsgivaren har skyldighet att utfärda ett intyg ännu tio år efter att anställningen upphört.
Du behöver vanligtvis inte skicka in dina arbetsintyg i förväg till arbetsgivaren, men det är bra att ta med dem till anställningsintervjun för det fall att arbetsgivaren vill se dem.
Det skulle vara bra att ha översättningar till finska eller svenska av alla intyg som du fått utomlands.
Mer information om detta finns på InfoFinlands sida Arbetsintyg.
Erkännande av examen
Det är lättare att söka jobb om du vet hur en examen som du avlagt utomlands motsvarar en finländsk examen.
Du kan ansöka om erkännande av utländsk examen vid Utbildningsstyrelsen.
Erkännande av examen är avgiftsbelagt.
Mer information om detta finns på InfoFinlands sida Utländsk examen i Finland.
linkkiUtbildningsstyrelsen:
Erkännande av en examenfinska _ svenska _ engelska
Öppen ansökan
Du kan ta direkt kontakt med en arbetsplats som du är intresserad av.
Du kan skicka in en öppen ansökan eller ringa arbetsgivaren, trots att de inte har några lediga jobb just nu.
I den öppna ansökan ska du berätta vad du kan och hurdana uppgifter du skulle kunna utföra.
Bifoga din meritförteckning, alltså CV, till ansökan.
Meritförteckning eller CV
En meritförteckning, eller ett CV, är en kortfattad och tydlig sammanfattning av ditt kunnande, din arbetserfarenhet och din utbildning.
Det finns olika CV-mallar.
I ett kompetensbaserat CV kan du gruppera dina färdigheter i olika kompetensområden.
CV:t kan även vara en video, en portfölj eller en webbsida.
Bekanta dig med olika CV-mallar och forma ditt eget CV såsom det passar dig.
Ett CV är vanligtvis 1–2 sidor långt.
Kom ihåg att uppdatera ditt CV för varje ny ansökan.
Vad innehåller ett CV?
Namn och kontaktuppgifter – Adress, e-postadress, telefonnummer
Arbetserfarenhet – Lista dina tidigare anställningar, den senaste först.
Ange också anställningens längd.
Beskriv dina arbetsuppgifter och de färdigheter som du lärt dig i arbetet.
Utbildning – Lista dina examina i kronologisk ordning, den senaste först.
Lägg till namnet på examen, utbildningsprogrammet och läroanstalten och när du tog examen.
Kurser – Lista kurserna i finska och andra kurser som du avlagt under en egen rubrik.
Övrigt kunnande – Språkkunskaper, IT-kunskaper, avlagda tillståndskort, till exempel hygienpass.
Publikationer eller andra arbetsprov
– Om du vill kan du även lista dina publikationer eller arbetsprov.
Fritidsintressen, förtroendeuppdrag
– Du kan även lyfta fram dina intressen.
Referenser – Du kan lägga till namnen på personer som har lovat att rekommendera dig för arbetsuppgiften.
Lägg till kontaktuppgifterna till dem.
Kom ihåg att be personen om tillstånd för detta.
I början av CV:t kan du tillfoga en sammanfattning eller profil där du beskriver din bakgrund och din kärnkompetens med några ord.
Du kan berätta vilka målsättningar du har med jobbsökningen eller vilken specialkompetens du besitter.
Du kan också lägga till ett fotografi.
linkkiArbets- och näringsministeriet:
Så här skriver du en jobbansökan och ett CVfinska _ svenska _ engelska
Kompetensbaserat CV
Ett kompetensbaserat CV lyfter fram ditt kunnande, dina färdigheter och dina erfarenheter.
Välj några kompetensområden och beskriv under rubrikerna dina erfarenheter, färdigheter och prestationer inom dem.
Du kan också lägga till sådant kunnande som du har införskaffat till exempel i frivilligarbete, fritidsintressen eller studier.
Dessutom kan du lista din arbetserfarenhet och utbildning i kronologisk ordning.
I början av CV:t kan du tillfoga en sammanfattning eller profil där du beskriver din bakgrund och din kärnkompetens med några ord.
Du kan berätta vilka målsättningar du har med jobbsökningen eller vilken specialkompetens du besitter.
Skriv ett eget CV för varje arbetsplats.
Lyft fram sådana färdigheter som behövs i uppgiften.
Fundera på vad arbetsgivaren bör veta om dina färdigheter och ditt kunnande.
Europass-CV
Europass är ett allmäneuropeiskt CV, alltså en allmäneuropeisk meritförteckning.
Det består av fem dokument som har till syfte att hjälpa arbetstagare och studerande att presentera sitt kunnande i Europa.
Dokumenten används i alla EU/EES-länderna.
Du kan använda Europass när du söker jobb eller studieplats.
Europass är särskilt nyttigt om du ansöker om ett jobb eller en utbildningsplats i Finland från ett annat EU-land.
linkkiEuropass.eu:
Information om CVfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Förbered dig på anställningsintervjun
Bekanta dig med arbetsgivaren i förväg till exempel med hjälp av webbplatsen.
Fundera på hur du ska lyfta fram ditt kunnande och din lämplighet för uppgiften.
Öva på att beskriva din bakgrund och din yrkeskunnighet med några meningar.
Fundera i förväg på vilka frågor arbetsgivaren kan ställa till dig.
Öva på att besvara allmänna frågor som ingår i en anställningsintervju.
Arbetsgivaren får inte fråga om din familj, vilken religion du har eller om du är politiskt aktiv.
Visa att du har bekantat dig med arbetsgivarens organisation och arbetsuppgiften i förväg och att du har ett äkta intresse för jobbet.
Fundera också på vilka frågor du vill ställa till arbetsgivaren.
linkkiArbets- och näringsministeriet:
Anvisningar för jobbintervjunfinska _ svenska _ engelska
Att börja på ett nytt jobb
Skriv alltid ett skriftligt anställningsavtal innan du börjar på ett nytt jobb.
Kom överens om anställningsavtalets innehåll med arbetsgivaren.
Läs avtalet noga innan du undertecknar det.
Läs mer på InfoFinlands sida Att komma överens om anställningsvillkoren.
När du börjar på ett nytt jobb ska du lämna ditt skattekort till arbetsgivaren.
Läs mer på InfoFinlands sida Skattekort.
Utlänningar som bor i Finland har nästan samma rättigheter och skyldigheter som finländarna.
Följande rättigheter och skyldigheter gäller även utlänningar som bor i Finland.
Rättigheter
Alla har rätt till likabehandling.
Ingen får särbehandlas till exempel på grund av kön, ålder, religion eller handikapp.
Var och en får fritt yttra sina åsikter i tal och skrift.
Människor får ordna möten och demonstrationer och delta i dem.
Demonstrationer ska anmälas till polisen på förhand.
Ingen får dömas till döden eller torteras.
Alla får själva välja sin bostadsort och röra sig fritt i Finland.
Alla har rätt till integritetsskydd.
Ett brev som tillhör en annan person får inte läsas och en annan persons telefonsamtal får inte avlyssnas.
Var och en får själv välja sin egen religion.
Om man inte vill behöver man inte välja någon religion alls.
Utlänningar som bor stadigvarande i Finland och som har fyllt 18 år har rätt att rösta i kommunalval.
Utlänningar som har rösträtt i kommunalval har även rätt att ställa upp som kandidat i kommunalval.
EU-medborgare som har hemort i Finland kan rösta i Europaparlamentsvalet om de har anmält sig till rösträttsregistret (äänioikeusrekisteri).
EU-medborgare som är i det finska rösträttsregistret kan också ställa upp som kandidat i Finlands Europaparlamentsval.
Läs mer om utlänningars rösträtt i Finland på InfoFinlands sida Val i Finland.
Skyldigheter
Alla som bor eller vistas i Finland måste följa Finlands lagar.
7–17-åringar har läroplikt (oppivelvollisuus), d.v.s. skyldighet att avlägga grundskolans (peruskoulu) lärokurs.
Ofta måste de som arbetar i Finland betalar skatt på sin lön i Finland.
Alla har skyldighet att vittna inför domstol om de blir kallade.
Föräldrar är skyldiga att ta hand om sina barn.
Alla har skyldighet att hjälpa vid en olycka.
Läs mer om beskattningen på InfoFinlands sida Beskattning.
Finska medborgares rättigheter och skyldigheter
Finska medborgare har utöver de ovannämnda också några ytterligare rättigheter och skyldigheter som utlänningar bosatta i Finland inte har.
Läs mer om finska medborgarnas rättigheter och skyldigheter på InfoFinlands sida Finskt medborgarskap.
Finlands grundlagfinska _ svenska _ engelska
Information om demokratin i Finlandfinska _ svenska _ engelska
Val i Finlandfinska _ svenska _ engelska
Flytta till Finland
Fortsatt uppehållstillstånd
Studera finska språket
Arbete och studier
Äktenskap och samboförhållande
Social trygghet
Tjänster för barnfamiljer
Hälsa
Flytta till Finland
Om du inte är medborgare i ett nordiskt land, EU-medborgare eller familjemedlem till en EU-medborgare som är bosatt i Finland, behöver du ett uppehållstillstånd.
Läs mer på InfoFinlands sida Familjen till Finland.
Om du är EU-medborgare behöver du inte uppehållstillstånd i Finland.
Om du vistas i Finland mer än tre månader, behöver du ett registreringsintyg för EU-medborgare (Unionin kansalaisen rekisteröintitodistus).
Om du inte är EU-medborgare, men din familjemedlem som är bosatt i Finland är EU-medborgare, behöver du ett uppehållskort för familjemedlem (perheenjäsenen oleskelukortti).
Läs mer på InfoFinlands sida EU-medborgare.
Om du är medborgare i ett nordiskt land behöver du inte uppehållstillstånd i Finland.
Läs mer på InfoFinlands sida Medborgare i nordiska länder.
På InfoFinlands sida Komihåglista för dig som flyttar till Finland hittar du nyttig information om vilka andra saker du bör ta hand om innan du flyttar till Finland.
När du flyttar till Finland ska du besöka magistraten (maistraatti)på orten där du är bosatt.
Vid magistraten kan du få en finsk personbeteckning, om du inte fick den redan i samband med att du beviljades uppehållstillstånd eller din uppehållsrätt för EU-medborgare registrerades vid Migrationsverket.
På magistraten utreder man även om det är möjligt att registrera en hemkommun i Finland för dig.
När du har en hemkommun kan du använda kommunens tjänster, såsom till exempel hälsovårdstjänster.
Läs mer på InfoFinlands sida Hemkommun i Finland.
Till Finland på grund av familjebandfinska _ svenska _ engelska
Registrering av uppehållsrätt för EU-medborgarefinska _ svenska _ engelska
Registrering av utlänningarfinska _ svenska _ engelska
Fortsatt uppehållstillstånd
Om du har ett uppehållstillstånd ska du komma ihåg att ansöka om fortsatt uppehållstillstånd i god tid innan giltigheten för det första tillståndet tar slut.
Ansök om fortsatt uppehållstillstånd elektroniskt i tjänsten Enter Finland eller på Migrationsverkets tjänsteställe.
Tillståndsbeslutet är avgiftsbelagt.
Du måste betala avgiften samtidigt som du ansöker om fortsatt uppehållstillstånd.
Mer information om att ansöka om fortsatt uppehållstillstånd hittar du på InfoFinlands sida Fortsatt uppehållstillstånd.
Om du är EU-medborgare kan du ansöka om permanent uppehållsrätt när du har bott i Finland fem år.
Att förlänga uppehållstillståndetfinska _ svenska _ engelska
Studera finska språket
Information om studier i finska språket hittar du på InfoFinlands sida Finska och svenska språket.
Om du bor i Helsingforsregionen, Tammerforsregionen eller Åboregionen kan du leta efter en kurs i finska språket som passar dig genom tjänsten Finnishcourses.fi.
Kurser i finska och svenska språketfinska _ engelska _ ryska
Arbete och studier
Om du har uppehållstillstånd på grund av familjeband, har du rätt att arbeta och studera i Finland.
Även medborgare i EU-länder och nordiska länder och deras familjemedlemmar har rätt att arbeta och studera.
Notera att om du har ansökt om ditt första uppehållstillstånd i Finland så har du inte rätt att arbeta innan tillståndet har beviljats.
Om du är intresserad av att grunda ett eget företag, gå in på InfoFinlands sida Att grunda ett företag.
Information om studier i Finland hittar du på InfoFinlands sida Utbildning.
Äktenskap och samboförhållande
Om du ska gifta dig i Finland hittar du nyttig information på InfoFinlands sida Äktenskap.
Information om att leva i ett samboförhållande i Finland hittar du på InfoFinlands sida Samboförhållande.
Du hittar information om skilsmässa på InfoFinlands sida Skilsmässa.
Notera att om du har ett uppehållstillstånd som beviljats på basis av familjeband, så kan förändringar i familjeförhållandena, såsom till exempel skilsmässa, påverka ditt uppehållstillstånd.
Läs mer på InfoFinlands sida Kan jag förlora mitt uppehållstillstånd?
På InfoFinlands sida Problem i äktenskap och parförhållande hittar du information om var du kan söka hjälp för problem i förhållandet.
Social trygghet
De flesta av FPA:s förmåner är sådana att du har rätt till dem endast om du flyttar ditt stadigvarande boende till Finland.
Social trygghet för dig som flyttar till Finlandfinska _ svenska _ engelska
Tjänster för barnfamiljer
Information om de tjänster och stöd som samhället erbjuder barnfamiljer hittar du på InfoFinlands sida Ekonomiskt stöd till familjer och Vård av barnet.
Hälsa
I Finland finns både offentliga och privata hälsovårdstjänster.
De offentliga hälsovårdstjänsterna är förmånligare än de privata.
Om du har en hemkommun i Finland kan du använda offentliga hälsovårdstjänster.
Om du flyttar till Finland av familjeskäl får du vanligen en hemkommun i Finland.
Magistraten fattar beslut om registrering av hemkommun.
Läs mer på InfoFinlands sida Hälsovårdstjänster i Finland och Hemkommun i Finland.
Lediga jobb
Sök lediga jobb på jobbförmedlingssidor på internet, i tidningar eller på sociala medier (till exempel Facebook och LinkedIn).
Du hittar jobbförmedlingssidor när du skriver "avoimet työpaikat" (lediga jobb) i sökmotorns sökfält.
linkkiArbets- och näringsministeriet:
Lediga jobbfinska _ svenska
linkkiArbets- och näringsförvaltningen:
Länkar till jobbsajterfinska _ svenska _ engelska
linkkiArbets- och näringsministeriet:
Yrkesbarometern finska _ svenska _ engelska
linkkiEures-portalen:
information om arbetsplatser i Europafinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiArbets- och näringsministeriet:
Tips för jobbsökningenfinska _ svenska _ engelska
Skapa nätverk och upprätthåll ditt kunnande
Du har nytta av nätverk när du söker jobb.
Identifiera och dra nytta av dina nätverk.
Lärare, studiekamrater, bekanta, tidigare kollegor och chefer kan också ingå i ditt nätverk.
Be om tips till jobbsökningen och hjälp med att skriva ansökningar av andra.
Fundera också på om du har någon i ditt nätverk som kan berätta om jobbtillfällen eller rekommendera dig.
Var aktiv.
Upprätthåll ditt kunnande, följ aktuella händelser och nyheter i din bransch, delta i kompletteringsutbildning och utveckla tidigare kunskaper.
Upprätthåll och utvidga ditt nätverk.
Även korta anställningar eller en praktik kan hjälpa dig att bygga ut ditt nätverk.
Besök fackevenemang i din bransch, gör frivilligarbete eller sök till ett mentorprogram.
Tänk på att frivilligarbete kan påverka din arbetslöshetsförsäkring.
Läs mer om frivilligarbete på InfoFinlands sida Frivilligarbete.
Lär dig finska eller svenska
När du kan språket är det lättare för dig att hitta jobb och sköta dina ärenden i det finländska samhället.
Du kan studera finska och svenska på olika kurser eller på egen hand via internet.
Läs mer om språkstudier i InfoFinlands avsnitt Finska och svenska språket.
Utnyttja sociala medier i jobbsökningen
Sociala nätverk på internet, såsom Facebook och LinkedIn, är bra verktyg för jobbsökningen.
Många arbetsgivare använder även Twitter som kommunikationskanal.
I tjänsterna kan du söka information om lediga jobb och bygga upp fackliga nätverk.
Du kan få viktig information om olika organisationers verksamhet och aktuella händelser i olika branscher eller delta i diskussioner.
Kontakta arbetsgivarna direkt
Du kan kontakta intressanta organisationer direkt och fråga om de har lediga jobb.
De flesta jobben är dolda jobb.
De annonseras inte ut öppet, utan arbetsgivarna söker arbetstagare via sina egna nätverk.
Du kan ringa en arbetsgivare direkt eller skicka en öppen ansökan via e-post.
Ofta kan du även skicka in en öppen ansökan via företagets webbplats.
Arbetsförmedlingstjänster
Du kan även söka jobb via företag som erbjuder arbetsförmedlingstjänster.
Arbetet kan vara kortvarigt, men det kan ge dig värdefull erfarenhet och du kan utvidga dina nätverk.
Du ingår ett avtal med företaget och företaget skickar dig till arbete för en annan arbetsgivare.
Via dessa företag kan du även få en fast anställning.
linkkiArbets- och näringsministeriet:
Hyrarbetsguidefinska _ svenska _ engelska
linkkiFörbundet för personaltjänsteföretag:
Personalbranschens regler om rekrytering av utlänningarfinska _ engelska
Sysselsätt dig som freelancer eller företagare
Arbete som freelancer innebär att du arbetar för flera uppdragsgivare utan fast anställning.
En freelancer måste själv sköta beskattningen och pensionsbetalningar.
Du kan fakturera vi en faktureringstjänst utan att starta ett eget företag.
Det kallas för lättföretagande.
Du kan även starta ett eget företag.
Tänk på att arbete som freelancer eller företagare kan påverka din arbetslöshetsförsäkring.
linkkiFreelanceri.info:
Länkar för frilansarefinska
Arbets- och näringsbyrån stöttar dig i jobbsökningen
Arbets- och näringsbyrån eller TE-byrån (TE-toimisto) ger dig handledning i jobbsökningen och information om lediga jobb och tillgängliga utbildningar.
Om du inte har ett jobb eller om du blir arbetslös, anmäl dig på arbets- och näringsbyrån senast på din första dag som arbetslös.
Läs mer på InfoFinlands sida Om du blir arbetslös.
Att anmäla sig som kund
Du kan anmäla dig som kund vid TE-byrån antingen vid den lokala TE-byrån eller på TE-byråns webbplats.
Om du är arbetslös arbetssökande, upprättar ni en integrationsplan eller en sysselsättningsplan.
Om du arbetar deltid eller bara lite, bedömer TE-byrån om du kan få en arbetslöshetsförmån samtidigt.
TE-byrån ordnar
yrkesutbildning
integrationsutbildning
utbildningsförsök
arbetsförsök
arbete med lönebidrag
arbetsträning
yrkesvägledning och karriärvägledning
linkkiArbets- och näringsministeriet:
Anmälan till arbets- och näringsbyrån finska _ svenska
linkkiTE-tjänster:
Videoklipp och broschyrer för invandrarefinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska
Integrationsutbildning
Om du har flyttat till Finland nyligen och behöver stöd med integrationen, kan du få plats i en integrationsutbildning via TE-byrån.
Integrationsutbildningen kan omfatta studier i finska, andra studier eller arbetsförsök.
Du kan även ansöka till utbildningen själv.
Du måste avtala om utbildningen med TE-byrån innan du inleder utbildningen.
Läs mer på InfoFinlands sida Integration i Finland.
linkkiArbets- och näringsministeriet:
Integrationstjänster för invandrarefinska _ svenska _ engelska
Stöd med jobbsökningen för under 30-åringar vid Navigatorn
Om du är under 30 år kan du få information om arbete, studier och annat som hör vardagslivet till vid Navigatorn.
Ohjaamofinska _ svenska _ engelska
Utbildnings- och arbetslivsguide för unga(pdf, 26 MB)finska _ svenska _ engelska _ ryska _ estniska _ somaliska
Välkommen till arbetslivet finska
Arbetslivets ABC finska
linkkiFFC:
Arbetslivet i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ kinesiska _ arabiska
linkkiArbets- och näringsministeriet:
Hitta jobb med hjälp av sysselsättningsprogrammet Kotouttamisen SIB finska _ engelska
Om du måste sköta ärenden med finländska myndigheter, men inte kan finska eller svenska och det inte heller finns något annat språk som både du och myndigheten talar, kan du i vissa fall ha rätt till tolkning.
Då beställer myndigheten tolken och betalar för tolkningen.
Myndigheten kan ordna och betala tolkningen när det gäller skötsel av ärenden som behandlas på myndighetens initiativ.
Detta är dock inte alltid möjligt.
Om du behöver en tolk för den inledande kartläggningen och integrationsplanen, måste myndigheten beställa en tolk.
Du kan på förhand fråga myndigheten om detta.
Om du söker asyl i Finland har du rätt till tolkning i ärenden som rör behandlingen av din asylansökan.
Du har rätt att få information om ett beslut gällande dig på ditt modersmål eller ett annat språk som du förstår.
Information om beslutet ges genom tolkning eller översättning.
Om du själv bokar tolken och betalar tolkningen, kan du anlita en tolk när som helst.
Tolktjänsterfinska _ svenska _ engelska
Vad gör tolken?
Tolken är med på möten mellan dig och myndigheten.
Han eller hon tolkar det som du och myndigheten säger.
Tolken är antingen på plats eller också kan tolkningen ordnas via telefon eller video.
Tolken har som uppgift att tolka det som du och myndigheten säger.
Tolken sköter inga andra uppgifter utöver tolkningen.
Han eller hon kan således inte hjälpa dig med annat.
Tolken är en neutral, utomstående person som varken är på din eller på myndighetens sida.
Tolken har sekretessplikt och får inte berätta inte om dina angelägenheter för andra.
Var kan man beställa en tolk?
I Finland finns åtta kommunala tolkcentraler (tulkkikeskus).
Tolkcentralernas tjänster är främst avsedda för myndigheter som arbetar med invandrare.
Också många företag erbjuder tolktjänster.
linkkiFinlands översättar- och tolkförbund:
Sök tolk eller översättarefinska _ svenska _ engelska
Kommunala tolkcentraler
linkkiHelsingforsnejdens kontakttolkcentral:
Tolkningfinska
linkkiMellersta Finlands tolkcentral:
Tolkningfinska _ svenska _ engelska
Tolkningfinska
Tolkningfinska _ engelska
linkkiÖsterbottens tolkcentral:
Tolkningfinska
linkkiNorra Finlands tolktjänst:
Tolkningfinska
linkkiÅboregionens tolkcentral:
Tolkningfinska _ svenska
Tolkningfinska
Vem är asylsökande?
Asylsökandes uppehållsrätt
Social trygghet
Familjeåterförening
Hälsa
Vem är asylsökande?
En asylsökande (turvapaikanhakija) är en person som söker skydd och uppehållsrätt i en främmande stat.
Internationellt skydd kan beviljas om personen känner välgrundad fruktan för förföljelse (på grund av ras, religion, tillhörighet till en viss samhällsgrupp eller politisk samhörighet) eller om personen annars är utsatt för verklig fara i sitt hemland eller sitt permanenta bosättningsland.
En asylsökande är alltså inte en flykting (pakolainen).
Om en asylsökande beviljas flyktingstatus eller uppehållstillstånd på grund av skyddsbehov eller på någon annan grund får han eller hon stanna i Finland.
Broschyren Information till asylsökandefinska _ svenska _ engelska _ ryska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
Asylsökandes uppehållsrätt
Du får stanna i Finland om du beviljas asyl eller uppehållstillstånd på någon annan grund.
Om förhållandena i ditt hemland är sådana att du inte behöver asyl och det inte heller finns andra grunder att bevilja uppehållstillstånd, avslås din ansökan och du utvisas från Finland.
Om du får avslag på din asylansökan eller ansökan om uppehållstillstånd har du rätt att överklaga beslutet.
Läs mer på InfoFinlands sida Som asylsökande till Finland.
Att söka asyl i Finlandfinska _ svenska _ engelska
Social trygghet
Asylsökande har inte rätt till finskt socialskydd.
Detta innebär att de inte har rätt till FPA:s förmåner.
Mottagningscentralen betalar mottagningspenning till asylsökande.
Den utbetalas så länge som asylansökan behandlas.
Mottagningspenningen är ett litet belopp som är avsett för ofrånkomliga utgifter.
Om den asylsökande beviljas uppehållstillstånd och är fast bosatt i Finland har han eller hon rätt till finskt socialskydd.
Man kan ansöka om att omfattas av det finska socialskyddet av FPA då uppehållstillstånd har beviljats.
Familjeåterförening
Asylsökande har inte rätt till familjeåterförening.
Dina familjemedlemmar kan inte få uppehållstillstånd i Finland på grund av familjeband.
Om du får uppehållstillstånd i Finland kan dina familjemedlemmar ansöka om tillstånd på grund av familjeband.
Läs mer på InfoFinlands sida Till familjemedlem i Finland.
Att söka uppehållstillstånd på grund av familjebandfinska _ svenska _ engelska
Hälsa
Asylsökande har vanligtvis inte tillgång till offentlig hälsoåvård exempelvis på hälsocentraler.
Mottagningscentralen anordnar hälsovårdstjänster för asylsökande.
Hälsovårdare på mottagningscentralen ser till att asylsökande får den vård de behöver.
Fråga mer på din mottagningscentral.
Om du fått uppehållstillstånd och din hemkommun finns i Finland kan du använda tjänsterna inom den offentliga hälsovården på samma sätt som de övriga invånarna i kommunen.
Hälsovård för papperslösa
Global Clinic är en klinik där du kan få hjälp eller råd av en läkare eller sjukskötare om du vistas i Finland utan uppehållstillstånd.
Du kan besöka Global Clinic även om du inte behöver brådskande sjukvård.
Global Clinic bedriver verksamhet i följande städer:
Åbo
Tammerfors
Uleåborg
Joensuu
Du kan ringa eller skicka e-post.
En sjukskötare eller läkare besvarar ditt samtal.
Du hittar kontaktinformation på Global Clinic:s hemsidor.
Global Clinic:s tjänster är avgiftsfria för kunderna.
Global Clinic anmäler inte sina kunder till polisen eller andra myndigheter.
Klinikens adress eller öppettider meddelas inte offentligt.
Kontaktuppgifterfinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Anmäl flyttningen till myndigheterna
När du flyttar utomlands från Finland ska du göra en flyttanmälan till magistraten (maistraatti)
Du kan göra flyttanmälan på internet eller med en blankett som du får i magistraten eller på posten.
Om du flyttar permanent från Finland eller vistas utomlands två år utan avbrott återkallas ditt uppehållstillstånd.
Du kan ställa Migrationsverket (Maahanmuuttovirasto) en ansökan om att inte återkalla ditt uppehållstillstånd.
Ansökan ska göras innan du har vistats utomlands över två år.
Mer information om detta hittar du på InfoFinlands sida Kan jag förlora mitt uppehållstillstånd?.
Flyttning utomlands och social trygghet
När du flyttar utomlands för att bo där eller lämnar
Finland för en längre tid än för en kort semesterresa, ska du också anmäla detta till FPA (Kela) Om du omfattas av den sociala tryggheten i Finland och flyttar utomlands för högst ett år, bibehålls din rätt till den sociala tryggheten i Finland vanligen under din vistelse utomlands.
Om du flyttar till något EU- eller EES-land för att arbeta övergår du till den sociala tryggheten i det land där du arbetar, även om din vistelse varar under ett år.
Då kan du inte omfattas av den sociala tryggheten i Finland.
Om du flyttar utomlands för över ett år, betraktas flyttningen som permanent flyttning.
Då upphör din rätt till den sociala tryggheten i Finland när du flyttar bort från Finland.
I vissa fall kan du dock bibehålla din rätt till den sociala tryggheten i Finland även om du vistas utomlands över ett år.
Till exempel studerande har denna möjlighet.
Det gäller även arbetstagare som blivit utsända utomlands av sin finska arbetsgivare.
Detta förutsätter att du lämnar in en ansökan i ärendet inom ett år efter din flytt utomlands.
Om du flyttar till ett EU-land, ett EES-land eller Schweiz som utsänd arbetstagare (lähetetty työntekijä), ska din arbetsgivare hämta intyget E101/A1 för dig vid Pensionsskyddscentralen.
Intyget ska hämtas innan du åker utomlands.
Med intyget kan du bevisa att du omfattas av den sociala tryggheten i Finland även om du arbetar utomlands.
När du är utomlands kan din sociala trygghet påverkas till exempel av att du inleder studier eller börjar arbeta.
Anmäl alltid förändringar i omständigheterna till FPA.
Mer information om den sociala tryggheten i Finland hittar du på FPA:s webbplats och på InfoFinlands sida Den sociala tryggheten i Finland.
Frivillig återflyttning av flyktingar, asylsökande och emigranter
Om du vill återvända till ditt hemland kan du i vissa fall få stöd för frivilligt återvändande.
Stödet består antingen av pengar eller tjänster.
Penningsummans storlek beror på vilket land du återvänder till.
Tjänsten kan till exempel vara att du får hjälp med att leta efter en bostad eller arbetsplats i det land dit du återvänder.
Du kan få stöd om:
du är asylsökande och handläggningen av din ansökan är oavslutad
du har fått ett negativt beslut på din asylansökan
du är ett offer för människohandel och du inte har en hemkommun i Finland
du har ett tillfälligt uppehållstillstånd på grund av hinder för avlägsnande ur landet
du har fått tillfälligt skydd
din flyktingstatus i Finland har upphört eller återkallats eller det har fattats beslut om att avvisa dig.
Om du är kund hos en mottagningscentral kan du ansöka om stöd för frivilligt återvändande vid din egen mottagningscentral.
Om du inte är kund hos en mottagningscentral kan du ansöka om stöd hos Migrationsverket.
Flyttanmälanfinska _ svenska _ engelska
Återkallelse av uppehållstillståndfinska _ svenska _ engelska
Flytt utomlands och social trygghetfinska _ svenska _ engelska
Frivillig återflyttningfinska _ svenska _ engelska
Social- och hälsovårdsministeriet:
Ditt sociala skydd när du flyttar utomlands
Bankkonto
Du behöver ett bankkonto för att sköta din dagliga ekonomi.
Det lönar sig att jämföra tjänsterna och priserna som olika banker tillhandahåller så att du hittar det alternativ som är förmånligast för dig.
När du öppnar ett bankkonto behöver du ett pass, ett identitetskort för utlänningar eller någon annan officiell identitetshandling.
Om du saknar pass eller ett identitetskort för utlänningar kan du ta reda på vilken typ av identitetshandling banken kan godta.
Vissa banker godtar främlingspass, som de finska myndigheterna har utfärdat, resedokument för flykting eller någon annan identitetshandling som kan godtas som resedokument.
I vissa fall kan banken även kräva andra utredningar av identiteten, om du har en notering i din handling som anger att din identitet inte har kunnat fastställas.
Du kan inte identifiera dig med ett körkort.
När du öppnar ett bankkonto har banken en lagstadgad skyldighet att fråga vad ditt konto ska användas till.
Banken har även rätt att kontrollera om du har betalningsanmärkningar.
Banken behöver följande uppgifter från dig:
personnummer
adress i Finland eller i ett annat land
om du betalar skatt i ett annat land än Finland, din adress i det landet
samma uppgifter för de personer som har rätt att använda kontot.
När du öppnar ett bankkonto lönar det sig att även skaffa webbankkoder.
Med hjälp av webbankkoderna kan du till exempel uträtta många myndighetsärenden på nätet.
För dessa koder gäller dock hårdare krav än för öppning av ett bankkonto.
I vissa fall kan du alltså inte få webbankkoder även om du har ett bankkonto.
Vill du ha råd i bankfrågor kan du ringa till Försäkrings- och finansrådgivningen (Fine).
Tjänsten är kostnadsfri för kunderna, dvs. du betalar endast din egen samtalskostnad.
Tjänsten tillhandahålls på finska, svenska och engelska.
Försäkrings- och finansrådgivningen
tfn. 09 6850 120
linkkiFinansbranschens Centralförbund:
Utländska medborgares bankärendenfinska _ engelska
Identitetskort för utlänningar
Polisen kan utfärda dig ett identitetskort för utlänningar om du har identifierats och din identitet har verifierats på ett tillförlitligt sätt.
Din identitet kan verifieras från en handling som styrker identiteten.
Om du inte har en sådan handling, kan dina fingeravtryck jämföras med de fingeravtryck som lagrats i uppehållstillståndskortet eller uppehållskortet.
Dessutom krävs att:
du har ett giltigt uppehållstillstånd eller uppehållskort eller att din uppehållsrätt är registrerad,
du har hemkommun i Finland och
uppgifter om dig har registrerats i befolkningsdatasystemet.
Med ett identitetskort för utlänningar kan du styrka din identitet i Finland.
Du kan använda det till exempel när du ska öppna ett bankkonto i Finland.
Du kan emellertid inte använda det som resedokument på utlandsresor.
ID-kortfinska _ svenska _ engelska
Försäkringar
När du har en bostad är det bra att ta en hemförsäkring.
Hemförsäkringen ersätter till exempel skador på möbler och andra ägodelar.
Hemförsäkringar säljs av försäkringsbolag.
Om du använder en egen bil ska du enligt lagen ha en trafikförsäkring.
Om du vill ta en personförsäkring i ett finländskt försäkringsbolag ska du vanligtvis ha ett finländskt FPA-kort.
Personförsäkringar kan vara till exempel olycksfallsförsäkring, vårdkostnadsförsäkring och livförsäkring.
Försäkringsbolag i Finlandfinska
Telefon
När du tecknar ett telefonabonnemang i Finland får du ett finskt telefonnummer.
Många företag erbjuder telefonabonnemang.
För att teckna ett abonnemang behöver du ett finländskt identitetsnummer och du måste ha en adress i Finland.
Du ska vanligtvis även kunna visa ditt betalningsbeteende, dvs. uppgifter som visar att du har betalat dina räkningar och inte har några betalningsanmärkningar.
I annat fall måste du betala abonnemanget i förskott.
Du kan också köpa ett prepaid-abonnemang.
Då behöver du inte ha en finländsk identitetshandling eller adress i Finland.
Prepaid-kortet är i förväg laddat med en summa som man sedan kan ringa för.
Prepaid-abonnemang kan köpas till exempel i R-kiosker, en del snabbköp och på Internet.
När du ringer till utlandet med telefon lönar det sig att kontrollera vilket utlandsprefix du ringer förmånligast med.
Många företag erbjuder förmånliga utlandsprefix.
Observera att samtalspriset ändå alltid beror på vilket land du ringer till.
Kontrollera vilket alternativ som är förmånligast för dig.
Telefonoperatörer i Finlandfinska
linkkiTeleAle:
Förmånliga utlandssamtalfinska _ svenska _ engelska
Förmånliga utlandssamtalfinska _ engelska
linkkiSkype:
Förmånliga utlandssamtalfinska _ svenska _ engelska _ ryska _ estniska _ franska _ spanska _ turkiska _ kinesiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ ungerska _ japanska
Internet
I Finland kan du sköta många ärenden via Internet.
Man kan ofta uträtta ärenden hos myndigheter eller företag via deras webbsidor.
Det är bra att skaffa sig en Internetanslutning så fort som möjligt efter att du har flyttat till Finland.
Du får en Internetanslutning hem till dig genom att teckna ett avtal med en Internettjänsteleverantör.
Det lönar sig att jämföra olika tjänsteleverantörers priser innan man ingår ett avtal.
I Finland finns många företag som erbjuder olika typer av Internetanslutningar.
Dessa företag hittar till exempel genom sökning på nätet när du skriver ”internetliittymä” i sökmaskinens sökfält.
Anslutningarnas priser varierar mycket.
Om du har ett bibliotekskort kan du också använda internet gratis på biblioteken.
Ett bibliotekskort får du gratis på biblioteket.
Läs mer på InfoFinlands sida Bibliotek.
Det finns också caféer där kunderna har möjlighet att använda Internet.
linkkiKommunikationsverket:
Internet- och telefonabonnemangfinska _ svenska _ engelska
Prisnivån i Finland
Prisnivån är hög i Finland.
Till exempel mat och många typer av tjänster kostar i genomsnitt mer i Finland än i övriga Europa.
Boendekostnaderna varierar mycket.
I storstäderna kostar boendet mycket mer än på mindre orter.
Konsumentpriser i de Europeiska ländernafinska _ svenska
Priser på icke subventionerade hyresbostäderengelska
Priser på hyresbostäder med statliga stödengelska
Information om priser på sålda bostäderfinska _ svenska
Köp och konsumentens rättigheter
Alla som köper varor och tjänster är konsumenter.
Konsumentskyddslagen tryggar konsumentens rättigheter i Finland.
Du har rätt till gottgörelse till exempel då varan som du köpt har fel som inte du har orsakat.
Du kan till exempel ersättas med en felfri vara eller få dina pengar tillbaka.
Om en vara som du köpt har brister ska du först kontakt säljaren.
Om du inte kan komma överens om saken med säljaren, ta då kontakt med konsumentrådgivningen.
linkkiKonkurrens- och konsumentverket:
Konsumentrådgivningfinska _ svenska _ engelska
Information om konsumenträttigheterfinska _ svenska _ engelska
linkkiKonsumentförbundet:
Information om konsumenträttigheterfinska
Kollektivtrafik
Kollektivtrafiken fungerar väl i Finland.
Man kan resa nästan över allt i Finland med tåg eller buss.
Man kan också flyga till många städer.
I stora städer och deras näromgivning finns en välfungerande lokaltrafik.
Lokaltrafiken trafikeras vanligtvis med bussar.
Läs mer på InfoFinlands sida Trafiken i Finland.
Körkort
Du kan ta körkort i Finland när du har fyllt 18 år.
Om du har ett körkort som beviljats i ett annat land, beror det på situationen hur du ska gå tillväga.
Läs mer på InfoFinlands sida Trafiken i Finland.
Klimat och kläder
Klimatet i Finland är kallare än i många andra länder.
I Finland ligger medeltemperaturen på vintern under noll Celsiusgrader och på sommaren över +10 Celsiusgrader.
På våren och hösten ligger temperaturerna här emellan.
På vintern ska man klä sig varmt i Finland.
Läs mer om klimatet i Finland på InfoFinlands sida Klimatet i Finland.
Medier
I Finland utkommer nästan 200 tidningar.
Läs mer på InfoFinlands sida Medier i Finland.
Kulturen i Finland
Du hittar information om den finländska kulturen på InfoFinlands sidor Finländska seder och Den finländska arbetskulturen.
Vem är flykting?
Familjeåterförening
Eftersökning av försvunna anhöriga
Hälsa
Stöd för flyktingar
Vem är flykting?
En flykting är en person med flyktingstatus.
Flyktingstatus får de som beviljas asyl eller som tas till Finland i flyktingkvoten.
Kvotflyktingar
Man kan inte ansöka om att bli kvotflykting (kiintiöpakolainen) via myndigheterna i Finland.
Man kan inte heller föreslå en annan person, till exempel en släkting eller vän, som kvotflykting.
Finland tar som kvotflyktingar emot personer som har flyktingstatus enligt Förenta nationernas flyktingorganisation UNHCR.
Kvotflyktingarna väljs bland de personer som UNHCR föreslår till Finland.
De finländska myndigheterna intervjuar flyktingarna som UNHCR har föreslagit och väljer bland dem de personer som tas emot till Finland.
Intervjuerna görs i de länder där flyktingarna vistas, vanligen i flyktingläger eller i UNHCR:s lokaler.
Valet av kvotflyktingar påverkas till exempel av följande faktorer:
Flyktingen är i behov av internationellt skydd.
Flyktingens mänskliga rättigheter förverkligas inte i det land där han eller hon vistas.
Flyktingen utgör inget hot för Finlands säkerhet.
Flyktingen har förutsättningar att integreras i Finland.
En del flyktingar väljs utan intervju på basis av UNHCR:s dokument.
Dessa är vanligen nödfall, med andra ord flyktingar som är i ett brådskande behov av asyl till exempel av hälsorelaterade eller politiska orsaker.
Finlands riksdag beslutar hur många flyktingar som tas till landet.
Från och med år 2001 har Finlands flyktingkvot varit 750 personer per år.
Inrikesministeriet beslutar från vilka länder kvotflyktingarna tas.
Beviljande av flyktingstatus till asylsökande
En person kan erhålla flyktingstatus också genom att söka asyl i Finland.
Asylsökanden kan beviljas flyktingstatus om han eller hon har befogade skäl att frukta förföljelse i sitt hemland på grund av ras, religion, nationalitet, tillhörighet till en viss samhällsgrupp eller på grund av sin politiska uppfattning och då sökanden på grund av detta inte kan återvända till sitt hemland.
Asylsökande som inte beviljas flyktingstatus kan ändå få uppehållstillstånd i Finland på någon annan grund.
Läs mer på InfoFinlands sida Som asylsökande till Finland.
Information om val av kvotflyktingarfinska _ svenska _ engelska
Familjeåterförening
Också flyktingens familjemedlemmar kan få uppehållstillstånd i Finland.
Vilka som är familjemedlemmar definieras i lagen.
Endast dessa familjemedlemmar kan få uppehållstillstånd på grund av familjeband.
I Finland betraktas som familjemedlemmar
registrerad partner
sambo
vårdnadshavaren till ett barn under 18 år.
För att familjemedlemmarna ska kunna få uppehållstillstånd, krävs det i vissa fall att flyktingen har en tillräcklig inkomst för att försörja sina familjemedlemmar i Finland.
Mer information om familjeåterförening finns på InfoFinlands sida Till familjemedlem i Finland.
Hjälp med familjeåterföreningen
Om du har kommit till Finland som kvotflykting, kan Migrationsverket ersätta kostnaderna för en familjemedlems inresa.
Kostnaderna ersätts dock endast i de fall där familjebandet har funnits redan före du fick ditt första uppehållstillstånd i Finland.
Andra anhörigas resekostnader ersätts inte.
Endast kvotflyktingar kan få ersättning för familjemedlemmarnas resekostnader.
Finlands Rösa Kors hjälper med researrangemangen för kvotflyktingar
Migrationsverket ersätter resekostnaderna endast i det fall att familjemedlemmen reser till Finland på en resa som arrangeras av Finlands Röda Kors och Internationella organisationen för migration.
Finlands Röda Kors hjälper med att ordna resan till Finland för kvotflyktingens familjemedlemmar när dessa fått uppehållstillstånd.
Röda Korset ger också rådgivning om reglerna för familjeåterförening och därom, hur familjemedlemmarna ska gå tillväga för att ansöka om familjeåterförening.
När Migrationsverket har gett ett positivt beslut på din ansökan om återförening på grund av familjeband och anser att staten kan bekosta resan för dina familjemedlemmar, skickar det sitt beslut till Röda Korset.
Om du har kommit till Finland som kvotflykting och vill att finska staten bekostar resan för dina familjemedlemmar ska du ta kontakt med Röda Korsets beredskapsenhet som sätter igång researrangemangen.
Finlands Röda Kors kan inte bistå familjemedlemmarnas flygresor eller andra resor ekonomiskt.
Att söka uppehållstillstånd på grund av familjebandfinska _ svenska _ engelska
Familjemedlem till en flyktingfinska _ svenska _ engelska
Eftersökning av försvunna anhöriga
Om du vill ha kontakt med en anhörig som försvunnit kan du be om hjälp vid personefterforskningen vid Finlands Röda Kors.
Röda Korset hjälper familjer som skilts åt vid olika katastrofer eller kriser.
Röda Korset söker försvunna anhöriga och förmedlar meddelanden på krisområden.
linkkiFinlands Röda Kors:
Efterforskning av anhörigafinska _ svenska _ engelska _ franska _ somaliska
linkkiFinlands Röda Kors:
Efterforskning av anhörigafinska _ svenska _ engelska _ ryska _ somaliska _ spanska _ persiska _ arabiska _ portugisiska
Hälsa
Om du har kommit till Finland som kvotflykting, har du hemkommun i Finland och då kan du använda de offentliga hälsovårdstjänsterna.
Stöd för flyktingar
Flyktingar och asylsökande kan söka hjälp och rådgivning i juridiska frågor bland annat vid Flyktingrådgivningen r.f. eller rättshjälpsbyråerna (oikeusaputoimisto).
Flyktingrådgivningen ger asylsökande rättshjälp i asylprocessens första skede.
Flyktingrådgivningen ger också andra utlänningar allmän rättshjälp.
Rättshjälpsbyråerna ger personer som är bosatta i Finland expertråd i skötseln av juridiska ärenden.
För att sköta ett juridiskt ärende kan man få ett rättsbiträde bekostat antingen helt eller delvis med statliga medel.
Finlands flyktinghjälp r.f. är en organisation som arbetar för att främja flyktingarnas grundläggande rättigheter.
Organisationens verksamhet i Finland omfattar informering, utbildning och socialarbete.
Flyktinghjälpen hjälper flyktingar och invandrare till exempel i frågor som rör integrationen, boendet och grundandet av egna organisationer.
linkkiFinlands flyktinghjälp r.f.:
Stöd till flyktingarfinska _ svenska _ engelska
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Många länder har en beskickning i Finland.
Beskickningen kan antingen vara en ambassad eller ett konsulat.
Ambassaderna finns i Helsingfors.
Vissa länder har också konsulat i andra städer.
Om du behöver sköta ett ärende med myndigheterna i ditt hemland ska du ta kontakt med ditt lands beskickning.
Via beskickningen kan du ofta uträtta till exempel följande ärenden:
Få en födelseattest
Ansöka om medborgarskap i ditt hemland om du har förlorat det eller avstått från det
Anmäla födelsen av ditt barn till myndigheterna i ditt hemland om barnet föds i Finland
Ansöka om medborgarskap i ditt hemland för ditt barn om barnet har fötts i Finland
Registrera ett äktenskap i ditt hemland om du har gift dig i Finland
Rösta i val i ditt hemland
Observera att alla beskickningar inte erbjuder samma tjänster.
Det är inte nödvändigtvis möjligt att sköta alla ovannämnda ärenden i alla beskickningar.
Vilka tjänster ditt lands beskickning tillhandahåller beror på lagen i ditt hemland.
Mer information får du från ditt hemlands beskickning.
Alla länder har inte en beskickning i Finland.
I detta fall betjänas du ofta av ditt hemlands beskickning i något av Finlands grannländer.
På det finska utrikesministeriets webbplats finns en förteckning över andra länders beskickningar i Finland.
Där hittar du även kontaktuppgifterna till beskickningarna.
Andra länders beskickningar i Finlandfinska _ svenska _ engelska
Med integration (kotoutuminen) avses att du bosätter dig i Finland och skaffar kunskaper och färdigheter som du behöver i det finländska samhället.
Integrationen underlättas t.ex. av att
du lär dig språket,
hittar en arbetsplats eller studieplats,
får kontakter till det finländska samhället.
I Finland finns det olika tjänster som främjar din integration, hjälper dig att hitta sysselsättning och lära dig språket.
Också dina familjemedlemmar kan ha rätt till dessa tjänster om de flyttar till Finland tillsammans med dig.
Det är viktigt att du även själv aktivt främjar din integration.
Integrationsfrämjande tjänster
Grundläggande information om Finland
Alla invandrare har rätt att få grundläggande information om Finland.
När du får uppehållstillstånd eller registrerar din uppehållsrätt, får du samtidigt skriftlig information om
det finländska samhället och arbetslivet,
dina rättigheter och skyldigheter
tjänster som främjar din integration.
Invandrarrådgivning
Arbets- och näringsbyråerna och kommunerna tillhandahåller invandrarrådgivning.
De hjälper dig att integrera dig i Finland.
integration och integrationsfrämjande tjänster
arbetslivet
utbildning och studier.
Inledande kartläggning
Vid den inledande kartläggningen görs en utvärdering av det tjänster som kan främja din integration.
Vid den inledande kartläggningen utreds t.ex. din utbildning, din arbetserfarenhet och dina språkkunskaper.
Den inledande kartläggningen görs vid arbets- och näringsbyrån eller vid kommunen.
Den kan också göras på ett annat ställe, t.ex. vid en läroinrättning.
Detta beror på vilken kommun du bor i.
Du kan framföra en begäran om en inledande kartläggning av din situation t.ex. till arbets- och näringsbyrån eller socialbyrån i din kommun.
Invandrarrådgivningen ger dig närmare information om den inledande kartläggningen och hur den ordnas i din hemkommun.
Om du behöver stöd för din integration, utarbetas en integrationsplan för dig efter den inledande kartläggningen.
En integrationsplan utarbetas för dig åtminstone om
du är arbetslös arbetssökande eller
får utkomststöd eller
du inte fyllt 18 år och inte har en vårdnadshavare i Finland.
I integrationsplanen antecknas åtgärder som främjar din integration.
Planen kan omfatta t.ex. studier i finska, andra studier eller arbetspraktik.
Du kan utarbeta en integrationsplan t.ex. med en arbetskraftsrådgivare vid arbets- och näringsbyrån, alltså TE-byrån (TE-toimisto), eller med en socialarbetare på socialbyrån.
Integrationsplanen ska utarbetas senast tre år efter att du fått ditt första uppehållstillstånd eller din uppehållsrätt registrerades.
Integrationsplanens längd beror på hur lång tid du behöver stöd för din integration.
Integrationsplanen gäller vanligen i högst tre år.
I vissa specialfall kan den gälla i fem år.
När en integrationsplan har utarbetats för dig, är det viktigt att du följer planen.
TE-byrån eller kommunen anvisar dig vid behov till integrationsutbildning.
I utbildningen ingår studier i finska eller svenska och introduktion i det finländska samhället och arbetslivet samt den finländska kulturen.
I utbildningen kan även andra studier och praktik ingå.
TE-byrån, FPA eller kommunen utreder din rätt till arbetslöshetstförmån eller utkomststöd under integrationsplanen.
Om du har en arbetsplats kan din arbetsgivare eventuellt stöda din integration.
Arbetsgivaren kan t.ex. betala avgifter för en kurs i finska för din räkning.
Ibland kan arbetsgivaren också hjälpa dig med praktiska ärenden, t.ex. leta efter en bostad åt dig.
Fråga mer om detta av din arbetsgivare.
linkkiArbets- och näringsministeriet:
Inledande kartläggning och integrationsplanfinska _ svenska _ engelska
Stöd till arbetslösa invandrarefinska _ svenska _ engelska
Integrationsutbildning
När en integrationsplan utarbetats kan du få integrationsutbildning.
Integrationsutbildning ordnas av kommuner, arbets- och näringsbyråer och många läroanstalter.
Arbets- och näringsbyrån eller kommunen hänvisar dig till integrationsutbildningen.
Integrationsutbildningen omfattar vanligen studier i finska eller svenska. I utbildningen bekantar du dig med det finländska samhället och arbetslivet och den finländska kulturen.
Studier i finska och svenska
På InfoFinlands sida Finska och svenska språket hittar du information om möjligheterna att studera finska eller svenska.
Din kultur i Finland
Din kultur, ditt språk och din religion kan fortfarande utgöra en viktig del av ditt liv också i Finland.
En invandrarförening kan hjälpa dig att bevara och utveckla din kultur.
I Finland finns många föreningar för invandrare.
Du hitar mer information om föreningar på InfoFinlands sida Föreningar.
Barn med invandrarbakgrund kan få undervisning i det egna modersmålet.
Du hitar mer information på InfoFinlands sida Grundläggande utbildning.
I Finland råder religionsfrihet (uskonnonvapaus).
Var och en har alltså rätt att bekänna och utöva sin religion.
Var och en får själv välja sin religion.
Om du vill, kan du låta att bli att välja en religion.
Du hittar mer information om religionsutövning i Finland på InfoFinlands sida Kulturer och religioner i Finland.
linkkiArbets- och näringsministeriet:
Guiden Välkommen till Finland(pdf, 3,40 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
linkkiArbets- och näringsbyrån:
Information om integrationfinska _ svenska _ engelska
linkkiArbets- och näringsbyrån:
Broschyren Jobba i Finland(pdf, 5,51 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ polska
Uppehållstillstånd
Studier i Finland
Boende
Arbete
Hälsa
Den sociala tryggheten
Utländsk examen i Finland
Uppehållstillstånd
Om du är medborgare i något av de nordiska länderna, ett EU-land, ett EES-land eller i Schweiz och kommer till Finland för att studera, måste du registrera din uppehållsrätt.
Läs mer på InfoFinlands sida EU-medborgare och Nordisk medborgare.
Om du är medborgare i något annat land behöver du ett uppehållstillstånd för studier.
Om dina studier i Finland pågår högst tre månader behöver du inget uppehållstillstånd.
Du kan ändå behöva ett visum.
Läs mer på InfoFinlands sida Att studera i Finland.
Information för utländska studerandeengelska
Studier i Finland
Du kan studera i Finland som utbytesstudent eller avlägga hela examen här.
Om du vill komma till Finland som utbytesstudent ska du kontakta till exempel studentexpeditionen eller den internationella enheten vid din egen läroanstalt.
På InfoFinlands sida Ansökan till utbildning hittar du information om hur du ansöker som examensstuderande till gymnasier, yrkesläroanstalter eller högskolor i Finland.
I Finland kan du studera på finska, svenska och ibland på engelska.
Högskolor ordnar engelskspråkig undervisning i vissa utbildningsprogram.
Läs mer på InfoFinlands sida Utländska studerande i Finland.
Boende
Om du är studerande kan du söka hyresbostäder som är speciellt avsedda för studerande.
Studentbostäder har ofta lägre hyra än vanliga bostäder.
Studentbostäder hyrs ut av studentbostadsstiftelser, universitetens studentkårer, nationer och vissa andra stiftelser.
Dessutom har vissa läroanstalter egna studenthem.
Fråga på din studieort var du kan söka en studentbostad.
Du kan söka bostad direkt när du blivit antagen till studier.
I de största städerna kan det ta flera veckor eller månader innan man får en bostad.
På InfoFinlands sida Boende hittar du mer information om hur du söker bostad och andra frågor i anslutning till boende.
Studentbostäderfinska _ engelska
Arbete
Om du är medborgare i ett EU-land, ett EES-land, Schweiz eller i något av de nordiska länderna, har du rätt att arbeta obegränsat under din studietid och du behöver inget särskilt tillstånd för det.
Arbete kan ge dig rätt till den sociala tryggheten i Finland.
Om du är medborgare i något annat land har du med ditt uppehållstillstånd för studerande rätt att arbeta i begränsad omfattning, om arbetet är
arbetspraktik som ingår i examen eller ett slutarbete eller
ett deltidsarbete, i genomsnitt högst 25 timmar per vecka under terminen
ett heltidsarbete under de tider då ingen undervisning ordnas vid läroanstalten, vanligen under sommar- och vinterlov.
På InfoFinlands sida Var hittar jag jobb? får du information om hur du söker arbete i Finland.
Studerandes rätt att arbetafinska _ svenska _ engelska
Hälsa
Om du kommer från ett annat nordiskt land till Finland för att studera har du rätt till sjukvård i Finland.
Du får vård på samma villkor och till samma kostnad som finländarna.
Ta med dig ett officiellt identitetsbevis när du använder hälsovårdstjänsterna.
Om du kommer från ett EU-land, ett EES-land eller Schweiz till Finland för att studera har du rätt till nödvändig sjukvård med det europeiska sjukvårdskortet.
Skaffa det europeiska sjukvårdskortet i ditt hemland innan du kommer till Finland.
Om du kommer från något annat land till Finland för att studera behöver du en omfattande sjukförsäkring innan du kan få uppehållstillstånd i Finland.
Mer information om uppehållstillstånd för studerande och om den sjukförsäkring som krävs för att få uppehållstillstånd får du på InfoFinlands sida Att studera i Finland eller på Migrationsverkets (Maahanmuuttovirasto) webbplats.
I Finland omfattas högskolestuderande av studerandehälsovården.
Fråga mer vid din egen läroanstalt.
Mer information om studerandehälsovården får du på Studenternas hälsovårdsstiftelses (SHVS) (YTHS) och social- och hälsovårdsministeriets (Sosiaali- ja terveysministeriö) webbplatser.
Du får information om hälsovårdstjänster i Finland på InfoFinlands sida Hälsa.
linkkiSHVS:
Hälsovård för högskolestuderandefinska _ svenska _ engelska
linkkiSocial- och hälsovårdsministeriet:
Studerandehälsovårdfinska _ svenska
Den sociala tryggheten
De flesta av FPA:s förmåner är sådana att du har rätt till dem endast om du flyttar ditt stadigvarande boende till Finland.
En studerande från ett land utanför EU/EES kan ha rätt till vissa av FPA:s förmåner, till exempel de förmåner som ingår i sjukförsäkringen.
Läs mer på InfoFinlands sida Den sociala tryggheten i Finland.
Social trygghet för dig som flyttar till Finlandfinska _ svenska _ engelska
Utländsk examen i Finland
Om du har avlagt en examen utomlands kan du ha nytta av jämställande av examen, erkännande av yrkeskompetens eller av att skaffa dig rätt till yrkesutövning eller en fristående examen.
På InfoFinlands sida Utländska examina i Finland hittar du information om hur du kan få din examen eller dina studier erkända i Finland.
linkkiUtbildningsstyrelsen:
Erkännande av en examenfinska _ svenska _ engelska
Finska medborgare har vissa rättigheter och skyldigheter som utlänningar bosatta i Finland inte nödvändigtvis har.
Rättigheter
rätt att få finskt pass
rätt att resa till Finland och vägra att bli utlämnad till ett annat land
rätt att rösta i presidentval, riksdagsval och folkomröstningar då man fyllt 18 år.
rätt att ställa upp som kandidat i riksdagsval då man fyllt 18 år.
möjlighet att bli utnämnd till sådana statliga ämbeten för vilka det krävs finskt medborgarskap
EU-medborgarnas rättigheter som rätten att fritt röra sig och arbeta inom EU:s område och rätten att rösta och ställa upp som kandidat i EU-val
Skyldigheter
Skyldighet att delta i landets försvar eller bistå i det.
Män som har fyllt 18 år har värnplikt (asevelvollisuus).
Skyldighet att följa Finlands lagar även annanstans än i Finland.
Finska medborgare kan i Finland dömas för brott som begåtts utomlands.
Observera att dessa är rättigheter och skyldigheter som ingår i det finska medborgarskapet.
Information om rättigheter och skyldigheter som gäller alla som är bosatta i Finland finns på InfoFinlands sida Dina rättigheter och skyldigheter i Finland.
Finska medborgares rättigheter och skyldigheterfinska _ svenska _ engelska
linkkiFörsvarsmakten:
Värnpliktfinska _ svenska _ engelska
Att ansöka om finskt passfinska _ svenska _ engelska
Att ansöka om finskt pass utomlandsfinska _ svenska _ engelska
Flytta till Finland
Fortsatt uppehållstillstånd
Studera finska språket
Arbete och studier
Äktenskap och samboförhållande
Social trygghet
Tjänster för barnfamiljer
Hälsa
Flytta till Finland
Om du inte är medborgare i ett nordiskt land, EU-medborgare eller familjemedlem till en EU-medborgare som är bosatt i Finland, behöver du ett uppehållstillstånd.
Läs mer på InfoFinlands sida Familjen till Finland.
Om du är EU-medborgare behöver du inte uppehållstillstånd i Finland.
Om du vistas i Finland mer än tre månader, behöver du ett registreringsintyg för EU-medborgare (Unionin kansalaisen rekisteröintitodistus).
Om du inte är EU-medborgare, men din familjemedlem som är bosatt i Finland är EU-medborgare, behöver du ett uppehållskort för familjemedlem (perheenjäsenen oleskelukortti).
Läs mer på InfoFinlands sida EU-medborgare.
Om du är medborgare i ett nordiskt land behöver du inte uppehållstillstånd i Finland.
Läs mer på InfoFinlands sida Medborgare i nordiska länder.
På InfoFinlands sida Komihåglista för dig som flyttar till Finland hittar du nyttig information om vilka andra saker du bör ta hand om innan du flyttar till Finland.
När du flyttar till Finland ska du besöka magistraten (maistraatti)på orten där du är bosatt.
Vid magistraten kan du få en finsk personbeteckning, om du inte fick den redan i samband med att du beviljades uppehållstillstånd eller din uppehållsrätt för EU-medborgare registrerades vid Migrationsverket.
På magistraten utreder man även om det är möjligt att registrera en hemkommun i Finland för dig.
När du har en hemkommun kan du använda kommunens tjänster, såsom till exempel hälsovårdstjänster.
Läs mer på InfoFinlands sida Hemkommun i Finland.
Till Finland på grund av familjebandfinska _ svenska _ engelska
Registrering av uppehållsrätt för EU-medborgarefinska _ svenska _ engelska
Registrering av utlänningarfinska _ svenska _ engelska
Fortsatt uppehållstillstånd
Om du har ett uppehållstillstånd ska du komma ihåg att ansöka om fortsatt uppehållstillstånd i god tid innan giltigheten för det första tillståndet tar slut.
Ansök om fortsatt uppehållstillstånd elektroniskt i tjänsten Enter Finland eller på Migrationsverkets tjänsteställe.
Tillståndsbeslutet är avgiftsbelagt.
Du måste betala avgiften samtidigt som du ansöker om fortsatt uppehållstillstånd.
Mer information om att ansöka om fortsatt uppehållstillstånd hittar du på InfoFinlands sida Fortsatt uppehållstillstånd.
Om du är EU-medborgare kan du ansöka om permanent uppehållsrätt när du har bott i Finland fem år.
Att förlänga uppehållstillståndetfinska _ svenska _ engelska
Studera finska språket
Information om studier i finska språket hittar du på InfoFinlands sida Finska och svenska språket.
Om du bor i Helsingforsregionen, Tammerforsregionen eller Åboregionen kan du leta efter en kurs i finska språket som passar dig genom tjänsten Finnishcourses.fi.
Kurser i finska och svenska språketfinska _ engelska _ ryska
Arbete och studier
Om du har uppehållstillstånd på grund av familjeband, har du rätt att arbeta och studera i Finland.
Även medborgare i EU-länder och nordiska länder och deras familjemedlemmar har rätt att arbeta och studera.
Notera att om du har ansökt om ditt första uppehållstillstånd i Finland så har du inte rätt att arbeta innan tillståndet har beviljats.
Om du är intresserad av att grunda ett eget företag, gå in på InfoFinlands sida Att grunda ett företag.
Information om studier i Finland hittar du på InfoFinlands sida Utbildning.
Äktenskap och samboförhållande
Om du ska gifta dig i Finland hittar du nyttig information på InfoFinlands sida Äktenskap.
Information om att leva i ett samboförhållande i Finland hittar du på InfoFinlands sida Samboförhållande.
Du hittar information om skilsmässa på InfoFinlands sida Skilsmässa.
Notera att om du har ett uppehållstillstånd som beviljats på basis av familjeband, så kan förändringar i familjeförhållandena, såsom till exempel skilsmässa, påverka ditt uppehållstillstånd.
Läs mer på InfoFinlands sida Kan jag förlora mitt uppehållstillstånd?
På InfoFinlands sida Problem i äktenskap och parförhållande hittar du information om var du kan söka hjälp för problem i förhållandet.
Social trygghet
De flesta av FPA:s förmåner är sådana att du har rätt till dem endast om du flyttar ditt stadigvarande boende till Finland.
Social trygghet för dig som flyttar till Finlandfinska _ svenska _ engelska
Tjänster för barnfamiljer
Information om de tjänster och stöd som samhället erbjuder barnfamiljer hittar du på InfoFinlands sida Ekonomiskt stöd till familjer och Vård av barnet.
Hälsa
I Finland finns både offentliga och privata hälsovårdstjänster.
De offentliga hälsovårdstjänsterna är förmånligare än de privata.
Om du har en hemkommun i Finland kan du använda offentliga hälsovårdstjänster.
Om du flyttar till Finland av familjeskäl får du vanligen en hemkommun i Finland.
Magistraten fattar beslut om registrering av hemkommun.
Läs mer på InfoFinlands sida Hälsovårdstjänster i Finland och Hemkommun i Finland.
Uppehållstillstånd
Fortsatt uppehållstillstånd
Arbete och företagande i Finland
Finska och svenska språket
Studier
Den sociala tryggheten
Hälsan
Uppehållstillstånd
Om du är medborgare i något av de nordiska länderna, ett EU-land, ett EES-land eller i Schweiz och kommer till Finland för att arbeta, behöver du inget uppehållstillstånd.
Läs mer på InfoFinlands sida Nordisk medborgare eller EU-medborgare.
Om du är medborgare i något annat land behöver du ett uppehållstillstånd för arbetstagare.
Om du redan befinner dig i Finland på någon annan grund kan du ha rätt att arbeta även om du inte har ansökt om ett uppehållstillstånd på grund av arbete.
Läs mer på InfoFinlands sida Till Finland för att arbeta.
Om du inte är medborgare i något av Europeiska unionens medlemsländer, ett EES-land eller i Schweiz och vill driva ett företag i Finland, behöver du ett uppehållstillstånd för företagare.
Mer information om uppehållstillstånd för företagare hittar du på InfoFinlands sida Bli företagare i Finland.
Arbete i Finlandfinska _ svenska _ engelska
Uppehållstillstånd för företagarefinska _ svenska _ engelska
Fortsatt uppehållstillstånd
Ansök om fortsatt uppehållstillstånd på internet i tjänsten Enter Finland eller på Migrationsverkets tjänsteställe.
Gör en ansökan innan ditt föregående uppehållstillstånd går ut.
Du får mer information om att ansöka om fortsatt uppehållstillstånd på InfoFinlands sida Fortsatt uppehållstillstånd.
Att förlänga uppehållstillståndetfinska _ svenska _ engelska
Arbete och företagande i Finland
I InfoFinlands avsnitt Arbete och företagande hittar du mycket information om arbetslivet och företagandet i Finland.
Finska och svenska språket
En del arbetsgivare ordnar undervisning i det finska språket för sina anställda.
Fråga din arbetsgivare som det ordnas undervisning i det finska språket på din arbetsplats.
Information om andra möjligheter att studera finska eller svenska hittar du i InfoFinlands avsnitt Finska och svenska språket.
Studier
Om du vill avlägga examen eller fortbilda dig kan du delta i fortbildning.
Fortbildning ordnas bland annat av läroanstalter, fackförbund och Institutet för Yrkenas befrämjande.
Också många arbetsplatser utbildar sina anställda till exempel i användningen av nya apparater eller program.
Studierna är inte alltid inriktade på att skaffa ett yrke.
Du kan också ha studier som hobby.
Läs mer på InfoFinlands sida Studier som hobby.
Grundläggande information om fortbildningfinska _ svenska
Den sociala tryggheten
Du kan omfattas av den finländska sociala tryggheten endera på basis av stadigvarande bosättning eller på basis av arbete.
De flesta av FPA:s förmåner är sådana att du har rätt till dem endast om du flyttar ditt stadigvarande boende till Finland.
Dessutom måste du uppfylla samma villkor för att få förmånen som alla andra som bor i Finland.
Om du flyttar till Finland för att arbeta, har du vanligtvis rätt till FPA:s förmåner under din anställning också när din anställning endast är kortvarig.
Om din lön uppgår till minst 696,60 € i månaden, har du rätt till de flesta av FPA:s förmåner.
Hur många timmar per vecka du arbetar eller hur lång din anställning är spelar ingen roll.
Om du har anställning i Finland, är det skäl för dig att ansluta dig till en finländsk arbetslöshetskassa.
Om du är medlem av en arbetslöshetskassa kan du få inkomstrelaterad arbetslöshetsersättning, om du blir arbetslös.
Läs mer på InfoFinlands sidor Fackförbund och Arbetslöshetsförsäkring.
Social trygghet för dig som flyttar till Finlandfinska _ svenska _ engelska
Hälsan
Hälsovård för anställda och företagare
Om du har kommit till Finland för att arbeta har du vanligen rätt att använda de offentliga hälsovårdstjänsterna i Finland.
Detta beror på hurdant och hur långt arbetsavtal du har samt från vilket land du har kommit till Finland.
Du kan begära att FPA utreder din rätt till de offentliga hälsovårdstjänsterna.
Du hittar mer information om den offentliga hälso- och sjukvården på InfoFinlands sida Hälsovårdstjänster i Finland.
I Finland är arbetsgivare skyldiga att ordna förebyggande företagshälsovård för sina anställda.
Företagare kan ordna sin egen företagshälsovård om de vill.
Företagare måste alltså inte ordna företagshälsovård för sig.
Företagare måste ändå ordna företagshälsovård för sina anställda.
Företagshälsovården kan ordnas vid den lokala hälsovårdscentralen eller till exempel på en privat läkarcentral.
Mer information får du på InfoFinlands sida Företagshälsovården och på social- och hälsovårdsministeriets webbplats.
linkkiSocial- och hälsovårdsministeriet:
Företagshälsovårdfinska _ svenska _ engelska
Om du förlorar ditt jobb
Om du har ett uppehållstillstånd för arbetstagare som endast gäller arbete för en viss arbetsgivare och du förlorar din arbetsplats, ska du ansöka om ett nytt uppehållstillstånd för arbetstagare eller ett uppehållstillstånd på andra grunder.
Om Migrationsverket har beviljat dig ett uppehållstillstånd för arbetstagare och din anställning upphör tidigare än uppehållstillståndet, måste du eller din arbetsgivare skriftligt meddela Migrationsverket att din anställning upphör.
Om ditt uppehållstillstånd för arbetstagare inte har begränsats att gälla arbete för en viss arbetsgivare, utan för en viss bransch och tillståndet är fortfarande giltigt, kan du byta jobb inom samma bransch.
Problem i arbetslivet
Om du råkar ut för problematiska situationer på arbetsplatsen ska du först kontakta din chef.
Om ärendet inte kan lösas på arbetsplatsen, ska du kontakta arbetarskyddsdistriktet (työsuojelupiiri) i ditt område eller ditt fackförbund.
Information och råd om var du kan få hjälp med olika slags problem i arbetslivet hittar du på InfoFinlands sida Problem i arbetslivet.
För att få finskt medborgarskap genom en medborgarskapsansökan krävs något av följande:
Du kan tillförlitligt intyga din identitet.
Du är minst 18 år gammal eller gift.
Du har bott i Finland tillräckligt länge.
Hur lång boendetid som krävs beror på din situation, vanligtvis ska du ha bott här minst 4–7 år.
Du har inte begått brott.
Du har inte lämnat till exempel skatter, böter, underhållsbidrag eller sjukhusavgifter obetalda.
Du kan redogöra för hur du försörjer dig i Finland.
Du kan finska, svenska eller det finska eller finlandssvenska teckenspråket åtminstone nöjaktigt.
Läs mer om att bevisa dina språkkunskaper på InfoFinlands sida Officiellt intyg över språkkunskaper.
Läs mer om att studera finska och svenska på InfoFinlands sida Finska och svenska språket.
Du kan ansöka om medborgarskap elektroniskt i tjänsten Enter Finland.
Fyll i en ansökan och lägg till bilagorna.
För en ansökan behöver du åtminstone följande dokument:
Ett giltigt identitetsbevis
En utredning om dina språkkunskaper
En utredning om ditt uppehälle.
Betala samtidigt också ansökningens handläggningsavgift.
När du fyllt i ansökningen i tjänsten har du tre månader på dig att styrka din identitet.
Boka en tid vid Migrationsverkets tjänsteställe på Migrationsverkets webbplats.
När du besöker tjänstestället för att styrka din identitet ska du ta med dig ditt identitetsbevis och ansökningsbilagorna i original.
Om du även ansöker om medborgarskap för ditt barn ska barnet följa med till tjänstestället för att styrka sin identitet.
När du fyllt i ansökningen, kom ihåg att följa ditt konto i Enter Finland-tjänsten.
Om Migrationsverket behöver ytterligare utredningar av dig, meddelas detta i Enter Finland-tjänsten.
Ansökningen kan avslås om du inte lämnar in begärda utredningar i tid.
När ett beslut har fattats får du ett meddelande.
Om du inte kan ansöka om medborgarskap elektroniskt eller inte vet hur man gör det kan du även ansöka om medborgarskap med en pappersblankett.
Skriv ut blanketten på Migrationsverkets webbplats och fyll i den färdigt.
Lämna den ifyllda ansökningen och ansökningsbilagorna personligen till Migrationsverkets tjänsteställe.
Mer information om medborgarskapsansökan och om annat som rör medborgarskap får du på Migrationsverkets webbplats.
Finskt medborgarskap är inte samma sak som uppehållstillstånd.
Om du först planerar att flytta till Finland, läs mer på InfoFinlands sida Flytta till Finland.
Att ansöka om finskt medborgarskapfinska _ svenska _ engelska
Barnets medborgarskapfinska _ svenska _ engelska
Medborgarskapsansökanfinska _ svenska _ engelska
Elektroniska tjänsterfinska _ svenska _ engelska
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Vem är asylsökande?
Asylsökandes uppehållsrätt
Social trygghet
Familjeåterförening
Hälsa
Vem är asylsökande?
En asylsökande (turvapaikanhakija) är en person som söker skydd och uppehållsrätt i en främmande stat.
Internationellt skydd kan beviljas om personen känner välgrundad fruktan för förföljelse (på grund av ras, religion, tillhörighet till en viss samhällsgrupp eller politisk samhörighet) eller om personen annars är utsatt för verklig fara i sitt hemland eller sitt permanenta bosättningsland.
En asylsökande är alltså inte en flykting (pakolainen).
Om en asylsökande beviljas flyktingstatus eller uppehållstillstånd på grund av skyddsbehov eller på någon annan grund får han eller hon stanna i Finland.
Broschyren Information till asylsökandefinska _ svenska _ engelska _ ryska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
Asylsökandes uppehållsrätt
Du får stanna i Finland om du beviljas asyl eller uppehållstillstånd på någon annan grund.
Om förhållandena i ditt hemland är sådana att du inte behöver asyl och det inte heller finns andra grunder att bevilja uppehållstillstånd, avslås din ansökan och du utvisas från Finland.
Om du får avslag på din asylansökan eller ansökan om uppehållstillstånd har du rätt att överklaga beslutet.
Läs mer på InfoFinlands sida Som asylsökande till Finland.
Att söka asyl i Finlandfinska _ svenska _ engelska
Social trygghet
Asylsökande har inte rätt till finskt socialskydd.
Detta innebär att de inte har rätt till FPA:s förmåner.
Mottagningscentralen betalar mottagningspenning till asylsökande.
Den utbetalas så länge som asylansökan behandlas.
Mottagningspenningen är ett litet belopp som är avsett för ofrånkomliga utgifter.
Om den asylsökande beviljas uppehållstillstånd och är fast bosatt i Finland har han eller hon rätt till finskt socialskydd.
Man kan ansöka om att omfattas av det finska socialskyddet av FPA då uppehållstillstånd har beviljats.
Familjeåterförening
Asylsökande har inte rätt till familjeåterförening.
Dina familjemedlemmar kan inte få uppehållstillstånd i Finland på grund av familjeband.
Om du får uppehållstillstånd i Finland kan dina familjemedlemmar ansöka om tillstånd på grund av familjeband.
Läs mer på InfoFinlands sida Till familjemedlem i Finland.
Att söka uppehållstillstånd på grund av familjebandfinska _ svenska _ engelska
Hälsa
Asylsökande har vanligtvis inte tillgång till offentlig hälsoåvård exempelvis på hälsocentraler.
Mottagningscentralen anordnar hälsovårdstjänster för asylsökande.
Hälsovårdare på mottagningscentralen ser till att asylsökande får den vård de behöver.
Fråga mer på din mottagningscentral.
Om du fått uppehållstillstånd och din hemkommun finns i Finland kan du använda tjänsterna inom den offentliga hälsovården på samma sätt som de övriga invånarna i kommunen.
Hälsovård för papperslösa
Global Clinic är en klinik där du kan få hjälp eller råd av en läkare eller sjukskötare om du vistas i Finland utan uppehållstillstånd.
Du kan besöka Global Clinic även om du inte behöver brådskande sjukvård.
Global Clinic bedriver verksamhet i följande städer:
Åbo
Tammerfors
Uleåborg
Joensuu
Du kan ringa eller skicka e-post.
En sjukskötare eller läkare besvarar ditt samtal.
Du hittar kontaktinformation på Global Clinic:s hemsidor.
Global Clinic:s tjänster är avgiftsfria för kunderna.
Global Clinic anmäler inte sina kunder till polisen eller andra myndigheter.
Klinikens adress eller öppettider meddelas inte offentligt.
Kontaktuppgifterfinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Arbetstagare, företagare, studerande, flykting, asylsökande eller en familjemedlem till en person bosatt i Finland hittar information speciellt om sin egen situation på dessa sidor i Infobanken.
Via dessa sidor hittar du snabbt den information som du behöver i kortfattade form.
Arbetstagare eller företagare
Studerande
Flykting
Asylsökande
Familjemedlem
Du kan få finskt medborgarskap
om du har en förälder som är finsk medborgare,
genom ansökan eller anmälan om medborgarskap.
I vissa undantagsfall kan man dessutom få medborgarskap på grundval av att man är född i Finland.
Ansöka om medborgarskap
Du kan ansöka om finskt medborgarskap när du har fyllt 18 år, har bott permanent i Finland i tillräckligt många år, har nöjaktiga muntliga och skriftliga kunskaper i finska eller svenska eller motsvarande kunskaper i finskt eller finlandssvenskt teckenspråk och din identitet är tillförlitligt utredd.
Det finns också andra villkor; till exempel måste du kunna visa hur du försörjer dig.
Du kan samtidigt ansöka om medborgarskap för ett minderårigt barn som du har vårdnaden om.
Om du har begått ett brott eller till exempel inte har betalat dina skatter, kan detta utgöra ett hinder för att få finskt medborgarskap.
Läs mer på InfoFinlands sida Hur kan man ansöka om finskt medborgarskap?
Finskt medborgarskap är inte samma sak som uppehållstillstånd.
Om du först planerar att flytta till Finland, läs mer på InfoFinlands sida Flytta till Finland.
Finskt medborgarskapfinska _ svenska _ engelska
Barnets medborgarskap
Samtidigt som du ansöker om medborgarskap för dig själv, kan du ansöka om det för ett minderårigt barn som du har vårdnaden om.
Läs mer på InfoFinlands sida Hur kan man ansöka om finskt medborgarskap?
Ett ofött barns medborgarskap
Barnet får automatiskt finskt medborgarskap vid födseln i följande fall:
Barnets mor är finsk medborgare.
Barnets far är finsk medborgare, men modern är inte det och föräldrarna är gifta med varandra.
Om föräldrarna inte är gifta, får barnet finskt medborgarskap av sin far enligt följande:
Vid födseln, då barnet föds i Finland och faderskapet bekräftas.
Genom medborgarskapsanmälan, då barnet föds i något annat land och faderskapet har bekräftats.
Också ett barn till utländska föräldrar som föds i Finland kan få finskt medborgarskap, om hen inte får medborgarskap i något annat land av sina föräldrar.
På InfoFinlands sida När ett barn föds i Finland finns mer information för föräldrar vars barn föds i Finland.
Barnets medborgarskapfinska _ svenska _ engelska
Finskt medborgarskap genom anmälan
Du kan få finskt medborgarskap genom medborgarskapsanmälan (kansalaisuusilmoitus) om du är
en före detta finska medborgare
utlänning och din far är finsk medborgare,
18–22 år och har bott i Finland i flera år
12–17 år och adoptivbarn till en finsk medborgare
medborgare i ett nordiskt land och har varit bosatt i Finland de senaste fem åren
Du kan göra en anmälan om medborgarskap på internet.
Fyll i blanketten i Enter Finland-tjänsten.
Lägg till bilagorna till ansökningen.
Betala samtidigt också ansökningens handläggningsavgift.
När du fyllt i anmälan, kom ihåg att följa ditt konto i tjänsten Enter Finland.
Du har tre månader på dig att styrka din identitet efter att du fyllt i blanketten i Enter Finland-tjänsten.
Du kan styrka din identitet vid Migrationsverkets tjänsteställe eller utomlands vid Finlands beskickning.
Fråga utrikesministeriet vilken beskickning du kan besöka för att styrka din identitet.
Boka en tid i förväg.
Ta med dig ett identitetsbevis och ansökningsbilagorna i original.
Om du inte kan göra din ansökan elektroniskt eller inte vet hur man gör det kan du också lämna in anmälan på en pappersblankett.
Mer information om hur du gör medborgarskapsanmälan hittar du på Migrationsverkets webbplats.
Medborgarskapsanmälanfinska _ svenska _ engelska
Flerfaldigt medborgarskap
Finland godkänner flerfaldigt medborgarskap, d.v.s. att du utöver ditt finska medborgarskap även har medborgarskap i ett annat land.
Alla stater godkänner dock inte flerfaldigt medborgarskap.
Innan du ansöker om finskt medborgarskap är det bra att ta reda på om flerfaldigt medborgarskap också är tillåtet i det land där du är medborgare.
Om denna stat inte tillåter flerfaldigt medborgarskap kan du förlora ditt nuvarande medborgarskap när du får finskt medborgarskap.
Flerfaldigt medborgarskap kan vara en fördel, men också en nackdel.
Det lönar sig att till exempel ta reda på om man tvingas göra värnplikten i flera medborgarskapsstater eller om det räcker med ett intyg över fullgjord värnplikt i ett land.
Flerfaldigt medborgarskap kan vara en fördel när man till exempel flyttar från ett land till ett annat.
Migrationsverket ger råd i frågor som rör medborgarskap:
Telefon 0295 419 626 tisdag, onsdag och fredag kl. 10.00–11.00
Barnets flerfaldiga medborgarskap
Barnet kan ha finskt medborgarskap och medborgarskap i något annat land.
Detta beror på huruvida det andra landet godkänner flerfaldigt medborgarskap för barnet.
Fråga mer om detta vid beskickningen för ditt eget land.
Kan man förlora sitt finska medborgarskap?
Man kan förlora sitt finska medborgarskap om man
är 22 år gammal, har medborgarskap också i en annan stat och saknar tillräcklig anknytning till Finland
har angett felaktiga uppgifter i medborgarskapsansökan eller medborgarskapsanmälan
har förvärvat sitt medborgarskap på grund av faderns finska medborgarskap och faderskapet upphävs.
Att förlora sitt finska medborgarskapfinska _ svenska _ engelska
Vem är flykting?
Familjeåterförening
Eftersökning av försvunna anhöriga
Hälsa
Stöd för flyktingar
Vem är flykting?
En flykting är en person med flyktingstatus.
Flyktingstatus får de som beviljas asyl eller som tas till Finland i flyktingkvoten.
Kvotflyktingar
Man kan inte ansöka om att bli kvotflykting (kiintiöpakolainen) via myndigheterna i Finland.
Man kan inte heller föreslå en annan person, till exempel en släkting eller vän, som kvotflykting.
Finland tar som kvotflyktingar emot personer som har flyktingstatus enligt
Förenta nationernas flyktingorganisation UNHCR. Kvotflyktingarna väljs bland de personer som UNHCR föreslår till Finland.
De finländska myndigheterna intervjuar flyktingarna som UNHCR har föreslagit och väljer bland dem de personer som tas emot till Finland.
Intervjuerna görs i de länder där flyktingarna vistas, vanligen i flyktingläger eller i UNHCR:s lokaler.
Valet av kvotflyktingar påverkas till exempel av följande faktorer:
Flyktingen är i behov av internationellt skydd.
Flyktingens mänskliga rättigheter förverkligas inte i det land där han eller hon vistas.
Flyktingen utgör inget hot för Finlands säkerhet.
Flyktingen har förutsättningar att integreras i Finland.
En del flyktingar väljs utan intervju på basis av UNHCR:s dokument.
Dessa är vanligen nödfall, med andra ord flyktingar som är i ett brådskande behov av asyl till exempel av hälsorelaterade eller politiska orsaker.
Finlands riksdag beslutar hur många flyktingar som tas till landet.
Från och med år 2001 har Finlands flyktingkvot varit 750 personer per år.
Inrikesministeriet beslutar från vilka länder kvotflyktingarna tas.
Beviljande av flyktingstatus till asylsökande
En person kan erhålla flyktingstatus också genom att söka asyl i Finland.
Asylsökanden kan beviljas flyktingstatus om han eller hon har befogade skäl att frukta förföljelse i sitt hemland på grund av ras, religion, nationalitet, tillhörighet till en viss samhällsgrupp eller på grund av sin politiska uppfattning och då sökanden på grund av detta inte kan återvända till sitt hemland.
Asylsökande som inte beviljas flyktingstatus kan ändå få uppehållstillstånd i Finland på någon annan grund.
Läs mer på InfoFinlands sida Som asylsökande till Finland.
Information om val av kvotflyktingarfinska _ svenska _ engelska
Familjeåterförening
Också flyktingens familjemedlemmar kan få uppehållstillstånd i Finland.
Vilka som är familjemedlemmar definieras i lagen.
Endast dessa familjemedlemmar kan få uppehållstillstånd på grund av familjeband.
I Finland betraktas som familjemedlemmar
registrerad partner
sambo
vårdnadshavaren till ett barn under 18 år.
För att familjemedlemmarna ska kunna få uppehållstillstånd, krävs det i vissa fall att flyktingen har en tillräcklig inkomst för att försörja sina familjemedlemmar i Finland.
Mer information om familjeåterförening finns på InfoFinlands sida Till familjemedlem i Finland.
Hjälp med familjeåterföreningen
Om du har kommit till Finland som kvotflykting, kan Migrationsverket ersätta kostnaderna för en familjemedlems inresa.
Kostnaderna ersätts dock endast i de fall där familjebandet har funnits redan före du fick ditt första uppehållstillstånd i Finland.
Andra anhörigas resekostnader ersätts inte.
Endast kvotflyktingar kan få ersättning för familjemedlemmarnas resekostnader.
Finlands Rösa Kors hjälper med researrangemangen för kvotflyktingar
Migrationsverket ersätter resekostnaderna endast i det fall att familjemedlemmen reser till Finland på en resa som arrangeras av Finlands Röda Kors och Internationella organisationen för migration.
Finlands Röda Kors hjälper med att ordna resan till Finland för kvotflyktingens familjemedlemmar när dessa fått uppehållstillstånd.
Röda Korset ger också rådgivning om reglerna för familjeåterförening och därom, hur familjemedlemmarna ska gå tillväga för att ansöka om familjeåterförening.
När Migrationsverket har gett ett positivt beslut på din ansökan om återförening på grund av familjeband och anser att staten kan bekosta resan för dina familjemedlemmar, skickar det sitt beslut till Röda Korset.
Om du har kommit till Finland som kvotflykting och vill att finska staten bekostar resan för dina familjemedlemmar ska du ta kontakt med Röda Korsets beredskapsenhet som sätter igång researrangemangen.
Finlands Röda Kors kan inte bistå familjemedlemmarnas flygresor eller andra resor ekonomiskt.
Att söka uppehållstillstånd på grund av familjebandfinska _ svenska _ engelska
Familjemedlem till en flyktingfinska _ svenska _ engelska
Eftersökning av försvunna anhöriga
Om du vill ha kontakt med en anhörig som försvunnit kan du be om hjälp vid personefterforskningen vid Finlands Röda Kors.
Röda Korset hjälper familjer som skilts åt vid olika katastrofer eller kriser.
Röda Korset söker försvunna anhöriga och förmedlar meddelanden på krisområden.
linkkiFinlands Röda Kors:
Efterforskning av anhörigafinska _ svenska _ engelska _ franska _ somaliska
linkkiFinlands Röda Kors:
Efterforskning av anhörigafinska _ svenska _ engelska _ ryska _ somaliska _ spanska _ persiska _ arabiska _ portugisiska
Hälsa
Om du har kommit till Finland som kvotflykting, har du hemkommun i Finland och då kan du använda de offentliga hälsovårdstjänsterna.
Stöd för flyktingar
Flyktingar och asylsökande kan söka hjälp och rådgivning i juridiska frågor bland annat vid Flyktingrådgivningen r.f. eller rättshjälpsbyråerna (oikeusaputoimisto).
Flyktingrådgivningen ger asylsökande rättshjälp i asylprocessens första skede.
Flyktingrådgivningen ger också andra utlänningar allmän rättshjälp.
Rättshjälpsbyråerna ger personer som är bosatta i Finland expertråd i skötseln av juridiska ärenden.
För att sköta ett juridiskt ärende kan man få ett rättsbiträde bekostat antingen helt eller delvis med statliga medel.
Finlands flyktinghjälp r.f. är en organisation som arbetar för att främja flyktingarnas grundläggande rättigheter.
Organisationens verksamhet i Finland omfattar informering, utbildning och socialarbete.
Flyktinghjälpen hjälper flyktingar och invandrare till exempel i frågor som rör integrationen, boendet och grundandet av egna organisationer.
linkkiFinlands flyktinghjälp r.f.:
Stöd till flyktingarfinska _ svenska _ engelska
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Före flytten till Finland
Efter flytten till Finland
Bekanta dig med innehållen i InfoFinland före flytten.
I InfoFinland hittar du pålitlig information på ditt eget språk om flytten till Finland, arbetslivet, boende, studier i finska eller svenska språket, utbildning, social trygghet, hälsotjänster, tjänster för familjer, problematiska situationer och fritid.
På sidorna finns nyttiga praktiska råd, kontaktuppgifter och länkar till tilläggsinformation.
Med hjälp av menyn Städer får du fram information om den kommun som du är intresserad av.
De olika språkversionerna av InfoFinlands är identiska.
Komihåglistan för dig som flyttar till Finland är avsedd att hjälpa dig med de viktigaste praktiska frågorna som har med flytten att göra.
Observera att listan inte nödvändigtvis innehåller allt som måste göras när du flyttar till Finland.
Före flytten till Finland
Uppehållstillstånd eller registrering av uppehållsrätt?
Om du ska vistas i Finland mer än 90 dagar och är EU-medborgare, måste du registrera din uppehållsrätt.
Om du är medborgare i ett land utanför EU, måste du ansöka om uppehållstillstånd i Finland.
Läs mer på InfoFinlands sida EU-medborgare eller Icke-EU-medborgare.
När du ansöker om uppehållstillstånd eller registrering av uppehållsrätten måste du bevisa att din utkomst i Finland är tryggad.
Om du kommer till Finland för att arbeta eller som företagare måste du bevisa att ditt arbete eller din företagsverksamhet inbringar dig en tillräcklig utkomst.
Om du flyttar till en familjemedlem i Finland, krävs det ofta även att den person som bor i Finland har tillräckliga medel för att försörja sig själv och den familjemedlem som flyttar till Finland.
Flyttsaker från EU-området
Om du flyttar till Finland från ett annat EU-land behöver du vanligen inte betala tull eller mervärdesskatt på dina flyttsaker, d.v.s. de personliga föremål som du tar med dig.
Du behöver inte heller anmäla dina flyttsaker i tullen (tulli).
Observera att tull- och skattefriheten för flyttsaker inte gäller alkohol eller tobaksprodukter.
För import av dessa gäller separata begränsningar.
Mer information får du på Tullrådgivningen +358 (0)295 5201 eller på tullens webbplats.
Tullrådgivningen betjänar på finska, svenska och engelska.
Flyttsaker från länder utanför EU
Om du flyttar till Finland från ett land som inte hör till EU behöver du vanligen inte betala tull eller mervärdesskatt på dina flyttsaker, d.v.s. de personliga föremål som du tar med dig.
Du måste dock göra en tullanmälan på flyttsakerna till de finländska tullmyndigheterna.
Som flyttsaker betraktas till exempel:
möbler och andra husgeråd
husdjur
cyklar och motorcyklar
bilar och släpvagnar avsedda för privat bruk.
Observera att tull- och skattefriheten för flyttsaker inte gäller alkohol eller tobaksprodukter.
För import av dessa gäller separata begränsningar.
linkkiTullen:
Införsel av flyttsaker till Finlandfinska _ svenska _ engelska _ ryska
Införsel av bil till Finland som flyttsak
När du tar med dig en bil till Finland som flyttsak, måste du tullanmäla den.
Om du tar med dig en bil till Finland måste du registrera den och betala bilskatt (autovero) för den innan du kan använda den i trafiken.
Man kan dock använda bilen tillfälligt innan bilskatten är betald.
Detta förutsätter att du har gjort en anmälan om ibruktagande av fordonet (auton käyttöönottoilmoitus) till skatteförvaltningen.
Du ska också ha en giltig trafikförsäkring (liikennevakuutus) för din bil i Finland.
Om du för in en bil från ett land utanför EES-området behöver du också ett förflyttningstillstånd innan du kan använda bilen.
Förflyttningstillstånd beviljas av besiktningskontor och vissa av Tullens verksamhetsställen.
Du får inte använda din bil i Finland förrän du har gjort en anmälan om ibruktagande av fordonet och skaffat ett förflyttningstillstånd.
Om du har frågor kring fordonsskatten eller anmälan om ibruktagande, kan du ringa skatteförvaltningens telefontjänst:
+358 (0)29 497 150 (finska)
+358 (0)29 497 151 (svenska)
+358 (0)29 497 152 (engelska)
linkkiTullen:
Fordon som flyttgodsfinska _ svenska _ engelska _ ryska
Införsel av sällskapsdjur
Mer information om reglerna i Finland ges av Livsmedelsverket (Ruokavirasto).
linkkiLivsmedelsverket:
Införsel av djur från EU-länderfinska _ svenska _ engelska
linkkiLivsmedelsverket:
Införsel av djur från länder utanför EUfinska _ svenska _ engelska
Flyttfirmor
En del företag som tillhandahåller flyttservice sköter också flytt från ett land till ett annat.
Du kan anlita dessa företag att transportera dina ägodelar från ett land till ett annat och också att packa dina saker och tillhandahålla förpackningsmaterial.
Flyttkostnaderna beror på varifrån du flyttar och hur mycket saker du har.
Tjänsterna och priserna i olika flyttfirmor kan variera stort och därför lönar det sig att jämföra.
Flyttjänsterfinska _ svenska _ engelska
linkkiViktor Ek:
Flyttjänsterfinska _ svenska _ engelska
Hjälp när du flyttarfinska _ svenska _ engelska _ norska
_ danska
Efter flytten till Finland
I den här listan har vi samlat de vanligaste ärendena som du måste ta hand om när du har kommit till Finland.
Bostad och hemförsäkring
De flesta invandrare bor först i en hyresbostad när de kommer till Finland.
Det är bra att reservera minst en månad för att söka hyresbostad.
Läs mer på InfoFinlands sida Boende.
När du har en bostad är det bra att också ta en hemförsäkring (kotivakuutus).
Hemförsäkringen ersätter till exempel skador på möbler och andra ägodelar.
Hemförsäkringar säljs av försäkringsbolag.Information om försäkringar finns på InfoFinlands sida Vardagslivet i Finland.
Finsk personbeteckning
Om du får ett uppehållstillstånd i Finland registreras du automatiskt i det finska befolkningsdatasystemet.
Du får samtidigt även en finsk personbeteckning.
I Finland kan du få personbeteckningen även vid magistraten eller skattebyrån på din hemort.
Läs mer på InfoFinlands sida Registrering som invånare.
Hemkommun i Finland
Om du flyttar till och blir stadigvarande bosatt i Finland registreras en hemkommun för dig i Finland.
Hemkommunen är den kommun där du bor.
När du har en hemkommun har du rätt att använda denna kommuns tjänster såsom till exempel offentliga hälsovårdstjänster.
Du kan ta reda på om det är möjligt att registrera en hemkommun i Finland för dig vid magistraten på din hemort.
Läs mer på InfoFinlands sida Hemkommun i Finland.
Registrering av utlänningarfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Registrering av utlänningar på skattebyrånfinska _ svenska _ engelska
Social trygghet
Du kan omfattas av den finländska sociala tryggheten endera på basis av stadigvarande bosättning eller på basis av arbete.
De flesta av FPA:s förmåner är sådana att du har rätt till dem endast om du flyttar ditt stadigvarande boende till Finland.
Dessutom måste du uppfylla samma villkor för att få förmånen som alla andra som bor i Finland.
Social trygghet för dig som flyttar till Finlandfinska _ svenska _ engelska
Bankkonto
Du behöver ett bankkonto för att sköta din dagliga ekonomi.
När du öppnar ett bankkonto behöver du ett pass eller någon annan officiell identitetshandling.
Det lönar sig att jämföra tjänsterna och priserna som olika banker tillhandahåller så att du hittar det alternativ som är förmånligast för dig.
Information om att öppna ett bankonto finns på InfoFinlands sida Vardagslivet i Finland.
linkkiFinansbranschens Centralförbund:
Utländska medborgares bankärendenfinska _ engelska
Skattekort
Om du arbetar och får lön eller är företagare behöver du ett finskt skattekort (verokortti).
Skattekortet får du vid skattebyrån.
Läs mer om beskattningen i Finland på InfoFinlands sida Beskattning.
Kollektivtrafik
Om du bor i en stad är det inte nödvändigt att äga en bil.
Kollektivtrafiken fungerar väl i Finland.
Man kan resa nästan över allt i Finland med tåg eller buss.
Man kan också flyga till många städer.
I stora städer och deras näromgivning finns en välfungerande lokaltrafik.
Lokaltrafiken trafikeras vanligtvis med bussar.
Läs mer på InfoFinlands sida Trafiken i Finland.
Körkort
Om du har ett körkort som utfärdats i ett av de nordiska länderna eller i ett EU-/EES-land, är det giltigt även i Finland.
Om du bor stadigvarande i Finland kan du byta ut kortet mot ett finländskt körkort.
Om du har ett körkort som utfärdats i ett land som är anslutet till Genève- eller Wien-konventionerna kan du köra med detta kort högst två år i Finland.
Du måste byta ut ditt körkort mot ett finländskt körkort inom två år efter att du flyttat till Finland.
Om du har ett körkort som utfärdats i ett land som inte är anslutet till Genève- eller Wien-konventionerna kan du köra bil med detta kort under ett års tid efter att ha registrerats i befolkningsregistret i Finland.
Du kan byta ut ditt körkort till ett finskt körkort på Ajovarmas serviceställe.
linkkiTrafiksäkerhetsverket:
Utländskt körkort i Finlandfinska _ svenska _ engelska
Internet
I Finland kan du sköta många ärenden via Internet.
Det är bra att skaffa sig en Internetuppkoppling så fort som möjligt efter att du har flyttat till Finland.
På InfoFinlands sida Vardagslivet i Finland finns mer information om att skaffa en internetuppkoppling.
linkkiKommunikationsverket:
Internet- och telefonabonnemangfinska _ svenska _ engelska
Telefon
När du köper ett telefonabonnemang i Finland får du ett finskt telefonnummer.
Många företag erbjuder telefonabonnemang.
Du kan också köpa ett prepaid-abonnemang.
Prepaid-kortet är i förväg laddat med en summa som man sedan kan ringa för.
Prepaid-abonnemang kan köpas till exempel i R-kiosker, en del snabbköp och på Internet.
linkkiSkype:
Förmånliga utlandssamtalfinska _ svenska _ engelska _ ryska _ estniska _ franska _ spanska _ turkiska _ kinesiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ rumänska _ ungerska _ japanska _ italienska
_ danska
_ bulgariska
_ grekiska
_ tjeckiska
Hälsa
I Finland finns offentliga och privata hälsovårdstjänster.
Du kan använda de offentliga hälsovårdstjänsterna om du har en hemkommun i Finland.
Till de offentliga hälsovårdstjänsterna hör till exempel hälsocentralerna.
De offentliga tjänsterna är förmånligare än de privata.
Om du vill reservera tid till en läkare ska du ta kontakt med hälsocentralen.
Om du inte har rätt att använda de offentliga hälsovårdstjänsterna kan du kontakta en privat läkarcentral.
Mer information om hälsovården i Finland får du på InfoFinlands sida Hälsa.
Språkstudier
Finlands officiella språk är finska och svenska.
Språkkunskaper hjälper dig att förstå det nya samhället och underlättar skötseln av ärenden.
Mer information hittar du på InfoFinlands sida Finska och svenska språket.
Jobbsökning
Arbets- och näringsbyrån hjälper dig i jobbsökningen.
Du kan söka jobb på Internet och via tidningar.
Du kan också hitta ett jobb genom att själv kontakta arbetsgivare som du är intresserad av.
Läs mer om jobbsökning i Finland på InfoFinlands sida Var hittar jag jobb?
Fritid och hobbyer
Information om möjligheter till fritidsaktiviteter hittar du på InfoFinlands sida Fritid.
linkkiExpat Finland:
Information om Finland för utlänningarengelska
På den här sidan finns information om den bosättningsbaserade sociala tryggheten som hör till FPA:s ansvarsområde.
På sidan finns information om de situationer då du betraktas ha rätt till den sociala trygghet som grundar sig på boende.
På InfoFinlands sida Utkomstskydd för arbetslösa får du mer information om vem som har rätt till utkomstskydd för arbetslösa.
FPA har bland annat hand om folkpensionen, barnbidrag, det grundläggande utkomstskyddet för arbetslösa, sjuk- och föräldradagpenningar, utkomststöd och rehabilitering.
FPA sköter även de sjukvårdsersättningar som betalas för privat sjukvård.
Grunderna för FPA:s bidrag definieras i lagen.
Du måste ansöka separat om att omfattas av den sociala tryggheten i Finland.
Du måste också separat söka de enskilda bidragen.
Varje sökandes livssituation behandlas individuellt när FPA fattar beslut om bidrag.
Sökandens livssituation och behov av understöd är ofta mycket olika.
Därför varierar även bidragens belopp och grunder.
Du ska alltid utreda din egen situation individuellt.
Offentliga hälso- och sjukvårdstjänster samt socialtjänster är kommunernas ansvar i Finland.
Läs mer på InfoFinlands sida Hälsovårdstjänster i Finland.
Mer information om rätten till hemkommun finns på InfoFinlands sida Hemkommun i Finland.
Information om social trygghetfinska _ svenska _ engelska
Social trygghet för dig som flyttar till Finland(pdf, 560 kb)finska _ svenska _ engelska _ ryska _ estniska
Information om sjukförsäkringfinska _ svenska _ engelska
linkkiSocial- och hälsovårdsministeriet:
Information om den sociala tryggheten i Finlandengelska
Att höra till den sociala tryggheten i Finland
Huvudregeln är att du omfattas av den sociala tryggheten i Finland och har rätt till FPA:s förmåner om du bor stadigvarande i Finland.
Vad stadigvarande boende betyder definieras i lagen.
Du kan också få rätt till den sociala tryggheten i Finland genom att arbeta i Finland.
Omfattas du av den sociala tryggheten och kan du få bidrag?
På detta inverkar om du flyttar till Finland från
ett nordiskt land
ett land inom Europeiska unionen (EU), ett land inom det Europeiska ekonomiska samarbetsområdet (EES) eller Schweiz eller
EES-länderna är Europeiska unionens medlemsländer samt Norge, Island och Liechtenstein.
Huruvida du omfattas du av den sociala tryggheten och kan få bidrag påverkas också av om du flyttar till Finland till exempel som
arbetstagare eller företagare
studerande
familjemedlem
utsänd arbetstagare.
Finland har ingått avtal om den sociala tryggheten med ett antal länder.
Dessa länder är de nordiska länderna (Sverige, Danmark, Norge och Island), USA, Kanada och Quebec, Chile, Israel, Indien och Australien.
Avtalen rör främst pensioner.
En del avtal gäller även sjukvård.
Om du kommer från ett av dessa länder ska du kontrollera hos FPA om avtalen påverkar din sociala trygghet.
Lag om hemkommunfinska _ svenska
Information om internationella socialskyddsavtalfinska _ svenska _ engelska
Information om den sociala tryggheten i Finland för EU-medborgarefinska _ svenska _ engelska
Stadigvarande flytt till Finland och stadigvarande boende i Finland
När du flyttar till Finland bedömer FPA alltid först om din flytt till Finland är stadigvarande boende i den mening som avses i lagarna om social trygghet.
(Det är bra att veta att stadigvarande boende definieras på olika sätt i olika lagar.
Här menas lagar om social trygghet.)
Om ditt boende i Finland inte anses stadigvarande, kan du ändå ha rätt att omfattas av den sociala tryggheten i Finland på grund av att du arbetar.
Din flytt till Finland kan betraktas som stadigvarande i följande situationer:
du är återflyttare, det vill säga återvänder till Finland från utlandet
du har ett arbetsavtal eller motsvarande avtal för ett arbete som du utför i Finland
du är gift eller annars i ett nära familjeförhållande till en person som redan bor stadigvarande i Finland.
Dessutom krävs det i allmänhet att ditt uppehållstillstånd har beviljats för minst ett år, om du är skyldig att ha ett uppehållstillstånd.
Din situation bedöms i sin helhet.
På basis av bedömningen beslutas om boendet är stadigvarande eller inte.
Om du flyttar till Finland tillfälligt har du vanligtvis inte rätt till den sociala tryggheten i Finland.
Till exempel befinner sig en studerande vars enda orsak till vistelsen i landet är studierna tillfälligt i Finland.
När ett beslut fattats att ditt boende i Finland är stadigvarande, anses du bo stadigvarande i Finland så länge som
du har din egentliga bostad och ditt hem här och så länge du huvudsakligen vistas här
eller
du har en annan grund för den stadigvarande vistelsen, till exempel ett familjeband eller arbete.
Om du emellertid börjar arbeta i ett annat land eller reser utomlands för över ett år, kan din rätt till den sociala tryggheten i Finland upphöra.
Mer information om sådana situationer får du vid FPA.
Det finns även bidrag som du inte kan få om du inte bor stadigvarande i Finland eller har gjort det tidigare.
Till exempel kan föräldrar få föräldradagpenning endast om de har bott i Finland minst 180 dagar före barnets beräknade födelsedatum.
Om du kommer från ett annat EU-land kan du i vissa fall utnyttja de försäkringsperioder som du har ackumulerat i andra EU-länder.
Fråga mer hos FPA.
Social trygghet för dig som flyttar till Finlandfinska _ svenska _ engelska
Flytt utomlands och social trygghetfinska _ svenska _ engelska
Kontaktuppgifter till FPAfinska _ svenska _ engelska
Arbete ger dig åtminstone delvis rätt till den sociala tryggheten i Finland
EU-länderna, EES-länderna och Schweiz
Om du flyttar till Finland för att arbeta från EU-området eller ett EES-land eller Schweiz, omfattas du vanligtvis av den sociala tryggheten i Finland under din anställning, även när din anställning är kortvarig.
Exempel:
Om du kommer till Finland för att arbeta under fyra månader, kan du ha rätt till hemvårdsstöd för barn och den offentliga hälsovården.
Om din anställning varar fyra månader eller längre, omfattas du av den sociala tryggheten i Finland under tiden för din anställning.
Övriga länder
Om du kommer till Finland som arbetstagare någon annanstans ifrån än ett EU-land, ett EES-land eller Schweiz påverkas din sociala trygghet av följande faktorer:
hur länge arbetet varar
från vilket land du flyttar till Finland.
De flesta av FPA:s förmåner är sådana att du har rätt till dem endast om du flyttar ditt stadigvarande boende till Finland eller om din anställning varar i minst fyra månader.
Dessutom måste du uppfylla samma villkor för att få förmånen som alla andra som bor i Finland.
Om du inte flyttar stadigvarande till Finland, omfattas du vanligen av den sociala tryggheten i Finland så länge din anställning varar.
Anställningen ska vara minst fyra månader lång och din arbetstid och lön ska vara tillräcklig.
Därtill behöver du ett uppehållstillstånd som omfattar rätt att arbeta.
Minimiarbetstiden är vanligtvis 18 timmar i veckan.
Lönen ska vara minst i enlighet med kollektivavtalet eller om inget kollektivavtal finns, uppgå till minst 1211 euro per månad (år 2019).
Arbetstagaren och den sociala tryggheten i Finlandfinska _ svenska _ engelska
Asylsökande
Asylsökande har inte rätt till finskt socialskydd.
Detta innebär att de inte har rätt till FPA:s förmåner.
Mottagningscentralen betalar mottagningspenning till asylsökande.
Den utbetalas så länge som asylansökan behandlas.
Mottagningspenningen är ett litet belopp som är avsett för ofrånkomliga utgifter.
Om den asylsökande beviljas uppehållstillstånd och är fast bosatt i Finland har han eller hon rätt till finskt socialskydd.
Man kan ansöka om att omfattas av det finska socialskyddet av FPA då uppehållstillstånd har beviljats.
Uppehållstillstånd
Studier i Finland
Boende
Arbete
Hälsa
Den sociala tryggheten
Utländsk examen i Finland
Uppehållstillstånd
Om du är medborgare i något av de nordiska länderna, ett EU-land, ett EES-land eller i Schweiz och kommer till Finland för att studera, måste du registrera din uppehållsrätt.
Läs mer på InfoFinlands sida EU-medborgare och Nordisk medborgare.
Om du är medborgare i något annat land behöver du ett uppehållstillstånd för studier.
Om dina studier i Finland pågår högst tre månader behöver du inget uppehållstillstånd.
Du kan ändå behöva ett visum.
Läs mer på InfoFinlands sida Att studera i Finland.
Information för utländska studerandeengelska
Studier i Finland
Du kan studera i Finland som utbytesstudent eller avlägga hela examen här.
Om du vill komma till Finland som utbytesstudent ska du kontakta till exempel studentexpeditionen eller den internationella enheten vid din egen läroanstalt.
På InfoFinlands sida Ansökan till utbildning hittar du information om hur du ansöker som examensstuderande till gymnasier, yrkesläroanstalter eller högskolor i Finland.
I Finland kan du studera på finska, svenska och ibland på engelska.
Högskolor ordnar engelskspråkig undervisning i vissa utbildningsprogram.
Läs mer på InfoFinlands sida Utländska studerande i Finland.
Boende
Om du är studerande kan du söka hyresbostäder som är speciellt avsedda för studerande.
Studentbostäder har ofta lägre hyra än vanliga bostäder.
Studentbostäder hyrs ut av studentbostadsstiftelser, universitetens studentkårer, nationer och vissa andra stiftelser.
Dessutom har vissa läroanstalter egna studenthem.
Fråga på din studieort var du kan söka en studentbostad.
Du kan söka bostad direkt när du blivit antagen till studier.
I de största städerna kan det ta flera veckor eller månader innan man får en bostad.
På InfoFinlands sida Boende hittar du mer information om hur du söker bostad och andra frågor i anslutning till boende.
Studentbostäderfinska _ engelska
Arbete
Om du är medborgare i ett EU-land, ett EES-land, Schweiz eller i något av de nordiska länderna, har du rätt att arbeta obegränsat under din studietid och du behöver inget särskilt tillstånd för det.
Arbete kan ge dig rätt till den sociala tryggheten i Finland.
Om du är medborgare i något annat land har du med ditt uppehållstillstånd för studerande rätt att arbeta i begränsad omfattning, om arbetet är
arbetspraktik som ingår i examen eller ett slutarbete eller
ett deltidsarbete, i genomsnitt högst 25 timmar per vecka under terminen
ett heltidsarbete under de tider då ingen undervisning ordnas vid läroanstalten, vanligen under sommar- och vinterlov.
På InfoFinlands sida Var hittar jag jobb? får du information om hur du söker arbete i Finland.
Studerandes rätt att arbetafinska _ svenska _ engelska
Hälsa
Om du kommer från ett annat nordiskt land till Finland för att studera har du rätt till sjukvård i Finland.
Du får vård på samma villkor och till samma kostnad som finländarna.
Ta med dig ett officiellt identitetsbevis när du använder hälsovårdstjänsterna.
Om du kommer från ett EU-land, ett EES-land eller Schweiz till Finland för att studera har du rätt till nödvändig sjukvård med det europeiska sjukvårdskortet.
Skaffa det europeiska sjukvårdskortet i ditt hemland innan du kommer till Finland.
Om du kommer från något annat land till Finland för att studera behöver du en omfattande sjukförsäkring innan du kan få uppehållstillstånd i Finland.
Mer information om uppehållstillstånd för studerande och om den sjukförsäkring som krävs för att få uppehållstillstånd får du på InfoFinlands sida Att studera i Finland eller på Migrationsverkets (Maahanmuuttovirasto) webbplats.
I Finland omfattas högskolestuderande av studerandehälsovården.
Fråga mer vid din egen läroanstalt.
Mer information om studerandehälsovården får du på Studenternas hälsovårdsstiftelses (SHVS) (YTHS) och social- och hälsovårdsministeriets (Sosiaali- ja terveysministeriö) webbplatser.
Du får information om hälsovårdstjänster i Finland på InfoFinlands sida Hälsa.
linkkiSHVS:
Hälsovård för högskolestuderandefinska _ svenska _ engelska
linkkiSocial- och hälsovårdsministeriet:
Studerandehälsovårdfinska _ svenska
Den sociala tryggheten
De flesta av FPA:s förmåner är sådana att du har rätt till dem endast om du flyttar ditt stadigvarande boende till Finland.
En studerande från ett land utanför EU/EES kan ha rätt till vissa av FPA:s förmåner, till exempel de förmåner som ingår i sjukförsäkringen.
Läs mer på InfoFinlands sida Den sociala tryggheten i Finland.
Social trygghet för dig som flyttar till Finlandfinska _ svenska _ engelska
Utländsk examen i Finland
Om du har avlagt en examen utomlands kan du ha nytta av jämställande av examen, erkännande av yrkeskompetens eller av att skaffa dig rätt till yrkesutövning eller en fristående examen.
På InfoFinlands sida Utländska examina i Finland hittar du information om hur du kan få din examen eller dina studier erkända i Finland.
linkkiUtbildningsstyrelsen:
Erkännande av en examenfinska _ svenska _ engelska
Kommunerna tillhandahåller många tjänster för sina invånare.
Till kommunens tjänster hör till exempel hälsovård och barndagvård.
Om du har en hemkommun (kotikunta) i Finland, har du vanligen rätt att använda dig av den kommunens tjänster.
Det lönar sig för dig att utreda om du och de andra medlemmarna i din familj har rätt till en hemkommun i Finland.
Rätten till en hemkommun i Finland bestäms enligt hemkommunslagen.
Vid magistraten (maistraatti) på din egen boningsort kan du ta reda på om du har rätt till en hemkommun i Finland.
Hur kan du få en hemkommun i Finland
För att du ska kunna få en hemkommun i Finland måste du flytta till och vara stadigvarande bosatt i Finland.
Om du bor i Finland tillfälligt, till exempel om du flyttar till Finland för studier eller jobb under högst ett år, kan du vanligen inte få en hemkommun i Finland.
Du har möjlighet att få en hemkommun i Finland om:
du är finsk medborgare
du är medborgare i ett nordiskt land
du är medborgare i EU, Schweiz eller Liechtenstein och du har registrerat din uppehållsrätt i Finland
du har permanent (P) eller kontinuerligt (A) uppehållstillstånd som är i kraft
du är familjemedlem till en person som har en hemkommun i Finland
Om du har ett tillfälligt uppehållstillstånd (B-tillstånd) som är i kraft kan du få en hemkommun om du kan påvisa att det är din avsikt att bo stadigvarande i Finland.
Stadigvarande boende kan påvisas till exempel genom följande omständigheter:
du har en arbetsplats i Finland och ditt arbetskontrakt är i kraft minst två år
du studerar i Finland och dina studier räcker minst två år
du är av finländsk härkomst
du har tidigare haft en hemkommun i Finland
du har varit fortlöpande bosatt i Finland under minst ett års tid.
Din hemkommun är vanligen den kommun du bor i.
Om du inte har en bostad eller om du har bostäder på flera kommuners område är din hemkommun den kommun som du själv uppfattar som din hemkommun och som du har någon fast förbindelse till, till exempel genom familjeförhållanden eller arbetsplats.
Kontaktuppgifter till magistratfinska _ svenska _ engelska
Lag om hemkommunfinska _ svenska
Utlänningar som bor i Finland har nästan samma rättigheter och skyldigheter som finländarna.
Följande rättigheter och skyldigheter gäller även utlänningar som bor i Finland.
Rättigheter
Alla har rätt till likabehandling.
Ingen får särbehandlas till exempel på grund av kön, ålder, religion eller handikapp.
Var och en får fritt yttra sina åsikter i tal och skrift.
Människor får ordna möten och demonstrationer och delta i dem.
Demonstrationer ska anmälas till polisen på förhand.
Ingen får dömas till döden eller torteras.
Alla får själva välja sin bostadsort och röra sig fritt i Finland.
Alla har rätt till integritetsskydd.
Ett brev som tillhör en annan person får inte läsas och en annan persons telefonsamtal får inte avlyssnas.
Var och en får själv välja sin egen religion.
Om man inte vill behöver man inte välja någon religion alls.
Utlänningar som bor stadigvarande i Finland och som har fyllt 18 år har rätt att rösta i kommunalval.
Utlänningar som har rösträtt i kommunalval har även rätt att ställa upp som kandidat i kommunalval.
EU-medborgare som har hemort i Finland kan rösta i Europaparlamentsvalet om de har anmält sig till rösträttsregistret (äänioikeusrekisteri).
EU-medborgare som är i det finska rösträttsregistret kan också ställa upp som kandidat i Finlands Europaparlamentsval.
Läs mer om utlänningars rösträtt i Finland på InfoFinlands sida Val i Finland.
Skyldigheter
Alla som bor eller vistas i Finland måste följa Finlands lagar.
7–17-åringar har läroplikt (oppivelvollisuus), d.v.s. skyldighet att avlägga grundskolans (peruskoulu) lärokurs.
Ofta måste de som arbetar i Finland betalar skatt på sin lön i Finland.
Alla har skyldighet att vittna inför domstol om de blir kallade.
Föräldrar är skyldiga att ta hand om sina barn.
Alla har skyldighet att hjälpa vid en olycka.
Läs mer om beskattningen på InfoFinlands sida Beskattning.
Finska medborgares rättigheter och skyldigheter
Finska medborgare har utöver de ovannämnda också några ytterligare rättigheter och skyldigheter som utlänningar bosatta i Finland inte har.
Läs mer om finska medborgarnas rättigheter och skyldigheter på InfoFinlands sida Finskt medborgarskap.
Finlands grundlagfinska _ svenska _ engelska
Information om demokratin i Finlandfinska _ svenska _ engelska
Val i Finlandfinska _ svenska _ engelska
Uppehållstillstånd
Fortsatt uppehållstillstånd
Arbete och företagande i Finland
Finska och svenska språket
Studier
Den sociala tryggheten
Hälsan
Uppehållstillstånd
Om du är medborgare i något av de nordiska länderna, ett EU-land, ett EES-land eller i Schweiz och kommer till Finland för att arbeta, behöver du inget uppehållstillstånd.
Läs mer på InfoFinlands sida Nordisk medborgare eller EU-medborgare.
Om du är medborgare i något annat land behöver du ett uppehållstillstånd för arbetstagare.
Om du redan befinner dig i Finland på någon annan grund kan du ha rätt att arbeta även om du inte har ansökt om ett uppehållstillstånd på grund av arbete.
Läs mer på InfoFinlands sida Till Finland för att arbeta.
Om du inte är medborgare i något av Europeiska unionens medlemsländer, ett EES-land eller i Schweiz och vill driva ett företag i Finland, behöver du ett uppehållstillstånd för företagare.
Mer information om uppehållstillstånd för företagare hittar du på InfoFinlands sida Bli företagare i Finland.
Arbete i Finlandfinska _ svenska _ engelska
Uppehållstillstånd för företagarefinska _ svenska _ engelska
Fortsatt uppehållstillstånd
Ansök om fortsatt uppehållstillstånd på internet i tjänsten Enter Finland eller på Migrationsverkets tjänsteställe.
Gör en ansökan innan ditt föregående uppehållstillstånd går ut.
Du får mer information om att ansöka om fortsatt uppehållstillstånd på InfoFinlands sida Fortsatt uppehållstillstånd.
Att förlänga uppehållstillståndetfinska _ svenska _ engelska
Arbete och företagande i Finland
I InfoFinlands avsnitt Arbete och företagande hittar du mycket information om arbetslivet och företagandet i Finland.
Finska och svenska språket
En del arbetsgivare ordnar undervisning i det finska språket för sina anställda.
Fråga din arbetsgivare som det ordnas undervisning i det finska språket på din arbetsplats.
Information om andra möjligheter att studera finska eller svenska hittar du i InfoFinlands avsnitt Finska och svenska språket.
Studier
Om du vill avlägga examen eller fortbilda dig kan du delta i fortbildning.
Fortbildning ordnas bland annat av läroanstalter, fackförbund och Institutet för Yrkenas befrämjande.
Också många arbetsplatser utbildar sina anställda till exempel i användningen av nya apparater eller program.
Studierna är inte alltid inriktade på att skaffa ett yrke.
Du kan också ha studier som hobby.
Läs mer på InfoFinlands sida Studier som hobby.
Grundläggande information om fortbildningfinska _ svenska
Den sociala tryggheten
Du kan omfattas av den finländska sociala tryggheten endera på basis av stadigvarande bosättning eller på basis av arbete.
De flesta av FPA:s förmåner är sådana att du har rätt till dem endast om du flyttar ditt stadigvarande boende till Finland.
Dessutom måste du uppfylla samma villkor för att få förmånen som alla andra som bor i Finland.
Om du flyttar till Finland för att arbeta, har du vanligtvis rätt till FPA:s förmåner under din anställning också när din anställning endast är kortvarig.
Om din lön uppgår till minst 696,60 € i månaden, har du rätt till de flesta av FPA:s förmåner.
Hur många timmar per vecka du arbetar eller hur lång din anställning är spelar ingen roll.
Om du har anställning i Finland, är det skäl för dig att ansluta dig till en finländsk arbetslöshetskassa.
Om du är medlem av en arbetslöshetskassa kan du få inkomstrelaterad arbetslöshetsersättning, om du blir arbetslös.
Läs mer på InfoFinlands sidor Fackförbund och Arbetslöshetsförsäkring.
Social trygghet för dig som flyttar till Finlandfinska _ svenska _ engelska
Hälsan
Hälsovård för anställda och företagare
Om du har kommit till Finland för att arbeta har du vanligen rätt att använda de offentliga hälsovårdstjänsterna i Finland.
Detta beror på hurdant och hur långt arbetsavtal du har samt från vilket land du har kommit till Finland.
Du kan begära att FPA utreder din rätt till de offentliga hälsovårdstjänsterna.
Du hittar mer information om den offentliga hälso- och sjukvården på InfoFinlands sida Hälsovårdstjänster i Finland.
I Finland är arbetsgivare skyldiga att ordna förebyggande företagshälsovård för sina anställda.
Företagare kan ordna sin egen företagshälsovård om de vill.
Företagare måste alltså inte ordna företagshälsovård för sig.
Företagare måste ändå ordna företagshälsovård för sina anställda.
Företagshälsovården kan ordnas vid den lokala hälsovårdscentralen eller till exempel på en privat läkarcentral.
Mer information får du på InfoFinlands sida Företagshälsovården och på social- och hälsovårdsministeriets webbplats.
linkkiSocial- och hälsovårdsministeriet:
Företagshälsovårdfinska _ svenska _ engelska
Om du förlorar ditt jobb
Om du har ett uppehållstillstånd för arbetstagare som endast gäller arbete för en viss arbetsgivare och du förlorar din arbetsplats, ska du ansöka om ett nytt uppehållstillstånd för arbetstagare eller ett uppehållstillstånd på andra grunder.
Om Migrationsverket har beviljat dig ett uppehållstillstånd för arbetstagare och din anställning upphör tidigare än uppehållstillståndet, måste du eller din arbetsgivare skriftligt meddela Migrationsverket att din anställning upphör.
Om ditt uppehållstillstånd för arbetstagare inte har begränsats att gälla arbete för en viss arbetsgivare, utan för en viss bransch och tillståndet är fortfarande giltigt, kan du byta jobb inom samma bransch.
Problem i arbetslivet
Om du råkar ut för problematiska situationer på arbetsplatsen ska du först kontakta din chef.
Om ärendet inte kan lösas på arbetsplatsen, ska du kontakta arbetarskyddsdistriktet (työsuojelupiiri) i ditt område eller ditt fackförbund.
Information och råd om var du kan få hjälp med olika slags problem i arbetslivet hittar du på InfoFinlands sida Problem i arbetslivet.
När du har flyttat till Finland ska du besöka magistraten på din hemort för att registrera dig som invånare.
Innan du besöker magistraten kan du fylla i Registreringsanmälan för utlänningar som finns på adressen maistraatti.fi.
Du kan även fylla i anmälan på magistraten.
Magistraten registrerar dina uppgifter i det finska befolkningsdatasystemet.
Dessa uppgifter är bland annat namn, födelsedatum, medborgarskap, kön och adress.
Om du flyttar till Finland för att bo här stadigvarande i ett år eller längre kan du ha rätt till hemkommun i Finland.
Du behöver en hemkommun för att kunna använda kommunala tjänster, såsom hälso- och sjukvården eller dagvården.
Magistraten utreder om du kan få en hemkommun registrerad.
När du besöker magistraten, ta med dig minst följande handlingar:
Om du är EU-medborgare eller nordisk medborgare:
Giltigt pass eller annan identitetshandling som styrker ditt medborgarskap
Arbetsavtal, intyg om studier eller någon annan utredning över registreringsbehovet (om du är EU-medborgare och ännu inte har registrerat din uppehållsrätt vid Migrationsverket)
Äktenskapsintyget i original (om du är gift)
Dina barns födelseattester i original (om du har barn under 18 år som flyttar till Finland)
Observera att du måste legalisera handlingar som har utfärdats av myndigheter utanför EU eller Norden.
Det gäller till exempel äktenskapsintyg som utfärdats i USA.
Om du är medborgare i något annat land:
Giltigt pass
Uppehållstillstånd (om du behöver uppehållstillstånd i Finland)
Vid behov utredning över arbete eller studier i Finland (t.ex. arbetsavtal eller närvarointyg som utfärdats av din läroanstalt) eller någon annan utredning över orsakerna till registreringen
Legaliserat äktenskapsintyg i original (om du är gift)
Legaliserade födelseattester för dina barn i original (om du har barn under 18 år som flyttar till Finland)
Legalisering av handlingar
På magistraten ska du visa upp originalhandlingen eller en vidimerad kopia av den.
Kopian kan pålitligt vidimeras av den myndighet som utfärdat handlingen eller notarius publicus i det land där handlingen utfärdades.
Handlingen ska vara legaliserad för att magistraten ska kunna föra in dina uppgifter i befolkningsdatasystemet.
Om ditt land har tillträtt Haagkonventionen ska du begära om ett så kallat Apostille-intyg för din handling.
Du behöver inget Apostille-intyg om du har en allmän handling som utfärdats av en myndighet i ett EU-land.
Du kan emellertid behöva en standardblankett som används som översättningsstöd som bilaga till en allmän handling.
Du får mer information om dessa standardblanketter hos myndigheterna i det land där du begär intyget.
Ett annat alternativ är att handlingen översätts av en auktoriserad översättare som godkänts av ett EU-land.
Observera att handlingarna ska vara på finska, svenska eller engelska.
Om din handling är på något annat språk måste du se till att få den översatt till finska, svenska eller engelska.
En auktoriserad översättare kan översätta handlingen åt dig.
Om översättningen görs utomlands måste även översättningen vara legaliserad.
Om du behöver mer information om legalisering av handlingar, kontakta magistraten eller utrikesministeriet i ditt eget land.
Finsk personbeteckning
Du får en personbeteckning av Migrationsverket när du beviljas uppehållstillstånd i Finland eller när din uppehållsrätt för EU-medborgare registreras.
Du kan även få en finsk personbeteckning vid:
skattebyrån, om du behöver personbeteckningen för beskattningen.
Den finska personbeteckningen är en nummerserie med elva siffror som bildas baserat på ditt födelsedatum och ditt kön.
Du behöver personbeteckningen till exempel för din arbetsgivare eller läroanstalt.
Den underlättar även skötseln av många officiella ärenden.
Om du har fått din personbeteckning någon annanstans än vid magistraten och vill ha en hemkommun, måste du även besöka magistraten.
Läs mer på InfoFinlands sida Hemkommun i Finland.
Registrering av utlänningarfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Registrering av utlänningar på skattebyrånfinska _ svenska _ engelska
Om du måste sköta ärenden med finländska myndigheter, men inte kan finska eller svenska och det inte heller finns något annat språk som både du och myndigheten talar, kan du i vissa fall ha rätt till tolkning.
Då beställer myndigheten tolken och betalar för tolkningen.
Myndigheten kan ordna och betala tolkningen när det gäller skötsel av ärenden som behandlas på myndighetens initiativ.
Detta är dock inte alltid möjligt.
Om du behöver en tolk för den inledande kartläggningen och integrationsplanen, måste myndigheten beställa en tolk.
Du kan på förhand fråga myndigheten om detta.
Om du söker asyl i Finland har du rätt till tolkning i ärenden som rör behandlingen av din asylansökan.
Du har rätt att få information om ett beslut gällande dig på ditt modersmål eller ett annat språk som du förstår.
Information om beslutet ges genom tolkning eller översättning.
Om du själv bokar tolken och betalar tolkningen, kan du anlita en tolk när som helst.
Tolktjänsterfinska _ svenska _ engelska
Vad gör tolken?
Tolken är med på möten mellan dig och myndigheten.
Han eller hon tolkar det som du och myndigheten säger.
Tolken är antingen på plats eller också kan tolkningen ordnas via telefon eller video.
Tolken har som uppgift att tolka det som du och myndigheten säger.
Tolken sköter inga andra uppgifter utöver tolkningen.
Han eller hon kan således inte hjälpa dig med annat.
Tolken är en neutral, utomstående person som varken är på din eller på myndighetens sida.
Tolken har sekretessplikt och får inte berätta inte om dina angelägenheter för andra.
Var kan man beställa en tolk?
I Finland finns åtta kommunala tolkcentraler (tulkkikeskus).
Tolkcentralernas tjänster är främst avsedda för myndigheter som arbetar med invandrare.
Också många företag erbjuder tolktjänster.
linkkiFinlands översättar- och tolkförbund:
Sök tolk eller översättarefinska _ svenska _ engelska
Kommunala tolkcentraler
linkkiHelsingforsnejdens kontakttolkcentral:
Tolkningfinska
linkkiMellersta Finlands tolkcentral:
Tolkningfinska _ svenska _ engelska
Tolkningfinska
Tolkningfinska _ engelska
linkkiÖsterbottens tolkcentral:
Tolkningfinska
linkkiNorra Finlands tolktjänst:
Tolkningfinska
linkkiÅboregionens tolkcentral:
Tolkningfinska _ svenska
Tolkningfinska
Arbetstagare, företagare, studerande, flykting, asylsökande eller en familjemedlem till en person bosatt i Finland hittar information speciellt om sin egen situation på dessa sidor i Infobanken.
Via dessa sidor hittar du snabbt den information som du behöver i kortfattade form.
Arbetstagare eller företagare
Studerande
Flykting
Asylsökande
Familjemedlem
Om du är medborgare i något nordiskt land behöver du inte uppehållstillstånd i Finland.
Du har rätt att jobba, fungera som företagare och studera i Finland.
När du flyttar till Finland måste du göra en flyttanmälan och gå och registrera dig vid magistraten (maistraatti) på din egen hemort.
Notera att du måste besöka magistraten personligen.
Gör flyttanmälan senast inom en vecka från din flyttningsdag.
För registreringen behöver du ett officiellt identitetskort där ditt medborgarskap framgår eller pass som är i kraft.
Familjemedlemmar till nordiska medborgare
Om en av dina familjemedlemmar, som flyttar med dig till Finland, inte är medborgare i ett nordiskt land, kan han/hon behöva uppehållstillstånd eller ett registreringsintyg över uppehållsrätt för EU-medborgare.
Läs mer på InfoFinlands sidor EU-medborgare eller Icke-EU-medborgare.
Finsk personbeteckning
När du registrerar dig vid magistraten kan du på samma gång få en finsk personbeteckning (henkilötunnus).
Du behöver en personbeteckning när du sköter ärenden hos myndigheter, och dessutom underlättar den skötandet av ärenden i till exempel banker och med din arbetsgivare.
Läs mer på InfoFinlands sidor Registrering som invånare.
Registrering av utlänningarfinska _ svenska _ engelska
Information för nordiska medborgarefinska _ svenska _ engelska _ norska
_ danska
_ isländska
Rådgivningstjänst för nordiska medborgarefinska _ engelska _ norska
_ danska
_ isländska
Bankkonto
Du behöver ett bankkonto för att sköta din dagliga ekonomi.
Det lönar sig att jämföra tjänsterna och priserna som olika banker tillhandahåller så att du hittar det alternativ som är förmånligast för dig.
När du öppnar ett bankkonto behöver du ett pass, ett identitetskort för utlänningar eller någon annan officiell identitetshandling.
Om du saknar pass eller ett identitetskort för utlänningar kan du ta reda på vilken typ av identitetshandling banken kan godta.
Vissa banker godtar främlingspass, som de finska myndigheterna har utfärdat, resedokument för flykting eller någon annan identitetshandling som kan godtas som resedokument.
I vissa fall kan banken även kräva andra utredningar av identiteten, om du har en notering i din handling som anger att din identitet inte har kunnat fastställas.
Du kan inte identifiera dig med ett körkort.
När du öppnar ett bankkonto har banken en lagstadgad skyldighet att fråga vad ditt konto ska användas till.
Banken har även rätt att kontrollera om du har betalningsanmärkningar.
Banken behöver följande uppgifter från dig:
personnummer
adress i Finland eller i ett annat land
om du betalar skatt i ett annat land än Finland, din adress i det landet
samma uppgifter för de personer som har rätt att använda kontot.
När du öppnar ett bankkonto lönar det sig att även skaffa webbankkoder.
Med hjälp av webbankkoderna kan du till exempel uträtta många myndighetsärenden på nätet.
För dessa koder gäller dock hårdare krav än för öppning av ett bankkonto.
I vissa fall kan du alltså inte få webbankkoder även om du har ett bankkonto.
Vill du ha råd i bankfrågor kan du ringa till Försäkrings- och finansrådgivningen (Fine).
Tjänsten är kostnadsfri för kunderna, dvs. du betalar endast din egen samtalskostnad.
Tjänsten tillhandahålls på finska, svenska och engelska.
Försäkrings- och finansrådgivningen
tfn. 09 6850 120
linkkiFinansbranschens Centralförbund:
Utländska medborgares bankärendenfinska _ engelska
Identitetskort för utlänningar
Polisen kan utfärda dig ett identitetskort för utlänningar om du har identifierats och din identitet har verifierats på ett tillförlitligt sätt.
Din identitet kan verifieras från en handling som styrker identiteten.
Om du inte har en sådan handling, kan dina fingeravtryck jämföras med de fingeravtryck som lagrats i uppehållstillståndskortet eller uppehållskortet.
Dessutom krävs att:
du har ett giltigt uppehållstillstånd eller uppehållskort eller att din uppehållsrätt är registrerad,
du har hemkommun i Finland och
uppgifter om dig har registrerats i befolkningsdatasystemet.
Med ett identitetskort för utlänningar kan du styrka din identitet i Finland.
Du kan använda det till exempel när du ska öppna ett bankkonto i Finland.
Du kan emellertid inte använda det som resedokument på utlandsresor.
ID-kortfinska _ svenska _ engelska
Försäkringar
När du har en bostad är det bra att ta en hemförsäkring.
Hemförsäkringen ersätter till exempel skador på möbler och andra ägodelar.
Hemförsäkringar säljs av försäkringsbolag.
Om du använder en egen bil ska du enligt lagen ha en trafikförsäkring.
Om du vill ta en personförsäkring i ett finländskt försäkringsbolag ska du vanligtvis ha ett finländskt FPA-kort.
Personförsäkringar kan vara till exempel olycksfallsförsäkring, vårdkostnadsförsäkring och livförsäkring.
Försäkringsbolag i Finlandfinska
Telefon
När du tecknar ett telefonabonnemang i Finland får du ett finskt telefonnummer.
Många företag erbjuder telefonabonnemang.
För att teckna ett abonnemang behöver du ett finländskt identitetsnummer och du måste ha en adress i Finland.
Du ska vanligtvis även kunna visa ditt betalningsbeteende, dvs. uppgifter som visar att du har betalat dina räkningar och inte har några betalningsanmärkningar.
I annat fall måste du betala abonnemanget i förskott.
Du kan också köpa ett prepaid-abonnemang.
Då behöver du inte ha en finländsk identitetshandling eller adress i Finland.
Prepaid-kortet är i förväg laddat med en summa som man sedan kan ringa för.
Prepaid-abonnemang kan köpas till exempel i R-kiosker, en del snabbköp och på Internet.
När du ringer till utlandet med telefon lönar det sig att kontrollera vilket utlandsprefix du ringer förmånligast med.
Många företag erbjuder förmånliga utlandsprefix.
Observera att samtalspriset ändå alltid beror på vilket land du ringer till.
Kontrollera vilket alternativ som är förmånligast för dig.
Telefonoperatörer i Finlandfinska
linkkiTeleAle:
Förmånliga utlandssamtalfinska _ svenska _ engelska
Förmånliga utlandssamtalfinska _ engelska
linkkiSkype:
Förmånliga utlandssamtalfinska _ svenska _ engelska _ ryska _ estniska _ franska _ spanska _ turkiska _ kinesiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ ungerska _ japanska
Internet
I Finland kan du sköta många ärenden via Internet.
Man kan ofta uträtta ärenden hos myndigheter eller företag via deras webbsidor.
Det är bra att skaffa sig en Internetanslutning så fort som möjligt efter att du har flyttat till Finland.
Du får en Internetanslutning hem till dig genom att teckna ett avtal med en Internettjänsteleverantör.
Det lönar sig att jämföra olika tjänsteleverantörers priser innan man ingår ett avtal.
I Finland finns många företag som erbjuder olika typer av Internetanslutningar.
Dessa företag hittar till exempel genom sökning på nätet när du skriver ”internetliittymä” i sökmaskinens sökfält.
Anslutningarnas priser varierar mycket.
Om du har ett bibliotekskort kan du också använda internet gratis på biblioteken.
Ett bibliotekskort får du gratis på biblioteket.
Läs mer på InfoFinlands sida Bibliotek.
Det finns också caféer där kunderna har möjlighet att använda Internet.
linkkiKommunikationsverket:
Internet- och telefonabonnemangfinska _ svenska _ engelska
Prisnivån i Finland
Prisnivån är hög i Finland.
Till exempel mat och många typer av tjänster kostar i genomsnitt mer i Finland än i övriga Europa.
Boendekostnaderna varierar mycket.
I storstäderna kostar boendet mycket mer än på mindre orter.
Konsumentpriser i de Europeiska ländernafinska _ svenska
Priser på icke subventionerade hyresbostäderengelska
Priser på hyresbostäder med statliga stödengelska
Information om priser på sålda bostäderfinska _ svenska
Köp och konsumentens rättigheter
Alla som köper varor och tjänster är konsumenter.
Konsumentskyddslagen tryggar konsumentens rättigheter i Finland.
Du har rätt till gottgörelse till exempel då varan som du köpt har fel som inte du har orsakat.
Du kan till exempel ersättas med en felfri vara eller få dina pengar tillbaka.
Om en vara som du köpt har brister ska du först kontakt säljaren.
Om du inte kan komma överens om saken med säljaren, ta då kontakt med konsumentrådgivningen.
linkkiKonkurrens- och konsumentverket:
Konsumentrådgivningfinska _ svenska _ engelska
Information om konsumenträttigheterfinska _ svenska _ engelska
linkkiKonsumentförbundet:
Information om konsumenträttigheterfinska
Kollektivtrafik
Kollektivtrafiken fungerar väl i Finland.
Man kan resa nästan över allt i Finland med tåg eller buss.
Man kan också flyga till många städer.
I stora städer och deras näromgivning finns en välfungerande lokaltrafik.
Lokaltrafiken trafikeras vanligtvis med bussar.
Läs mer på InfoFinlands sida Trafiken i Finland.
Körkort
Du kan ta körkort i Finland när du har fyllt 18 år.
Om du har ett körkort som beviljats i ett annat land, beror det på situationen hur du ska gå tillväga.
Läs mer på InfoFinlands sida Trafiken i Finland.
Klimat och kläder
Klimatet i Finland är kallare än i många andra länder.
I Finland ligger medeltemperaturen på vintern under noll Celsiusgrader och på sommaren över +10 Celsiusgrader.
På våren och hösten ligger temperaturerna här emellan.
På vintern ska man klä sig varmt i Finland.
Läs mer om klimatet i Finland på InfoFinlands sida Klimatet i Finland.
Medier
I Finland utkommer nästan 200 tidningar.
Läs mer på InfoFinlands sida Medier i Finland.
Kulturen i Finland
Du hittar information om den finländska kulturen på InfoFinlands sidor Finländska seder och Den finländska arbetskulturen.
Före flytten till Finland
Efter flytten till Finland
Bekanta dig med innehållen i InfoFinland före flytten.
I InfoFinland hittar du pålitlig information på ditt eget språk om flytten till Finland, arbetslivet, boende, studier i finska eller svenska språket, utbildning, social trygghet, hälsotjänster, tjänster för familjer, problematiska situationer och fritid.
På sidorna finns nyttiga praktiska råd, kontaktuppgifter och länkar till tilläggsinformation.
Med hjälp av menyn Städer får du fram information om den kommun som du är intresserad av.
De olika språkversionerna av InfoFinlands är identiska.
Komihåglistan för dig som flyttar till Finland är avsedd att hjälpa dig med de viktigaste praktiska frågorna som har med flytten att göra.
Observera att listan inte nödvändigtvis innehåller allt som måste göras när du flyttar till Finland.
Före flytten till Finland
Uppehållstillstånd eller registrering av uppehållsrätt?
Om du ska vistas i Finland mer än 90 dagar och är EU-medborgare, måste du registrera din uppehållsrätt.
Om du är medborgare i ett land utanför EU, måste du ansöka om uppehållstillstånd i Finland.
Läs mer på InfoFinlands sida EU-medborgare eller Icke-EU-medborgare.
När du ansöker om uppehållstillstånd eller registrering av uppehållsrätten måste du bevisa att din utkomst i Finland är tryggad.
Om du kommer till Finland för att arbeta eller som företagare måste du bevisa att ditt arbete eller din företagsverksamhet inbringar dig en tillräcklig utkomst.
Om du flyttar till en familjemedlem i Finland, krävs det ofta även att den person som bor i Finland har tillräckliga medel för att försörja sig själv och den familjemedlem som flyttar till Finland.
Flyttsaker från EU-området
Om du flyttar till Finland från ett annat EU-land behöver du vanligen inte betala tull eller mervärdesskatt på dina flyttsaker, d.v.s. de personliga föremål som du tar med dig.
Du behöver inte heller anmäla dina flyttsaker i tullen (tulli).
Observera att tull- och skattefriheten för flyttsaker inte gäller alkohol eller tobaksprodukter.
För import av dessa gäller separata begränsningar.
Mer information får du på Tullrådgivningen +358 (0)295 5201 eller på tullens webbplats.
Tullrådgivningen betjänar på finska, svenska och engelska.
Flyttsaker från länder utanför EU
Om du flyttar till Finland från ett land som inte hör till EU behöver du vanligen inte betala tull eller mervärdesskatt på dina flyttsaker, d.v.s. de personliga föremål som du tar med dig.
Du måste dock göra en tullanmälan på flyttsakerna till de finländska tullmyndigheterna.
Som flyttsaker betraktas till exempel:
möbler och andra husgeråd
husdjur
cyklar och motorcyklar
bilar och släpvagnar avsedda för privat bruk.
Observera att tull- och skattefriheten för flyttsaker inte gäller alkohol eller tobaksprodukter.
För import av dessa gäller separata begränsningar.
linkkiTullen:
Införsel av flyttsaker till Finlandfinska _ svenska _ engelska _ ryska
Införsel av bil till Finland som flyttsak
När du tar med dig en bil till Finland som flyttsak, måste du tullanmäla den.
Om du tar med dig en bil till Finland måste du registrera den och betala bilskatt (autovero) för den innan du kan använda den i trafiken.
Man kan dock använda bilen tillfälligt innan bilskatten är betald.
Detta förutsätter att du har gjort en anmälan om ibruktagande av fordonet (auton käyttöönottoilmoitus) till skatteförvaltningen.
Du ska också ha en giltig trafikförsäkring (liikennevakuutus) för din bil i Finland.
Om du för in en bil från ett land utanför EES-området behöver du också ett förflyttningstillstånd innan du kan använda bilen.
Förflyttningstillstånd beviljas av besiktningskontor och vissa av Tullens verksamhetsställen.
Du får inte använda din bil i Finland förrän du har gjort en anmälan om ibruktagande av fordonet och skaffat ett förflyttningstillstånd.
Om du har frågor kring fordonsskatten eller anmälan om ibruktagande, kan du ringa skatteförvaltningens telefontjänst:
+358 (0)29 497 150 (finska)
+358 (0)29 497 151 (svenska)
+358 (0)29 497 152 (engelska)
linkkiTullen:
Fordon som flyttgodsfinska _ svenska _ engelska _ ryska
Införsel av sällskapsdjur
Mer information om reglerna i Finland ges av Livsmedelsverket (Ruokavirasto).
linkkiLivsmedelsverket:
Införsel av djur från EU-länderfinska _ svenska _ engelska
linkkiLivsmedelsverket:
Införsel av djur från länder utanför EUfinska _ svenska _ engelska
Flyttfirmor
En del företag som tillhandahåller flyttservice sköter också flytt från ett land till ett annat.
Du kan anlita dessa företag att transportera dina ägodelar från ett land till ett annat och också att packa dina saker och tillhandahålla förpackningsmaterial.
Flyttkostnaderna beror på varifrån du flyttar och hur mycket saker du har.
Tjänsterna och priserna i olika flyttfirmor kan variera stort och därför lönar det sig att jämföra.
Flyttjänsterfinska _ svenska _ engelska
linkkiViktor Ek:
Flyttjänsterfinska _ svenska _ engelska
Hjälp när du flyttarfinska _ svenska _ engelska _ norska
_ danska
Efter flytten till Finland
I den här listan har vi samlat de vanligaste ärendena som du måste ta hand om när du har kommit till Finland.
Bostad och hemförsäkring
De flesta invandrare bor först i en hyresbostad när de kommer till Finland.
Det är bra att reservera minst en månad för att söka hyresbostad.
Läs mer på InfoFinlands sida Boende.
När du har en bostad är det bra att också ta en hemförsäkring (kotivakuutus).
Hemförsäkringen ersätter till exempel skador på möbler och andra ägodelar.
Hemförsäkringar säljs av försäkringsbolag.Information om försäkringar finns på InfoFinlands sida Vardagslivet i Finland.
Finsk personbeteckning
Om du får ett uppehållstillstånd i Finland registreras du automatiskt i det finska befolkningsdatasystemet.
Du får samtidigt även en finsk personbeteckning.
I Finland kan du få personbeteckningen även vid magistraten eller skattebyrån på din hemort.
Läs mer på InfoFinlands sida Registrering som invånare.
Hemkommun i Finland
Om du flyttar till och blir stadigvarande bosatt i Finland registreras en hemkommun för dig i Finland.
Hemkommunen är den kommun där du bor.
När du har en hemkommun har du rätt att använda denna kommuns tjänster såsom till exempel offentliga hälsovårdstjänster.
Du kan ta reda på om det är möjligt att registrera en hemkommun i Finland för dig vid magistraten på din hemort.
Läs mer på InfoFinlands sida Hemkommun i Finland.
Registrering av utlänningarfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Registrering av utlänningar på skattebyrånfinska _ svenska _ engelska
Social trygghet
Du kan omfattas av den finländska sociala tryggheten endera på basis av stadigvarande bosättning eller på basis av arbete.
De flesta av FPA:s förmåner är sådana att du har rätt till dem endast om du flyttar ditt stadigvarande boende till Finland.
Dessutom måste du uppfylla samma villkor för att få förmånen som alla andra som bor i Finland.
Social trygghet för dig som flyttar till Finlandfinska _ svenska _ engelska
Bankkonto
Du behöver ett bankkonto för att sköta din dagliga ekonomi.
När du öppnar ett bankkonto behöver du ett pass eller någon annan officiell identitetshandling.
Det lönar sig att jämföra tjänsterna och priserna som olika banker tillhandahåller så att du hittar det alternativ som är förmånligast för dig.
Information om att öppna ett bankonto finns på InfoFinlands sida Vardagslivet i Finland.
linkkiFinansbranschens Centralförbund:
Utländska medborgares bankärendenfinska _ engelska
Skattekort
Om du arbetar och får lön eller är företagare behöver du ett finskt skattekort (verokortti).
Skattekortet får du vid skattebyrån.
Läs mer om beskattningen i Finland på InfoFinlands sida Beskattning.
Kollektivtrafik
Om du bor i en stad är det inte nödvändigt att äga en bil.
Kollektivtrafiken fungerar väl i Finland.
Man kan resa nästan över allt i Finland med tåg eller buss.
Man kan också flyga till många städer.
I stora städer och deras näromgivning finns en välfungerande lokaltrafik.
Lokaltrafiken trafikeras vanligtvis med bussar.
Läs mer på InfoFinlands sida Trafiken i Finland.
Körkort
Om du har ett körkort som utfärdats i ett av de nordiska länderna eller i ett EU-/EES-land, är det giltigt även i Finland.
Om du bor stadigvarande i Finland kan du byta ut kortet mot ett finländskt körkort.
Om du har ett körkort som utfärdats i ett land som är anslutet till Genève- eller Wien-konventionerna kan du köra med detta kort högst två år i Finland.
Du måste byta ut ditt körkort mot ett finländskt körkort inom två år efter att du flyttat till Finland.
Om du har ett körkort som utfärdats i ett land som inte är anslutet till Genève- eller Wien-konventionerna kan du köra bil med detta kort under ett års tid efter att ha registrerats i befolkningsregistret i Finland.
Du kan byta ut ditt körkort till ett finskt körkort på Ajovarmas serviceställe.
linkkiTrafiksäkerhetsverket:
Utländskt körkort i Finlandfinska _ svenska _ engelska
Internet
I Finland kan du sköta många ärenden via Internet.
Det är bra att skaffa sig en Internetuppkoppling så fort som möjligt efter att du har flyttat till Finland.
På InfoFinlands sida Vardagslivet i Finland finns mer information om att skaffa en internetuppkoppling.
linkkiKommunikationsverket:
Internet- och telefonabonnemangfinska _ svenska _ engelska
Telefon
När du köper ett telefonabonnemang i Finland får du ett finskt telefonnummer.
Många företag erbjuder telefonabonnemang.
Du kan också köpa ett prepaid-abonnemang.
Prepaid-kortet är i förväg laddat med en summa som man sedan kan ringa för.
Prepaid-abonnemang kan köpas till exempel i R-kiosker, en del snabbköp och på Internet.
linkkiSkype:
Förmånliga utlandssamtalfinska _ svenska _ engelska _ ryska _ estniska _ franska _ spanska _ turkiska _ kinesiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ ungerska _ japanska
Hälsa
I Finland finns offentliga och privata hälsovårdstjänster.
Du kan använda de offentliga hälsovårdstjänsterna om du har en hemkommun i Finland.
Till de offentliga hälsovårdstjänsterna hör till exempel hälsocentralerna.
De offentliga tjänsterna är förmånligare än de privata.
Om du vill reservera tid till en läkare ska du ta kontakt med hälsocentralen.
Om du inte har rätt att använda de offentliga hälsovårdstjänsterna kan du kontakta en privat läkarcentral.
Mer information om hälsovården i Finland får du på InfoFinlands sida Hälsa.
Språkstudier
Finlands officiella språk är finska och svenska.
Språkkunskaper hjälper dig att förstå det nya samhället och underlättar skötseln av ärenden.
Mer information hittar du på InfoFinlands sida Finska och svenska språket.
Jobbsökning
Arbets- och näringsbyrån hjälper dig i jobbsökningen.
Du kan söka jobb på Internet och via tidningar.
Du kan också hitta ett jobb genom att själv kontakta arbetsgivare som du är intresserad av.
Läs mer om jobbsökning i Finland på InfoFinlands sida Var hittar jag jobb?
Fritid och hobbyer
Information om möjligheter till fritidsaktiviteter hittar du på InfoFinlands sida Fritid.
linkkiExpat Finland:
Information om Finland för utlänningarengelska
Om du behöver visum eller uppehållstillstånd för att vistas i Finland, men inte har det, vistas du illegalt i Finland.
Asylsökande har rätt att uppehålla dig i Finland även utan visum eller uppehållstillstånd under den tid som det tar att handlägga asylansökan.
Även om du har kommit lagligt till Finland kan din vistelse i landet bli illegal till exempel om du stannar kvar i landet fastän du inte beviljas ett uppehållstillstånd eller om ditt visum eller uppehållstillstånd har gått ut.
Information om hur du kan få ett uppehållstillstånd i Finland finns på InfoFinlands sida Flytta till Finland.
Hjälp och rådgivning
Mathjälp och inkvartering
Du har rätt till nödinkvartering och mathjälp om du inte har pengar till mat eller någonstans att övernatta.
Kommuner, församlingar och vissa organisationer ordnar nödinkvartering.
Juridisk rådgivning
Flyktingrådgivningen r.f. ger kostnadsfri juridisk rådgivning för papperslösa invandrare.
Rådgivningen betjänar telefonledes på numret 045-237 7104 (måndagar kl. 14–16).
Rådgivningen ges av en jurist.
Fler kontaktuppgifter hittar du på Flyktingrådgivningens webbplats.
Sjukvård
Om du blir sjuk eller skadas, har du rätt till brådskande vård inom den offentliga hälso- och sjukvården, till exempel på en hälsostation eller ett sjukhus.
Du måste i regel själv betala kostnaderna för vården.
I Helsingfors, Åbo, Tammerfors och Esbo får barn och gravida kvinnor samma hälso- och sjukvårdstjänster som övriga invånare.
De måste betala samma avgifter för vården som övriga invånare.
Global Clinic är en klinik där du kan få hjälp eller råd av en läkare eller sjukskötare om du vistas i Finland utan uppehållstillstånd.
Du kan besöka Global Clinic även om du inte behöver brådskande sjukvård.
Global Clinic bedriver verksamhet i följande städer:
Åbo
Tammerfors
Uleåborg
Joensuu
Du kan ringa eller skicka e-post.
En sjukskötare eller läkare besvarar ditt samtal.
Du hittar kontaktinformation på Global Clinic:s hemsidor.
Global Clinic:s tjänster är avgiftsfria för kunderna.
Global Clinic anmäler inte sina kunder till polisen eller andra myndigheter.
Klinikens adress eller öppettider meddelas inte offentligt.
linkkiFlyktingrådgivningen rf:
Juridisk rådgivningfinska _ engelska _ franska _ arabiska
Kontaktuppgifterfinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Med integration (kotoutuminen) avses att du bosätter dig i Finland och skaffar kunskaper och färdigheter som du behöver i det finländska samhället.
Integrationen underlättas t.ex. av att
du lär dig språket,
hittar en arbetsplats eller studieplats,
får kontakter till det finländska samhället.
I Finland finns det olika tjänster som främjar din integration, hjälper dig att hitta sysselsättning och lära dig språket.
Också dina familjemedlemmar kan ha rätt till dessa tjänster om de flyttar till Finland tillsammans med dig.
Det är viktigt att du även själv aktivt främjar din integration.
Integrationsfrämjande tjänster
Grundläggande information om Finland
Alla invandrare har rätt att få grundläggande information om Finland.
När du får uppehållstillstånd eller registrerar din uppehållsrätt, får du samtidigt skriftlig information om
det finländska samhället och arbetslivet,
dina rättigheter och skyldigheter
tjänster som främjar din integration.
Invandrarrådgivning
Arbets- och näringsbyråerna och kommunerna tillhandahåller invandrarrådgivning.
De hjälper dig att integrera dig i Finland.
integration och integrationsfrämjande tjänster
arbetslivet
utbildning och studier.
Inledande kartläggning
Vid den inledande kartläggningen görs en utvärdering av det tjänster som kan främja din integration.
Vid den inledande kartläggningen utreds t.ex. din utbildning, din arbetserfarenhet och dina språkkunskaper.
Den inledande kartläggningen görs vid arbets- och näringsbyrån eller vid kommunen.
Den kan också göras på ett annat ställe, t.ex. vid en läroinrättning.
Detta beror på vilken kommun du bor i.
Du kan framföra en begäran om en inledande kartläggning av din situation t.ex. till arbets- och näringsbyrån eller socialbyrån i din kommun.
Invandrarrådgivningen ger dig närmare information om den inledande kartläggningen och hur den ordnas i din hemkommun.
Om du behöver stöd för din integration, utarbetas en integrationsplan för dig efter den inledande kartläggningen.
En integrationsplan utarbetas för dig åtminstone om
du är arbetslös arbetssökande eller
får utkomststöd eller
du inte fyllt 18 år och inte har en vårdnadshavare i Finland.
I integrationsplanen antecknas åtgärder som främjar din integration.
Planen kan omfatta t.ex. studier i finska, andra studier eller arbetspraktik.
Du kan utarbeta en integrationsplan t.ex. med en arbetskraftsrådgivare vid arbets- och näringsbyrån, alltså TE-byrån (TE-toimisto), eller med en socialarbetare på socialbyrån.
Integrationsplanen ska utarbetas senast tre år efter att du fått ditt första uppehållstillstånd eller din uppehållsrätt registrerades.
Integrationsplanens längd beror på hur lång tid du behöver stöd för din integration.
Integrationsplanen gäller vanligen i högst tre år.
I vissa specialfall kan den gälla i fem år.
När en integrationsplan har utarbetats för dig, är det viktigt att du följer planen.
TE-byrån eller kommunen anvisar dig vid behov till integrationsutbildning.
I utbildningen ingår studier i finska eller svenska och introduktion i det finländska samhället och arbetslivet samt den finländska kulturen.
I utbildningen kan även andra studier och praktik ingå.
TE-byrån, FPA eller kommunen utreder din rätt till arbetslöshetstförmån eller utkomststöd under integrationsplanen.
Om du har en arbetsplats kan din arbetsgivare eventuellt stöda din integration.
Arbetsgivaren kan t.ex. betala avgifter för en kurs i finska för din räkning.
Ibland kan arbetsgivaren också hjälpa dig med praktiska ärenden, t.ex. leta efter en bostad åt dig.
Fråga mer om detta av din arbetsgivare.
linkkiArbets- och näringsministeriet:
Inledande kartläggning och integrationsplanfinska _ svenska _ engelska
Stöd till arbetslösa invandrarefinska _ svenska _ engelska
Integrationsutbildning
När en integrationsplan utarbetats kan du få integrationsutbildning.
Integrationsutbildning ordnas av kommuner, arbets- och näringsbyråer och många läroanstalter.
Arbets- och näringsbyrån eller kommunen hänvisar dig till integrationsutbildningen.
Integrationsutbildningen omfattar vanligen studier i finska eller svenska. I utbildningen bekantar du dig med det finländska samhället och arbetslivet och den finländska kulturen.
Studier i finska och svenska
På InfoFinlands sida Finska och svenska språket hittar du information om möjligheterna att studera finska eller svenska.
Din kultur i Finland
Din kultur, ditt språk och din religion kan fortfarande utgöra en viktig del av ditt liv också i Finland.
En invandrarförening kan hjälpa dig att bevara och utveckla din kultur.
I Finland finns många föreningar för invandrare.
Du hitar mer information om föreningar på InfoFinlands sida Föreningar.
Barn med invandrarbakgrund kan få undervisning i det egna modersmålet.
Du hitar mer information på InfoFinlands sida Grundläggande utbildning.
I Finland råder religionsfrihet (uskonnonvapaus).
Var och en har alltså rätt att bekänna och utöva sin religion.
Var och en får själv välja sin religion.
Om du vill, kan du låta att bli att välja en religion.
Du hittar mer information om religionsutövning i Finland på InfoFinlands sida Kulturer och religioner i Finland.
linkkiArbets- och näringsministeriet:
Guiden Välkommen till Finland(pdf, 3,40 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
linkkiArbets- och näringsbyrån:
Information om integrationfinska _ svenska _ engelska
linkkiArbets- och näringsbyrån:
Broschyren Jobba i Finland(pdf, 5,51 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ polska
Kommunerna tillhandahåller många tjänster för sina invånare.
Till kommunens tjänster hör till exempel hälsovård och barndagvård.
Om du har en hemkommun (kotikunta) i Finland, har du vanligen rätt att använda dig av den kommunens tjänster.
Det lönar sig för dig att utreda om du och de andra medlemmarna i din familj har rätt till en hemkommun i Finland.
Rätten till en hemkommun i Finland bestäms enligt hemkommunslagen.
Vid magistraten (maistraatti) på din egen boningsort kan du ta reda på om du har rätt till en hemkommun i Finland.
Hur kan du få en hemkommun i Finland
För att du ska kunna få en hemkommun i Finland måste du flytta till och vara stadigvarande bosatt i Finland.
Om du bor i Finland tillfälligt, till exempel om du flyttar till Finland för studier eller jobb under högst ett år, kan du vanligen inte få en hemkommun i Finland.
Du har möjlighet att få en hemkommun i Finland om:
du är finsk medborgare
du är medborgare i ett nordiskt land
du är medborgare i EU, Schweiz eller Liechtenstein och du har registrerat din uppehållsrätt i Finland
du har permanent (P) eller kontinuerligt (A) uppehållstillstånd som är i kraft
du är familjemedlem till en person som har en hemkommun i Finland
Om du har ett tillfälligt uppehållstillstånd (B-tillstånd) som är i kraft kan du få en hemkommun om du kan påvisa att det är din avsikt att bo stadigvarande i Finland.
Stadigvarande boende kan påvisas till exempel genom följande omständigheter:
du har en arbetsplats i Finland och ditt arbetskontrakt är i kraft minst två år
du studerar i Finland och dina studier räcker minst två år
du är av finländsk härkomst
du har tidigare haft en hemkommun i Finland
du har varit fortlöpande bosatt i Finland under minst ett års tid.
Din hemkommun är vanligen den kommun du bor i.
Om du inte har en bostad eller om du har bostäder på flera kommuners område är din hemkommun den kommun som du själv uppfattar som din hemkommun och som du har någon fast förbindelse till, till exempel genom familjeförhållanden eller arbetsplats.
Kontaktuppgifter till magistratfinska _ svenska _ engelska
Lag om hemkommunfinska _ svenska
Återkallande av uppehållstillstånd
Om du flyttar utomlands
Om ditt äktenskap eller registrerade parförhållande upphör
Om du förlorar ditt jobb
Återkallande av uppehållstillstånd
Ditt permanenta eller tidsbegränsade uppehållstillstånd återkallas om
du flyttar permanent från Finland
du har vistats två år utomlands utan avbrott.
Ditt permanenta eller tidsbegränsade uppehållstillstånd kan också återkallas om
du har uppgett felaktiga uppgifter i din ansökan om tillstånd
du har hemlighållit information som hade kunnat förhindra att tillståndet beviljas
ett annat Schengen-land begär att Finland återkallar ditt uppehållstillstånd.
Ett tidsbegränsat uppehållstillstånd kan också återkallas om de grunder på vilka tillståndet beviljades inte längre gäller.
Beslut om återkallelse av uppehållstillstånd fattas av Migrationsverket.
Om du flyttar utomlands
Om du ämnar flytta utomlands från Finland för två år, till exempel på grund av arbete eller studier, kan du ansöka hos Migrationsverket om att ditt uppehållstillstånd inte återkallas.
Ansökan är fritt formulerad men datum, underskrift och dina personuppgifter ska finnas med.
Ur ansökan bör även framgå hur länge och varför du studerar utomlands.
I din ansökning ska du motivera varför ditt uppehållstillstånd inte bör återkallas.
Ansökan ska göras innan du har vistats utomlands två år.
Om din finländska arbetsgivare har sänt dig utomlands för att arbeta förlorar du inte ditt uppehållstillstånd i Finland även om du vistas utomlands på grund av arbetet i över två år.
Om ditt äktenskap eller registrerade parförhållande upphör
Om du har ett tidsbestämt uppehållstillstånd med familjeband som grund kan det faktum att äktenskapet eller det registrerade parförhållandet upphör påverka uppehållstillståndet.
Om familjebandet inte längre existerar kan det hända att uppehållstillståndet inte förlängs.
Det är även möjligt att ett existerande tillstånd upphävs.
Uppehållstillståndet kan dock förlängas om du fortsättningsvis har starka band till Finland.
Exempel på sådana är:
barn eller andra familjemedlemmar i Finland
arbetsplats eller eget företag i Finland
studieplats i Finland
Om du skiljer dig på grund av att din make/maka varit våldsam mot dig kan ditt uppehållstillstånd förlängas trots skilsmässan.
Du ska lämna in en redovisning, exempelvis läkarintyg eller utlåtande från familjerådgivning.
Bifoga även till ansökan om uppehållstillstånd din egen redovisning av situationen.
Mer information om skilsmässa och upplösande av ett registrerat parförhållande hittar du på InfoFinlands sidor Skilsmässa.
Om du förlorar ditt jobb
Om du har ett uppehållstillstånd för arbetstagare som endast gäller arbete för en viss arbetsgivare och du förlorar din arbetsplats, ska du ansöka om ett nytt uppehållstillstånd för arbetstagare eller ett uppehållstillstånd på andra grunder.
Om Migrationsverket har beviljat dig ett uppehållstillstånd för arbetstagare och din anställning upphör tidigare än uppehållstillståndet, måste du eller din arbetsgivare skriftligt meddela Migrationsverket att din anställning upphör.
Om ditt uppehållstillstånd för arbetstagare inte har begränsats att gälla arbete för en viss arbetsgivare, utan för en viss bransch och tillståndet är fortfarande giltigt, kan du byta jobb inom samma bransch.
Mer information om arbete och företagande i Finland hittar du på InfoFinlands sida Arbete och entreprenörskap.
Mer information om uppehållstillstånd för arbetstagare och företagare hittar du på sidan Arbeta i Finland och Till Finland som företagare.
Om du redan har haft ett uppehållstillstånd i Finland, men tillståndet inte förlängs, fattar Migrationsverket beslut om utvisning.
Om du begår brott i Finland, kan du även utvisas på grund av brotten.
Om du blir utvisad, förfaller ditt eventuella giltiga uppehållstillstånd och du måste lämna landet.
Vanligtvis får du en tidsfrist inom vilken du måste lämna Finland.
Om du inte lämnar Finland inom tidsfristen avlägsnar polisen eller gränsbevakningsväsendet dig ur landet.
Enligt lag kan du inte utvisas om du hotas av dödsstraff, tortyr, förföljelse eller någon annan behandling som är omänsklig eller kränker människovärdet i ditt hemland.
Återkallelse av uppehållstillståndfinska _ svenska _ engelska
Avvisning och utvisningfinska _ svenska _ engelska
Flytta till Finland
Fortsatt uppehållstillstånd
Studera finska språket
Arbete och studier
Äktenskap och samboförhållande
Social trygghet
Tjänster för barnfamiljer
Hälsa
Flytta till Finland
Om du inte är medborgare i ett nordiskt land, EU-medborgare eller familjemedlem till en EU-medborgare som är bosatt i Finland, behöver du ett uppehållstillstånd.
Läs mer på InfoFinlands sida Familjen till Finland.
Om du är EU-medborgare behöver du inte uppehållstillstånd i Finland.
Om du vistas i Finland mer än tre månader, behöver du ett registreringsintyg för EU-medborgare (Unionin kansalaisen rekisteröintitodistus).
Läs mer på InfoFinlands sida EU-medborgare.
Om du inte är EU-medborgare, men din familjemedlem som är bosatt i Finland är EU-medborgare, behöver du ett uppehållskort för familjemedlem (perheenjäsenen oleskelukortti).
Läs mer på InfoFinlands sida EU-medborgare.
Om du är medborgare i ett nordiskt land behöver du inte uppehållstillstånd i Finland.
Läs mer på InfoFinlands sida Medborgare i nordiska länder.
På InfoFinlands sida Komihåglista för dig som flyttar till Finland hittar du nyttig information om vilka andra saker du bör ta hand om innan du flyttar till Finland.
När du flyttar till Finland ska du besöka magistraten (maistraatti)på orten där du är bosatt.
Vid magistraten kan du få en finsk personbeteckning, om du inte har ansökt om detta samtidigt som du ansökte om uppehållstillstånd.
På magistraten utreder man även om det är möjligt att registrera en hemkommun i Finland för dig.
När du har en hemkommun kan du använda kommunens tjänster, såsom till exempel hälsovårdstjänster.
Läs mer på InfoFinlands sida Hemkommun i Finland.
Till Finland på grund av familjebandfinska _ svenska _ engelska
Registrering av uppehållsrätt för EU-medborgarefinska _ svenska _ engelska
Registrering av utlänningarfinska _ svenska _ engelska
Fortsatt uppehållstillstånd
Om du har ett uppehållstillstånd ska du komma ihåg att ansöka om fortsatt uppehållstillstånd i god tid innan giltigheten för det första tillståndet tar slut.
Ansök om fortsatt uppehållstillstånd elektroniskt i tjänsten Enter Finland eller på Migrationsverkets tjänsteställe.
Tillståndsbeslutet är avgiftsbelagt.
Du måste betala avgiften samtidigt som du ansöker om fortsatt uppehållstillstånd.
Mer information om att ansöka om fortsatt uppehållstillstånd hittar du på InfoFinlands sida Fortsatt uppehållstillstånd.
Om du är EU-medborgare kan du ansöka om permanent uppehållsrätt när du har bott i Finland fem år.
Att förlänga uppehållstillståndetfinska _ svenska _ engelska
Studera finska språket
Information om studier i finska språket hittar du på InfoFinlands sida Finska och svenska språket.
Om du bor i Helsingforsregionen, Tammerforsregionen eller Åboregionen kan du leta efter en kurs i finska språket som passar dig genom tjänsten Finnishcourses.fi.
Kurser i finska och svenska språketfinska _ engelska _ ryska
Arbete och studier
Om du har uppehållstillstånd på grund av familjeband, har du rätt att arbeta och studera i Finland.
Även medborgare i EU-länder och nordiska länder och deras familjemedlemmar har rätt att arbeta och studera.
Notera att om du har ansökt om ditt första uppehållstillstånd i Finland så har du inte rätt att arbeta innan tillståndet har beviljats.
På InfoFinlands sida Var hittar jag jobb? hittar du information om jobbsökning i Finland.
Om du är intresserad av att grunda ett eget företag, gå in på InfoFinlands sida Att grunda ett företag.
Information om studier i Finland hittar du på InfoFinlands sida Utbildning.
Äktenskap och samboförhållande
Om du ska gifta dig i Finland hittar du nyttig information på InfoFinlands sida Äktenskap.
Information om att leva i ett samboförhållande i Finland hittar du på InfoFinlands sida Samboförhållande.
Du hittar information om skilsmässa på InfoFinlands sida Skilsmässa.
Notera att om du har ett uppehållstillstånd som beviljats på basis av familjeband, så kan förändringar i familjeförhållandena, såsom till exempel skilsmässa, påverka ditt uppehållstillstånd.
Läs mer på InfoFinlands sida Kan jag förlora mitt uppehållstillstånd?
På InfoFinlands sida Problem i äktenskap och parförhållande hittar du information om var du kan söka hjälp för problem i förhållandet.
Social trygghet
Om du flyttar till Finland av familjeskäl omfattas du vanligen av det finländska socialskyddet.
Detta är ändå inte alltid fallet.
Du kan kontrollera saken vid Fpa.
Social trygghet för dig som flyttar till Finlandfinska _ svenska _ engelska
Tjänster för barnfamiljer
Information om de tjänster och stöd som samhället erbjuder barnfamiljer hittar du på InfoFinlands sida Ekonomiskt stöd till familjer och Vård av barnet.
Hälsa
I Finland finns både offentliga och privata hälsovårdstjänster.
De offentliga hälsovårdstjänsterna är förmånligare än de privata.
Om du har en hemkommun i Finland kan du använda offentliga hälsovårdstjänster.
Om du flyttar till Finland av familjeskäl får du vanligen en hemkommun i Finland.
Magistraten fattar beslut om registrering av hemkommun.
Läs mer på InfoFinlands sida Hälsovårdstjänster i Finland och Hemkommun i Finland.
När du har flyttat till Finland ska du besöka magistraten på din hemort för att registrera dig som invånare.
Innan du besöker magistraten kan du fylla i Registreringsanmälan för utlänningar som finns på adressen maistraatti.fi.
Du kan även fylla i anmälan på magistraten.
Magistraten registrerar dina uppgifter i det finska befolkningsdatasystemet.
Dessa uppgifter är bland annat namn, födelsedatum, medborgarskap, kön och adress.
Om du flyttar till Finland för att bo här stadigvarande i ett år eller längre kan du ha rätt till hemkommun i Finland.
Du behöver en hemkommun för att kunna använda kommunala tjänster, såsom hälso- och sjukvården eller dagvården.
Magistraten utreder om du kan få en hemkommun registrerad.
När du besöker magistraten, ta med dig minst följande handlingar:
Om du är EU-medborgare eller nordisk medborgare:
Giltigt pass eller annan identitetshandling som styrker ditt medborgarskap
Arbetsavtal, intyg om studier eller någon annan utredning över registreringsbehovet (om du är EU-medborgare och ännu inte har registrerat din uppehållsrätt vid Migrationsverket)
Äktenskapsintyget i original (om du är gift)
Dina barns födelseattester i original (om du har barn under 18 år som flyttar till Finland)
Observera att du måste legalisera handlingar som har utfärdats av myndigheter utanför EU eller Norden.
Det gäller till exempel äktenskapsintyg som utfärdats i USA.
Om du är medborgare i något annat land:
Giltigt pass
Uppehållstillstånd (om du behöver uppehållstillstånd i Finland)
Vid behov utredning över arbete eller studier i Finland (t.ex. arbetsavtal eller närvarointyg som utfärdats av din läroanstalt) eller någon annan utredning över orsakerna till registreringen
Legaliserat äktenskapsintyg i original (om du är gift)
Legaliserade födelseattester för dina barn i original (om du har barn under 18 år som flyttar till Finland)
Legalisering av handlingar
På magistraten ska du visa upp originalhandlingen eller en vidimerad kopia av den.
Kopian kan pålitligt vidimeras av den myndighet som utfärdat handlingen eller notarius publicus i det land där handlingen utfärdades.
Handlingen ska vara legaliserad för att magistraten ska kunna föra in dina uppgifter i befolkningsdatasystemet.
Om ditt land har tillträtt Haagkonventionen ska du begära om ett så kallat Apostille-intyg för din handling.
Du behöver inget Apostille-intyg om du har en allmän handling som utfärdats av en myndighet i ett EU-land.
Du kan emellertid behöva en standardblankett som används som översättningsstöd som bilaga till en allmän handling.
Du får mer information om dessa standardblanketter hos myndigheterna i det land där du begär intyget.
Ett annat alternativ är att handlingen översätts av en auktoriserad översättare som godkänts av ett EU-land.
Observera att handlingarna ska vara på finska, svenska eller engelska.
Om din handling är på något annat språk måste du se till att få den översatt till finska, svenska eller engelska.
En auktoriserad översättare kan översätta handlingen åt dig.
Om översättningen görs utomlands måste även översättningen vara legaliserad.
Om du behöver mer information om legalisering av handlingar, kontakta magistraten eller utrikesministeriet i ditt eget land.
Finsk personbeteckning
Du får en personbeteckning av Migrationsverket när du beviljas uppehållstillstånd i Finland eller när din uppehållsrätt för EU-medborgare registreras.
Du kan även få en finsk personbeteckning vid:
skattebyrån, om du behöver personbeteckningen för beskattningen.
Den finska personbeteckningen är en nummerserie med elva siffror som bildas baserat på ditt födelsedatum och ditt kön.
Du behöver personbeteckningen till exempel för din arbetsgivare eller läroanstalt.
Den underlättar även skötseln av många officiella ärenden.
Om du har fått din personbeteckning någon annanstans än vid magistraten och vill ha en hemkommun, måste du även besöka magistraten.
Läs mer på InfoFinlands sida Hemkommun i Finland.
Registrering av utlänningarfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Registrering av utlänningar på skattebyrånfinska _ svenska _ engelska
Om du redan är i Finland och får ett negativt beslut om uppehållstillstånd från Migrationsverket (Maahanmuuttovirasto), måste du antingen lämna Finland eller överklaga beslutet.
Du får vistas i Finland så länge som behandlingen av besvären pågår.
Du kan överklaga också om du har ansökt om uppehållstillstånd utomlands.
Då måste du vänta på behandlingen av besvären utomlands.
Om du är asylsökande i Finland eller offer för människohandel, har du rätt att få stöd för frivillig återresa (vapaaehtoisen paluun tuki), om du beslutar att återvända till ditt hemland.
Läs mer under rubriken Stöd för frivillig återresa.
Att överklaga ett beslut om uppehållstillstånd
En besvärsanvisning om hur beslutet får överklagas bifogas alltid beslutet.
Besvären behandlas av förvaltningsdomstolen (hallinto-oikeus).
Förvaltningsdomstolen kan antingen avslå besvären eller sända ärendet till Migrationsverket för ny behandling.
Avslag innebär att Migrationsverkets beslut förblir gällande.
Om förvaltningsdomstolen avslår besvären kan du i vissa fall ansöka om besvärstillstånd hos högsta förvaltningsdomstolen (korkein hallinto-oikeus).
Om högsta förvaltningsdomstolen beviljar besvärstillstånd, behandlar den besvären.
Du kan få hjälp med att överklaga av antingen en privat jurist, en statlig rättshjälpsbyrå (valtion oikeusaputoimisto) eller Flyktingrådgivningen rf (Pakolaisneuvonta) (endast asylsökande).
På InfoFinlands sida Behöver du en jurist? finns mer information om hur du kan få hjälp i juridiska ärenden.
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Att lämna Finland
Om du får avslag på din ansökan om uppehållstillstånd eller om förvaltningsrätten avslår ditt överklagande, måste du lämna Finland.
Du ges möjlighet att lämna landet frivilligt.
Tidsfristen är vanligtvis 30 dagar.
Om du inte lämnar landet inom tidsfristen, avlägsnar polisen eller gränsbevakningsväsendet dig ur landet.
Du får inreseförbud till Schengenområdet om:
Du har brutit mot inresereglerna och din ansökan har avslagits, till exempel på grund av skenäktenskap.
Du har begått brott och du anses utgöra ett hot mot den allmänna ordningen och säkerheten.
Din asylansökan avslås i ett påskyndat förfarande.
Du inte lämnar landet frivilligt inom den tidsfrist som meddelats för dig.
När du har inreseförbud kan du inte besöka Finland eller något annat Schengenland.
Avvisning och utvisningfinska _ svenska _ engelska
Stöd för frivillig återresa
Om du vill återvända till ditt hemland kan du i vissa fall få stöd för frivilligt återvändande.
Stödet består antingen av pengar eller tjänster.
Penningsummans storlek beror på vilket land du återvänder till.
Tjänsten kan till exempel vara att du får hjälp med att leta efter en bostad eller arbetsplats i det land dit du återvänder.
Du kan få stöd om:
du har fått ett negativt beslut på din asylansökan
du återkallar din asylansökan
du är ett offer för människohandel och du inte har en hemkommun i Finland
du har ett tillfälligt uppehållstillstånd på grund av hinder för avlägsnande ur landet
du har fått tillfälligt skydd
din flyktingstatus i Finland har upphört eller återkallats eller det har fattats beslut om att avvisa dig
du har fått humanitärt skydd, men ditt uppehållstillstånd löper ut eller har redan löpt ut.
Om du är kund hos en mottagningscentral kan du ansöka om stöd för frivilligt återvändande vid din egen mottagningscentral.
Om du inte är kund hos en mottagningscentral kan du ansöka om stöd hos Migrationsverket.
Frivillig återflyttningfinska _ svenska _ engelska
Stöd för frivilligt återvändandefinska _ svenska _ engelska _ persiska _ arabiska
Vem är asylsökande?
Asylsökandes uppehållsrätt
Social trygghet
Familjeåterförening
Hälsa
Vem är asylsökande?
En asylsökande (turvapaikanhakija) är en person som söker skydd och uppehållsrätt i en främmande stat.
Internationellt skydd kan beviljas om personen känner välgrundad fruktan för förföljelse (på grund av ras, religion, tillhörighet till en viss samhällsgrupp eller politisk samhörighet) eller om personen annars är utsatt för verklig fara i sitt hemland eller sitt permanenta bosättningsland.
En asylsökande är alltså inte en flykting (pakolainen).
Om en asylsökande beviljas flyktingstatus eller uppehållstillstånd på grund av skyddsbehov eller på någon annan grund får han eller hon stanna i Finland.
Broschyren Information till asylsökandefinska _ svenska _ engelska _ ryska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
Asylsökandes uppehållsrätt
Du får stanna i Finland om du beviljas asyl eller uppehållstillstånd på någon annan grund.
Om förhållandena i ditt hemland är sådana att du inte behöver asyl och det inte heller finns andra grunder att bevilja uppehållstillstånd, avslås din ansökan och du utvisas från Finland.
Om du får avslag på din asylansökan eller ansökan om uppehållstillstånd har du rätt att överklaga beslutet.
Läs mer på InfoFinlands sida Som asylsökande till Finland.
Att söka asyl i Finlandfinska _ svenska _ engelska
Social trygghet
Asylsökande har inte rätt till finskt socialskydd.
Detta innebär att de inte har rätt till FPA:s förmåner.
Mottagningscentralen betalar mottagningspenning till asylsökande.
Den utbetalas så länge som asylansökan behandlas.
Mottagningspenningen är ett litet belopp som är avsett för ofrånkomliga utgifter.
Om den asylsökande beviljas uppehållstillstånd och är fast bosatt i Finland har han eller hon rätt till finskt socialskydd.
Man kan ansöka om att omfattas av det finska socialskyddet av FPA då uppehållstillstånd har beviljats.
Familjeåterförening
Asylsökande har inte rätt till familjeåterförening.
Dina familjemedlemmar kan inte få uppehållstillstånd i Finland på grund av familjeband.
Om du får uppehållstillstånd i Finland kan dina familjemedlemmar ansöka om tillstånd på grund av familjeband.
Läs mer på InfoFinlands sida Till familjemedlem i Finland.
Att söka uppehållstillstånd på grund av familjebandfinska _ svenska _ engelska
Hälsa
Asylsökande har vanligtvis inte tillgång till offentlig hälsoåvård exempelvis på hälsocentraler.
Mottagningscentralen anordnar hälsovårdstjänster för asylsökande.
Hälsovårdare på mottagningscentralen ser till att asylsökande får den vård de behöver.
Fråga mer på din mottagningscentral.
Om du fått uppehållstillstånd och din hemkommun finns i Finland kan du använda tjänsterna inom den offentliga hälsovården på samma sätt som de övriga invånarna i kommunen.
Hälsovård för papperslösa
Global Clinic är en klinik där du kan få hjälp eller råd av en läkare eller sjukskötare om du vistas i Finland utan uppehållstillstånd.
Du kan besöka Global Clinic även om du inte behöver brådskande sjukvård.
Global Clinic bedriver verksamhet i följande städer:
Åbo
Tammerfors
Uleåborg
Joensuu
Du kan ringa eller skicka e-post.
En sjukskötare eller läkare besvarar ditt samtal.
Du hittar kontaktinformation på Global Clinic:s hemsidor.
Global Clinic:s tjänster är avgiftsfria för kunderna.
Global Clinic anmäler inte sina kunder till polisen eller andra myndigheter.
Klinikens adress eller öppettider meddelas inte offentligt.
Kontaktuppgifterfinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Om du är medborgare i något nordiskt land behöver du inte uppehållstillstånd i Finland.
Du har rätt att jobba, fungera som företagare och studera i Finland.
När du flyttar till Finland måste du göra en flyttanmälan och gå och registrera dig vid magistraten (maistraatti) på din egen hemort.
Notera att du måste besöka magistraten personligen.
Gör flyttanmälan senast inom en vecka från din flyttningsdag.
För registreringen behöver du ett officiellt identitetskort där ditt medborgarskap framgår eller pass som är i kraft.
Familjemedlemmar till nordiska medborgare
Om en av dina familjemedlemmar, som flyttar med dig till Finland, inte är medborgare i ett nordiskt land, kan han/hon behöva uppehållstillstånd eller ett registreringsintyg över uppehållsrätt för EU-medborgare.
Läs mer på InfoFinlands sidor EU-medborgare eller Icke-EU-medborgare.
Finsk personbeteckning
När du registrerar dig vid magistraten kan du på samma gång få en finsk personbeteckning (henkilötunnus).
Du behöver en personbeteckning när du sköter ärenden hos myndigheter, och dessutom underlättar den skötandet av ärenden i till exempel banker och med din arbetsgivare.
Läs mer på InfoFinlands sidor Registrering som invånare.
Registrering av utlänningarfinska _ svenska _ engelska
Information för nordiska medborgarefinska _ svenska _ engelska _ norska
_ danska
_ isländska
Rådgivningstjänst för nordiska medborgarefinska _ engelska _ norska
_ danska
_ isländska
Rådgivning i uppehållstillståndsärenden
Om du har problem eller oklarheter med uppehållstillståndet, kan du ta kontakt med följande instanser för att be om råd:
Finlands beskickningar utomlands
Invandrarrådgivarna i din kommun i Finland
På Migrationsverkets webbplats finns mycket information om uppehållstillstånd.
Migrationsverket ger rådgivning angående tillstånd också per telefon.
Finlands beskickningar utomlands betjänar personer som ansöker om uppehållstillstånd i utlandet.
Många städer har rådgivningstjänster för invandrare med rådgivare som specialiserat sig på invandringsfrågor.
Flyktingsrådgivningen bistår asylsökande juridiskt i asylprocessen.
Dessutom tillhandahåller Flyktingrådgivningen allmän juridisk rådgivning för andra utlänningar.
Vänligen observera att endast Migrationsverket kan fatta beslut om uppehållstillstånd.
Information om uppehållstillståndfinska _ svenska _ engelska
linkkiFlyktingrådgivningen rf:
Juridisk rådgivningfinska _ engelska _ franska _ arabiska
Vem är flykting?
Familjeåterförening
Eftersökning av försvunna anhöriga
Hälsa
Stöd för flyktingar
Vem är flykting?
En flykting är en person med flyktingstatus.
Flyktingstatus får de som beviljas asyl eller som tas till Finland i flyktingkvoten.
Kvotflyktingar
Man kan inte ansöka om att bli kvotflykting (kiintiöpakolainen) via myndigheterna i Finland.
Man kan inte heller föreslå en annan person, till exempel en släkting eller vän, som kvotflykting.
Finland tar som kvotflyktingar emot personer som har flyktingstatus enligt
Förenta nationernas flyktingorganisation UNHCR. Kvotflyktingarna väljs bland de personer som UNHCR föreslår till Finland.
De finländska myndigheterna intervjuar flyktingarna som UNHCR har föreslagit och väljer bland dem de personer som tas emot till Finland.
Intervjuerna görs i de länder där flyktingarna vistas, vanligen i flyktingläger eller i UNHCR:s lokaler.
Valet av kvotflyktingar påverkas till exempel av följande faktorer:
Flyktingen är i behov av internationellt skydd.
Flyktingens mänskliga rättigheter förverkligas inte i det land där han eller hon vistas.
Flyktingen utgör inget hot för Finlands säkerhet.
Flyktingen har förutsättningar att integreras i Finland.
En del flyktingar väljs utan intervju på basis av UNHCR:s dokument.
Dessa är vanligen nödfall, med andra ord flyktingar som är i ett brådskande behov av asyl till exempel av hälsorelaterade eller politiska orsaker.
Finlands riksdag beslutar hur många flyktingar som tas till landet.
Från och med år 2001 har Finlands flyktingkvot varit 750 personer per år.
Inrikesministeriet beslutar från vilka länder kvotflyktingarna tas.
Beviljande av flyktingstatus till asylsökande
En person kan erhålla flyktingstatus också genom att söka asyl i Finland.
Asylsökanden kan beviljas flyktingstatus om han eller hon har befogade skäl att frukta förföljelse i sitt hemland på grund av ras, religion, nationalitet, tillhörighet till en viss samhällsgrupp eller på grund av sin politiska uppfattning och då sökanden på grund av detta inte kan återvända till sitt hemland.
Asylsökande som inte beviljas flyktingstatus kan ändå få uppehållstillstånd i Finland på någon annan grund.
Läs mer på InfoFinlands sida Som asylsökande till Finland.
Information om val av kvotflyktingarfinska _ svenska _ engelska
Familjeåterförening
Också flyktingens familjemedlemmar kan få uppehållstillstånd i Finland.
Vilka som är familjemedlemmar definieras i lagen.
Endast dessa familjemedlemmar kan få uppehållstillstånd på grund av familjeband.
I Finland betraktas som familjemedlemmar
registrerad partner
sambo
vårdnadshavaren till ett barn under 18 år.
För att familjemedlemmarna ska kunna få uppehållstillstånd, krävs det i vissa fall att flyktingen har en tillräcklig inkomst för att försörja sina familjemedlemmar i Finland.
Mer information om familjeåterförening finns på InfoFinlands sida Till familjemedlem i Finland.
Hjälp med familjeåterföreningen
Om du har kommit till Finland som kvotflykting, kan Migrationsverket ersätta kostnaderna för en familjemedlems inresa.
Kostnaderna ersätts dock endast i de fall där familjebandet har funnits redan före du fick ditt första uppehållstillstånd i Finland.
Andra anhörigas resekostnader ersätts inte.
Endast kvotflyktingar kan få ersättning för familjemedlemmarnas resekostnader.
Finlands Rösa Kors hjälper med researrangemangen för kvotflyktingar
Migrationsverket ersätter resekostnaderna endast i det fall att familjemedlemmen reser till Finland på en resa som arrangeras av Finlands Röda Kors och Internationella organisationen för migration.
Finlands Röda Kors hjälper med att ordna resan till Finland för kvotflyktingens familjemedlemmar när dessa fått uppehållstillstånd.
Röda Korset ger också rådgivning om reglerna för familjeåterförening och därom, hur familjemedlemmarna ska gå tillväga för att ansöka om familjeåterförening.
När Migrationsverket har gett ett positivt beslut på din ansökan om återförening på grund av familjeband och anser att staten kan bekosta resan för dina familjemedlemmar, skickar det sitt beslut till Röda Korset.
Om du har kommit till Finland som kvotflykting och vill att finska staten bekostar resan för dina familjemedlemmar ska du ta kontakt med Röda Korsets beredskapsenhet som sätter igång researrangemangen.
Finlands Röda Kors kan inte bistå familjemedlemmarnas flygresor eller andra resor ekonomiskt.
Att söka uppehållstillstånd på grund av familjebandfinska _ svenska _ engelska
Familjemedlem till en flyktingfinska _ svenska _ engelska
Eftersökning av försvunna anhöriga
Om du vill ha kontakt med en anhörig som försvunnit kan du be om hjälp vid personefterforskningen vid Finlands Röda Kors.
Röda Korset hjälper familjer som skilts åt vid olika katastrofer eller kriser.
Röda Korset söker försvunna anhöriga och förmedlar meddelanden på krisområden.
linkkiFinlands Röda Kors:
Efterforskning av anhörigafinska _ svenska _ engelska _ franska _ somaliska
linkkiFinlands Röda Kors:
Efterforskning av anhörigafinska _ svenska _ engelska _ ryska _ somaliska _ spanska _ persiska _ arabiska _ portugisiska
Hälsa
Om du har kommit till Finland som kvotflykting, har du hemkommun i Finland och då kan du använda de offentliga hälsovårdstjänsterna.
Stöd för flyktingar
Flyktingar och asylsökande kan söka hjälp och rådgivning i juridiska frågor bland annat vid Flyktingrådgivningen r.f. eller rättshjälpsbyråerna (oikeusaputoimisto).
Flyktingrådgivningen ger asylsökande rättshjälp i asylprocessens första skede.
Flyktingrådgivningen ger också andra utlänningar allmän rättshjälp.
Rättshjälpsbyråerna ger personer som är bosatta i Finland expertråd i skötseln av juridiska ärenden.
För att sköta ett juridiskt ärende kan man få ett rättsbiträde bekostat antingen helt eller delvis med statliga medel.
Finlands flyktinghjälp r.f. är en organisation som arbetar för att främja flyktingarnas grundläggande rättigheter.
Organisationens verksamhet i Finland omfattar informering, utbildning och socialarbete.
Flyktinghjälpen hjälper flyktingar och invandrare till exempel i frågor som rör integrationen, boendet och grundandet av egna organisationer.
linkkiFinlands flyktinghjälp r.f.:
Stöd till flyktingarfinska _ svenska _ engelska
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Om du behöver visum eller uppehållstillstånd för att vistas i Finland, men inte har det, vistas du illegalt i Finland.
Asylsökande har rätt att uppehålla dig i Finland även utan visum eller uppehållstillstånd under den tid som det tar att handlägga asylansökan.
Även om du har kommit lagligt till Finland kan din vistelse i landet bli illegal till exempel om du stannar kvar i landet fastän du inte beviljas ett uppehållstillstånd eller om ditt visum eller uppehållstillstånd har gått ut.
Information om hur du kan få ett uppehållstillstånd i Finland finns på InfoFinlands sida Flytta till Finland.
Hjälp och rådgivning
Mathjälp och inkvartering
Du har rätt till nödinkvartering och mathjälp om du inte har pengar till mat eller någonstans att övernatta.
Kommuner, församlingar och vissa organisationer ordnar nödinkvartering.
Juridisk rådgivning
Flyktingrådgivningen r.f. ger kostnadsfri juridisk rådgivning för papperslösa invandrare.
Rådgivningen betjänar telefonledes på numret 045-237 7104 (måndagar kl. 14–16).
Rådgivningen ges av en jurist.
Fler kontaktuppgifter hittar du på Flyktingrådgivningens webbplats.
Sjukvård
Om du blir sjuk eller skadas, har du rätt till brådskande vård inom den offentliga hälso- och sjukvården, till exempel på en hälsostation eller ett sjukhus.
Du måste i regel själv betala kostnaderna för vården.
I Helsingfors, Åbo, Tammerfors och Esbo får barn och gravida kvinnor samma hälso- och sjukvårdstjänster som övriga invånare.
De måste betala samma avgifter för vården som övriga invånare.
Global Clinic är en klinik där du kan få hjälp eller råd av en läkare eller sjukskötare om du vistas i Finland utan uppehållstillstånd.
Du kan besöka Global Clinic även om du inte behöver brådskande sjukvård.
Global Clinic bedriver verksamhet i följande städer:
Åbo
Tammerfors
Uleåborg
Joensuu
Du kan ringa eller skicka e-post.
En sjukskötare eller läkare besvarar ditt samtal.
Du hittar kontaktinformation på Global Clinic:s hemsidor.
Global Clinic:s tjänster är avgiftsfria för kunderna.
Global Clinic anmäler inte sina kunder till polisen eller andra myndigheter.
Klinikens adress eller öppettider meddelas inte offentligt.
linkkiFlyktingrådgivningen rf:
Juridisk rådgivningfinska _ engelska _ franska _ arabiska
Kontaktuppgifterfinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Du kan få permanent uppehållstillstånd (pysyvä oleskelulupa) (P), om
du bott i Finland i minst fyra år med A-tillstånd och
inte under tiden har bott utomlands i över två år och
grunden för de tidigare uppehållstillstånden fortfarande existerar
Om du hade A-tillstånd då du kom till Finland beräknas de fyra åren från den dag du anlände till Finland Om du fått A-tillstånd i Finland beräknas de fyra åren från den dag då det första A-tillståndet trädde i kraft.
Om du har fått internationellt skydd i Finland beräknas de fyra åren från att du anlände till Finland.
Permanent uppehållstillstånd kan eventuellt inte beviljas om:
du har begått ett brott som är belagt med fängelsestraff
du är misstänkt för ett brott som är belagt med fängelsestraff
du har begått två eller flera brott
du misstänks för två eller flera brott
Permanen uppehållstillstånd gäller tills vidare.
Tillstånet kan dras tillbaka om du permanent flyttar från Finland, uppehåller dig utomlands kontinuerligt i minst två år eller har lämnar felaktiga uppgifter då du ansökt om tillståndet.
EU-uppehållstillstånd för tredjelandsmedborgare som uppehållit sig länge i landet
Tredjelandsmedborgare äe medborgare i annat land än de nordiska länderna, EU-länderna, Liechtenstein eller Schweiz.
Du kan beviljas EU-uppehållstillstånd (P-EU) för tredjelandsmedborgare om:
du har bott i Finland i minst fem år med A-tillstånd och
inte under denna tid har bott utomlands längre än 10 månader och
grunden för de tidigare uppehållstillstånden fortfarande existerar
P-EU-tillstånd ansöks om på samma sätt som permanent uppehållstillstånd.
P-EU-tillstånd gäller tills vidare.
P-EU-tillståndsansökan kan även avslås på samma grunder som permanent uppehållstillstånd.
Ansökan
Du kan ansöka om permanent uppehållstillstånd på internet i tjänsten Enter Finland.
När du ställt ansökan ska du besöka Migrationsverkets tjänsteställe för att styrka din identitet.
Ta med dig en identitetshandling och originalexemplaren av ansökningsbilagorna.
Det är bra att boka en tid hos Migrationsverkets tjänsteställe i förväg.
Du kan boka tiden via Migrationsverkets elektroniska tidsbokningssystem.
Om du gjort ansökningen på internet, kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan, kommer detta att meddelas via ditt Enter Finland-konto.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du ansöka om tillståndet med en pappersblankett vid Migrationsverkets tjänsteställe.
Du kan skriva ut blanketten på Migrationsverkets webbplats.
Boka en tid vid tjänstestället och ta med dig den ifyllda ansökningen, bilagorna och en identitetshandling.
Handläggning av ansökan är avgiftsbelagd.
Avgiften ska betalas då ansökan ställs.
I tjänsten Enter Finland kan du betala med nätbankskoderna för en finsk bank eller med kreditkort.
Permanent uppehållstillståndfinska _ svenska _ engelska
Ansökningsblankettfinska _ svenska _ engelska
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Uppehållstillstånd
Studier i Finland
Boende
Arbete
Hälsa
Den sociala tryggheten
Utländsk examen i Finland
Uppehållstillstånd
Om du är medborgare i något av de nordiska länderna, ett EU-land, ett EES-land eller i Schweiz och kommer till Finland för att studera, måste du registrera din uppehållsrätt.
Läs mer på InfoFinlands sida EU-medborgare och Nordisk medborgare.
Om du är medborgare i något annat land behöver du ett uppehållstillstånd för studier.
Om dina studier i Finland pågår högst tre månader behöver du inget uppehållstillstånd.
Du kan ändå behöva ett visum.
Läs mer på InfoFinlands sida Att studera i Finland.
Information för utländska studerandeengelska
Studier i Finland
Du kan studera i Finland som utbytesstudent eller avlägga hela examen här.
Om du vill komma till Finland som utbytesstudent ska du kontakta till exempel studentexpeditionen eller den internationella enheten vid din egen läroanstalt.
På InfoFinlands sida Ansökan till utbildning hittar du information om hur du ansöker som examensstuderande till gymnasier, yrkesläroanstalter eller högskolor i Finland.
I Finland kan du studera på finska, svenska och ibland på engelska.
Högskolor ordnar engelskspråkig undervisning i vissa utbildningsprogram.
Läs mer på InfoFinlands sida Utländska studerande i Finland.
Boende
Om du är studerande kan du söka hyresbostäder som är speciellt avsedda för studerande.
Studentbostäder har ofta lägre hyra än vanliga bostäder.
Studentbostäder hyrs ut av studentbostadsstiftelser, universitetens studentkårer, nationer och vissa andra stiftelser.
Dessutom har vissa läroanstalter egna studenthem.
Fråga på din studieort var du kan söka en studentbostad.
Du kan söka bostad direkt när du blivit antagen till studier.
I de största städerna kan det ta flera veckor eller månader innan man får en bostad.
På InfoFinlands sida Boende hittar du mer information om hur du söker bostad och andra frågor i anslutning till boende.
Studentbostäderfinska _ engelska
Arbete
Om du är medborgare i ett EU-land, ett EES-land, Schweiz eller i något av de nordiska länderna, har du rätt att arbeta obegränsat under din studietid och du behöver inget särskilt tillstånd för det.
Arbete kan ge dig rätt till den sociala tryggheten i Finland.
Om du är medborgare i något annat land har du med ditt uppehållstillstånd för studerande rätt att arbeta i begränsad omfattning, om arbetet är
arbetspraktik som ingår i examen eller ett slutarbete eller
ett deltidsarbete, i genomsnitt högst 25 timmar per vecka under terminen
ett heltidsarbete under de tider då ingen undervisning ordnas vid läroanstalten, vanligen under sommar- och vinterlov.
På InfoFinlands sida Var hittar jag jobb? får du information om hur du söker arbete i Finland.
Studerandes rätt att arbetafinska _ svenska _ engelska
Hälsa
Om du kommer från ett annat nordiskt land till Finland för att studera har du rätt till sjukvård i Finland.
Du får vård på samma villkor och till samma kostnad som finländarna.
Ta med dig ett officiellt identitetsbevis när du använder hälsovårdstjänsterna.
Om du kommer från ett EU-land, ett EES-land eller Schweiz till Finland för att studera har du rätt till nödvändig sjukvård med det europeiska sjukvårdskortet.
Skaffa det europeiska sjukvårdskortet i ditt hemland innan du kommer till Finland.
Om du kommer från något annat land till Finland för att studera behöver du en omfattande sjukförsäkring innan du kan få uppehållstillstånd i Finland.
Mer information om uppehållstillstånd för studerande och om den sjukförsäkring som krävs för att få uppehållstillstånd får du på InfoFinlands sida Att studera i Finland eller på Migrationsverkets (Maahanmuuttovirasto) webbplats.
I Finland omfattas högskolestuderande av studerandehälsovården.
Fråga mer vid din egen läroanstalt.
Mer information om studerandehälsovården får du på Studenternas hälsovårdsstiftelses (SHVS) (YTHS) och social- och hälsovårdsministeriets (Sosiaali- ja terveysministeriö) webbplatser.
Du får information om hälsovårdstjänster i Finland på InfoFinlands sida Hälsa.
linkkiSHVS:
Hälsovård för högskolestuderandefinska _ svenska _ engelska
linkkiSocial- och hälsovårdsministeriet:
Studerandehälsovårdfinska _ svenska
Den sociala tryggheten
Om du flyttar till Finland tillfälligt har du vanligtvis inte rätt till den sociala tryggheten i Finland.
Till exempel befinner sig en studerande vars enda orsak till vistelsen i landet är studierna tillfälligt i Finland.
Arbete kan ge dig partiell rätt till social trygghet i Finland.
Läs mer på InfoFinlands sida Den sociala tryggheten i Finland.
Social trygghet för dig som flyttar till Finlandfinska _ svenska _ engelska
Utländsk examen i Finland
Om du har avlagt en examen utomlands kan du ha nytta av jämställande av examen, erkännande av yrkeskompetens eller av att skaffa dig rätt till yrkesutövning eller en fristående examen.
På InfoFinlands sida Utländska examina i Finland hittar du information om hur du kan få din examen eller dina studier erkända i Finland.
linkkiUtbildningsstyrelsen:
Erkännande av en examenfinska _ svenska _ engelska
Återkallande av uppehållstillstånd
Om du flyttar utomlands
Om ditt äktenskap eller registrerade parförhållande upphör
Om du förlorar ditt jobb
Återkallande av uppehållstillstånd
Ditt permanenta eller tidsbegränsade uppehållstillstånd återkallas om
du flyttar permanent från Finland
du har vistats två år utomlands utan avbrott.
Ditt permanenta eller tidsbegränsade uppehållstillstånd kan också återkallas om
du har uppgett felaktiga uppgifter i din ansökan om tillstånd
du har hemlighållit information som hade kunnat förhindra att tillståndet beviljas
ett annat Schengen-land begär att Finland återkallar ditt uppehållstillstånd.
Ett tidsbegränsat uppehållstillstånd kan också återkallas om de grunder på vilka tillståndet beviljades inte längre gäller.
Beslut om återkallelse av uppehållstillstånd fattas av Migrationsverket.
Om du flyttar utomlands
Om du ämnar flytta utomlands från Finland för två år, till exempel på grund av arbete eller studier, kan du ansöka hos Migrationsverket om att ditt uppehållstillstånd inte återkallas.
Ansökan är fritt formulerad men datum, underskrift och dina personuppgifter ska finnas med.
Ur ansökan bör även framgå hur länge och varför du studerar utomlands.
I din ansökning ska du motivera varför ditt uppehållstillstånd inte bör återkallas.
Ansökan ska göras innan du har vistats utomlands två år.
Om din finländska arbetsgivare har sänt dig utomlands för att arbeta förlorar du inte ditt uppehållstillstånd i Finland även om du vistas utomlands på grund av arbetet i över två år.
Om ditt äktenskap eller registrerade parförhållande upphör
Om du har ett tidsbestämt uppehållstillstånd med familjeband som grund kan det faktum att äktenskapet eller det registrerade parförhållandet upphör påverka uppehållstillståndet.
Om familjebandet inte längre existerar kan det hända att uppehållstillståndet inte förlängs.
Det är även möjligt att ett existerande tillstånd upphävs.
Uppehållstillståndet kan dock förlängas om du fortsättningsvis har starka band till Finland.
Exempel på sådana är:
barn eller andra familjemedlemmar i Finland
arbetsplats eller eget företag i Finland
studieplats i Finland
Om du skiljer dig på grund av att din make/maka varit våldsam mot dig kan ditt uppehållstillstånd förlängas trots skilsmässan.
Du ska lämna in en redovisning, exempelvis läkarintyg eller utlåtande från familjerådgivning.
Bifoga även till ansökan om uppehållstillstånd din egen redovisning av situationen.
Mer information om skilsmässa och upplösande av ett registrerat parförhållande hittar du på InfoFinlands sidor Skilsmässa.
Om du förlorar ditt jobb
Om du har ett uppehållstillstånd för arbetstagare som endast gäller arbete för en viss arbetsgivare och du förlorar din arbetsplats, ska du ansöka om ett nytt uppehållstillstånd för arbetstagare eller ett uppehållstillstånd på andra grunder.
Om Migrationsverket har beviljat dig ett uppehållstillstånd för arbetstagare och din anställning upphör tidigare än uppehållstillståndet, måste du eller din arbetsgivare skriftligt meddela Migrationsverket att din anställning upphör.
Om ditt uppehållstillstånd för arbetstagare inte har begränsats att gälla arbete för en viss arbetsgivare, utan för en viss bransch och tillståndet är fortfarande giltigt, kan du byta jobb inom samma bransch.
Mer information om arbete och företagande i Finland hittar du på InfoFinlands sida Arbete och entreprenörskap.
Mer information om uppehållstillstånd för arbetstagare och företagare hittar du på sidan Arbeta i Finland och Till Finland som företagare.
Om du redan har haft ett uppehållstillstånd i Finland, men tillståndet inte förlängs, fattar Migrationsverket beslut om utvisning.
Om du begår brott i Finland, kan du även utvisas på grund av brotten.
Om du blir utvisad, förfaller ditt eventuella giltiga uppehållstillstånd och du måste lämna landet.
Vanligtvis får du en tidsfrist inom vilken du måste lämna Finland.
Om du inte lämnar Finland inom tidsfristen avlägsnar polisen eller gränsbevakningsväsendet dig ur landet.
Enligt lag kan du inte utvisas om du hotas av dödsstraff, tortyr, förföljelse eller någon annan behandling som är omänsklig eller kränker människovärdet i ditt hemland.
Återkallelse av uppehållstillståndfinska _ svenska _ engelska
Avvisning och utvisningfinska _ svenska _ engelska
Om du har ett tillfälligt uppehållstillstånd (A- eller B-tillstånd) och orsaken för din vistelse i Finland ändras måste du ansöka om ett nytt uppehållstillstånd på den nya grunden.
Om du har ett permanent uppehållstillstånd (P) i Finland behöver du inte ändra grunden för ditt uppehållstillstånd även om orsaken till din vistelse ändras.
Du kan ansöka om uppehållstillstånd på något av följande grunder:
arbete
studier
familjeband
återflyttning
finländsk härkomst
internationellt skydd
annan orsak
Det är bra att komma ihåg att grunden för uppehållstillståndet kan påverka vilka rättigheter du har i Finland.
Till exempel ger ett uppehållstillstånd på grund av familjeband mer omfattande rätt att arbeta än ett tillstånd som beviljats på grund av studier.
Hur får jag ett tillfälligt uppehållstillstånd ändrat till ett kontinuerligt tillstånd?
Om du har ett tillfälligt uppehållstillstånd (B-tillstånd) kan du ansöka om ett kontinuerligt uppehållstillstånd (A-tillstånd) om grunden för vistelsen i Finland har ändrats från tillfällig till kontinuerlig.
Om du har ett tillfälligt uppehållstillstånd på grund av familjeband kan du ansöka om ett kontinuerligt uppehållstillstånd när en familjemedlem till dig ansöker om ett kontinuerligt uppehållstillstånd.
Du kan ansöka om ett kontinuerligt uppehållstillstånd också på någon annan grund om grunden är kontinuerlig.
Om du har ett tillfälligt uppehållstillstånd på grund av studier kan du få ett kontinuerligt tillstånd endast i det fall att grunden för din vistelse i Finland ändras.
Du kan inte få ett kontinuerligt tillstånd på basis av studier.
Grunden för din vistelse kan ändras till exempel om du får en arbetsplats i Finland eller gifter dig med en finsk medborgare eller en person som har kontinuerligt eller fortsatt tillstånd i Finland.
Om du har ett tillfälligt uppehållstillstånd för arbete eller näringsidkande kan du ansöka om ett kontinuerligt uppehållstillstånd när du har vistats i Finland två år utan avbrott.
Hur söker jag ett uppehållstillstånd på nya grunder?
Välj ansökningsblankett utifrån grunden för din ansökan om nytt tillstånd.
Lämna in din ansökan på internet i tjänsten Enter Finland eller vid Migrationsverkets tjänsteställe.
Mer information om ansökningsproceduren hittar du på InfoFinlands sida Fortsatt uppehållstillstånd.
Från studerande till anställd
Om du har avlagt en examen i Finland kan du få ett uppehållstillstånd för att söka arbete.
När du är klar med dina studier och ditt uppehållstillstånd för studerande går ut, kan du ansöka om fortsatt tillstånd (jatkolupa) för att söka arbete.
Tillståndet är i kraft ett år.
Detta tillstånd kan endast fås en gång och det kan inte förnyas.
När du får en arbetsplats kan du få uppehållstillstånd på grund av arbete.
Uppehållstillstånd på en ny grundfinska _ svenska _ engelska
Uppehållstillstånd för sökande av arbetefinska _ svenska _ engelska
Uppehållstillstånd
Fortsatt uppehållstillstånd
Arbete och företagande i Finland
Finska och svenska språket
Studier
Den sociala tryggheten
Hälsan
Uppehållstillstånd
Om du är medborgare i något av de nordiska länderna, ett EU-land, ett EES-land eller i Schweiz och kommer till Finland för att arbeta eller driva ett företag, måste du registrera din uppehållsrätt.
Läs mer på InfoFinlands sida EU-medborgare.
Om du är medborgare i något annat land behöver du ett uppehållstillstånd för arbetstagare.
Om du redan befinner dig i Finland på någon annan grund kan du ha rätt att arbeta även om du inte har ansökt om ett uppehållstillstånd på grund av arbete.
Läs mer på InfoFinlands sida Till Finland för att arbeta.
Om du inte är medborgare i något av Europeiska unionens medlemsländer, ett EES-land eller i Schweiz och vill driva ett företag i Finland, behöver du ett uppehållstillstånd för företagare.
Mer information om uppehållstillstånd för företagare hittar du på InfoFinlands sida Bli företagare i Finland.
Arbete i Finlandfinska _ svenska _ engelska
Uppehållstillstånd för företagarefinska _ svenska _ engelska
Fortsatt uppehållstillstånd
Ansök om fortsatt uppehållstillstånd på internet i tjänsten Enter Finland eller på Migrationsverkets tjänsteställe.
Gör en ansökan innan ditt föregående uppehållstillstånd går ut.
Du får mer information om att ansöka om fortsatt uppehållstillstånd på InfoFinlands sida Fortsatt uppehållstillstånd.
Att förlänga uppehållstillståndetfinska _ svenska _ engelska
Arbete och företagande i Finland
I InfoFinlands avsnitt Arbete och företagande hittar du mycket information om arbetslivet och företagandet i Finland.
Finska och svenska språket
En del arbetsgivare ordnar undervisning i det finska språket för sina anställda.
Fråga din arbetsgivare som det ordnas undervisning i det finska språket på din arbetsplats.
Information om andra möjligheter att studera finska eller svenska hittar du i InfoFinlands avsnitt Finska och svenska språket.
Studier
Om du vill avlägga examen eller fortbilda dig kan du delta i fortbildning.
Fortbildning ordnas bland annat av läroanstalter, fackförbund och Institutet för Yrkenas befrämjande.
Också många arbetsplatser utbildar sina anställda till exempel i användningen av nya apparater eller program.
Studierna är inte alltid inriktade på att skaffa ett yrke.
Du kan också ha studier som hobby.
Läs mer på InfoFinlands sida Studier som hobby.
Grundläggande information om fortbildningfinska _ svenska
Den sociala tryggheten
Om du flyttar till Finland för att arbeta från EU-området eller ett EES-land eller Schweiz, omfattas du vanligtvis delvis av den sociala tryggheten i Finland också när din anställning endast är kortvarig.
Om du kommer till Finland som arbetstagare någon annanstans ifrån än ett EU-land, ett EES-land eller Schweiz påverkas din sociala trygghet av följande faktorer:
hur länge arbetet varar
från vilket land du flyttar till Finland.
De flesta av FPA:s förmåner är sådana att du har rätt till dem endast om du flyttar ditt stadigvarande boende till Finland.
Dessutom måste du uppfylla samma villkor för att få förmånen som alla andra som bor i Finland.
Om du inte flyttar stadigvarande till Finland, kan du i vissa situationer ändå ha rätt att åtminstone delvis omfattas av den sociala tryggheten i Finland medan du arbetar här.
Detta förutsätter att din arbetstid och lön uppfyller minimikraven.
Om du har anställning i Finland, är det skäl för dig att ansluta dig till en finländsk arbetslöshetskassa.
Om du är medlem av en arbetslöshetskassa kan du få inkomstrelaterad arbetslöshetsersättning, om du blir arbetslös.
Läs mer på InfoFinlands sidor Fackförbund och Arbetslöshetsförsäkring.
Social trygghet för dig som flyttar till Finlandfinska _ svenska _ engelska
Hälsan
Hälsovård för anställda och företagare
Om du har kommit till Finland för att arbeta har du vanligen rätt att använda de offentliga hälsovårdstjänsterna i Finland.
Detta beror på hurdant och hur långt arbetsavtal du har samt från vilket land du har kommit till Finland.
Du kan begära att FPA utreder din rätt till de offentliga hälsovårdstjänsterna.
Du hittar mer information om den offentliga hälso- och sjukvården på InfoFinlands sida Hälsovårdstjänster i Finland.
I Finland är arbetsgivare skyldiga att ordna förebyggande företagshälsovård för sina anställda.
Företagare kan ordna sin egen företagshälsovård om de vill.
Företagare måste alltså inte ordna företagshälsovård för sig.
Företagare måste ändå ordna företagshälsovård för sina anställda.
Företagshälsovården kan ordnas vid den lokala hälsovårdscentralen eller till exempel på en privat läkarcentral.
Mer information får du på InfoFinlands sida Företagshälsovården och på social- och hälsovårdsministeriets webbplats.
linkkiSocial- och hälsovårdsministeriet:
Företagshälsovårdfinska _ svenska _ engelska
Om du förlorar ditt jobb
Om du har ett uppehållstillstånd för arbetstagare som endast gäller arbete för en viss arbetsgivare och du förlorar din arbetsplats, ska du ansöka om ett nytt uppehållstillstånd för arbetstagare eller ett uppehållstillstånd på andra grunder.
Om Migrationsverket har beviljat dig ett uppehållstillstånd för arbetstagare och din anställning upphör tidigare än uppehållstillståndet, måste du eller din arbetsgivare skriftligt meddela Migrationsverket att din anställning upphör.
Om ditt uppehållstillstånd för arbetstagare inte har begränsats att gälla arbete för en viss arbetsgivare, utan för en viss bransch och tillståndet är fortfarande giltigt, kan du byta jobb inom samma bransch.
Problem i arbetslivet
Om du råkar ut för problematiska situationer på arbetsplatsen ska du först kontakta din chef.
Om ärendet inte kan lösas på arbetsplatsen, ska du kontakta arbetarskyddsdistriktet (työsuojelupiiri) i ditt område eller ditt fackförbund.
Information och råd om var du kan få hjälp med olika slags problem i arbetslivet hittar du på InfoFinlands sida Problem i arbetslivet.
Om du redan är i Finland och får ett negativt beslut om uppehållstillstånd från Migrationsverket (Maahanmuuttovirasto), måste du antingen lämna Finland eller överklaga beslutet.
Du får vistas i Finland så länge som behandlingen av besvären pågår.
Du kan överklaga också om du har ansökt om uppehållstillstånd utomlands.
Då måste du vänta på behandlingen av besvären utomlands.
Om du är asylsökande i Finland eller offer för människohandel, har du rätt att få stöd för frivillig återresa (vapaaehtoisen paluun tuki), om du beslutar att återvända till ditt hemland.
Läs mer under rubriken Stöd för frivillig återresa.
Att överklaga ett beslut om uppehållstillstånd
En besvärsanvisning om hur beslutet får överklagas bifogas alltid beslutet.
Besvären behandlas av förvaltningsdomstolen (hallinto-oikeus).
Förvaltningsdomstolen kan antingen avslå besvären eller sända ärendet till Migrationsverket för ny behandling.
Avslag innebär att Migrationsverkets beslut förblir gällande.
Om förvaltningsdomstolen avslår besvären kan du i vissa fall ansöka om besvärstillstånd hos högsta förvaltningsdomstolen (korkein hallinto-oikeus).
Om högsta förvaltningsdomstolen beviljar besvärstillstånd, behandlar den besvären.
Du kan få hjälp med att överklaga av antingen en privat jurist, en statlig rättshjälpsbyrå (valtion oikeusaputoimisto) eller Flyktingrådgivningen rf (Pakolaisneuvonta) (endast asylsökande).
På InfoFinlands sida Behöver du en jurist? finns mer information om hur du kan få hjälp i juridiska ärenden.
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Att lämna Finland
Om du får avslag på din ansökan om uppehållstillstånd eller om förvaltningsrätten avslår ditt överklagande, måste du lämna Finland.
Du ges möjlighet att lämna landet frivilligt.
Tidsfristen är vanligtvis 30 dagar.
Om du inte lämnar landet inom tidsfristen, avlägsnar polisen eller gränsbevakningsväsendet dig ur landet.
Du får inreseförbud till Schengenområdet om:
Du har brutit mot inresereglerna och din ansökan har avslagits, till exempel på grund av skenäktenskap.
Du har begått brott och du anses utgöra ett hot mot den allmänna ordningen och säkerheten.
Din asylansökan avslås i ett påskyndat förfarande.
Du inte lämnar landet frivilligt inom den tidsfrist som meddelats för dig.
När du har inreseförbud kan du inte besöka Finland eller något annat Schengenland.
Avvisning och utvisningfinska _ svenska _ engelska
Stöd för frivillig återresa
Om du vill återvända till ditt hemland kan du i vissa fall få stöd för frivilligt återvändande.
Stödet består antingen av pengar eller tjänster.
Penningsummans storlek beror på vilket land du återvänder till.
Tjänsten kan till exempel vara att du får hjälp med att leta efter en bostad eller arbetsplats i det land dit du återvänder.
Du kan få stöd om:
du har fått ett negativt beslut på din asylansökan
du återkallar din asylansökan
du är ett offer för människohandel och du inte har en hemkommun i Finland
du har ett tillfälligt uppehållstillstånd på grund av hinder för avlägsnande ur landet
du har fått tillfälligt skydd
din flyktingstatus i Finland har upphört eller återkallats eller det har fattats beslut om att avvisa dig
du har fått humanitärt skydd, men ditt uppehållstillstånd löper ut eller har redan löpt ut.
Om du är kund hos en mottagningscentral kan du ansöka om stöd för frivilligt återvändande vid din egen mottagningscentral.
Om du inte är kund hos en mottagningscentral kan du ansöka om stöd hos Migrationsverket.
Frivillig återflyttningfinska _ svenska _ engelska
Stöd för frivilligt återvändandefinska _ svenska _ engelska _ persiska _ arabiska
Det är viktigt att du ansöker om fortsatt uppehållstillstånd innan ditt tidigare uppehållstillstånd går ut.
Om ditt tidigare uppehållstillstånd går ut under behandlingen av ansökan får du uppehålla dig i Finland och har vanligtvis även rätt att arbeta under den tid som ansökan behandlas.
Om du ansöker om fortsatt uppehållstillstånd först efter att ditt tidigare uppehållstillstånd gått ut, får du uppehålla dig i Finland under tiden då ansökan behandlas men har inte rätt att arbeta innan du erhållit fortsatt uppehållstillstånd.
Att ansöka
Du kan ansöka om tillståndet på internet i tjänsten Enter Finland.
När du ställt ansökan ska du besöka Migrationsverkets tjänsteställe för att styrka din identitet.
Du ska besöka tjänstestället inom tre månader efter att ha gjort ansökan.
Ta med dig pass, passfoto och originalexemplaren av ansökningsbilagorna.
Det är bra att boka en tid hos Migrationsverkets tjänsteställe i förväg.
Du kan boka tiden via Migrationsverkets elektroniska tidsbokningssystem.
Om du gjort ansökningen på internet, kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan, kommer detta att meddelas via ditt Enter Finland-konto.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du ansöka om tillståndet med en pappersblankett vid Migrationsverkets tjänsteställe.
Skriv ut blanketten på Migrationsverkets webbplats och fyll i den färdigt.
Boka en tid vid tjänstestället.
När du ska besöka tjänstestället, ta med dig din ifyllda ansökan, bilagorna och kopior på bilagor samt pass och passfoto.
Migrationsverket beviljar dig fortsatt uppehållstillstånd om grunden för det tidigare uppehållstillståndet fortfarande existerar.
Du kan även ansöka om fortsatt uppehållstillstånd på annan grund än för det tidigare tillståndet
Hanteringen av ansökan är avgiftsbelagd. Avgiften ska betalas då ansökan görs.
I tjänsten Enter Finland kan du betala med nätbankskoderna för en finsk bank eller med kreditkort.
Att förlänga uppehållstillståndetfinska _ svenska _ engelska
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Blanketter för ansökan om uppehållstillståndfinska _ svenska _ engelska
Migrationsverket:
Presentation av e-tjänsten Enter Finland
Arbetstagare, företagare, studerande, flykting, asylsökande eller en familjemedlem till en person bosatt i Finland hittar information speciellt om sin egen situation på dessa sidor i Infobanken.
Via dessa sidor hittar du snabbt den information som du behöver i kortfattade form.
Arbetstagare eller företagare
Studerande
Flykting
Asylsökande
Familjemedlem
Rådgivning i uppehållstillståndsärenden
Om du har problem eller oklarheter med uppehållstillståndet, kan du ta kontakt med följande instanser för att be om råd:
Finlands beskickningar utomlands
Invandrarrådgivarna i din kommun i Finland
På Migrationsverkets webbplats finns mycket information om uppehållstillstånd.
Migrationsverket ger rådgivning angående tillstånd också per telefon.
Finlands beskickningar utomlands betjänar personer som ansöker om uppehållstillstånd i utlandet.
Många städer har rådgivningstjänster för invandrare med rådgivare som specialiserat sig på invandringsfrågor.
Flyktingsrådgivningen bistår asylsökande juridiskt i asylprocessen.
Dessutom tillhandahåller Flyktingrådgivningen allmän juridisk rådgivning för andra utlänningar.
Vänligen observera att endast Migrationsverket kan fatta beslut om uppehållstillstånd.
Information om uppehållstillståndfinska _ svenska _ engelska
linkkiFlyktingrådgivningen rf:
Juridisk rådgivningfinska _ engelska _ franska _ arabiska
Finland tillhör Schengenområdet.
Länderna som tillhör Schengenområdet har enhetlig visering.
Utlänningar som vill resa till Finland för en kort tid, till exempel på semester, affärsresa eller på besök hos släktingar, behöver ett visum om de inte är medborgare i ett viseringsfritt land.
Ett visum är ett inresetillstånd för en kortvarig och tillfällig, högst tre månader lång vistelse.
På utrikesministeriets webbplats eller vid den närmast belägna finländska beskickningen kan du kontrollera om du behöver ett visum i Schengenområdet.
Visumbehovet till Schengenområdet och av
Finland accepterade resedokumentfinska _ svenska _ engelska
Information för viseringsfria personer
Du kan resa till Finland och de övriga Schengenländerna om du har ett giltigt pass eller något annat resedokument som godkänns i Finland.
Du får vistas högst tre månader under en period på sex månader i Finland och de övriga Schengenländerna räknat från den dag du reste in till Schengenområdet.
Information för viseringsskyldiga personer
Du ska alltid ha ett visum när du kommer till Finland eller något annat land i Schengenområdet.
Du får vistas i Finland eller något annat land i Schengenområdet utan uppehållstillstånd så länge som ditt visum är i kraft.
Om du har ett visum eller uppehållstillstånd i något Schengenland kan du resa inom Schengenområdet utan att behöva skaffa ett separat visum för de andra Schengenländerna.
Så här ansöker du om Schengenvisum
Du ansöker om visum i den närmast belägna finländska beskickningen eller visumcentralen.
Du ska vistas lagligt i det land där du ansöker om visum. I länder där
Finland inte har en beskickning kan något annat land representera Finland i visumärenden.
I detta fall kan du ansöka om visum i detta lands beskickning.
På utrikesministeriets webbplats finns en förteckning över de länder där ett annat land representerar Finland i visumärenden.
Du ansöker om visum med en visumansökningsblankett.
Blanketten får du på utrikesministeriets webbplats och från beskickningar i Schengenländer.
Antalet bilagor som krävs till visumansökan kan variera beroende på i vilket land du söker visum.
Hos beskickningen kan du kontrollera vilka bilagor du behöver för din visumansökan.
Lämna din ansökning till den beskickning eller visumcentral dit du ställer din ansökan.
Du kan inte skicka din ansökning via e-post eller fax.
Förlängning av visum i Finland
Polisen kan förlänga uppehållstiden för ditt visum eller visumets utgångstid om du av motiverade skäl inte kan lämna Finland när ditt visum utgår.
Motiverade skäl för förlängning av visum kan till exempel vara:
en akut, svår sjukdom som hindrar dig från att resa,
en släkting som är bosatt i Finland har plötsligt insjuknat svårt eller avlidit,
inställt flyg på grund av strejk eller väderförhållanden,
viktiga affärsförhandlingar som pågår längre än väntat.
Information till medborgare från viseringsskyldiga länderfinska _ svenska _ engelska
Ansökan om Schengenvisumfinska _ svenska _ engelska
Länder där en annan Schengenstat representerar Finlandfinska _ svenska _ engelska
Förlängning av visum i Finlandfinska _ svenska _ engelska
Hjälp i nödsituationer
Beskickningarna hjälper sitt lands medborgare som hamnat i nödläge i Finland.
De kan till exempel hjälpa dig om du har råkat ut för en olycka, blivit sjuk eller fallit offer för ett brott.
Beskickningen kan bevilja dig ett nytt pass om ditt pass har gått förlorat eller stulits.
Om du är turist i Finland och hamnar i en svår situation, ska du kontakta ditt hemlands beskickning.
linkkiVisitFinland.com:
Information om Finland till turistersvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ japanska _ italienska
Före flytten till Finland
Efter flytten till Finland
Bekanta dig med innehållen i InfoFinland före flytten.
I InfoFinland hittar du pålitlig information på ditt eget språk om flytten till Finland, arbetslivet, boende, studier i finska eller svenska språket, utbildning, social trygghet, hälsotjänster, tjänster för familjer, problematiska situationer och fritid.
På sidorna finns nyttiga praktiska råd, kontaktuppgifter och länkar till tilläggsinformation.
Med hjälp av menyn Städer får du fram information om den kommun som du är intresserad av.
De olika språkversionerna av InfoFinlands är identiska.
Komihåglistan för dig som flyttar till Finland är avsedd att hjälpa dig med de viktigaste praktiska frågorna som har med flytten att göra.
Observera att listan inte nödvändigtvis innehåller allt som måste göras när du flyttar till Finland.
Före flytten till Finland
Uppehållstillstånd eller registrering av uppehållsrätt?
Om du ska vistas i Finland mer än 90 dagar och är EU-medborgare, måste du registrera din uppehållsrätt.
Om du är medborgare i ett land utanför EU, måste du ansöka om uppehållstillstånd i Finland.
Läs mer på InfoFinlands sida EU-medborgare eller Icke-EU-medborgare.
När du ansöker om uppehållstillstånd eller registrering av uppehållsrätten måste du bevisa att din utkomst i Finland är tryggad.
Om du kommer till Finland för att arbeta eller som företagare måste du bevisa att ditt arbete eller din företagsverksamhet inbringar dig en tillräcklig utkomst.
Om du flyttar till en familjemedlem i Finland, krävs det ofta även att den person som bor i Finland har tillräckliga medel för att försörja sig själv och den familjemedlem som flyttar till Finland.
Flyttsaker från EU-området
Om du flyttar till Finland från ett annat EU-land behöver du vanligen inte betala tull eller mervärdesskatt på dina flyttsaker, d.v.s. de personliga föremål som du tar med dig.
Du behöver inte heller anmäla dina flyttsaker i tullen (tulli).
Observera att tull- och skattefriheten för flyttsaker inte gäller alkohol eller tobaksprodukter.
För import av dessa gäller separata begränsningar.
Mer information får du på Tullrådgivningen +358 (0)295 5201 eller på tullens webbplats.
Tullrådgivningen betjänar på finska, svenska och engelska.
Flyttsaker från länder utanför EU
Om du flyttar till Finland från ett land som inte hör till EU behöver du vanligen inte betala tull eller mervärdesskatt på dina flyttsaker, d.v.s. de personliga föremål som du tar med dig.
Du måste dock göra en tullanmälan på flyttsakerna till de finländska tullmyndigheterna.
Som flyttsaker betraktas till exempel:
möbler och andra husgeråd
husdjur
cyklar och motorcyklar
bilar och släpvagnar avsedda för privat bruk.
Observera att tull- och skattefriheten för flyttsaker inte gäller alkohol eller tobaksprodukter.
För import av dessa gäller separata begränsningar.
linkkiTullen:
Införsel av flyttsaker till Finlandfinska _ svenska _ engelska _ ryska
Införsel av bil till Finland som flyttsak
När du tar med dig en bil till Finland som flyttsak, måste du tullanmäla den.
Om du tar med dig en bil till Finland måste du registrera den och betala bilskatt (autovero) för den innan du kan använda den i trafiken.
Man kan dock använda bilen tillfälligt innan bilskatten är betald.
Detta förutsätter att du har gjort en anmälan om ibruktagande av fordonet (auton käyttöönottoilmoitus) till skatteförvaltningen.
Du ska också ha en giltig trafikförsäkring (liikennevakuutus) för din bil i Finland.
Om du för in en bil från ett land utanför EES-området behöver du också ett förflyttningstillstånd innan du kan använda bilen.
Förflyttningstillstånd beviljas av besiktningskontor och vissa av Tullens verksamhetsställen.
Du får inte använda din bil i Finland förrän du har gjort en anmälan om ibruktagande av fordonet och skaffat ett förflyttningstillstånd.
Om du har frågor kring fordonsskatten eller anmälan om ibruktagande, kan du ringa skatteförvaltningens telefontjänst:
+358 (0)29 497 150 (finska)
+358 (0)29 497 151 (svenska)
+358 (0)29 497 152 (engelska)
linkkiTullen:
Fordon som flyttgodsfinska _ svenska _ engelska _ ryska
Införsel av sällskapsdjur
Om du vill ta med dig ett husdjur till Finland är det bra att på förhand bekanta sig med reglerna som gäller införsel av djur.
Ofta krävs till exempel att djuren har fått vissa vaccinationer.
Mer information om reglerna i Finland ges av Livsmedelssäkerhetsverket Evira.
linkkiEvira:
Införsel av djur från EU-länderfinska _ svenska _ engelska
linkkiEvira:
Införsel av djur från länder utanför EUfinska _ svenska _ engelska _ ryska
Flyttfirmor
En del företag som tillhandahåller flyttservice sköter också flytt från ett land till ett annat.
Du kan anlita dessa företag att transportera dina ägodelar från ett land till ett annat och också att packa dina saker och tillhandahålla förpackningsmaterial.
Flyttkostnaderna beror på varifrån du flyttar och hur mycket saker du har.
Tjänsterna och priserna i olika flyttfirmor kan variera stort och därför lönar det sig att jämföra.
Flyttjänsterfinska _ svenska _ engelska
linkkiViktor Ek:
Flyttjänsterfinska _ svenska _ engelska
Hjälp när du flyttarfinska _ svenska _ engelska _ norska
_ danska
Efter flytten till Finland
I den här listan har vi samlat de vanligaste ärendena som du måste ta hand om när du har kommit till Finland.
Bostad och hemförsäkring
De flesta invandrare bor först i en hyresbostad när de kommer till Finland.
Det är bra att reservera minst en månad för att söka hyresbostad.
Läs mer på InfoFinlands sida Boende.
När du har en bostad är det bra att också ta en hemförsäkring (kotivakuutus).
Hemförsäkringen ersätter till exempel skador på möbler och andra ägodelar.
Hemförsäkringar säljs av försäkringsbolag.Information om försäkringar finns på InfoFinlands sida Vardagslivet i Finland.
Finsk personbeteckning
När du ansöker om ditt första uppehållstillstånd i Finland eller om registrering av uppehållsrätten för EU-medborgare kan du samtidigt ansöka om en finsk personbeteckning.
Du kan även ansöka om en personbeteckning i Finland vid magistraten eller skattebyrån på din hemort.
Mer information hittar du på InfoFinlands sida Registrering som invånare.
Hemkommun i Finland
Om du flyttar till och blir stadigvarande bosatt i Finland registreras en hemkommun för dig i Finland.
Hemkommunen är den kommun där du bor.
När du har en hemkommun har du rätt att använda denna kommuns tjänster såsom till exempel offentliga hälsovårdstjänster.
Du kan ta reda på om det är möjligt att registrera en hemkommun i Finland för dig vid magistraten på din hemort.
Läs mer på InfoFinlands sida Hemkommun i Finland.
Registrering av utlänningarfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Registrering av utlänningar på skattebyrånfinska _ svenska _ engelska
Social trygghet
Huvudregeln är att du omfattas av den sociala tryggheten i Finland och har rätt till FPA:s förmåner om du bor stadigvarande i Finland.
Vad stadigvarande boende betyder definieras i lagen.
Du kan också ha rätt till den sociala tryggheten i Finland om du arbetar i Finland.
Det finns dock fler omständigheter som påverkar den sociala tryggheten, till exempel vilket land du kommer ifrån.
Social trygghet för dig som flyttar till Finlandfinska _ svenska _ engelska
Bankkonto
Du behöver ett bankkonto för att sköta din dagliga ekonomi.
När du öppnar ett bankkonto behöver du ett pass eller någon annan officiell identitetshandling.
Det lönar sig att jämföra tjänsterna och priserna som olika banker tillhandahåller så att du hittar det alternativ som är förmånligast för dig.
Information om att öppna ett bankonto finns på InfoFinlands sida Vardagslivet i Finland.
linkkiFinansbranschens Centralförbund:
Utländska medborgares bankärendenfinska _ engelska
Skattekort
Om du arbetar och får lön eller är företagare behöver du ett finskt skattekort (verokortti).
Skattekortet får du vid skattebyrån.
Läs mer om beskattningen i Finland på InfoFinlands sida Beskattning.
Kollektivtrafik
Om du bor i en stad är det inte nödvändigt att äga en bil.
Kollektivtrafiken fungerar väl i Finland.
Man kan resa nästan över allt i Finland med tåg eller buss.
Man kan också flyga till många städer.
I stora städer och deras näromgivning finns en välfungerande lokaltrafik.
Lokaltrafiken trafikeras vanligtvis med bussar.
Läs mer på InfoFinlands sida Trafiken i Finland.
Körkort
Om du har ett körkort som utfärdats i ett av de nordiska länderna eller i ett EU-/EES-land, är det giltigt även i Finland.
Om du bor stadigvarande i Finland kan du byta ut kortet mot ett finländskt körkort.
Om du har ett körkort som utfärdats i ett land som är anslutet till Genève- eller Wien-konventionerna kan du köra med detta kort högst två år i Finland.
Du måste byta ut ditt körkort mot ett finländskt körkort inom två år efter att du flyttat till Finland.
Om du har ett körkort som utfärdats i ett land som inte är anslutet till Genève- eller Wien-konventionerna kan du köra bil med detta kort under ett års tid efter att ha registrerats i befolkningsregistret i Finland.
Du kan byta ut ditt körkort till ett finskt körkort på Ajovarmas serviceställe.
linkkiTrafiksäkerhetsverket:
Utländskt körkort i Finlandfinska _ svenska _ engelska
Internet
I Finland kan du sköta många ärenden via Internet.
Det är bra att skaffa sig en Internetuppkoppling så fort som möjligt efter att du har flyttat till Finland.
På InfoFinlands sida Vardagslivet i Finland finns mer information om att skaffa en internetuppkoppling.
linkkiKommunikationsverket:
Internet- och telefonabonnemangfinska _ svenska _ engelska
Telefon
När du köper ett telefonabonnemang i Finland får du ett finskt telefonnummer.
Många företag erbjuder telefonabonnemang.
Du kan också köpa ett prepaid-abonnemang.
Prepaid-kortet är i förväg laddat med en summa som man sedan kan ringa för.
Prepaid-abonnemang kan köpas till exempel i R-kiosker, en del snabbköp och på Internet.
linkkiSkype:
Förmånliga utlandssamtalfinska _ svenska _ engelska _ ryska _ estniska _ franska _ spanska _ turkiska _ kinesiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ ungerska _ japanska
Hälsa
I Finland finns offentliga och privata hälsovårdstjänster.
Du kan använda de offentliga hälsovårdstjänsterna om du har en hemkommun i Finland.
Till de offentliga hälsovårdstjänsterna hör till exempel hälsocentralerna.
De offentliga tjänsterna är förmånligare än de privata.
Om du vill reservera tid till en läkare ska du ta kontakt med hälsocentralen.
Om du inte har rätt att använda de offentliga hälsovårdstjänsterna kan du kontakta en privat läkarcentral.
Mer information om hälsovården i Finland får du på InfoFinlands sida Hälsa.
Språkstudier
Finlands officiella språk är finska och svenska.
Språkkunskaper hjälper dig att förstå det nya samhället och underlättar skötseln av ärenden.
Mer information hittar du på InfoFinlands sida Finska och svenska språket.
Jobbsökning
Arbets- och näringsbyrån hjälper dig i jobbsökningen.
Du kan söka jobb på Internet och via tidningar.
Du kan också hitta ett jobb genom att själv kontakta arbetsgivare som du är intresserad av.
Läs mer om jobbsökning i Finland på InfoFinlands sida Var hittar jag jobb?
Fritid och hobbyer
Information om möjligheter till fritidsaktiviteter hittar du på InfoFinlands sida Fritid.
linkkiExpat Finland:
Information om Finland för utlänningarengelska
Du kan få permanent uppehållstillstånd (pysyvä oleskelulupa) (P), om
du bott i Finland i minst fyra år med A-tillstånd och
inte under tiden har bott utomlands i över två år och
grunden för de tidigare uppehållstillstånden fortfarande existerar
Om du hade A-tillstånd då du kom till Finland beräknas de fyra åren från den dag du anlände till Finland Om du fått A-tillstånd i Finland beräknas de fyra åren från den dag då det första A-tillståndet trädde i kraft.
Om du har fått internationellt skydd i Finland beräknas de fyra åren från att du anlände till Finland.
Permanent uppehållstillstånd kan eventuellt inte beviljas om:
du har begått ett brott som är belagt med fängelsestraff
du är misstänkt för ett brott som är belagt med fängelsestraff
du har begått två eller flera brott
du misstänks för två eller flera brott
Permanen uppehållstillstånd gäller tills vidare.
Tillstånet kan dras tillbaka om du permanent flyttar från Finland, uppehåller dig utomlands kontinuerligt i minst två år eller har lämnar felaktiga uppgifter då du ansökt om tillståndet.
EU-uppehållstillstånd för tredjelandsmedborgare som uppehållit sig länge i landet
Tredjelandsmedborgare äe medborgare i annat land än de nordiska länderna, EU-länderna, Liechtenstein eller Schweiz.
Du kan beviljas EU-uppehållstillstånd (P-EU) för tredjelandsmedborgare om:
du har bott i Finland i minst fem år med A-tillstånd och
inte under denna tid har bott utomlands längre än 10 månader och
grunden för de tidigare uppehållstillstånden fortfarande existerar
P-EU-tillstånd ansöks om på samma sätt som permanent uppehållstillstånd.
P-EU-tillstånd gäller tills vidare.
P-EU-tillståndsansökan kan även avslås på samma grunder som permanent uppehållstillstånd.
Ansökan
Du kan ansöka om permanent uppehållstillstånd på internet i tjänsten Enter Finland.
När du ställt ansökan ska du besöka Migrationsverkets tjänsteställe för att styrka din identitet.
Ta med dig en identitetshandling och originalexemplaren av ansökningsbilagorna.
Det är bra att boka en tid hos Migrationsverkets tjänsteställe i förväg.
Du kan boka tiden via Migrationsverkets elektroniska tidsbokningssystem.
Om du gjort ansökningen på internet, kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan, kommer detta att meddelas via ditt Enter Finland-konto.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du ansöka om tillståndet med en pappersblankett vid Migrationsverkets tjänsteställe.
Du kan skriva ut blanketten på Migrationsverkets webbplats.
Boka en tid vid tjänstestället och ta med dig den ifyllda ansökningen, bilagorna och en identitetshandling.
Handläggning av ansökan är avgiftsbelagd.
Avgiften ska betalas då ansökan ställs.
I tjänsten Enter Finland kan du betala med nätbankskoderna för en finsk bank eller med kreditkort.
Permanent uppehållstillståndfinska _ svenska _ engelska
Ansökningsblankettfinska _ svenska _ engelska
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Om du är av finländsk härkomst eller har en nära kontakt med Finland kan du beviljas uppehållstillstånd i Finland på grund av detta.
Då är du återflyttare (paluumuuttaja).
Huruvida du beviljas uppehållstillstånd beror på hur starka och nära släktband du har till Finland.
För att få tillståndet krävs inga andra skäl, som till exempel arbete eller studier.
Personer som aldrig själv har varit finska medborgare men vars ena förälder eller mor- eller farförälder är eller har varit infödd finsk medborgare betraktas som återflyttare (paluumuuttaja) av finsk härkomst.
Också före detta finska medborgare räknas som återflyttare.
Uppehållstillstånd för återflyttarefinska _ svenska _ engelska
Avkomlingar till infödda finska medborgare
Du kan beviljas uppehållstillstånd i Finland om minst en av dina föräldrar eller mor- eller farföräldrar är eller har varit infödd finsk medborgare.
Med infödd finsk medborgare avses en person som har fått finskt medborgarskap vid födseln.
När du ansöker om tillstånd måste du ge en tillförlitlig bild av din härkomst, som till exempel uppvisa den ursprungliga födelseattesten av en förälder eller en mor- eller farförälder samt ett intyg över ert släktskap.
Du krävs inte på redogörelse över din utkomst.
Före detta finska medborgare
Om du är en före detta finsk medborgare kan du på denna grund få uppehållstillstånd i Finland.
Förutsättningen är inte att du är en infödd finsk medborgare, utan du kan också ha fått det finska medborgarskapet på ansökan.
Du krävs inte på redogörelse över din utkomst.
Om du är en före detta finsk medborgare kan du återfå ditt finska medborgarskap genom att göra en medborgarskapsanmälan (kansalaisuusilmoitus).
Läs mer på InfoFinlands sida Finskt medborgarskap.
Ansökan om uppehållstillstånd
Du kan ansöka om uppehållstillstånd antingen utomlands innan du kommer till Finland eller i Finland.
Utomlands kan du ansöka om tillstånd vid den närmaste av Finlands ambassader, i Finland vid Migrationsverkets tjänsteställe.
Du måste personligen gå och lämna in ansökan om uppehållstillstånd.
Ta med dig originalexemplaren av de bilagor som krävs för ansökan när du lämnar in din ansökan vid ambassaden eller Migrationsverkets tjänsteställe.
När du ansöker om uppehållstillstånd måste du ha med dig ett pass för att kunna styrka din identitet.
När du ansöker om tillstånd tas dina fingeravtryck för det biometriska uppehållstillståndskortet.
Ansökan om uppehållstillstånd är avgiftsbelagd.
Avgiften måste betalas i samband med att man lämnar in sin tillståndsansökan.
Finsk personbeteckning
Om du får ett uppehållstillstånd i Finland registreras du automatiskt i det finska befolkningsdatasystemet.
Du får samtidigt även en finsk personbeteckning.
När du har flyttat till Finland ska du besöka magistraten på din hemort för att registrera dig som invånare.
Läs mer på InfoFinlands sida Registrering som invånare.
Uppehållstillstånd för avkomlingar till infödda finländarefinska _ svenska _ engelska
Uppehållstillstånd för före detta finska medborgarefinska _ svenska _ engelska
linkkiFinland-Samfundet:
Utlandsfinländarnas intresseorganisationfinska _ svenska _ engelska
Kommunerna tillhandahåller många tjänster för sina invånare.
Till kommunens tjänster hör till exempel hälsovård och barndagvård.
Om du har en hemkommun (kotikunta) i Finland, har du vanligen rätt att använda dig av den kommunens tjänster.
Det lönar sig för dig att utreda om du och de andra medlemmarna i din familj har rätt till en hemkommun i Finland.
Rätten till en hemkommun i Finland bestäms enligt hemkommunslagen.
Vid magistraten (maistraatti) på din egen boningsort kan du ta reda på om du har rätt till en hemkommun i Finland.
Hur kan du få en hemkommun i Finland
För att du ska kunna få en hemkommun i Finland måste du flytta till och vara stadigvarande bosatt i Finland.
Om du bor i Finland tillfälligt, till exempel om du flyttar till Finland för studier eller jobb under högst ett år, kan du vanligen inte få en hemkommun i Finland.
Du har möjlighet att få en hemkommun i Finland om:
du är finsk medborgare
du är medborgare i ett nordiskt land
du är medborgare i EU, Schweiz eller Liechtenstein och du har registrerat din uppehållsrätt i Finland
du har permanent (P) eller kontinuerligt (A) uppehållstillstånd som är i kraft
du är familjemedlem till en person som har en hemkommun i Finland
Om du har ett tillfälligt uppehållstillstånd (B-tillstånd) som är i kraft kan du få en hemkommun om du kan påvisa att det är din avsikt att bo stadigvarande i Finland.
Stadigvarande boende kan påvisas till exempel genom följande omständigheter:
du har en arbetsplats i Finland och ditt arbetskontrakt är i kraft minst två år
du studerar i Finland och dina studier räcker minst två år
du är av finländsk härkomst
du har tidigare haft en hemkommun i Finland
du har varit fortlöpande bosatt i Finland under minst ett års tid.
Din hemkommun är vanligen den kommun du bor i.
Om du inte har en bostad eller om du har bostäder på flera kommuners område är din hemkommun den kommun som du själv uppfattar som din hemkommun och som du har någon fast förbindelse till, till exempel genom familjeförhållanden eller arbetsplats.
Kontaktuppgifter till magistratfinska _ svenska _ engelska
Lag om hemkommunfinska _ svenska
Om du har ett tillfälligt uppehållstillstånd (A- eller B-tillstånd) och orsaken för din vistelse i Finland ändras måste du ansöka om ett nytt uppehållstillstånd på den nya grunden.
Om du har ett permanent uppehållstillstånd (P) i Finland behöver du inte ändra grunden för ditt uppehållstillstånd även om orsaken till din vistelse ändras.
Du kan ansöka om uppehållstillstånd på något av följande grunder:
arbete
studier
familjeband
återflyttning
finländsk härkomst
internationellt skydd
annan orsak
Det är bra att komma ihåg att grunden för uppehållstillståndet kan påverka vilka rättigheter du har i Finland.
Till exempel ger ett uppehållstillstånd på grund av familjeband mer omfattande rätt att arbeta än ett tillstånd som beviljats på grund av studier.
Hur får jag ett tillfälligt uppehållstillstånd ändrat till ett kontinuerligt tillstånd?
Om du har ett tillfälligt uppehållstillstånd (B-tillstånd) kan du ansöka om ett kontinuerligt uppehållstillstånd (A-tillstånd) om grunden för vistelsen i Finland har ändrats från tillfällig till kontinuerlig.
Om du har ett tillfälligt uppehållstillstånd på grund av familjeband kan du ansöka om ett kontinuerligt uppehållstillstånd när en familjemedlem till dig ansöker om ett kontinuerligt uppehållstillstånd.
Du kan ansöka om ett kontinuerligt uppehållstillstånd också på någon annan grund om grunden är kontinuerlig.
Om du har ett tillfälligt uppehållstillstånd på grund av studier kan du få ett kontinuerligt tillstånd endast i det fall att grunden för din vistelse i Finland ändras.
Du kan inte få ett kontinuerligt tillstånd på basis av studier.
Grunden för din vistelse kan ändras till exempel om du får en arbetsplats i Finland eller gifter dig med en finsk medborgare eller en person som har kontinuerligt eller fortsatt tillstånd i Finland.
Om du har ett tillfälligt uppehållstillstånd för arbete eller näringsidkande kan du ansöka om ett kontinuerligt uppehållstillstånd när du har vistats i Finland två år utan avbrott.
Hur söker jag ett uppehållstillstånd på nya grunder?
Välj ansökningsblankett utifrån grunden för din ansökan om nytt tillstånd.
Lämna in din ansökan på internet i tjänsten Enter Finland eller vid Migrationsverkets tjänsteställe.
Mer information om ansökningsproceduren hittar du på InfoFinlands sida Fortsatt uppehållstillstånd.
Från studerande till anställd
Om du har avlagt en examen i Finland kan du få ett uppehållstillstånd för att söka arbete.
När du är klar med dina studier och ditt uppehållstillstånd för studerande går ut, kan du ansöka om fortsatt tillstånd (jatkolupa) för att söka arbete.
Tillståndet är i kraft ett år.
Detta tillstånd kan endast fås en gång och det kan inte förnyas.
När du får en arbetsplats kan du få uppehållstillstånd på grund av arbete.
Uppehållstillstånd på en ny grundfinska _ svenska _ engelska
Uppehållstillstånd för sökande av arbetefinska _ svenska _ engelska
På denna sida finns information riktad till kvotflyktingar.
Information om att ansöka om asyl hittar du på InfoFinlands sida Till Finland som asylsökande.
Kvotflyktingar
Man kan inte ansöka om att bli kvotflykting via myndigheterna i Finland.
Man kan inte heller föreslå en annan person, till exempel en släkting eller vän, som kvotflykting.
Finland tar som kvotflyktingar emot personer som har flyktingstatus enligt
Förenta nationernas flyktingorganisation UNHCR.
Intervjuerna görs i de länder där flyktingarna vistas, vanligen i flyktingläger eller i UNHCR:s lokaler.
Information om val av kvotflyktingarfinska _ svenska _ engelska
Flytta till Finland
På webbsidan Movingtofinland.fi finns mycket information avsedd för kvotflyktingar om att flytta till Finland och om livet i Finland.
Information för flyktingarfinska _ engelska _ franska _ persiska _ arabiska _ kurdiska
Stöd till flyktingar
Finlands röda kors (FRK) hjälper kvotflyktingar när de flyttar till Finland.
När flyktingarna anländer till Finland kommer en anställd från röda korset till flygplatsen och tar emot dem.
Röda korsets frivilligarbetare hjälper även flyktingar att bosätta sig och integreras i Finland.
Flyktingar kan be om hjälp och rådgivning i rättsliga frågor bland annat från flyktingrådgivningen r.f. eller från rättshjälpsbyråer.
Finlands flyktinghjälp r.f. är en organisation som strävar efter att främja de grundläggande rättigheterna för flyktingar.
Organisationen utför informations-, utbildnings och socialarbete i Finland.
Flyktinghjälpen hjälper flyktingar och invandrare till exempel med ärenden som gäller integrering, boende och grundande av egna organisationer.
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ engelska
linkkiFinlands flyktinghjälp r.f.:
Stöd till flyktingarfinska _ svenska _ engelska
linkkiFinlands röda kors:
Stöd till flyktingarfinska _ svenska _ engelska
Rehabiliteringscentret för tortyrofferfinska _ engelska
Som flykting i Finland
På InfoFinlands sida Flykting hittar du mer information avsedd för flyktingar.
När du har flyttat till Finland, måste du besöka magistraten (maistraatti) på din hemort.
Innan du besöker magistraten kan du fylla i en registreringsanmälan som du kan ladda ned på adressen maistraatti.fi.
Du kan även fylla i anmälan i magistraten.
På magistraten kan du, under förutsättning att villkoren för detta uppfylls, även få en finsk personbeteckning, om du inte redan fick en sådan då du beviljades uppehållstillstånd eller din uppehållsrätt för EU-medborgare registrerades.
Om du behöver en personbeteckning för arbete, kan du få en personbeteckning även på skattebyrån.
På magistraten utreder man om det är möjligt att registrera en hemkommun (kotikunta)för dig.
När du går till magistraten ska du ta med dig åtminstone följande handlingar:
pass eller
annat identitetsbevis där ditt medborgarskap framgår (om du är medborgare i ett EU-land eller ett nordiskt land)
legaliserat äktenskapsintyg (om du är gift)
legaliserade födelseattester för barnen (om du har barn under 18 år)
uppehållstillstånd (om du behöver ett uppehållstillstånd i Finland)
Registreringsintyg över uppehållsrätt för EU-medborgare (om du är EU-medborgare och din uppehållsrätt måste registreras)
arbetskontrakt eller intyg om studier (om din uppehållsrätt som EU-medborgare inte har registrerats)
Notera att utländska handlingar måste vara legaliserade för att man utgående från dem ska kunna föra in personuppgifter i befolkningsdatasystemet.
Du måste även låta översätta handlingarna till finska, svenska eller engelska om de är på något annat språk.
Om du behöver mer information om legalisering av handlingar, kontakta magistraten eller utrikesministeriet i ditt hemland.
Registrering av utlänningarfinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Registrering av utlänningar på skattebyrånfinska _ svenska _ engelska
Finsk personbeteckning
Personbeteckningen (henkilötunnus) är en 11 tecken lång sifferserie som bildas på basis av ditt födelsedatum och ditt kön.
Du behöver en personbeteckning till för din arbetsgivare eller läroanstalt.
Det underlättar även skötandet av många officiella ärenden.
För att du ska kunna få en finsk personbeteckning måste dina uppgifter registreras i Finlands befolkningsdatasystem.
Det innebär att grundinformation om dig förs in i befolkningsdatasystemet.
Dessa uppgifter är till exempel namn, födelsedatum, nationalitet, kön och adress.
När du ansöker om uppehållstillstånd, kan du samtidigt även ansöka om en finsk personbeteckning.
Då måste du i din ansökan be om att din information registreras i Finlands befolkningsdatasystem.
Om du är EU-medborgare kan du ansöka om personbeteckning samtidigt som du ansöker om registrering av uppehållsrätt.
I registreringsblanketten finns en punkt där du kan be om att dina uppgifter registreras i befolkningsdatasystemet.
Läs mer på InfoFinlands sida Hemkommun i Finland.
Det är viktigt att du ansöker om fortsatt uppehållstillstånd innan ditt tidigare uppehållstillstånd går ut.
Om ditt tidigare uppehållstillstånd går ut under behandlingen av ansökan får du uppehålla dig i Finland och har vanligtvis även rätt att arbeta under den tid som ansökan behandlas.
Om du ansöker om fortsatt uppehållstillstånd först efter att ditt tidigare uppehållstillstånd gått ut, får du uppehålla dig i Finland under tiden då ansökan behandlas men har inte rätt att arbeta innan du erhållit fortsatt uppehållstillstånd.
Att ansöka
Du kan ansöka om tillståndet på internet i tjänsten Enter Finland.
När du ställt ansökan ska du besöka Migrationsverkets tjänsteställe för att styrka din identitet.
Du ska besöka tjänstestället inom tre månader efter att ha gjort ansökan.
Ta med dig pass, passfoto och originalexemplaren av ansökningsbilagorna.
Det är bra att boka en tid hos Migrationsverkets tjänsteställe i förväg.
Du kan boka tiden via Migrationsverkets elektroniska tidsbokningssystem.
Om du gjort ansökningen på internet, kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan, kommer detta att meddelas via ditt Enter Finland-konto.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du ansöka om tillståndet med en pappersblankett vid Migrationsverkets tjänsteställe.
Skriv ut blanketten på Migrationsverkets webbplats och fyll i den färdigt.
Boka en tid vid tjänstestället.
När du ska besöka tjänstestället, ta med dig din ifyllda ansökan, bilagorna och kopior på bilagor samt pass och passfoto.
Migrationsverket beviljar dig fortsatt uppehållstillstånd om grunden för det tidigare uppehållstillståndet fortfarande existerar.
Du kan även ansöka om fortsatt uppehållstillstånd på annan grund än för det tidigare tillståndet
Hanteringen av ansökan är avgiftsbelagd. Avgiften ska betalas då ansökan görs.
I tjänsten Enter Finland kan du betala med nätbankskoderna för en finsk bank eller med kreditkort.
Att förlänga uppehållstillståndetfinska _ svenska _ engelska
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Blanketter för ansökan om uppehållstillståndfinska _ svenska _ engelska
Migrationsverket:
Presentation av e-tjänsten Enter Finland
Söka asyl
Asylsökande från Europeiska unionens område
Minderåriga asylsökande
Handläggning av asylansökan
Asylsamtal
Positivt beslut
Negativt beslut
Rättshjälp för asylsökande
Asylsökandes rätt att arbeta
Du kan söka asyl i Finland om du har välgrundad fruktan för förföljelse i ditt hemland.
Orsaker till förföljelse kan vara etniskt ursprung, religion, medborgarskap, tillhörighet till en viss grupp i samhället eller politiska åsikter.
Migrationsverket utreder om det finns asylskäl och fattar ett beslut.
Du kan endast söka asyl för dig själv.
Broschyren Information till asylsökandefinska _ svenska _ engelska _ ryska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
Söka asyl
Du kan endast söka asyl i Finland på det finska territoriet.
Det finns ingen särskild asylansökningsblankett som du skulle kunna fylla i förväg.
När du kommer till Finland, meddela gränskontrollmyndigheten eller polisen genast att du vill söka asyl.
Gränskontrollmyndigheten eller polisen registrerar dig som asylsökande, antecknar uppgifter om dig och tar dina fingeravtryck.
När myndigheten har mottagit din asylansökan, hänvisas du till ett mottagningscenter.
Där kan du bo under tiden då Migrationsverket behandlar din ansökan.
Du kan även bo någon annanstans, men då måste du själv bekosta boendet.
Att söka asyl i Finlandfinska _ svenska _ engelska
Asylsökande från Europeiska unionens område
Inom EU (och i Schweiz, Norge, Island och Liechtenstein) måste man söka asyl i det land, till vars territorium man kommer först.
Om du har sökt asyl eller vistats i något annat EU-land (eller i Schweiz, Norge, Island eller Liechtenstein) innan du kom till Finland, behandlas din ansökan inte i Finland.
I detta fall avvisas du tillbaka till det land där du var innan du kom till Finland.
Detta kallas för Dublinprocessen.
Om du är medborgare i ett EU-land, får du sannolikt inte asyl i Finland.
Finland anser att alla EU-länder är trygga för medborgarna.
Likväl utreds alla ansökningar som EU-medborgare skickar in.
På InfoFinlands sida EU-medborgare hittar du information om flytt till Finland av andra skäl än som asylsökande.
Att lämna asylansökan utan prövningfinska _ svenska _ engelska
Minderåriga asylsökande
Om du är under 18 år gammal och kommer till Finland som asylsökande utan vårdnadshavare, förordnas du ett ombud.
Ombudet är en pålitlig vuxen person som hjälper dig med olika ärenden under tiden då Migrationsverket behandlar din ansökan.
Ombudet följer med dig när du ska prata med myndigheter.
Dessutom utreder ditt ombud om du kan återförenas med din familj.
Du har rätt till boende, mat och hälsovård.
Du har även rätt att gå i skola.
Ensamkommande barn(pdf, 674)finska _ svenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ persiska _ arabiska _ kurdiska
Handläggning av asylansökan
Migrationsverket handlägger din ansökan och fattar ett beslut.
Migrationsverket utreder din identitet och resväg till Finland och bedömer om du kan beviljas asyl i Finland.
Det är vanligt att behandlingen av ansökan tar flera månader.
När du har sökt asyl har du rätt att vistas i Finland medan din ansökan behandlas.
Under denna tid kan du inte resa utomlands.
Om du reser kan myndigheterna besluta att din ansökan inte längre gäller.
Migrationsverket skickar dig en kallelse till asylsamtal.
I kallelsen anges tolkningsspråket, den exakta adressen till verksamhetsstället där samtalet hålls och klockslaget.
Handläggning av asylansökanfinska _ svenska _ engelska
Asylsamtal
Asylsamtalet (turvapaikkapuhuttelu) är den viktigaste händelsen under behandlingen av din ansökan.
Under samtalet ställs frågor om de händelser och orsaker som tvingade dig att lämna ditt hemland.
Det är viktigt att du beskriver allt som hänt så exakt som möjligt.
Migrationsverket beslutar baserat på din berättelse om du beviljas asyl i Finland.
Som asylsökande har du rätt att använda ett rättsbiträde under samtalet.
Biträdet deltar i asylsamtalet efter sitt eget omdöme.
Om du behöver en tolk, skaffar Migrationsverket tolken.
Positivt beslut
Du får stanna i Finland om du beviljas asyl eller uppehållstillstånd på andra grunder.
Du kan beviljas asyl i Finland om myndigheterna anser att du blir förföljd i ditt hemland på grund av
etniskt ursprung,
religion,
medborgarskap,
tillhörighet till en viss grupp i samhället eller
politiska åsikter.
Om du inte får asyl kan du i vissa fall beviljas uppehållstillstånd på grund av alternativt skydd.
Du kan beviljas uppehållstillstånd på grund av alternativt skydd om du hotas av:
dödsstraff eller avrättning,
tortyr eller någon annan behandling eller bestraffning som är omänsklig eller kränker människovärdet eller
om du utsätts för allvarlig personlig fara på grund av en väpnad konflikt.
När du söker asyl utreder Migrationsverket samtidigt om du kan få uppehållstillstånd på någon annan grund.
Asylfinska _ svenska _ engelska
Negativt beslut
Om du inte beviljas asyl eller uppehållstillstånd på någon annan grund blir du avvisad från Finland.
Du har även möjlighet att överklaga ett negativt beslut till förvaltningsdomstolen.
Bifogat till beslutet finns en anvisning om hur du överklagar.
På InfoFinlands sida Negativt beslut om uppehållstillstånd hittar du information om vad du kan göra om du får ett negativt beslut.
Ändringssökande i asylbeslutfinska _ svenska _ engelska
Avvisning av en asylsökandefinska _ svenska _ engelska
Rättshjälp för asylsökande
Under tiden då din ansökan behandlas kan du få rådgivning och rättshjälp vid den offentliga rättshjälpsbyrån.
Kontakta rättshjälpsbyrån om du vill ha ett rättsbiträde.
Vid behov hjälper mottagningscentret dig.
Rättshjälpsbyrån (oikeusaputoimisto) kan även hänvisa dig till en privat jurist eller en privat juristbyrå.
Du kan även få rådgivning hos Flyktingrådgivningen rf (Pakolaisneuvonta ry).
Flyktingrådgivningen ger rådgivning även till personer som vistas i Finland utan uppehållstillstånd.
linkkiRättsväsendet:
Rättshjälpsbyråerfinska _ svenska _ engelska
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Asylsökandes rätt att arbeta
Du får förvärvsarbeta i Finland om det har gått tre månader sedan du lämnade in din asylansökan och du har ett giltigt pass eller någon annan resehandling som du har företett till myndigheten när du sökte asyl.
Om du inte företedde en giltig resehandling till myndigheten i samband med din asylansökan får du förvärvsarbeta i Finland när det har gått sex månader sedan du lämnade in din asylansökan.
Du har rätt att arbeta tills du har fått ett lagakraftvunnet beslut på din asylansökan.
Om Migrationsverket ger dig ett positivt beslut på din asylansökan, får du uppehållstillstånd.
I det ingår nästan alltid rätt att arbeta.
Om Migrationsverket fattar ett negativt beslut på din asylansökan, har du rätt att arbeta under tiden då en eventuell överklagan behandlas.
För att arbeta måste du ha ett finländskt skattekort.
Hämta ett skattekort på den närmaste skattebyrån och lämna kortet till din arbetsgivare.
Läs mer på InfoFinlands sida Skattekort.
Om du arbetar permanent kan du även ansöka om uppehållstillstånd i Finland på grund av arbete.
På InfoFinlands sida Arbeta i Finland hittar du mer information om uppehållstillstånd för arbetstagare.
Asylsökandes rätt att arbetafinska _ svenska _ engelska
Uppehållstillstånd på andra grunderfinska _ svenska _ engelska
Om du är medborgare i något nordiskt land behöver du inte uppehållstillstånd i Finland.
Du har rätt att jobba, fungera som företagare och studera i Finland.
När du flyttar till Finland måste du göra en flyttanmälan och gå och registrera dig vid magistraten (maistraatti) på din egen hemort.
Notera att du måste besöka magistraten personligen.
Gör flyttanmälan senast inom en vecka från din flyttningsdag.
För registreringen behöver du ett officiellt identitetskort där ditt medborgarskap framgår eller pass som är i kraft.
Familjemedlemmar till nordiska medborgare
Om en av dina familjemedlemmar, som flyttar med dig till Finland, inte är medborgare i ett nordiskt land, kan han/hon behöva uppehållstillstånd eller ett registreringsintyg över uppehållsrätt för EU-medborgare.
Läs mer på InfoFinlands sidor EU-medborgare eller Icke-EU-medborgare.
Finsk personbeteckning
När du registrerar dig vid magistraten kan du på samma gång få en finsk personbeteckning (henkilötunnus).
Du behöver en personbeteckning när du sköter ärenden hos myndigheter, och dessutom underlättar den skötandet av ärenden i till exempel banker och med din arbetsgivare.
Läs mer på InfoFinlands sidor Registrering som invånare.
Registrering av utlänningarfinska _ svenska _ engelska
Information för nordiska medborgarefinska _ svenska _ engelska _ norska
_ danska
_ isländska
Rådgivningstjänst för nordiska medborgarefinska _ engelska _ norska
_ danska
_ isländska
Information om den sociala tryggheten i de nordiska ländernafinska _ svenska _ engelska _ norska
Finland tillhör Schengenområdet.
Länderna som tillhör Schengenområdet har enhetlig visering.
Utlänningar som vill resa till Finland för en kort tid, till exempel på semester, affärsresa eller på besök hos släktingar, behöver ett visum om de inte är medborgare i ett viseringsfritt land.
Ett visum är ett inresetillstånd för en kortvarig och tillfällig, högst tre månader lång vistelse.
På utrikesministeriets webbplats eller vid den närmast belägna finländska beskickningen kan du kontrollera om du behöver ett visum i Schengenområdet.
Visumbehovet till Schengenområdet och av
Finland accepterade resedokumentfinska _ svenska _ engelska
Information för viseringsfria personer
Du kan resa till Finland och de övriga Schengenländerna om du har ett giltigt pass eller något annat resedokument som godkänns i Finland.
Du får vistas högst tre månader under en period på sex månader i Finland och de övriga Schengenländerna räknat från den dag du reste in till Schengenområdet.
Information för viseringsskyldiga personer
Du ska alltid ha ett visum när du kommer till Finland eller något annat land i Schengenområdet.
Du får vistas i Finland eller något annat land i Schengenområdet utan uppehållstillstånd så länge som ditt visum är i kraft.
Om du har ett visum eller uppehållstillstånd i något Schengenland kan du resa inom Schengenområdet utan att behöva skaffa ett separat visum för de andra Schengenländerna.
Så här ansöker du om Schengenvisum
Du ansöker om visum i den närmast belägna finländska beskickningen eller visumcentralen.
Du ska vistas lagligt i det land där du ansöker om visum. I länder där
Finland inte har en beskickning kan något annat land representera Finland i visumärenden.
I detta fall kan du ansöka om visum i detta lands beskickning.
På utrikesministeriets webbplats finns en förteckning över de länder där ett annat land representerar Finland i visumärenden.
Du ansöker om visum med en visumansökningsblankett.
Blanketten får du på utrikesministeriets webbplats och från beskickningar i Schengenländer.
Antalet bilagor som krävs till visumansökan kan variera beroende på i vilket land du söker visum.
Hos beskickningen kan du kontrollera vilka bilagor du behöver för din visumansökan.
Lämna din ansökning till den beskickning eller visumcentral dit du ställer din ansökan.
Du kan inte skicka din ansökning via e-post eller fax.
Förlängning av visum i Finland
Polisen kan förlänga uppehållstiden för ditt visum eller visumets utgångstid om du av motiverade skäl inte kan lämna Finland när ditt visum utgår.
Motiverade skäl för förlängning av visum kan till exempel vara:
en akut, svår sjukdom som hindrar dig från att resa,
en släkting som är bosatt i Finland har plötsligt insjuknat svårt eller avlidit,
inställt flyg på grund av strejk eller väderförhållanden,
viktiga affärsförhandlingar som pågår längre än väntat.
Information till medborgare från viseringsskyldiga länderfinska _ svenska _ engelska
Ansökan om Schengenvisumfinska _ svenska _ engelska
Länder där en annan Schengenstat representerar Finlandfinska _ svenska _ engelska
Förlängning av visum i Finlandfinska _ svenska _ engelska
Hjälp i nödsituationer
Beskickningarna hjälper sitt lands medborgare som hamnat i nödläge i Finland.
De kan till exempel hjälpa dig om du har råkat ut för en olycka, blivit sjuk eller fallit offer för ett brott.
Beskickningen kan bevilja dig ett nytt pass om ditt pass har gått förlorat eller stulits.
Om du är turist i Finland och hamnar i en svår situation, ska du kontakta ditt hemlands beskickning.
linkkiVisitFinland.com:
Information om Finland till turistersvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ japanska _ italienska
Också andra anhöriga till finska medborgare än en make/maka, en sambo, föräldrar till minderåriga barn eller minderåriga barn kan i vissa fall få uppehållstillstånd i Finland på grund av familjeband.
Även andra anhöriga till en person som har ett uppehållstillstånd på grund av internationellt skydd kan beviljas uppehållstillstånd.
Om uppehållstillståndet beviljats på någon annan grund än internationellt skydd, kan andra anhöriga inte få uppehållstillstånd.
En annan anhörig kan få uppehållstillstånd om han eller hon är helt beroende av den anhöriga som bor i Finland.
På denna grund kan uppehållstillstånd beviljas till exempel för en förälder till en myndig (18 år gammal) person.
Enbart ekonomiskt beroende eller svag hälsa räcker ändå inte för att beviljas uppehållstillstånd.
En annan anhörig kan få uppehållstillstånd också om han eller hon levt tillsammans som en familjemedlem till den anhöriga som är bosatt i Finland, innan denna person kom till Finland.
Dessutom krävs det att familjelivet upphört på grund av ett tvingande skäl, till exempel för att man blivit flyktingar.
Annan anhörig till en finsk medborgarefinska _ svenska _ engelska
Annan anhörig till en person som fått internationellt skyddfinska _ svenska _ engelska
Att ansöka om uppehållstillstånd
Vanligtvis måste du ansöka om ditt första uppehållstillstånd innan du kommer till Finland.
Ansök om tillståndet i ditt hemland eller i ett annat land där du vistas lagligt.
Du kan ansöka om tillståndet på internet via tjänsten Enter Finland.
När du ställt ansökan ska du besöka Finlands beskickning närmast dig eller Migrationsverkets tjänsteställe för att styrka din identitet och visa upp originalexemplaren av ansökningsbilagorna.
Du ska besöka beskickningen eller tjänstestället inom tre månader efter att ha gjort ansökan på internet.
Ansökningen kan tas för behandling först när du besökt beskickningen eller tjänstestället.
Vanligtvis måste du boka en tid hos beskickningen eller tjänstestället i förväg.
Kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan, kommer detta att meddelas via ditt Enter Finland-konto.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du också lämna in en pappersansökan jämte bilagor vid Finlands beskickning närmast dig eller på Migrationsverkets tjänsteställe i Finland.
Du kan skriva ut ansökningsblanketten på Migrationsverkets webbplats.
Ansökan om uppehållstillstånd är avgiftsbelagd.
Avgiften ska betalas då ansökan ställs.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Finlands beskickningar utomlandsfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Finsk personbeteckning
Om du får ett uppehållstillstånd i Finland registreras du automatiskt i det finska befolkningsdatasystemet.
Du får samtidigt även en finsk personbeteckning.
När du har flyttat till Finland ska du besöka magistraten på din hemort för att registrera dig som invånare.
Läs mer på InfoFinlands sida Registrering som invånare.
Om du behöver visum eller uppehållstillstånd för att vistas i Finland, men inte har det, vistas du illegalt i Finland.
Asylsökande har rätt att uppehålla dig i Finland även utan visum eller uppehållstillstånd under den tid som det tar att handlägga asylansökan.
Även om du har kommit lagligt till Finland kan din vistelse i landet bli illegal till exempel om du stannar kvar i landet fastän du inte beviljas ett uppehållstillstånd eller om ditt visum eller uppehållstillstånd har gått ut.
Information om hur du kan få ett uppehållstillstånd i Finland finns på InfoFinlands sida Flytta till Finland.
Hjälp och rådgivning
Mathjälp och inkvartering
Du har rätt till nödinkvartering och mathjälp om du inte har pengar till mat eller någonstans att övernatta.
Kommuner, församlingar och vissa organisationer ordnar nödinkvartering.
Juridisk rådgivning
Flyktingrådgivningen r.f. ger kostnadsfri juridisk rådgivning för papperslösa invandrare.
Rådgivningen betjänar telefonledes på numret 045-237 7104 (måndagar kl. 14–16).
Rådgivningen ges av en jurist.
Fler kontaktuppgifter hittar du på Flyktingrådgivningens webbplats.
Sjukvård
Om du blir sjuk eller skadas, har du rätt till brådskande vård inom den offentliga hälso- och sjukvården, till exempel på en hälsostation eller ett sjukhus.
Du måste i regel själv betala kostnaderna för vården.
I Helsingfors, Åbo, Tammerfors och Esbo får barn och gravida kvinnor samma hälso- och sjukvårdstjänster som övriga invånare.
De måste betala samma avgifter för vården som övriga invånare.
Global Clinic är en klinik där du kan få hjälp eller råd av en läkare eller sjukskötare om du vistas i Finland utan uppehållstillstånd.
Du kan besöka Global Clinic även om du inte behöver brådskande sjukvård.
Global Clinic bedriver verksamhet i följande städer:
Åbo
Tammerfors
Uleåborg
Joensuu
Du kan ringa eller skicka e-post.
En sjukskötare eller läkare besvarar ditt samtal.
Du hittar kontaktinformation på Global Clinic:s hemsidor.
Global Clinic:s tjänster är avgiftsfria för kunderna.
Global Clinic anmäler inte sina kunder till polisen eller andra myndigheter.
Klinikens adress eller öppettider meddelas inte offentligt.
linkkiFlyktingrådgivningen rf:
Juridisk rådgivningfinska _ engelska _ franska _ arabiska
Kontaktuppgifterfinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Om du är av finländsk härkomst eller har en nära kontakt med Finland kan du beviljas uppehållstillstånd i Finland på grund av detta.
Då är du återflyttare (paluumuuttaja).
Huruvida du beviljas uppehållstillstånd beror på hur starka och nära släktband du har till Finland.
För att få tillståndet krävs inga andra skäl, som till exempel arbete eller studier.
Personer som aldrig själv har varit finska medborgare men vars ena förälder eller mor- eller farförälder är eller har varit infödd finsk medborgare betraktas som återflyttare (paluumuuttaja) av finsk härkomst.
Också före detta finska medborgare räknas som återflyttare.
Uppehållstillstånd för återflyttarefinska _ svenska _ engelska
Avkomlingar till infödda finska medborgare
Du kan beviljas uppehållstillstånd i Finland om minst en av dina föräldrar eller mor- eller farföräldrar är eller har varit infödd finsk medborgare.
Med infödd finsk medborgare avses en person som har fått finskt medborgarskap vid födseln.
När du ansöker om tillstånd måste du ge en tillförlitlig bild av din härkomst, som till exempel uppvisa den ursprungliga födelseattesten av en förälder eller en mor- eller farförälder samt ett intyg över ert släktskap.
Du krävs inte på redogörelse över din utkomst.
Före detta finska medborgare
Om du är en före detta finsk medborgare kan du på denna grund få uppehållstillstånd i Finland.
Förutsättningen är inte att du är en infödd finsk medborgare, utan du kan också ha fått det finska medborgarskapet på ansökan.
Du krävs inte på redogörelse över din utkomst.
Om du är en före detta finsk medborgare kan du återfå ditt finska medborgarskap genom att göra en medborgarskapsanmälan (kansalaisuusilmoitus).
Läs mer på InfoFinlands sida Finskt medborgarskap.
Ansökan om uppehållstillstånd
Du kan ansöka om uppehållstillstånd antingen utomlands innan du kommer till Finland eller i Finland.
Utomlands kan du ansöka om tillstånd vid den närmaste av Finlands ambassader, i Finland vid Migrationsverkets tjänsteställe.
Du måste personligen gå och lämna in ansökan om uppehållstillstånd.
Ta med dig originalexemplaren av de bilagor som krävs för ansökan när du lämnar in din ansökan vid ambassaden eller Migrationsverkets tjänsteställe.
När du ansöker om uppehållstillstånd måste du ha med dig ett pass för att kunna styrka din identitet.
När du ansöker om tillstånd tas dina fingeravtryck för det biometriska uppehållstillståndskortet.
Ansökan om uppehållstillstånd är avgiftsbelagd.
Avgiften måste betalas i samband med att man lämnar in sin tillståndsansökan.
Finsk personbeteckning
Om du får ett uppehållstillstånd i Finland registreras du automatiskt i det finska befolkningsdatasystemet.
Du får samtidigt även en finsk personbeteckning.
När du har flyttat till Finland ska du besöka magistraten på din hemort för att registrera dig som invånare.
Läs mer på InfoFinlands sida Registrering som invånare.
Uppehållstillstånd för avkomlingar till infödda finländarefinska _ svenska _ engelska
Uppehållstillstånd för före detta finska medborgarefinska _ svenska _ engelska
linkkiFinland-Samfundet:
Utlandsfinländarnas intresseorganisationfinska _ svenska _ engelska
Barn till en finsk medborgare
Barnet kan få uppehållstillstånd på grund av familjeband om hans/hennes förälder är finsk medborgare eller gift med en finsk medborgare och bor i Finland.
Barnet måste vara under 18 år gammalt och ogift den dag då beslutet om uppehållstillstånd fattas.
Den förälder till barnet som är bosatt i Finland måste vara barnets vårdnadshavare för att barnet ska kunna få uppehållstillstånd.
Om båda föräldrarna är vårdnadshavare måste även den andra föräldern ge sitt samtycke till att barnet flyttar till Finland.
En myndighet, till exempel en notaries publicus, måste verifiera överenskommelsen.
Familjebandet mellan föräldern och barnet måste bevisas, till exempel med en födelseattest med föräldrarnas namn.
Barnets vårdnadshavare gör ansökan för det minderåriga barnets del.
Även barnet måste vara närvarande när tillståndsansökan lämnas in.
Barn till en finsk medborgarefinska _ svenska _ engelska
Barn till en utländsk medborgare
Barnet kan få uppehållstillstånd på grund av familjeband om hans/hennes föräldrar har uppehållstillstånd i Finland och en förälder bor i Finland.
Barnet måste vara under 18 år gammalt och ogift den dag då beslutet om uppehållstillstånd fattas.
Även ett barn som föds i Finland behöver ett uppehållstillstånd i Finland.
Tillståndet måste sökas inom tre månader från barnets födelse.
Den förälder till barnet som är bosatt i Finland måste vara barnets vårdnadshavare för att barnet ska kunna få uppehållstillstånd.
Om båda föräldrarna är vårdnadshavare måste även den andra föräldern ge sitt samtycke till att barnet flyttar till Finland.
En myndighet, till exempel en notaries publicus, måste verifiera överenskommelsen.
Familjebandet mellan föräldern och barnet måste bevisas till exempel med en födelseattest med föräldrarnas namn.
För att barnet ska kunna få uppehållstillstånd måste hans/hennes uppehälle i Finland vara tryggat, till exempel genom förälderns löneinkomster.
Kravet på tillräcklig inkomst tillämpas dock inte på föräldern om barnet fötts innan föräldern anlänt till Finland och föräldern har flyktingstatus i Finland.
Om föräldern har fått flyktingstatus den 1.7.2016 eller senare, ska man ansöka om uppehållstillstånd för barnet inom tre månader från att föräldern fått flyktingstatus.
Ansökan kan även göras senare, men då tillämpas kravet på tillräcklig inkomst.
Om barnets förälder har uppehållstillstånd på grund av internetionellt skydd, men inte flyktingstatus, krävs att föräldern har en tillräcklig inkomst för att barnet ska kunna få uppehållstillstånd.
Barnets vårdnadshavare gör ansökan för det minderåriga barnets del.
Även barnet måste vara närvarande när tillståndsansökan lämnas in.
Barn till en utländsk medborgarefinska _ svenska _ engelska
Utkomstförutsättningfinska _ svenska _ engelska
Barn till en person som fått internationellt skyddfinska _ svenska _ engelska
Förälder eller annan vårdnadshavare
Om barnet inte är finsk medborgare måste han/hon ha uppehållstillstånd i Finland.
Barnet måste vara under 18 år gammalt och ogift den dag då beslutet om uppehållstillstånd fattas.
För att få uppehållstillstånd på grund av familjeband måste du vara barnets vårdnadshavare.
Vanligtvis är barnets mor eller far vårdnadshavare.
Vårdnadshavaren kan dock även vara någon annan, till exempel en mor- eller farförälder.
Familjebandet mellan barnet och föräldern måste bevisas till exempel med en födelseattest med föräldrarnas namn.
Om en annan vårdnadshavare än barnets mor eller far ansöker om uppehållstillstånd måste vårdnaden bevisas till exempel genom uppvisande av ett domstolsbeslut.
För att du ska kunna få uppehållstillstånd måste du ha tillräckliga medel för att leva i Finland.
Kravet på tillräcklig inkomst tillämpas dock inte på dig om ditt barn är en finsk medborgare.
Kravet på tillräcklig inkomst tillämpas inte heller om du varit barnets vårdnadshavare redan innan barnet anlänt till Finland och barnet har flyktingstatus i Finland.
Om barnet fått flyktingstatus den 1.7.2016 eller senare, ska du ansöka om uppehållstillstånd inom tre månader från att barnet fått flyktingstatus i Finland.
Ansökan kan även göras senare, men då tillämpas kravet på tillräcklig inkomst.
Vårdnadshavare till en finsk medborgarefinska _ svenska _ engelska
Vårdnadshavare till en utländsk medborgarefinska _ svenska _ engelska
Utkomstförutsättningfinska _ svenska _ engelska
Vårdnadshavare till en person som fått internationellt skyddfinska _ svenska _ engelska
Att ansöka om uppehållstillstånd
Vanligtvis måste du ansöka om ditt första uppehållstillstånd innan du kommer till Finland.
Ansök om tillståndet i ditt hemland eller i ett annat land där du vistas lagligt.
Du kan också ansöka om ditt första visum i Finland, om din familjemedlem är finsk medborgare och du själv är medborgare i ett visumfritt land, det vill säga du inte behöver visum för att komma till Finland.
Du kan ansöka om tillståndet på internet via tjänsten Enter Finland.
När du ställt ansökan ska du besöka Finlands beskickning närmast dig eller Migrationsverkets tjänsteställe för att styrka din identitet och visa upp originalexemplaren av ansökningsbilagorna.
Du ska besöka beskickningen eller tjänstestället inom tre månader efter att ha gjort ansökan på internet.
Ansökningen kan tas för behandling först när du besökt beskickningen eller tjänstestället.
Det är bra att boka en tid hos beskickningen eller tjänstestället i förväg.
Kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan, kommer detta att meddelas via ditt Enter Finland-konto.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du också lämna in en pappersansökan jämte bilagor vid Finlands beskickning närmast dig eller på Migrationsverkets tjänsteställe i Finland.
Du kan skriva ut ansökningsblanketten på Migrationsverkets webbplats.
Ansökan om uppehållstillstånd är avgiftsbelagd.
Avgiften ska betalas då ansökan ställs.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Finlands beskickningar utomlandsfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Finsk personbeteckning
Om du får ett uppehållstillstånd i Finland registreras du automatiskt i det finska befolkningsdatasystemet.
Du får samtidigt även en finsk personbeteckning.
När du har flyttat till Finland ska du besöka magistraten på din hemort för att registrera dig som invånare.
Läs mer på InfoFinlands sida Registrering som invånare.
Återkallande av uppehållstillstånd
Om du flyttar utomlands
Om ditt äktenskap eller registrerade parförhållande upphör
Om du förlorar ditt jobb
Återkallande av uppehållstillstånd
Ditt permanenta eller tidsbegränsade uppehållstillstånd återkallas om
du flyttar permanent från Finland
du har vistats två år utomlands utan avbrott.
Ditt permanenta eller tidsbegränsade uppehållstillstånd kan också återkallas om
du har uppgett felaktiga uppgifter i din ansökan om tillstånd
du har hemlighållit information som hade kunnat förhindra att tillståndet beviljas
ett annat Schengen-land begär att Finland återkallar ditt uppehållstillstånd.
Ett tidsbegränsat uppehållstillstånd kan också återkallas om de grunder på vilka tillståndet beviljades inte längre gäller.
Beslut om återkallelse av uppehållstillstånd fattas av Migrationsverket.
Om du flyttar utomlands
Om du ämnar flytta utomlands från Finland för två år, till exempel på grund av arbete eller studier, kan du ansöka hos Migrationsverket om att ditt uppehållstillstånd inte återkallas.
Ansökan är fritt formulerad men datum, underskrift och dina personuppgifter ska finnas med.
Ur ansökan bör även framgå hur länge och varför du studerar utomlands.
I din ansökning ska du motivera varför ditt uppehållstillstånd inte bör återkallas.
Ansökan ska göras innan du har vistats utomlands två år.
Om din finländska arbetsgivare har sänt dig utomlands för att arbeta förlorar du inte ditt uppehållstillstånd i Finland även om du vistas utomlands på grund av arbetet i över två år.
Om ditt äktenskap eller registrerade parförhållande upphör
Om du har ett tidsbestämt uppehållstillstånd med familjeband som grund kan det faktum att äktenskapet eller det registrerade parförhållandet upphör påverka uppehållstillståndet.
Om familjebandet inte längre existerar kan det hända att uppehållstillståndet inte förlängs.
Det är även möjligt att ett existerande tillstånd upphävs.
Uppehållstillståndet kan dock förlängas om du fortsättningsvis har starka band till Finland.
Exempel på sådana är:
barn eller andra familjemedlemmar i Finland
arbetsplats eller eget företag i Finland
studieplats i Finland
Om du skiljer dig på grund av att din make/maka varit våldsam mot dig kan ditt uppehållstillstånd förlängas trots skilsmässan.
Du ska lämna in en redovisning, exempelvis läkarintyg eller utlåtande från familjerådgivning.
Bifoga även till ansökan om uppehållstillstånd din egen redovisning av situationen.
Mer information om skilsmässa och upplösande av ett registrerat parförhållande hittar du på InfoFinlands sidor Skilsmässa.
Om du förlorar ditt jobb
Om du har ett uppehållstillstånd för arbetstagare som endast gäller arbete för en viss arbetsgivare och du förlorar din arbetsplats, ska du ansöka om ett nytt uppehållstillstånd för arbetstagare eller ett uppehållstillstånd på andra grunder.
Om Migrationsverket har beviljat dig ett uppehållstillstånd för arbetstagare och din anställning upphör tidigare än uppehållstillståndet, måste du eller din arbetsgivare skriftligt meddela Migrationsverket att din anställning upphör.
Om ditt uppehållstillstånd för arbetstagare inte har begränsats att gälla arbete för en viss arbetsgivare, utan för en viss bransch och tillståndet är fortfarande giltigt, kan du byta jobb inom samma bransch.
Mer information om arbete och företagande i Finland hittar du på InfoFinlands sida Arbete och entreprenörskap.
Mer information om uppehållstillstånd för arbetstagare och företagare hittar du på sidan Arbeta i Finland och Till Finland som företagare.
Om du redan har haft ett uppehållstillstånd i Finland, men tillståndet inte förlängs, fattar Migrationsverket beslut om utvisning.
Om du begår brott i Finland, kan du även utvisas på grund av brotten.
Om du blir utvisad, förfaller ditt eventuella giltiga uppehållstillstånd och du måste lämna landet.
Vanligtvis får du en tidsfrist inom vilken du måste lämna Finland.
Om du inte lämnar Finland inom tidsfristen avlägsnar polisen eller gränsbevakningsväsendet dig ur landet.
Enligt lag kan du inte utvisas om du hotas av dödsstraff, tortyr, förföljelse eller någon annan behandling som är omänsklig eller kränker människovärdet i ditt hemland.
Återkallelse av uppehållstillståndfinska _ svenska _ engelska
Avvisning och utvisningfinska _ svenska _ engelska
På denna sida finns information riktad till kvotflyktingar.
Information om att ansöka om asyl hittar du på InfoFinlands sida Till Finland som asylsökande.
Kvotflyktingar
Man kan inte ansöka om att bli kvotflykting via myndigheterna i Finland.
Man kan inte heller föreslå en annan person, till exempel en släkting eller vän, som kvotflykting.
Finland tar som kvotflyktingar emot personer som har flyktingstatus enligt
Förenta nationernas flyktingorganisation UNHCR.
Intervjuerna görs i de länder där flyktingarna vistas, vanligen i flyktingläger eller i UNHCR:s lokaler.
Information om val av kvotflyktingarfinska _ svenska _ engelska
Flytta till Finland
På webbsidan Movingtofinland.fi finns mycket information avsedd för kvotflyktingar om att flytta till Finland och om livet i Finland.
Information för flyktingarfinska _ engelska _ franska _ persiska _ arabiska _ kurdiska
Stöd till flyktingar
Finlands röda kors (FRK) hjälper kvotflyktingar när de flyttar till Finland.
När flyktingarna anländer till Finland kommer en anställd från röda korset till flygplatsen och tar emot dem.
Röda korsets frivilligarbetare hjälper även flyktingar att bosätta sig och integreras i Finland.
Flyktingar kan be om hjälp och rådgivning i rättsliga frågor bland annat från flyktingrådgivningen r.f. eller från rättshjälpsbyråer.
Finlands flyktinghjälp r.f. är en organisation som strävar efter att främja de grundläggande rättigheterna för flyktingar.
Organisationen utför informations-, utbildnings och socialarbete i Finland.
Flyktinghjälpen hjälper flyktingar och invandrare till exempel med ärenden som gäller integrering, boende och grundande av egna organisationer.
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
linkkiFinlands flyktinghjälp r.f.:
Stöd till flyktingarfinska _ svenska _ engelska
linkkiFinlands röda kors:
Stöd till flyktingarfinska _ svenska _ engelska
Rehabiliteringscentret för tortyrofferfinska _ engelska
Som flykting i Finland
På InfoFinlands sida Flykting hittar du mer information avsedd för flyktingar.
Make/maka till en finsk medborgare
Make/maka till en utländsk medborgare
Make/maka till en flykting
Partner
Att ansöka om uppehållstillstånd
Om maken/makan/sambon/partnern inte får uppehållstillstånd
Make/maka till en finsk medborgare
Om du har ingått äktenskap med en finländsk medborgare som är bosatt i Finland kan du få uppehållstillstånd i Finland på grund av familjeband.
Även en maka/make av samma kön kan få uppehållstillstånd, om ni är gifta eller i ett registrerat parförhållande.
Sambo med en finsk medborgare
Om du är sambo med en finsk medborgare som bor i Finland kan du få uppehållstillstånd på grund av familjeband.
Tillståndet kan beviljas om:
du har bott tillsammans med din sambo minst två år eller
du har ett gemensamt barn med din sambo (då uteblir kravet på gemensamt boende under två års tid) eller
det finns något annat vägande skäl för att bevilja tillståndet
Ifall du ansöker om tillstånd på dessa grunder måste du och din sambo bevisa att ni har bott tillsammans två år.
Som bevis godtas till exempel ett utdrag ur boenderegistret eller ett hyreskontrakt med bådas namn.
Om du och din sambo är bosatta i olika stater anses gemensamt boende till exempel under semesterresor inte som en tillräcklig grund för beviljande av uppehållstillstånd.
Varken du eller din sambo får vara gift med någon annan.
Försörjningsförutsättning för make/maka till en finsk medborgare
Om du är familjemedlem till en finsk medborgare, behöver din försörjning inte vara tryggad.
Du har obegränsad rätt att arbeta.
Du får börja arbeta först när du har fått ett uppehållstillstånd.
Information om hur du ansöker om tillståndet finns under rubriken Att ansöka om uppehållstillstånd.
Make eller maka till en finsk medborgarefinska _ svenska _ engelska
Sambo till en finsk medborgarefinska _ svenska _ engelska
Make/maka till en utländsk medborgare
Även en make/maka av samma kön kan få uppehållstillstånd.
Sambo med en utländsk medborgare
Om din sambo har uppehållstillstånd i Finland och bor i Finland kan du få uppehållstillstånd i Finland på grund av familjeband.
Du kan få tillståndet om:
du har bott tillsammans med din sambo minst två år eller
du har ett gemensamt barn tillsammans med din sambo (då uteblir kravet på gemensamt boende under två års tid)
Ifall du ansöker om tillstånd på dessa grunder måste du och din sambo bevisa att ni har bott tillsammans två år.
Som bevis duger till exempel ett utdrag ur boenderegistret eller ett hyreskontrakt med bådas namn.
Om du och din sambo är bosatta i olika stater anses gemensamt boende till exempel under semesterresor inte som en tillräcklig grund för beviljande av uppehållstillstånd.
Varken du eller din sambo får vara gift med någon annan.
Försörjningsförutsättning för make/maka till en utländsk medborgare
För att du ska få uppehållstillstånd i Finland måste du eller din make/maka ha tillräcklig inkomst även för din försörjning.
På Migrationsverkets sidor kan du kontrollera hur stor inkomst ni måste ha.
Om din maka/make fått uppehållstillstånd på grund av internationellt skydd, tillämpas kravet på tillräcklig inkomst på er.
Det är möjligt att i enskilda fall avvika från försörjningsförutsättningen, om det finns exceptionellt vägande skäl eller om barnets bästa kräver detta.
Information om hur du ansöker om tillståndet finns under rubriken Att ansöka om uppehållstillstånd.
Make eller maka till en utländsk medborgarefinska _ svenska _ engelska
Sambo till en utländsk medborgarefinska _ svenska _ engelska
Utkomstförutsättningfinska _ svenska _ engelska
Make/maka till en flykting
Om din maka/make har uppehållstillstånd i Finland på grund av internationellt skydd och flyktingstatus, kan du få uppehållstillstånd i Finland på grund av familjeband.
Sambo med flykting
Om din sambo har uppehållstillstånd i Finland på grund av internationellt skydd och flyktingstatus, kan du få uppehållstillstånd i Finland på grund av familjeband.
Du kan få tillståndet om:
du har bott tillsammans med din sambo minst två år eller
du har ett gemensamt barn tillsammans med din sambo (då uteblir kravet på gemensamt boende under två års tid)
Ifall du ansöker om tillstånd på dessa grunder måste du och din sambo bevisa att ni har bott tillsammans två år.
Som bevis duger till exempel ett utdrag ur boenderegistret eller ett hyreskontrakt med bådas namn.
Om du och din sambo är bosatta i olika stater anses gemensamt boende till exempel under semesterresor inte som en tillräcklig grund för beviljande av uppehållstillstånd.
Varken du eller din sambo får vara gift med någon annan.
Försörjningsförutsättning för make/maka/sambo/partner till en flykting
Försörjningsförutsättningen tillämpas på er på olika sätt, om din make/maka/sambo/partner har fått uppehållstillstånd på grund av internationellt skydd och har flyktingstatus i Finland.
Din försörjning behöver inte vara tryggad i följande fall:
Om din make/maka/sambo/partner har beviljats asyl eller godkänts som kvotflykting före den 1 juli 2016 och familjen har bildats före hen kom till Finland.
Om din make/maka/sambo/partner har fått flyktingstatus den 1 juli 2016 eller efter detta ska ansökan om uppehållstillstånd lämnas in inom tre månader efter att hen fått beslut på sin ansökan.
De tre månaderna räknas från den dag då din maka/make/sambo/partner delgivits beslutet.
Om du, av anledningar som du inte själv kan påverka, inte hinner ansöka om uppehållstillstånd inom tre månader, kan du ändå ansöka om familjeåterförening.
I din ansökan ska du ange varför tidsfristen på tre månader överskreds.
Du kan ansöka om familjeåterförening även senare, men då tillämpas kravet på tillräcklig inkomst på er.
Försörjningsförutsättningen gäller er även i det fall att ni gifte er efter att din make/maka kom till Finland.
I vissa enskilda fall kan man avvika från försörjningsförutsättningen om det finns exceptionellt vägande skäl eller om barnets bästa kräver detta.
Information om hur du ansöker om tillståndet finns under rubriken Att ansöka om uppehållstillstånd.
Maka eller make till en person som fått internationellt skyddfinska _ svenska _ engelska
Sambo till en person som fått internationellt skyddfinska _ svenska _ engelska
Försörjningsförutsättning för familjemedlemmar till personer som får internationellt skyddfinska _ svenska _ engelska
Partner
Man kan vanligen inte få uppehållstillstånd på grund av sällskapande.
I Finland är en person man sällskapar med inte en familjemedlem enligt lagen.
I vissa fall kan du ändå få ett tillfälligt (B) uppehållstillstånd i Finland på grund av sällskapande.
För att du ska kunna beviljas uppehållstillstånd i Finland måste ditt och din partners förhållande vara stadigt.
Ett bevis på stadigt sällskapande kan till exempel vara att er avsikt är att ingå äktenskap i Finland.
Varken du eller din partner får vara gift med någon annan.
För att du ska kunna få uppehållstillstånd måste du ha tillräckliga medel för ditt uppehälle.
Dessa medel bör vara fritt tillgängliga för dig till exempel på ditt eget bankkonto.
Inkomsterna för din partner som är bosatt i Finland beaktas inte.
Flick- eller pojkvän till en finsk medborgarefinska _ svenska _ engelska
Att ansöka om uppehållstillstånd
Vanligtvis måste du ansöka om ditt första uppehållstillstånd innan du kommer till Finland.
Ansök om tillståndet i ditt hemland eller i ett annat land där du vistas lagligt. Du kan också ansöka om ditt första uppehållstillstånd i Finland om din make eller maka är finsk medborgare och du själv är medborgare i ett visumfritt land, det vill säga du inte behöver visum för att komma till Finland.
Du kan ansöka om tillståndet på internet via tjänsten Enter Finland.
När du ställt ansökan ska du besöka Finlands beskickning närmast dig eller Migrationsverkets tjänsteställe för att styrka din identitet och visa upp originalexemplaren av ansökningsbilagorna.
Du ska besöka beskickningen eller tjänstestället inom tre månader efter att ha gjort ansökan på internet.
Ansökningen kan tas för behandling först när du besökt beskickningen eller tjänstestället.
Vanligtvis måste du boka en tid hos beskickningen eller tjänstestället i förväg.
Kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan, kommer detta att meddelas via ditt Enter Finland-konto.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du också lämna in en pappersansökan jämte bilagor vid Finlands beskickning närmast dig eller på Migrationsverkets tjänsteställe i Finland.
Du kan skriva ut ansökningsblanketten på Migrationsverkets webbplats.
Ansökan om uppehållstillstånd är avgiftsbelagd.
Avgiften ska betalas då ansökan ställs.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Finlands beskickningar utomlandsfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Handläggningstider för tillståndsansökningarfinska _ svenska _ engelska
Finsk personbeteckning
Om du får ett uppehållstillstånd i Finland registreras du automatiskt i det finska befolkningsdatasystemet.
Du får samtidigt även en finsk personbeteckning.
När du har flyttat till Finland ska du besöka magistraten på din hemort för att registrera dig som invånare.
Läs mer på InfoFinlands sida Registrering som invånare.
Om maken/makan/sambon/partnern inte får uppehållstillstånd
En make/maka/sambo/partner beviljas inte uppehållstillstånd om förutsättningarna för uppehållstillstånd inte uppfylls.
Man kan låta bli att bevilja tillståndet även då de finländska myndigheterna anser att parterna har ingått äktenskap endast för uppehållstillståndets skull och att makarna inte avser att leva tillsammans som en familj.
Myndigheterna kan misstänka att parterna ingått äktenskap endast för uppehållstillståndets skull till exempel om ni har ingått äktenskap efter endast en kort bekantskap, om det är stor åldersskillnad mellan er eller om den ena av er har haft flera korta äktenskap.
Om du får ett nekande beslut på din tillståndsansökan kan du överklaga den till förvaltningsdomstolen.
Du får instruktioner för detta bifogade till tillståndsbeslutet.
Läs mer om problem med uppehållstillståndet på InfoFinlands sida Problem med uppehållstillståndet.
Om du redan är i Finland och får ett negativt beslut om uppehållstillstånd från Migrationsverket (Maahanmuuttovirasto), måste du antingen lämna Finland eller överklaga beslutet.
Du får vistas i Finland så länge som behandlingen av besvären pågår.
Du kan överklaga också om du har ansökt om uppehållstillstånd utomlands.
Då måste du vänta på behandlingen av besvären utomlands.
Om du är asylsökande i Finland eller offer för människohandel, har du rätt att få stöd för frivillig återresa (vapaaehtoisen paluun tuki), om du beslutar att återvända till ditt hemland.
Läs mer under rubriken Stöd för frivillig återresa.
Att överklaga ett beslut om uppehållstillstånd
En besvärsanvisning om hur beslutet får överklagas bifogas alltid beslutet.
Besvären behandlas av förvaltningsdomstolen (hallinto-oikeus).
Förvaltningsdomstolen kan antingen avslå besvären eller sända ärendet till Migrationsverket för ny behandling.
Avslag innebär att Migrationsverkets beslut förblir gällande.
Om förvaltningsdomstolen avslår besvären kan du i vissa fall ansöka om besvärstillstånd hos högsta förvaltningsdomstolen (korkein hallinto-oikeus).
Om högsta förvaltningsdomstolen beviljar besvärstillstånd, behandlar den besvären.
Du kan få hjälp med att överklaga av antingen en privat jurist, en statlig rättshjälpsbyrå (valtion oikeusaputoimisto) eller Flyktingrådgivningen rf (Pakolaisneuvonta) (endast asylsökande).
På InfoFinlands sida Behöver du en jurist? finns mer information om hur du kan få hjälp i juridiska ärenden.
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Att lämna Finland
Om du får avslag på din ansökan om uppehållstillstånd eller om förvaltningsrätten avslår ditt överklagande, måste du lämna Finland.
Du ges möjlighet att lämna landet frivilligt.
Tidsfristen är vanligtvis 30 dagar.
Om du inte lämnar landet inom tidsfristen, avlägsnar polisen eller gränsbevakningsväsendet dig ur landet.
Du får inreseförbud till Schengenområdet om:
Du har brutit mot inresereglerna och din ansökan har avslagits, till exempel på grund av skenäktenskap.
Du har begått brott och du anses utgöra ett hot mot den allmänna ordningen och säkerheten.
Din asylansökan avslås i ett påskyndat förfarande.
Du inte lämnar landet frivilligt inom den tidsfrist som meddelats för dig.
När du har inreseförbud kan du inte besöka Finland eller något annat Schengenland.
Avvisning och utvisningfinska _ svenska _ engelska
Stöd för frivillig återresa
Om du vill återvända till ditt hemland kan du i vissa fall få stöd för frivilligt återvändande.
Stödet består antingen av pengar eller tjänster.
Penningsummans storlek beror på vilket land du återvänder till.
Tjänsten kan till exempel vara att du får hjälp med att leta efter en bostad eller arbetsplats i det land dit du återvänder.
Du kan få stöd om:
du har fått ett negativt beslut på din asylansökan
du återkallar din asylansökan
du är ett offer för människohandel och du inte har en hemkommun i Finland
du har ett tillfälligt uppehållstillstånd på grund av hinder för avlägsnande ur landet
du har fått tillfälligt skydd
din flyktingstatus i Finland har upphört eller återkallats eller det har fattats beslut om att avvisa dig
du har fått humanitärt skydd, men ditt uppehållstillstånd löper ut eller har redan löpt ut.
Om du är kund hos en mottagningscentral kan du ansöka om stöd för frivilligt återvändande vid din egen mottagningscentral.
Om du inte är kund hos en mottagningscentral kan du ansöka om stöd hos Migrationsverket.
Frivillig återflyttningfinska _ svenska _ engelska
Söka asyl
Asylsökande från Europeiska unionens område
Minderåriga asylsökande
Handläggning av asylansökan
Asylsamtal
Positivt beslut
Negativt beslut
Rättshjälp för asylsökande
Asylsökandes rätt att arbeta
Du kan söka asyl i Finland om du har välgrundad fruktan för förföljelse i ditt hemland.
Orsaker till förföljelse kan vara etniskt ursprung, religion, medborgarskap, tillhörighet till en viss grupp i samhället eller politiska åsikter.
Migrationsverket utreder om det finns asylskäl och fattar ett beslut.
Du kan endast söka asyl för dig själv.
Broschyren Information till asylsökandefinska _ svenska _ engelska _ ryska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
Söka asyl
Du kan endast söka asyl i Finland på det finska territoriet.
Det finns ingen särskild asylansökningsblankett som du skulle kunna fylla i förväg.
När du kommer till Finland, meddela gränskontrollmyndigheten eller polisen genast att du vill söka asyl.
Gränskontrollmyndigheten eller polisen registrerar dig som asylsökande, antecknar uppgifter om dig och tar dina fingeravtryck.
När myndigheten har mottagit din asylansökan, hänvisas du till ett mottagningscenter.
Där kan du bo under tiden då Migrationsverket behandlar din ansökan.
Du kan även bo någon annanstans, men då måste du själv bekosta boendet.
Att söka asyl i Finlandfinska _ svenska _ engelska
Asylsökande från Europeiska unionens område
Inom EU (och i Schweiz, Norge, Island och Liechtenstein) måste man söka asyl i det land, till vars territorium man kommer först.
Om du har sökt asyl eller vistats i något annat EU-land (eller i Schweiz, Norge, Island eller Liechtenstein) innan du kom till Finland, behandlas din ansökan inte i Finland.
I detta fall avvisas du tillbaka till det land där du var innan du kom till Finland.
Detta kallas för Dublinprocessen.
Om du är medborgare i ett EU-land, får du sannolikt inte asyl i Finland.
Finland anser att alla EU-länder är trygga för medborgarna.
Likväl utreds alla ansökningar som EU-medborgare skickar in.
På InfoFinlands sida EU-medborgare hittar du information om flytt till Finland av andra skäl än som asylsökande.
Att lämna asylansökan utan prövningfinska _ svenska _ engelska
Minderåriga asylsökande
Om du är under 18 år gammal och kommer till Finland som asylsökande utan vårdnadshavare, förordnas du ett ombud.
Ombudet är en pålitlig vuxen person som hjälper dig med olika ärenden under tiden då Migrationsverket behandlar din ansökan.
Ombudet följer med dig när du ska prata med myndigheter.
Dessutom utreder ditt ombud om du kan återförenas med din familj.
Du har rätt till boende, mat och hälsovård.
Du har även rätt att gå i skola.
Ensamkommande barn(pdf, 674)finska _ svenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ persiska _ arabiska _ kurdiska
Handläggning av asylansökan
Migrationsverket handlägger din ansökan och fattar ett beslut.
Migrationsverket utreder din identitet och resväg till Finland och bedömer om du kan beviljas asyl i Finland.
Det är vanligt att behandlingen av ansökan tar flera månader.
När du har sökt asyl har du rätt att vistas i Finland medan din ansökan behandlas.
Under denna tid kan du inte resa utomlands.
Om du reser kan myndigheterna besluta att din ansökan inte längre gäller.
Migrationsverket skickar dig en kallelse till asylsamtal.
I kallelsen anges tolkningsspråket, den exakta adressen till verksamhetsstället där samtalet hålls och klockslaget.
Handläggning av asylansökanfinska _ svenska _ engelska
Asylsamtal
Asylsamtalet (turvapaikkapuhuttelu) är den viktigaste händelsen under behandlingen av din ansökan.
Under samtalet ställs frågor om de händelser och orsaker som tvingade dig att lämna ditt hemland.
Det är viktigt att du beskriver allt som hänt så exakt som möjligt.
Migrationsverket beslutar baserat på din berättelse om du beviljas asyl i Finland.
Som asylsökande har du rätt att använda ett rättsbiträde under samtalet.
Biträdet deltar i asylsamtalet efter sitt eget omdöme.
Om du behöver en tolk, skaffar Migrationsverket tolken.
Positivt beslut
Du får stanna i Finland om du beviljas asyl eller uppehållstillstånd på andra grunder.
Du kan beviljas asyl i Finland om myndigheterna anser att du blir förföljd i ditt hemland på grund av
etniskt ursprung,
religion,
medborgarskap,
tillhörighet till en viss grupp i samhället eller
politiska åsikter.
Om du inte får asyl kan du i vissa fall beviljas uppehållstillstånd på grund av alternativt skydd.
Du kan beviljas uppehållstillstånd på grund av alternativt skydd om du hotas av:
dödsstraff eller avrättning,
tortyr eller någon annan behandling eller bestraffning som är omänsklig eller kränker människovärdet eller
om du utsätts för allvarlig personlig fara på grund av en väpnad konflikt.
När du söker asyl utreder Migrationsverket samtidigt om du kan få uppehållstillstånd på någon annan grund.
Asylfinska _ svenska _ engelska
Negativt beslut
Om du inte beviljas asyl eller uppehållstillstånd på någon annan grund blir du avvisad från Finland.
Du har även möjlighet att överklaga ett negativt beslut till förvaltningsdomstolen.
Bifogat till beslutet finns en anvisning om hur du överklagar.
På InfoFinlands sida Negativt beslut om uppehållstillstånd hittar du information om vad du kan göra om du får ett negativt beslut.
Ändringssökande i asylbeslutfinska _ svenska _ engelska
Avvisning av en asylsökandefinska _ svenska _ engelska
Rättshjälp för asylsökande
Under tiden då din ansökan behandlas kan du få rådgivning och rättshjälp vid den offentliga rättshjälpsbyrån.
Kontakta rättshjälpsbyrån om du vill ha ett rättsbiträde.
Vid behov hjälper mottagningscentret dig.
Rättshjälpsbyrån (oikeusaputoimisto) kan även hänvisa dig till en privat jurist eller en privat juristbyrå.
Du kan även få rådgivning hos Flyktingrådgivningen rf (Pakolaisneuvonta ry).
Flyktingrådgivningen ger rådgivning även till personer som vistas i Finland utan uppehållstillstånd.
linkkiRättsväsendet:
Rättshjälpsbyråerfinska _ svenska _ engelska
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Asylsökandes rätt att arbeta
Du får förvärvsarbeta i Finland om det har gått tre månader sedan du lämnade in din asylansökan och du har ett giltigt pass eller någon annan resehandling som du har företett till myndigheten när du sökte asyl.
Om du inte företedde en giltig resehandling till myndigheten i samband med din asylansökan får du förvärvsarbeta i Finland när det har gått sex månader sedan du lämnade in din asylansökan.
Du har rätt att arbeta tills du har fått ett lagakraftvunnet beslut på din asylansökan.
Om Migrationsverket ger dig ett positivt beslut på din asylansökan, får du uppehållstillstånd.
I det ingår nästan alltid rätt att arbeta.
Om Migrationsverket fattar ett negativt beslut på din asylansökan, har du rätt att arbeta under tiden då en eventuell överklagan behandlas.
För att arbeta måste du ha ett finländskt skattekort.
Hämta ett skattekort på den närmaste skattebyrån och lämna kortet till din arbetsgivare.
Läs mer på InfoFinlands sida Skattekort.
Om du arbetar permanent kan du även ansöka om uppehållstillstånd i Finland på grund av arbete.
På InfoFinlands sida Arbeta i Finland hittar du mer information om uppehållstillstånd för arbetstagare.
Asylsökandes rätt att arbetafinska _ svenska _ engelska
Uppehållstillstånd på andra grunderfinska _ svenska _ engelska
Om du vill flytta till en familjemedlem som bor i Finland behöver du ett uppehållstillstånd.
Om du bara vill hälsa på hos din familjemedlem i Finland hittar du mer information på InfoFinlands sida Kort vistelse i Finland.
Alla familjemedlemmar kan inte få uppehållstillstånd.
Vanligen kan man få tillstånd om man är make/maka, sambo, minderårigt barn eller förälder till minderårigt barn till personen bosatt i Finland.
Ofta krävs det även att personen bosatt i Finland ska ha tillräckliga medel för att försörja en familjemedlem som flyttar till Finland.
Notera att separata regler gäller för familjemedlemmar till EU-medborgare (inte finländska medborgare).
Om du är familjemedlem till en EU-medborgare bosatt i Finland hittar du mer information om tillståndsärenden på InfoFinlands sidan EU-medborgare.
Mer information om hur familjemedlemmar kan få uppehållstillstånd finns på InfoFinlands sidor Uppehållstillstånd för make eller maka, Uppehållstillstånd för barn eller förälder, Uppehållstillstånd för övriga anhöriga.
På InfoFinlands sida Familjemedlem hittar du mer information avsedd för personer som flyttar av familjeskäl.
Till Finland på grund av familjebandfinska _ svenska _ engelska
Rådgivning i uppehållstillståndsärenden
Om du har problem eller oklarheter med uppehållstillståndet, kan du ta kontakt med följande instanser för att be om råd:
Finlands beskickningar utomlands
Invandrarrådgivarna i din kommun i Finland
På Migrationsverkets webbplats finns mycket information om uppehållstillstånd.
Migrationsverket ger rådgivning angående tillstånd också per telefon.
Finlands beskickningar utomlands betjänar personer som ansöker om uppehållstillstånd i utlandet.
Många städer har rådgivningstjänster för invandrare med rådgivare som specialiserat sig på invandringsfrågor.
Flyktingsrådgivningen bistår asylsökande juridiskt i asylprocessen.
Dessutom tillhandahåller Flyktingrådgivningen allmän juridisk rådgivning för andra utlänningar.
Vänligen observera att endast Migrationsverket kan fatta beslut om uppehållstillstånd.
Information om uppehållstillståndfinska _ svenska _ engelska
linkkiFlyktingrådgivningen rf:
Juridisk rådgivningfinska _ engelska _ franska _ arabiska
Också andra anhöriga till finska medborgare än en make/maka, en sambo, föräldrar till minderåriga barn eller minderåriga barn kan i vissa fall få uppehållstillstånd i Finland på grund av familjeband.
Även andra anhöriga till en person som har ett uppehållstillstånd på grund av internationellt skydd kan beviljas uppehållstillstånd.
Om uppehållstillståndet beviljats på någon annan grund än internationellt skydd, kan andra anhöriga inte få uppehållstillstånd.
En annan anhörig kan få uppehållstillstånd om han eller hon är helt beroende av den anhöriga som bor i Finland.
På denna grund kan uppehållstillstånd beviljas till exempel för en förälder till en myndig (18 år gammal) person.
Enbart ekonomiskt beroende eller svag hälsa räcker ändå inte för att beviljas uppehållstillstånd.
En annan anhörig kan få uppehållstillstånd också om han eller hon levt tillsammans som en familjemedlem till den anhöriga som är bosatt i Finland, innan denna person kom till Finland.
Dessutom krävs det att familjelivet upphört på grund av ett tvingande skäl, till exempel för att man blivit flyktingar.
Annan anhörig till en finsk medborgarefinska _ svenska _ engelska
Annan anhörig till en person som fått internationellt skyddfinska _ svenska _ engelska
Att ansöka om uppehållstillstånd
Vanligtvis måste du ansöka om ditt första uppehållstillstånd innan du kommer till Finland.
Ansök om tillståndet i ditt hemland eller i ett annat land där du vistas lagligt.
Du kan ansöka om tillståndet på internet via tjänsten Enter Finland.
När du ställt ansökan ska du besöka Finlands beskickning närmast dig eller Migrationsverkets tjänsteställe för att styrka din identitet och visa upp originalexemplaren av ansökningsbilagorna.
Du ska besöka beskickningen eller tjänstestället inom tre månader efter att ha gjort ansökan på internet.
Ansökningen kan tas för behandling först när du besökt beskickningen eller tjänstestället.
Vanligtvis måste du boka en tid hos beskickningen eller tjänstestället i förväg.
Kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan, kommer detta att meddelas via ditt Enter Finland-konto.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du också lämna in en pappersansökan jämte bilagor vid Finlands beskickning närmast dig eller på Migrationsverkets tjänsteställe i Finland.
Du kan skriva ut ansökningsblanketten på Migrationsverkets webbplats.
Ansökan om uppehållstillstånd är avgiftsbelagd.
Avgiften ska betalas då ansökan ställs.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Finlands beskickningar utomlandsfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Finsk personbeteckning
Om du får ett uppehållstillstånd i Finland registreras du automatiskt i det finska befolkningsdatasystemet.
Du får samtidigt även en finsk personbeteckning.
När du har flyttat till Finland ska du besöka magistraten på din hemort för att registrera dig som invånare.
Läs mer på InfoFinlands sida Registrering som invånare.
Ansök om studieplats
Teckna en tillräckligt omfattande sjukförsäkring i ditt hemland
Reservera tillräckliga medel för din försörjning
Ansök om uppehållstillstånd för studerande
Uppehållstillstånd för studerande från andra EU-länder
Fortsatt uppehållstillstånd för studerande
När du avslutar dina studier
För praktik till Finland
Den här sidan är avsedd för dig som är medborgare i något annat land än ett EU-land, Norge, Island, Schweiz eller Liechtenstein.
Om du ska studera i Finland längre än 90 dagar behöver du ett uppehållstillstånd på grund av studier.
Du kan studera mindre än 90 dagar i Finland utan uppehållstillstånd.
Om du ska flytta till Finland för studier måste du ta hand om följande:
Ansök om studieplats
Innan du kan ansöka om uppehållstillstånd måste du skaffa dig en studieplats i Finland.
Godkända läroanstalter är läroanstalter efter grundskolan, till exempel universitet, högskolor och yrkesläroanstalter.
Studieplatsen ska uppfylla ett av följande villkor:
studierna leder till yrke eller examen
du deltar i ett utbytesprogram mellan läroanstalter eller något annat utbytesprogram
du avlägger en kompletterande utbildning eller en specialutbildning som hör till din examen.
Du kan ansöka om studieplats i skolornas gemensamma ansökan på våren eller hösten.
Till vissa utbildningar är den gemensamma ansökan (yhteishaku) redan i januari.
Ta i god tid reda på när du kan ansöka om en studieplats.
Fyll i ansökan i tjänsten Opintopolku.fi.
På InfoFinlands sida Ansökan till utbildning hittar du mer information om hur du ansöker om en studieplats i Finland.
Teckna en tillräckligt omfattande sjukförsäkring i ditt hemland
Som studerande betalar du själv vårdkostnaderna om du insjuknar i Finland.
För ditt uppehållstillstånd behöver du en privat försäkring som täcker kostnaderna för sjukdom och läkemedel.
Du kan teckna en försäkring hos ett försäkringsbolag i ditt hemland eller fråga om en lämplig försäkring hos internationella försäkringsbolag.
Alla försäkringar ska uppfylla följande villkor:
Försäkringens självrisk får inte överstiga 300 euro.
Försäkringen ska gälla under hela din vistelse i Finland.
Försäkringen ska gälla när du kommer till Finland.
Försäkringen får inte vara en vanlig reseförsäkring.
Säg inte upp din försäkring.
Om du insjuknar måste du själv betala läkar- och sjukhuskostnaderna.
Hur stora vårdkostnader som försäkringen måste täcka beror på hur länge dina studier varar.
Om dina studier i Finland till exempel varar mindre än två år, ska försäkringen täcka sjukvårdskostnader upp till minst 120 000 euro.
Om du har det europeiska sjukvårdskortet (European Health Insurance Card, EHIC), behöver du ingen separat försäkring.
Sjukvårdskortet ska vara giltigt under hela din vistelse i Finland.
Försäkring för studerandefinska _ svenska _ engelska
Reservera tillräckliga medel för din försörjning
Du måste också själv ansvara för levnadskostnaderna i Finland.
Du behöver ha minst 560 euro disponibla medel i månaden för att kunna betala för boende, mat och andra utgifter.
För en vistelse som varar ett år ska du alltså ha 6 720 euro i disponibla medel.
Försörjningsförutsättningen kan i vissa fall undgås.
Om till exempel läroanstalten ordnar dig en gratis bostad och även gratis måltider behöver du ha en mindre summa i disponibla medel.
Om studierna är avgiftsbelagda måste du även se till att du har tillräckliga medel för din försörjning efter att du har betalat läsårsavgiften.
Beloppet som krävs ska finnas på ditt bankkonto eller också ska du ha ett intyg över ett stipendium som beviljats av en officiell instans.
Sådana stipendier är till exempel de som beviljats av staten, läroanstalter eller organisationer.
Sponsringslöften eller kontoutdrag från privatpersoner, såsom släktingar, bekanta eller arbetsgivare, godkänns inte.
Försörjningsförutsättning för studerandefinska _ svenska _ engelska
Ansök om uppehållstillstånd för studerande
Du måste ansöka om ditt första uppehållstillstånd innan du kommer till Finland.
Du kan ansöka om tillståndet på internet via tjänsten Enter Finland.
När du ställt ansökan ska du besöka Finlands beskickning närmast dig för att styrka din identitet och visa upp originalexemplaren av ansökningsbilagorna.
Du ska besöka beskickningen inom tre månader efter att ha gjort ansökan på internet.
Ansökningen kan tas för behandling först när du besökt beskickningen.
Vanligtvis måste du boka en tid hos beskickningen i förväg.
Kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan kommer detta att meddelas via ditt konto.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du också lämna in en pappersansökan jämte bilagor vid Finlands beskickning närmast dig.
Du kan skriva ut ansökningsblanketten på Migrationsverkets webbplats.
Handläggningen av ansökan är avgiftsbelagd.
Du måste betala avgiften när du lämnar in ansökan om uppehållstillstånd.
Du ska bifoga följande handlingar till din ansökan om uppehållstillstånd för studerande:
Giltigt pass
Passfoto (anvisningar för fotot finns på Migrationsverkets webbplats)
Närvarointyg (intyg över att du är studerande vid en läroanstalt som är godkänd i Finland)
En utredning över att du har tillräckliga medel för din försörjning
Ett försäkringsintyg eller en kopia av det europeiska sjukvårdskortet
En utredning över att du har betalat läsårsavgiften eller har ett stipendium
Tidigare examensbetyg (om du inte ska avlägga examen eller är en utbytesstudent)
Eventuella arbetsintyg (om du inte ska avlägga examen eller är en utbytesstudent)
Information om uppehållstillstånd för studierfinska _ svenska _ engelska
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Finlands beskickningar utomlandsfinska _ svenska _ engelska
Uppehållstillstånd för studerande från andra EU-länder
Du behöver inget uppehållstillstånd i Finland om du har ett uppehållstillstånd som beviljats i ett annat EU-land och om du studerar vid en högskola.
Dessutom måste dina studier:
innefatta internationell rörlighet i ett EU-program eller ett mångformigt program eller
omfattas av ett avtal mellan två eller fler högskolor.
I detta fall måste du göra en underrättelse om rörlighet till Migrationsverket.
Du får studera i Finland högst 360 dagar när du gör en underrättelse om rörlighet.
Underrättelse om rörlighet i Finlandfinska _ svenska _ engelska
Finsk personbeteckning
Om du får ett uppehållstillstånd i Finland registreras du automatiskt i det finska befolkningsdatasystemet.
Du får samtidigt även en finsk personbeteckning.
När du har flyttat till Finland ska du besöka magistraten på din hemort för att registrera dig som invånare.
Läs mer på InfoFinlands sida Registrering som invånare.
Fortsatt uppehållstillstånd för studerande
Uppehållstillstånd för studerande beviljas högst för två år i taget.
Om dina studier fortsätter men uppehållstillståndet håller på att gå ut ska du ansöka om fortsatt uppehållstillstånd.
Kom ihåg att ansöka om fortsatt uppehållstillstånd för studerande i god tid innan giltighetstiden för det första tillståndet går ut.
Observera att Migrationsverket (Maahanmuuttovirasto) även kontrollerar om grunden för din vistelse i Finland verkligen har varit studier.
Om du till exempel avlägger en grundexamen vid universitet, högskola eller yrkeshögskola bör du avlägga 45 studiepoäng under ett läsår för att uppfylla villkoren för fortsatt uppehållstillstånd.
Du ska bifoga ett studieregisterutdrag till din ansökan om fortsatt uppehållstillstånd.
Fortsatt uppehållstillstånd för studerandefinska _ svenska _ engelska
När du avslutar dina studier
Om du har avlagt en examen i Finland kan du få ett tillfälligt uppehållstillstånd för arbetssökande.
Detta tillstånd kan beviljas endast som ett fortsatt tillstånd till ett uppehållstillstånd för studerande.
Du ska ansöka om tillståndet innan ditt uppehållstillstånd för studerande går ut.
Uppehållstillstånd för arbetssökande kan beviljas för högst ett år.
Om du får ett jobb kan du börja arbeta direkt.
Du måste ansöka om ett nytt uppehållstillstånd på grund av arbete innan ditt uppehållstillstånd för arbetssökande går ut.
Uppehållstillstånd för sökande av arbetefinska _ svenska _ engelska
Till Finland som praktikant
Om du studerar utomlands och vill komma till Finland för arbetspraktik behöver du ett uppehållstillstånd på grund av praktik.
Mer information hittar du på Migrationsverkets webbplats.
Praktik i Finlandfinska _ svenska _ engelska
InfoFinlands sida Utländska studerande i Finland innehåller viktig information om studielivet i Finland.
Information för utländska studerandeengelska
Migrationsverket:
Presentation av e-tjänsten Enter Finland
Du kan få permanent uppehållstillstånd (pysyvä oleskelulupa) (P), om
du bott i Finland i minst fyra år med A-tillstånd och
inte under tiden har bott utomlands i över två år och
grunden för de tidigare uppehållstillstånden fortfarande existerar
Om du hade A-tillstånd då du kom till Finland beräknas de fyra åren från den dag du anlände till Finland Om du fått A-tillstånd i Finland beräknas de fyra åren från den dag då det första A-tillståndet trädde i kraft.
Om du har fått internationellt skydd i Finland beräknas de fyra åren från att du anlände till Finland.
Permanent uppehållstillstånd kan eventuellt inte beviljas om:
du har begått ett brott som är belagt med fängelsestraff
du är misstänkt för ett brott som är belagt med fängelsestraff
du har begått två eller flera brott
du misstänks för två eller flera brott
Permanen uppehållstillstånd gäller tills vidare.
Tillstånet kan dras tillbaka om du permanent flyttar från Finland, uppehåller dig utomlands kontinuerligt i minst två år eller har lämnar felaktiga uppgifter då du ansökt om tillståndet.
EU-uppehållstillstånd för tredjelandsmedborgare som uppehållit sig länge i landet
Tredjelandsmedborgare äe medborgare i annat land än de nordiska länderna, EU-länderna, Liechtenstein eller Schweiz.
Du kan beviljas EU-uppehållstillstånd (P-EU) för tredjelandsmedborgare om:
du har bott i Finland i minst fem år med A-tillstånd och
inte under denna tid har bott utomlands längre än 10 månader och
grunden för de tidigare uppehållstillstånden fortfarande existerar
P-EU-tillstånd ansöks om på samma sätt som permanent uppehållstillstånd.
P-EU-tillstånd gäller tills vidare.
P-EU-tillståndsansökan kan även avslås på samma grunder som permanent uppehållstillstånd.
Ansökan
Du kan ansöka om permanent uppehållstillstånd på internet i tjänsten Enter Finland.
När du ställt ansökan ska du besöka Migrationsverkets tjänsteställe för att styrka din identitet.
Ta med dig en identitetshandling och originalexemplaren av ansökningsbilagorna.
Det är bra att boka en tid hos Migrationsverkets tjänsteställe i förväg.
Du kan boka tiden via Migrationsverkets elektroniska tidsbokningssystem.
Om du gjort ansökningen på internet, kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan, kommer detta att meddelas via ditt Enter Finland-konto.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du ansöka om tillståndet med en pappersblankett vid Migrationsverkets tjänsteställe.
Du kan skriva ut blanketten på Migrationsverkets webbplats.
Boka en tid vid tjänstestället och ta med dig den ifyllda ansökningen, bilagorna och en identitetshandling.
Handläggning av ansökan är avgiftsbelagd.
Avgiften ska betalas då ansökan ställs.
I tjänsten Enter Finland kan du betala med nätbankskoderna för en finsk bank eller med kreditkort.
Permanent uppehållstillståndfinska _ svenska _ engelska
Ansökningsblankettfinska _ svenska _ engelska
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Barn till en finsk medborgare
Barnet kan få uppehållstillstånd på grund av familjeband om hans/hennes förälder är finsk medborgare eller gift med en finsk medborgare och bor i Finland.
Barnet måste vara under 18 år gammalt och ogift den dag då beslutet om uppehållstillstånd fattas.
Den förälder till barnet som är bosatt i Finland måste vara barnets vårdnadshavare för att barnet ska kunna få uppehållstillstånd.
Om båda föräldrarna är vårdnadshavare måste även den andra föräldern ge sitt samtycke till att barnet flyttar till Finland.
En myndighet, till exempel en notaries publicus, måste verifiera överenskommelsen.
Familjebandet mellan föräldern och barnet måste bevisas, till exempel med en födelseattest med föräldrarnas namn.
Barnets vårdnadshavare gör ansökan för det minderåriga barnets del.
Även barnet måste vara närvarande när tillståndsansökan lämnas in.
Barn till en finsk medborgarefinska _ svenska _ engelska
Barn till en utländsk medborgare
Barnet kan få uppehållstillstånd på grund av familjeband om hans/hennes föräldrar har uppehållstillstånd i Finland och en förälder bor i Finland.
Barnet måste vara under 18 år gammalt och ogift den dag då beslutet om uppehållstillstånd fattas.
Även ett barn som föds i Finland behöver ett uppehållstillstånd i Finland.
Tillståndet måste sökas inom tre månader från barnets födelse.
Den förälder till barnet som är bosatt i Finland måste vara barnets vårdnadshavare för att barnet ska kunna få uppehållstillstånd.
Om båda föräldrarna är vårdnadshavare måste även den andra föräldern ge sitt samtycke till att barnet flyttar till Finland.
En myndighet, till exempel en notaries publicus, måste verifiera överenskommelsen.
Familjebandet mellan föräldern och barnet måste bevisas till exempel med en födelseattest med föräldrarnas namn.
För att barnet ska kunna få uppehållstillstånd måste hans/hennes uppehälle i Finland vara tryggat, till exempel genom förälderns löneinkomster.
Kravet på tillräcklig inkomst tillämpas dock inte på föräldern om barnet fötts innan föräldern anlänt till Finland och föräldern har flyktingstatus i Finland.
Om föräldern har fått flyktingstatus den 1.7.2016 eller senare, ska man ansöka om uppehållstillstånd för barnet inom tre månader från att föräldern fått flyktingstatus.
Ansökan kan även göras senare, men då tillämpas kravet på tillräcklig inkomst.
Om barnets förälder har uppehållstillstånd på grund av internetionellt skydd, men inte flyktingstatus, krävs att föräldern har en tillräcklig inkomst för att barnet ska kunna få uppehållstillstånd.
Barnets vårdnadshavare gör ansökan för det minderåriga barnets del.
Även barnet måste vara närvarande när tillståndsansökan lämnas in.
Barn till en utländsk medborgarefinska _ svenska _ engelska
Utkomstförutsättningfinska _ svenska _ engelska
Barn till en person som fått internationellt skyddfinska _ svenska _ engelska
Förälder eller annan vårdnadshavare
Du kan få uppehållstillstånd på grund av familjeband om ditt barn bor i Finland.
Barnet måste vara under 18 år gammalt och ogift den dag då beslutet om uppehållstillstånd fattas.
För att få uppehållstillstånd på grund av familjeband måste du vara barnets vårdnadshavare.
Vanligtvis är barnets mor eller far vårdnadshavare.
Vårdnadshavaren kan dock även vara någon annan, till exempel en mor- eller farförälder.
Familjebandet mellan barnet och föräldern måste bevisas till exempel med en födelseattest med föräldrarnas namn.
Om en annan vårdnadshavare än barnets mor eller far ansöker om uppehållstillstånd måste vårdnaden bevisas till exempel genom uppvisande av ett domstolsbeslut.
För att du ska kunna få uppehållstillstånd måste du ha tillräckliga medel för att leva i Finland.
Kravet på tillräcklig inkomst tillämpas dock inte på dig om ditt barn är en finsk medborgare.
Kravet på tillräcklig inkomst tillämpas inte heller om du varit barnets vårdnadshavare redan innan barnet anlänt till Finland och barnet har flyktingstatus i Finland.
Om barnet fått flyktingstatus den 1.7.2016 eller senare, ska du ansöka om uppehållstillstånd inom tre månader från att barnet fått flyktingstatus i Finland.
Ansökan kan även göras senare, men då tillämpas kravet på tillräcklig inkomst.
Vårdnadshavare till en finsk medborgarefinska _ svenska _ engelska
Vårdnadshavare till en utländsk medborgarefinska _ svenska _ engelska
Utkomstförutsättningfinska _ svenska _ engelska
Vårdnadshavare till en person som fått internationellt skyddfinska _ svenska _ engelska
Att ansöka om uppehållstillstånd
Vanligtvis måste du ansöka om ditt första uppehållstillstånd innan du kommer till Finland.
Ansök om tillståndet i ditt hemland eller i ett annat land där du vistas lagligt.
Du kan också ansöka om ditt första visum i Finland, om din familjemedlem är finsk medborgare och du själv är medborgare i ett visumfritt land, det vill säga du inte behöver visum för att komma till Finland.
Du kan ansöka om tillståndet på internet via tjänsten Enter Finland.
När du ställt ansökan ska du besöka Finlands beskickning närmast dig eller Migrationsverkets tjänsteställe för att styrka din identitet och visa upp originalexemplaren av ansökningsbilagorna.
Du ska besöka beskickningen eller tjänstestället inom tre månader efter att ha gjort ansökan på internet.
Ansökningen kan tas för behandling först när du besökt beskickningen eller tjänstestället.
Det är bra att boka en tid hos beskickningen eller tjänstestället i förväg.
Kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan, kommer detta att meddelas via ditt Enter Finland-konto.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du också lämna in en pappersansökan jämte bilagor vid Finlands beskickning närmast dig eller på Migrationsverkets tjänsteställe i Finland.
Du kan skriva ut ansökningsblanketten på Migrationsverkets webbplats.
Ansökan om uppehållstillstånd är avgiftsbelagd.
Avgiften ska betalas då ansökan ställs.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Finlands beskickningar utomlandsfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Finsk personbeteckning
Om du får ett uppehållstillstånd i Finland registreras du automatiskt i det finska befolkningsdatasystemet.
Du får samtidigt även en finsk personbeteckning.
När du har flyttat till Finland ska du besöka magistraten på din hemort för att registrera dig som invånare.
Läs mer på InfoFinlands sida Registrering som invånare.
Uppehållstillstånd för företagare
Uppehållstillstånd för uppstartsföretagare
Att ansöka om uppehållstillstånd
Företagare i Finland
I Finland kan vem som helst med hemvist i ett land som hör till Europeiska ekonomiska samarbetsområdet (EES) starta ett företag.
Behovet av tillstånd är inte beroende av din nationalitet utan din bosättningsort.
Om du är medborgare i ett EU-land, EES-land, nordiskt land eller Schweiz och vill flytta till Finland för att starta ett företag, behöver du inget uppehållstillstånd.
Läs mer på InfoFinlands sida EU-medborgare.
Om du inte har hemvist inom EES och är medborgare i något annat land än ett medlemsland i den Europeiska unionen, ett EES-land eller Schweiz, behöver du ett uppehållstillstånd för att driva ett företag i Finland.
Din företagsverksamhet ska vara lönsam och dina inkomster från företagsverksamheten måste ge dig en tryggad försörjning.
Du måste ansöka om ditt första uppehållstillstånd innan du kommer till Finland.
Uppehållstillstånd för företagare
Om du vill arbeta som företagare i Finland behöver du ett uppehållstillstånd för företagare.
Som företagare betraktas:
Uppstartsföretagare
Privat näringsidkare, som driver en så kallad firma
Bolagsman i ett öppet bolag
Ansvarig bolagsman i kommanditbolag
Medlem i andelslag med obegränsad tillskottsplikt
Delägare som innehar en ledande ställning i ett aktiebolag (verkställande direktör eller styrelsemedlem) eller person som innehar en ledande ställning i någon annan sammanslutning
För att få uppehållstillstånd för företagare måste du själv arbeta i ditt företag i Finland.
Om du inte har hemvist i Finland eller något annat land inom EES, måste du registrera din företagsverksamhet i Patent- och registerstyrelsens handelsregister innan du ansöker om uppehållstillstånd för företagare.
Om du flyttar stadigvarande till Finland eller EES-området behöver du inte Patent- och registerstyrelsens tillstånd för att grunda företaget.
Tillståndet är alltså inte kopplat till din nationalitet utan till var du har din hemvist.
Ansökan om uppehållstillstånd behandlas i två steg.
Först bedömer NTM-centralen (Närings-, trafik- och miljöcentralen) ditt företags lönsamhet bland annat utifrån affärsverksamhetsplanen och finansieringen.
Därefter fattar Migrationsverket beslut om uppehållstillstånd.
På Migrationsverkets webbplats hittar du mer information om villkoren för att ansöka om uppehållstillstånd.
linkkiPatent- och registerstyrelsen:
Tillstånd för företagare som är bosatta utanför EES-områdetfinska _ svenska _ engelska
Uppehållstillstånd för företagarefinska _ svenska _ engelska
Chatbot-tjänst för utländska företagarefinska _ engelska
Uppehållstillstånd för uppstartsföretagare
Om du vill grunda ett uppstartsföretag i Finland kan du ansöka om uppehållstillstånd för uppstartsföretagare som är avsett för tillväxtföretagare.
För att få uppehållstillstånd för uppstartsföretagare måste du ha en konkret affärsverksamhetsplan.
Ansökan om uppehållstillstånd för uppstartsföretagare är indelat i två steg:
Du behöver ett utlåtande från Business Finland som bifaller verksamheten som tillväxtföretagare.
Ansök om uppehållstillstånd för uppstartsföretagare och besök Finlands beskickning eller Migrationsverkets serviceställe för att styrka din identitet.
Processen är mycket snabb och smidig.
Finland som stöder företag bedömer ditt företags affärsmodell, kunnande och förmåga att få verksamheten att växa.
Du kan skicka uppgifterna om din affärsverksamhetsplan och erforderliga handlingar till Business Finland på elektronisk väg.
När du har fått ett positivt utlåtande från Business Finland kan du ansöka om uppehållstillstånd för uppstartsföretagare hos Migrationsverket.
Bifoga utlåtandet till din ansökan om uppehållstillstånd för uppstartsföretagare som du skickar till Migrationsverket.
Du kan inte få uppehållstillstånd för uppstartsföretagare i Finland utan ett positivt utlåtande från Business Finland.
Du hittar anvisningar och mer information om ansökan om uppehållstillstånd för uppstartsföretagare på Migrationsverkets och Business Finlands webbplatser.
Uppehållstillstånd för uppstartsföretagarefinska _ svenska _ engelska
Uppehållstillstånd för uppstartsföretagareengelska
Att ansöka om uppehållstillstånd
Du kan ansöka om uppehållstillstånd för företagare eller uppehållstillstånd för uppstartsföretagare på internet via tjänsten Enter Finland.
När du ställt ansökan ska du besöka Finlands beskickning närmast dig för att styrka din identitet och visa upp originalexemplaren av ansökningsbilagorna.
Du ska besöka beskickningen inom tre månader efter att ha gjort ansökan på internet.
Ansökningen kan tas för behandling först när du har besökt beskickningen.
Vanligtvis måste du boka en tid hos beskickningen i förväg.
Kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan kommer detta att meddelas via ditt konto.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du också lämna in en pappersansökan jämte bilagor vid Finlands beskickning närmast dig.
Du kan skriva ut ansökningsblanketten på Migrationsverkets webbplats.
Handläggning av tillståndsansökan är avgiftsbelagd.
Du betalar avgiften när du lämnar in din tillståndsansökan.
Läs mer om att grunda ett företag på InfoFinlands sida Att grunda ett företag i Finland.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Finsk personbeteckning
Om du får ett uppehållstillstånd i Finland registreras du automatiskt i det finska befolkningsdatasystemet.
Du får samtidigt även en finsk personbeteckning.
När du har flyttat till Finland ska du besöka magistraten på din hemort för att registrera dig som invånare.
Läs mer på InfoFinlands sida Registrering som invånare.
Företagare i Finland
På InfoFinlands sida Arbete och entreprenörskap hittar du mer information avsedd för företagare och arbetstagare.
Guide om att grunda ett företagfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ turkiska _ kinesiska _ arabiska
Tjänster för företagare-Startup Kitengelska
Migrationsverket:Presentation av e-tjänsten Enter Finland
Om du har ett tillfälligt uppehållstillstånd (A- eller B-tillstånd) och orsaken för din vistelse i Finland ändras måste du ansöka om ett nytt uppehållstillstånd på den nya grunden.
Om du har ett permanent uppehållstillstånd (P) i Finland behöver du inte ändra grunden för ditt uppehållstillstånd även om orsaken till din vistelse ändras.
Du kan ansöka om uppehållstillstånd på något av följande grunder:
arbete
studier
familjeband
återflyttning
finländsk härkomst
internationellt skydd
annan orsak
Det är bra att komma ihåg att grunden för uppehållstillståndet kan påverka vilka rättigheter du har i Finland.
Till exempel ger ett uppehållstillstånd på grund av familjeband mer omfattande rätt att arbeta än ett tillstånd som beviljats på grund av studier.
Hur får jag ett tillfälligt uppehållstillstånd ändrat till ett kontinuerligt tillstånd?
Om du har ett tillfälligt uppehållstillstånd (B-tillstånd) kan du ansöka om ett kontinuerligt uppehållstillstånd (A-tillstånd) om grunden för vistelsen i Finland har ändrats från tillfällig till kontinuerlig.
Om du har ett tillfälligt uppehållstillstånd på grund av familjeband kan du ansöka om ett kontinuerligt uppehållstillstånd när en familjemedlem till dig ansöker om ett kontinuerligt uppehållstillstånd.
Du kan ansöka om ett kontinuerligt uppehållstillstånd också på någon annan grund om grunden är kontinuerlig.
Om du har ett tillfälligt uppehållstillstånd på grund av studier kan du få ett kontinuerligt tillstånd endast i det fall att grunden för din vistelse i Finland ändras.
Du kan inte få ett kontinuerligt tillstånd på basis av studier.
Grunden för din vistelse kan ändras till exempel om du får en arbetsplats i Finland eller gifter dig med en finsk medborgare eller en person som har kontinuerligt eller fortsatt tillstånd i Finland.
Om du har ett tillfälligt uppehållstillstånd för arbete eller näringsidkande kan du ansöka om ett kontinuerligt uppehållstillstånd när du har vistats i Finland två år utan avbrott.
Hur söker jag ett uppehållstillstånd på nya grunder?
Välj ansökningsblankett utifrån grunden för din ansökan om nytt tillstånd.
Lämna in din ansökan på internet i tjänsten Enter Finland eller vid Migrationsverkets tjänsteställe.
Mer information om ansökningsproceduren hittar du på InfoFinlands sida Fortsatt uppehållstillstånd.
Från studerande till anställd
Om du har avlagt en examen i Finland kan du få ett uppehållstillstånd för att söka arbete.
När du är klar med dina studier och ditt uppehållstillstånd för studerande går ut, kan du ansöka om fortsatt tillstånd (jatkolupa) för att söka arbete.
Tillståndet är i kraft ett år.
Detta tillstånd kan endast fås en gång och det kan inte förnyas.
När du får en arbetsplats kan du få uppehållstillstånd på grund av arbete.
Uppehållstillstånd på en ny grundfinska _ svenska _ engelska
Uppehållstillstånd för sökande av arbetefinska _ svenska _ engelska
Make/maka till en finsk medborgare
Make/maka till en utländsk medborgare
Make/maka till en flykting
Partner
Att ansöka om uppehållstillstånd
Om maken/makan/sambon/partnern inte får uppehållstillstånd
Make/maka till en finsk medborgare
Om du har ingått äktenskap med en finländsk medborgare som är bosatt i Finland kan du få uppehållstillstånd i Finland på grund av familjeband.
Även en maka/make av samma kön kan få uppehållstillstånd, om ni är gifta eller i ett registrerat parförhållande.
Sambo med en finsk medborgare
Om du är sambo med en finsk medborgare som bor i Finland kan du få uppehållstillstånd på grund av familjeband.
Tillståndet kan beviljas om:
du har bott tillsammans med din sambo minst två år eller
du har ett gemensamt barn med din sambo (då uteblir kravet på gemensamt boende under två års tid) eller
det finns något annat vägande skäl för att bevilja tillståndet
Ifall du ansöker om tillstånd på dessa grunder måste du och din sambo bevisa att ni har bott tillsammans två år.
Som bevis godtas till exempel ett utdrag ur boenderegistret eller ett hyreskontrakt med bådas namn.
Om du och din sambo är bosatta i olika stater anses gemensamt boende till exempel under semesterresor inte som en tillräcklig grund för beviljande av uppehållstillstånd.
Varken du eller din sambo får vara gift med någon annan.
Försörjningsförutsättning för make/maka till en finsk medborgare
Om du är familjemedlem till en finsk medborgare, behöver din försörjning inte vara tryggad.
Du har obegränsad rätt att arbeta.
Du får börja arbeta först när du har fått ett uppehållstillstånd.
Information om hur du ansöker om tillståndet finns under rubriken Att ansöka om uppehållstillstånd.
Make eller maka till en finsk medborgarefinska _ svenska _ engelska
Sambo till en finsk medborgarefinska _ svenska _ engelska
Make/maka till en utländsk medborgare
Även en make/maka av samma kön kan få uppehållstillstånd.
Sambo med en utländsk medborgare
Om din sambo har uppehållstillstånd i Finland och bor i Finland kan du få uppehållstillstånd i Finland på grund av familjeband.
Du kan få tillståndet om:
du har bott tillsammans med din sambo minst två år eller
du har ett gemensamt barn tillsammans med din sambo (då uteblir kravet på gemensamt boende under två års tid)
Ifall du ansöker om tillstånd på dessa grunder måste du och din sambo bevisa att ni har bott tillsammans två år.
Som bevis duger till exempel ett utdrag ur boenderegistret eller ett hyreskontrakt med bådas namn.
Om du och din sambo är bosatta i olika stater anses gemensamt boende till exempel under semesterresor inte som en tillräcklig grund för beviljande av uppehållstillstånd.
Varken du eller din sambo får vara gift med någon annan.
Försörjningsförutsättning för make/maka till en utländsk medborgare
För att du ska få uppehållstillstånd i Finland måste du eller din make/maka ha tillräcklig inkomst även för din försörjning.
På Migrationsverkets sidor kan du kontrollera hur stor inkomst ni måste ha.
Om din maka/make fått uppehållstillstånd på grund av internationellt skydd, tillämpas kravet på tillräcklig inkomst på er.
Det är möjligt att i enskilda fall avvika från försörjningsförutsättningen, om det finns exceptionellt vägande skäl eller om barnets bästa kräver detta.
Information om hur du ansöker om tillståndet finns under rubriken Att ansöka om uppehållstillstånd.
Make eller maka till en utländsk medborgarefinska _ svenska _ engelska
Sambo till en utländsk medborgarefinska _ svenska _ engelska
Utkomstförutsättningfinska _ svenska _ engelska
Make/maka till en flykting
Om din maka/make har uppehållstillstånd i Finland på grund av internationellt skydd och flyktingstatus, kan du få uppehållstillstånd i Finland på grund av familjeband.
Sambo med flykting
Om din sambo har uppehållstillstånd i Finland på grund av internationellt skydd och flyktingstatus, kan du få uppehållstillstånd i Finland på grund av familjeband.
Du kan få tillståndet om:
du har bott tillsammans med din sambo minst två år eller
du har ett gemensamt barn tillsammans med din sambo (då uteblir kravet på gemensamt boende under två års tid)
Ifall du ansöker om tillstånd på dessa grunder måste du och din sambo bevisa att ni har bott tillsammans två år.
Som bevis duger till exempel ett utdrag ur boenderegistret eller ett hyreskontrakt med bådas namn.
Om du och din sambo är bosatta i olika stater anses gemensamt boende till exempel under semesterresor inte som en tillräcklig grund för beviljande av uppehållstillstånd.
Varken du eller din sambo får vara gift med någon annan.
Försörjningsförutsättning för make/maka/sambo/partner till en flykting
Försörjningsförutsättningen tillämpas på er på olika sätt, om din make/maka/sambo/partner har fått uppehållstillstånd på grund av internationellt skydd och har flyktingstatus i Finland.
Din försörjning behöver inte vara tryggad i följande fall:
Om din make/maka/sambo/partner har beviljats asyl eller godkänts som kvotflykting före den 1 juli 2016 och familjen har bildats före hen kom till Finland.
Om din make/maka/sambo/partner har fått flyktingstatus den 1 juli 2016 eller efter detta ska ansökan om uppehållstillstånd lämnas in inom tre månader efter att hen fått beslut på sin ansökan.
De tre månaderna räknas från den dag då din maka/make/sambo/partner delgivits beslutet.
Om du, av anledningar som du inte själv kan påverka, inte hinner ansöka om uppehållstillstånd inom tre månader, kan du ändå ansöka om familjeåterförening.
I din ansökan ska du ange varför tidsfristen på tre månader överskreds.
Du kan ansöka om familjeåterförening även senare, men då tillämpas kravet på tillräcklig inkomst på er.
Försörjningsförutsättningen gäller er även i det fall att ni gifte er efter att din make/maka kom till Finland.
I vissa enskilda fall kan man avvika från försörjningsförutsättningen om det finns exceptionellt vägande skäl eller om barnets bästa kräver detta.
Information om hur du ansöker om tillståndet finns under rubriken Att ansöka om uppehållstillstånd.
Maka eller make till en person som fått internationellt skyddfinska _ svenska _ engelska
Sambo till en person som fått internationellt skyddfinska _ svenska _ engelska
Försörjningsförutsättning för familjemedlemmar till personer som får internationellt skyddfinska _ svenska _ engelska
Partner
Man kan vanligen inte få uppehållstillstånd på grund av sällskapande.
I Finland är en person man sällskapar med inte en familjemedlem enligt lagen.
I vissa fall kan du ändå få ett tillfälligt (B) uppehållstillstånd i Finland på grund av sällskapande.
För att du ska kunna beviljas uppehållstillstånd i Finland måste ditt och din partners förhållande vara stadigt.
Ett bevis på stadigt sällskapande kan till exempel vara att er avsikt är att ingå äktenskap i Finland.
Varken du eller din partner får vara gift med någon annan.
För att du ska kunna få uppehållstillstånd måste du ha tillräckliga medel för ditt uppehälle.
Dessa medel bör vara fritt tillgängliga för dig till exempel på ditt eget bankkonto.
Inkomsterna för din partner som är bosatt i Finland beaktas inte.
Flick- eller pojkvän till en finsk medborgarefinska _ svenska _ engelska
Att ansöka om uppehållstillstånd
Vanligtvis måste du ansöka om ditt första uppehållstillstånd innan du kommer till Finland.
Ansök om tillståndet i ditt hemland eller i ett annat land där du vistas lagligt. Du kan också ansöka om ditt första uppehållstillstånd i Finland om din make eller maka är finsk medborgare och du själv är medborgare i ett visumfritt land, det vill säga du inte behöver visum för att komma till Finland.
Du kan ansöka om tillståndet på internet via tjänsten Enter Finland.
När du ställt ansökan ska du besöka Finlands beskickning närmast dig eller Migrationsverkets tjänsteställe för att styrka din identitet och visa upp originalexemplaren av ansökningsbilagorna.
Du ska besöka beskickningen eller tjänstestället inom tre månader efter att ha gjort ansökan på internet.
Ansökningen kan tas för behandling först när du besökt beskickningen eller tjänstestället.
Vanligtvis måste du boka en tid hos beskickningen eller tjänstestället i förväg.
Kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan, kommer detta att meddelas via ditt Enter Finland-konto.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du också lämna in en pappersansökan jämte bilagor vid Finlands beskickning närmast dig eller på Migrationsverkets tjänsteställe i Finland.
Du kan skriva ut ansökningsblanketten på Migrationsverkets webbplats.
Ansökan om uppehållstillstånd är avgiftsbelagd.
Avgiften ska betalas då ansökan ställs.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Finlands beskickningar utomlandsfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Handläggningstider för tillståndsansökningarfinska _ svenska _ engelska
Finsk personbeteckning
Om du får ett uppehållstillstånd i Finland registreras du automatiskt i det finska befolkningsdatasystemet.
Du får samtidigt även en finsk personbeteckning.
När du har flyttat till Finland ska du besöka magistraten på din hemort för att registrera dig som invånare.
Läs mer på InfoFinlands sida Registrering som invånare.
Om maken/makan/sambon/partnern inte får uppehållstillstånd
En make/maka/sambo/partner beviljas inte uppehållstillstånd om förutsättningarna för uppehållstillstånd inte uppfylls.
Man kan låta bli att bevilja tillståndet även då de finländska myndigheterna anser att parterna har ingått äktenskap endast för uppehållstillståndets skull och att makarna inte avser att leva tillsammans som en familj.
Myndigheterna kan misstänka att parterna ingått äktenskap endast för uppehållstillståndets skull till exempel om ni har ingått äktenskap efter endast en kort bekantskap, om det är stor åldersskillnad mellan er eller om den ena av er har haft flera korta äktenskap.
Om du får ett nekande beslut på din tillståndsansökan kan du överklaga den till förvaltningsdomstolen.
Du får instruktioner för detta bifogade till tillståndsbeslutet.
Läs mer om problem med uppehållstillståndet på InfoFinlands sida Problem med uppehållstillståndet.
Uppehållstillstånd för arbetstagare
Andra uppehållstillstånd för förvärvsarbete
Uppehållstillstånd för säsongsarbete
Arbete med ett annat uppehållstillstånd
Ansökan om uppehållstillstånd
Arbete utan uppehållstillstånd
Arbetstagare i Finland
Den här sidan är avsedd för dig som är medborgare i något annat land är ett EU-land, Norge, Island, Schweiz eller Liechtenstein.
Om du kommer till Finland för att arbeta behöver du ett uppehållstillstånd.
Innan du kan få ett uppehållstillstånd måste du hitta ett jobb i Finland.
När du har hittat ett jobb kan du ansöka om uppehållstillstånd.
Du måste ansöka om uppehållstillstånd innan du kommer till Finland.
För att kunna arbeta i Finland behöver du vanligen antingen ett uppehållstillstånd för arbetstagare eller någon annan typ av uppehållstillstånd för förvärvsarbete.
Arten av det arbete du ska utföra påverkar typen av tillstånd.
Uppehållstillstånd för arbetstagare
Om du inte kan arbeta med stöd av ett annat uppehållstillstånd eller utan uppehållstillstånd behöver du ett uppehållstillstånd för arbetstagare (työntekijän oleskelulupa).
Uppehållstillstånd för arbetstagare är inte nödvändigt för alla arbetsuppgifter.
Du kan granska hurudant uppehållstillstånd du behöver från Migrationsverkets webbplats.
Du behöver uppehållstillstånd för arbetstagare om du arbetar till exempel som:
städare
hemvårdare eller barnskötare.
Migrationsverket beslutar om du ska beviljas uppehållstillstånd eller inte.
Ett delbeslut av arbets- och näringsbyrån behövs också för tillståndet.
Uppehållstillstånd för arbetstagarefinska _ svenska _ engelska
Andra uppehållstillstånd för förvärvsarbete
För vissa arbetsuppgifter behöver du inte ett uppehållstillstånd för arbetstagare, men du behöver dock ett uppehållstillstånd som beviljas för vissa uppdrag.
Dessa uppdrag kan vara till exempel:
uppdrag inom företagsledning
uppdrag som sakkunnig
forskaruppdrag
uppdrag inom vetenskap, kultur och konst
arbetspraktik.
Migrationsverket beslutar om du får uppehållstillstånd eller inte.
Ett delbeslut av arbets- och näringsbyrån behövs inte för tillståndet.
Arbete i Finlandfinska _ svenska _ engelska
Uppehållstillstånd för säsongsarbete
Om du ska utföra säsongsarbete i Finland behöver du ett säsongsarbetstillstånd.
Säsongsarbetet kan pågå högst nio månader.
Säsongsarbete är till exempel:
växtodling
skogsvårdsarbete
festivalarbete
Om du kommer från ett viseringspliktigt land och ska arbeta i under tre månader, måste du ansöka om ett säsongsarbetsvisum hos den finländska beskickningen.
Om ditt arbete pågår över tre månader ska du ansöka om ett säsongsarbetstillstånd hos Migrationsverket.
Tillstånd för säsongsarbetefinska _ svenska _ engelska
Arbete med ett annat uppehållstillstånd
Om du redan har uppehållstillstånd i Finland utifrån en annan grund, till exempel familjeband, kan du ha rätt att arbeta i Finland.
Då behöver du inte ett separat uppehållstillstånd för att arbeta.
Du kan kontrollera om du har rätt att arbeta i Finland från ditt uppehållstillståndskort eller beslut om uppehållstillstånd.
Rätt att arbetafinska _ svenska _ engelska
Om du har avlagt examen i Finland kan du få ett tillfälligt uppehållstillstånd för att söka arbete.
Detta tillstånd kan beviljas endast som ett fortsatt tillstånd till ett uppehållstillstånd för studerande.
Ansök om tillståndet innan ditt uppehållstillstånd för studerande löper ut.
Du kan få ett tillstånd för högst ett år.
Detta tillstånd kan man endast få en gång.
Om du hittar en arbetsplats, kan du börja arbeta genast.
Du måste ansöka om ett nytt uppehållstillstånd på grund av arbete innan ditt uppehållstillstånd för att söka arbete går ut.
Om du har avlagt examen i Finland, behövs inte ett delbeslut av arbets- och näringsbyrån för ditt tillstånd.
Uppehållstillstånd för sökande av arbetefinska _ svenska _ engelska
Ansökan om uppehållstillstånd
Du måste ansöka om ditt första uppehållstillstånd innan du kommer till Finland.
Du kan ansöka om tillståndet på internet via tjänsten Enter Finland.
När du ställt ansökan ska du besöka Finlands beskickning närmast dig för att styrka din identitet och visa upp originalexemplaren av ansökningsbilagorna.
Du ska besöka beskickningen inom tre månader efter att ha gjort ansökan på internet.
Ansökningen kan tas för behandling först när du besökt beskickningen.
Vanligtvis måste du boka en tid hos beskickningen i förväg.
Kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan kommer detta att meddelas via ditt konto.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du också lämna in en pappersansökan jämte bilagor vid Finlands beskickning närmast dig.
Du kan skriva ut ansökningsblanketten på Migrationsverkets webbplats.
Handläggningen av din ansökan om tillstånd är avgiftsbelagd.
Du måste betala avgiften när du lämnar in ansökan om uppehållstillstånd.
Till ansökan om uppehållstillstånd för arbetstagare ska du bifoga blanketten TEM054 som din arbetsgivare fyller i och undertecknar.
Arbetsgivaren kan lämna uppgifterna om arbetet och sitt företag själv samt följa handläggning av ansökan direkt via tjänsten Enter Finland.
Arbetsgivaren kan även betala handläggningsavgiften för arbetstagaren.
Fråga din arbetsgivare som hen använder tjänsten Enter Finland för arbetsgivare.
Kom ändå ihåg att arbetsgivaren inte kan ansöka om uppehållstillstånd för dig, utan hen kompletterar din ansökan för egen del i tjänsten Enter Finland.
Så länge handläggningen av din första ansökan om uppehållstillstånd pågår har du inte rätt att arbeta.
Om du har ansökt om uppehållstillstånd utomlands, kan du inte komma till Finland innan tillstånd har beviljats.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Handläggningstider för tillståndsansökningarfinska _ svenska _ engelska
Ansökan om uppehållstillstånd för specialist
Om du ska arbeta i Finland som specialist kan du även komma till Finland utan uppehållstillstånd.
Du måste dock ha visum eller rätt att vistas i Finland tre månader utan visum.
Du ska också ha en arbetsplats som uppfyller kraven.
Om du arbetar i Finland längre än tre månader måste du ansöka om uppehållstillstånd.
Du kan ansöka om tillståndet elektroniskt via tjänsten Enter Finland eller på Migrationsverkets tjänsteställe.
Finsk personbeteckning
Om du får ett uppehållstillstånd i Finland registreras du automatiskt i det finska befolkningsdatasystemet.
Du får samtidigt även en finsk personbeteckning.
När du har flyttat till Finland ska du besöka magistraten på din hemort för att registrera dig som invånare.
Läs mer på InfoFinlands sida Registrering som invånare.
Arbete utan uppehållstillstånd
Oberoende av vilket land du är medborgare i kan du i vissa fall arbeta i Finland utan uppehållstillstånd.
Du måste dock ha ett visum, om du behöver visum till Finland.
Du kan arbeta i Finland utan uppehållstillstånd till exempel om:
du kommer till Finland för att arbeta som tolk, lärare, sakkunnig eller idrottsdomare i högst tre månader utifrån en inbjudan eller ett avtal;
du är fast anställd vid ett företag som bedriver verksamhet i ett annat EU/EES-land och ska komma till Finland för att utföra tillfälligt leverans- eller underleveransarbete och ditt arbete pågår högst tre månader;
du är asylsökande i Finland och har ett giltigt resedokument som berättigar till gränsövergång.
Trots att du inte har uppehållstillstånd kan du börja arbeta tre månader efter att du har lämnat in din asylansökan;
du är asylsökande i Finland och har inte ett giltigt resedokument som berättigar till gränsövergång.
Trots att du inte har uppehållstillstånd kan du börja arbeta när du vistats i sex månader i landet.
Du kan granska om du har rätt att arbeta i Finland utan uppehållstillstånd från Migrationsverkets webbplats.
Arbete utan uppehållstillståndfinska _ svenska _ engelska
Arbetstagare i Finland
På InfoFinlands sida Var hittar jag jobb? finns information om hur du kan hitta ett jobb i Finland.
InfoFinlands sidor Arbete och entreprenörskap innehåller mer information för arbetstagare och företagare.
linkkiArbets- och näringsministeriet:
Arbeta i Finlandfinska _ svenska _ engelska
linkkiArbets- och näringsbyrån:
Broschyren Jobba i Finland(pdf, 5,51 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ polska
linkkiArbetshälsoinstitutet:
Handboken Jobba i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ kurdiska _ tyska _ thai _ vietnamesiska
Migrationsverket:
Presentation av e-tjänsten Enter Finland
Det är viktigt att du ansöker om fortsatt uppehållstillstånd innan ditt tidigare uppehållstillstånd går ut.
Om ditt tidigare uppehållstillstånd går ut under behandlingen av ansökan får du uppehålla dig i Finland och har vanligtvis även rätt att arbeta under den tid som ansökan behandlas.
Om du ansöker om fortsatt uppehållstillstånd först efter att ditt tidigare uppehållstillstånd gått ut, får du uppehålla dig i Finland under tiden då ansökan behandlas men har inte rätt att arbeta innan du erhållit fortsatt uppehållstillstånd.
Att ansöka
Du kan ansöka om tillståndet på internet i tjänsten Enter Finland.
När du ställt ansökan ska du besöka Migrationsverkets tjänsteställe för att styrka din identitet.
Du ska besöka tjänstestället inom tre månader efter att ha gjort ansökan.
Ta med dig pass, passfoto och originalexemplaren av ansökningsbilagorna.
Det är bra att boka en tid hos Migrationsverkets tjänsteställe i förväg.
Du kan boka tiden via Migrationsverkets elektroniska tidsbokningssystem.
Om du gjort ansökningen på internet, kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan, kommer detta att meddelas via ditt Enter Finland-konto.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du ansöka om tillståndet med en pappersblankett vid Migrationsverkets tjänsteställe.
Skriv ut blanketten på Migrationsverkets webbplats och fyll i den färdigt.
Boka en tid vid tjänstestället.
När du ska besöka tjänstestället, ta med dig din ifyllda ansökan, bilagorna och kopior på bilagor samt pass och passfoto.
Migrationsverket beviljar dig fortsatt uppehållstillstånd om grunden för det tidigare uppehållstillståndet fortfarande existerar.
Du kan även ansöka om fortsatt uppehållstillstånd på annan grund än för det tidigare tillståndet
Hanteringen av ansökan är avgiftsbelagd. Avgiften ska betalas då ansökan görs.
I tjänsten Enter Finland kan du betala med nätbankskoderna för en finsk bank eller med kreditkort.
Att förlänga uppehållstillståndetfinska _ svenska _ engelska
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Blanketter för ansökan om uppehållstillståndfinska _ svenska _ engelska
Migrationsverket:
Presentation av e-tjänsten Enter Finland
Om du vill flytta till en familjemedlem som bor i Finland behöver du ett uppehållstillstånd.
Om du bara vill hälsa på hos din familjemedlem i Finland hittar du mer information på InfoFinlands sida Kort vistelse i Finland.
Alla familjemedlemmar kan inte få uppehållstillstånd.
Vanligen kan man få tillstånd om man är make/maka, sambo, minderårigt barn eller förälder till minderårigt barn till personen bosatt i Finland.
Ofta krävs det även att personen bosatt i Finland ska ha tillräckliga medel för att försörja en familjemedlem som flyttar till Finland.
Notera att separata regler gäller för familjemedlemmar till EU-medborgare (inte finländska medborgare).
Om du är familjemedlem till en EU-medborgare bosatt i Finland hittar du mer information om tillståndsärenden på InfoFinlands sidan EU-medborgare.
Mer information om hur familjemedlemmar kan få uppehållstillstånd finns på InfoFinlands sidor Uppehållstillstånd för make eller maka, Uppehållstillstånd för barn eller förälder, Uppehållstillstånd för övriga anhöriga.
På InfoFinlands sida Familjemedlem hittar du mer information avsedd för personer som flyttar av familjeskäl.
Till Finland på grund av familjebandfinska _ svenska _ engelska
Hur ansöker jag?
Vad behövs för registreringen?
Kan jag bli av med uppehållsrätten?
Registrering av uppehållsrätten för EU-medborgare sker inte per automatik.
Du kan ansöka om registrering av uppehållsrätten om din försörjning i Finland är tryggad.
Den kan vara baserad på ett jobb, studier, företagsverksamhet, familjeband eller tillräckliga medel.
Om du avser att bo i Finland längre än tre månader, måste du registrera din uppehållsrätt hos Migrationsverket (Maahanmuuttovirasto).
Ansökan ska lämnas in senast inom tre månader från datumet för inresa.
Registreringen hos Migrationsverket är inte samma sak som registreringen av din bosättningsort i befolkningsdatasystemet (väestötietojärjestelmä) vid magistraten (maistraatti).
Om din sammanhängande vistelse i Finland är kortare än tre månader behöver du inte registrera vistelsen vid Migrationsverket.
Vistelsetiden på tre månader räknas alltid från det att du varit utanför Finlands gränser.
Läs mer om förutsättningarna på sidan EU-medborgare.
Hur ansöker jag?
Handläggning av ansökan om registrering av uppehållsrätt är avgiftsbelagd.
Du betalar avgiften när du lämnar in din ansökan.
Ansök om registrering av uppehållsrätten för EU-medborgare i tjänsten Enter Finland:
Fyll i ansökningsblanketten och bifoga erforderliga bilagor.
Du hittar information om vilka bilagor som behövs till ansökningen i avsnittet
Vad behövs för registreringen?
Besök Migrationsverkets tjänsteställe; du måste styrka din identitet och visa upp originalexemplaren av ansökningsbilagorna.
Ta med dig ett giltigt ID-kort eller pass.
Du ska besöka tjänstestället inom tre månader efter att ha gjort ansökan.
Det är bra att boka en tid på tjänstestället i förväg.
Boka tiden via Migrationsverkets elektroniska tidsbokningssystem.
Kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan, kommer detta att meddelas via ditt Enter Finland-konto.
Du får också ett meddelande när beslutet är klart.
Om du inte kan eller inte vet hur du ska göra ansökan på internet:
Gör registreringsansökan på en pappersblankett.
Du kan även göra det personligen på Migrationsverkets tjänsteställe.
Gör ansökan inom tre månader efter datumet för inresa.
Skriv ut registreringsblanketten på Migrationsverkets webbplats och fyll i den färdigt.
Var noga när du fyller i ansökan.
Felaktigt ifyllda ansökningar tas inte emot.
Boka en tid på Migrationsverkets tjänsteställe i det elektroniska tidsbokningssystemet.
Det är bra att boka en tid på tjänstestället i förväg.
Ta med dig den ifyllda registreringsblanketten, ett giltigt ID-kort eller pass och erforderliga bilagor.
Du hittar information om vilka bilagor som behövs till ansökningen i avsnittet
Vad behövs för registreringen?
Om kraven på grund och förutsättningar för vistelsen Finland uppfylls, kan du få ett intyg över registrering av uppehållsrätten för medborgare i Europeiska unionen från Migrationsverket.
Registreringen av uppehållsrätten gäller tillsvidare.
När du har bott lagligt och utan avbrott i Finland i fem år, har du permanent uppehållsrätt.
Permanent uppehållsrätt för EU-medborgare ansöks separat från Migrationsverket.
Registrering av uppehållsrätt för EU-medborgarefinska _ svenska _ engelska
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Permanent uppehållstillståndfinska _ svenska _ engelska
Om magistraten registrerar din uppehållsrätt, registreras dina personuppgifter automatiskt även i befolkningsdatasystemet.
Du får samtidigt även en finsk personbeteckning.
Du kan få en finsk personbeteckning även vid magistraten eller skattebyrån på din hemort.
Om du flyttar till Finland för att bo här stadigvarande i ett år eller längre, ska du också registrera dig i magistraten på din hemort.
Läs mer på InfoFinlands sida Registrering som invånare.
På InfoFinlands sida Komihåglista för dig som flyttar till Finland hittar du nyttig information om allt som du ska ta hand om när du flyttar till Finland.
Vad behövs för registreringen?
Arbetstagare eller företagare
Din uppehållsrätt kan registreras om du är anställd eller har ett eget företag i Finland.
Du behöver följande handlingar:
EU-registreringsblankett
Giltigt ID-kort eller pass
Anställningsavtal (om du är anställd)
En utredning över företagsverksamheten (om du är egenföretagare)
Studerande
Din uppehållsrätt kan registreras om du studerar vid en läroanstalt som är godkänd i Finland.
Du behöver följande handlingar:
EU-registreringsblankett
Giltigt ID-kort eller pass
Närvarointyg (intyg över att du är studerande vid en läroanstalt som är godkänd i Finland)
Du har en sjukförsäkring (t.ex. det europeiska sjukvårdskortet)
En utredning över din försörjning i Finland
Familjemedlem till en person bosatt i Finland
Din uppehållsrätt kan registreras om du har en familjemedlem som är stadigvarande bosatt i Finland.
Du behöver följande handlingar:
EU-registreringsblankett
Giltigt ID-kort eller pass
Intyg över äktenskap eller registrerat parförhållande
En utredning över att ni har bott tillsammans i två år eller har gemensam vårdnad om ett barn, om du är i ett samboförhållande
Barnets födelseattest om du har vårdnaden om ett barn
En utredning över grunden för att den person som ansöker om familjeförening vistas i Finland.
Om du inte själv är medborgare i ett EU-land, Liechtenstein eller Schweiz men avser att flytta till Finland till en familjemedlem som är EU-medborgare, måste du ansöka om uppehållskort för en familjemedlem till en EU-medborgare.
Du kan ansöka om uppehållskortet elektroniskt via tjänsten Enter Finland eller på Migrationsverkets (Maahanmuuttovirasto) tjänsteställe.
Handläggning av ansökan om uppehållskort är avgiftsbelagd.
Du betalar avgiften när du lämnar in din ansökan.
Du behöver följande handlingar:
Ansökan om uppehållskort
Giltigt pass
Intyg över äktenskap eller registrerat parförhållande
Registreringsintyget för den EU-medborgare, med vem du kommer till Finland
Utredning över släktskapsförhållandet (barn till EU-medborgaren eller andra släktingar som står under dennes vårdnad)
Utredning över samboskap (om du är sambo med EU-medborgaren och ni inte har gemensam vårdnad om barn)
Uppehållskortet för en familjemedlem till en EU-medborgare beviljas för fem år eller en kortare tid om boendet i Finland varar mindre än fem år.
Uppehållskort för EU-medborgares familjemedlemfinska _ svenska _ engelska
Tillräckliga medel
Om din uppehållsrätt inte kan registreras på någon av de ovan nämnda grunderna kan du ansöka om registrering om du har tillräckliga medel för din försörjning i Finland.
Också tillräckliga medel är en grund.
Du behöver följande handlingar:
EU-registreringsblankett
Giltigt ID-kort eller pass
En utredning över att du har tillräckliga medel för din försörjning i Finland.
Kan jag bli av med uppehållsrätten?
Registreringen av uppehållsrätten för en EU-medborgare och uppehållskortet för en familjemedlem till en EU-medborgare kan återkallas eller bli ogiltigt om:
du flyttar permanent från Finland
du har vistats utomlands utan avbrott i två år
du lämnade felaktiga uppgifter när du ansökte om registreringen eller om uppehållskortet för en familjemedlem till en EU-medborgare
du har undanhållit sådan information som skulle kunna ha hindrat dig från att få registreringen eller uppehållskortet
du utvisas från Finland
du får finskt medborgarskap.
Tänk på att ändringar i din livssituation kan påverka din uppehållsrätt.
Om din uppehållsrätt registrerades på basis av arbete, ett aktivt företag, en studieplats, familjeband eller tillräckliga medel, och detta skäl inte längre existerar, kan registreringen återkallas.
Beslut om återkallande eller upphörande av uppehållsrätten fattas av Migrationsverket.
Om du flyttar utomlands
Om du inte vill att ditt uppehållstillstånd eller uppehållskort ska återkallas ska du lämna in en ansökan om detta hos Migrationsverket senast inom två år efter att du har flyttat utomlands.
Återkallande av uppehållsrättfinska _ svenska _ engelska
Finland tillhör Schengenområdet.
Länderna som tillhör Schengenområdet har enhetlig visering.
Utlänningar som vill resa till Finland för en kort tid, till exempel på semester, affärsresa eller på besök hos släktingar, behöver ett visum om de inte är medborgare i ett viseringsfritt land.
Ett visum är ett inresetillstånd för en kortvarig och tillfällig, högst tre månader lång vistelse.
På utrikesministeriets webbplats eller vid den närmast belägna finländska beskickningen kan du kontrollera om du behöver ett visum i Schengenområdet.
Visumbehovet till Schengenområdet och av Finland accepterade resedokumentfinska _ svenska _ engelska
Information för viseringsfria personer
Du kan resa till Finland och de övriga Schengenländerna om du har ett giltigt pass eller något annat resedokument som godkänns i Finland.
Du får vistas högst tre månader under en period på sex månader i Finland och de övriga Schengenländerna räknat från den dag du reste in till Schengenområdet.
Information för viseringsskyldiga personer
Du ska alltid ha ett visum när du kommer till Finland eller något annat land i Schengenområdet.
Du får vistas i Finland eller något annat land i Schengenområdet utan uppehållstillstånd så länge som ditt visum är i kraft.
Om du har ett visum eller uppehållstillstånd i något Schengenland kan du resa inom Schengenområdet utan att behöva skaffa ett separat visum för de andra Schengenländerna.
Så här ansöker du om Schengenvisum
Du ansöker om visum i den närmast belägna finländska beskickningen eller visumcentralen.
Du ska vistas lagligt i det land där du ansöker om visum.
I länder där Finland inte har en beskickning kan något annat land representera Finland i visumärenden.
I detta fall kan du ansöka om visum i detta lands beskickning.
På utrikesministeriets webbplats finns en förteckning över de länder där ett annat land representerar Finland i visumärenden.
Du ansöker om visum med en visumansökningsblankett.
Blanketten får du på utrikesministeriets webbplats och från beskickningar i Schengenländer.
Antalet bilagor som krävs till visumansökan kan variera beroende på i vilket land du söker visum.
Hos beskickningen kan du kontrollera vilka bilagor du behöver för din visumansökan.
Lämna din ansökning till den beskickning eller visumcentral dit du ställer din ansökan.
Du kan inte skicka din ansökning via e-post eller fax.
Förlängning av visum i Finland
Polisen kan förlänga uppehållstiden för ditt visum eller visumets utgångstid om du av motiverade skäl inte kan lämna Finland när ditt visum utgår.
Motiverade skäl för förlängning av visum kan till exempel vara:
en akut, svår sjukdom som hindrar dig från att resa,
en släkting som är bosatt i Finland har plötsligt insjuknat svårt eller avlidit,
inställt flyg på grund av strejk eller väderförhållanden,
viktiga affärsförhandlingar som pågår längre än väntat.
Information till medborgare från viseringsskyldiga länderfinska _ svenska _ engelska
Ansökan om Schengenvisumfinska _ svenska _ engelska
Länder där en annan Schengenstat representerar Finlandfinska _ svenska _ engelska
Förlängning av visum i Finlandfinska _ svenska _ engelska
Hjälp i nödsituationer
Beskickningarna hjälper sitt lands medborgare som hamnat i nödläge i Finland.
De kan till exempel hjälpa dig om du har råkat ut för en olycka, blivit sjuk eller fallit offer för ett brott.
Beskickningen kan bevilja dig ett nytt pass om ditt pass har gått förlorat eller stulits.
Om du är turist i Finland och hamnar i en svår situation, ska du kontakta ditt hemlands beskickning.
linkkiVisitFinland.com:
Information om Finland till turistersvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ japanska _ italienska
Ansök om studieplats
Teckna en tillräckligt omfattande sjukförsäkring i ditt hemland
Reservera tillräckliga medel för din försörjning
Ansök om uppehållstillstånd för studerande
Uppehållstillstånd för studerande från andra EU-länder
Fortsatt uppehållstillstånd för studerande
När du avslutar dina studier
För praktik till Finland
Den här sidan är avsedd för dig som är medborgare i något annat land än ett EU-land, Norge, Island, Schweiz eller Liechtenstein.
Om du ska studera i Finland längre än 90 dagar behöver du ett uppehållstillstånd på grund av studier.
Du kan studera mindre än 90 dagar i Finland utan uppehållstillstånd.
Om du ska flytta till Finland för studier måste du ta hand om följande:
Ansök om studieplats
Innan du kan ansöka om uppehållstillstånd måste du skaffa dig en studieplats i Finland.
Godkända läroanstalter är läroanstalter efter grundskolan, till exempel universitet, högskolor och yrkesläroanstalter.
Studieplatsen ska uppfylla ett av följande villkor:
studierna leder till yrke eller examen
du deltar i ett utbytesprogram mellan läroanstalter eller något annat utbytesprogram
du avlägger en kompletterande utbildning eller en specialutbildning som hör till din examen.
Du kan ansöka om studieplats i skolornas gemensamma ansökan på våren eller hösten.
Till vissa utbildningar är den gemensamma ansökan (yhteishaku) redan i januari.
Ta i god tid reda på när du kan ansöka om en studieplats.
Fyll i ansökan i tjänsten Opintopolku.fi.
På InfoFinlands sida Ansökan till utbildning hittar du mer information om hur du ansöker om en studieplats i Finland.
Teckna en tillräckligt omfattande sjukförsäkring i ditt hemland
Som studerande betalar du själv vårdkostnaderna om du insjuknar i Finland.
För ditt uppehållstillstånd behöver du en privat försäkring som täcker kostnaderna för sjukdom och läkemedel.
Du kan teckna en försäkring hos ett försäkringsbolag i ditt hemland eller fråga om en lämplig försäkring hos internationella försäkringsbolag.
Alla försäkringar ska uppfylla följande villkor:
Försäkringens självrisk får inte överstiga 300 euro.
Försäkringen ska gälla under hela din vistelse i Finland.
Försäkringen ska gälla när du kommer till Finland.
Försäkringen får inte vara en vanlig reseförsäkring.
Säg inte upp din försäkring.
Om du insjuknar måste du själv betala läkar- och sjukhuskostnaderna.
Hur stora vårdkostnader som försäkringen måste täcka beror på hur länge dina studier varar.
Om dina studier i Finland till exempel varar mindre än två år, ska försäkringen täcka sjukvårdskostnader upp till minst 120 000 euro.
Om du har det europeiska sjukvårdskortet (European Health Insurance Card, EHIC), behöver du ingen separat försäkring.
Sjukvårdskortet ska vara giltigt under hela din vistelse i Finland.
Försäkring för studerandefinska _ svenska _ engelska
Reservera tillräckliga medel för din försörjning
Du måste också själv ansvara för levnadskostnaderna i Finland.
Du behöver ha minst 560 euro disponibla medel i månaden för att kunna betala för boende, mat och andra utgifter.
För en vistelse som varar ett år ska du alltså ha 6 720 euro i disponibla medel.
Försörjningsförutsättningen kan i vissa fall undgås.
Om till exempel läroanstalten ordnar dig en gratis bostad och även gratis måltider behöver du ha en mindre summa i disponibla medel.
Om studierna är avgiftsbelagda måste du även se till att du har tillräckliga medel för din försörjning efter att du har betalat läsårsavgiften.
Beloppet som krävs ska finnas på ditt bankkonto eller också ska du ha ett intyg över ett stipendium som beviljats av en officiell instans.
Sådana stipendier är till exempel de som beviljats av staten, läroanstalter eller organisationer.
Sponsringslöften eller kontoutdrag från privatpersoner, såsom släktingar, bekanta eller arbetsgivare, godkänns inte.
Försörjningsförutsättning för studerandefinska _ svenska _ engelska
Ansök om uppehållstillstånd för studerande
Du måste ansöka om ditt första uppehållstillstånd innan du kommer till Finland.
Du kan ansöka om tillståndet på internet via tjänsten Enter Finland.
När du ställt ansökan ska du besöka Finlands beskickning närmast dig för att styrka din identitet och visa upp originalexemplaren av ansökningsbilagorna.
Du ska besöka beskickningen inom tre månader efter att ha gjort ansökan på internet.
Ansökningen kan tas för behandling först när du besökt beskickningen.
Vanligtvis måste du boka en tid hos beskickningen i förväg.
Kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan kommer detta att meddelas via ditt konto.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du också lämna in en pappersansökan jämte bilagor vid Finlands beskickning närmast dig.
Du kan skriva ut ansökningsblanketten på Migrationsverkets webbplats.
Handläggningen av ansökan är avgiftsbelagd.
Du måste betala avgiften när du lämnar in ansökan om uppehållstillstånd.
Du ska bifoga följande handlingar till din ansökan om uppehållstillstånd för studerande:
Giltigt pass
Passfoto (anvisningar för fotot finns på Migrationsverkets webbplats)
Närvarointyg (intyg över att du är studerande vid en läroanstalt som är godkänd i Finland)
En utredning över att du har tillräckliga medel för din försörjning
Ett försäkringsintyg eller en kopia av det europeiska sjukvårdskortet
En utredning över att du har betalat läsårsavgiften eller har ett stipendium
Tidigare examensbetyg (om du inte ska avlägga examen eller är en utbytesstudent)
Eventuella arbetsintyg (om du inte ska avlägga examen eller är en utbytesstudent)
Information om uppehållstillstånd för studierfinska _ svenska _ engelska
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Finlands beskickningar utomlandsfinska _ svenska _ engelska
Uppehållstillstånd för studerande från andra EU-länder
Du behöver inget uppehållstillstånd i Finland om du har ett uppehållstillstånd som beviljats i ett annat EU-land och om du studerar vid en högskola.
Dessutom måste dina studier:
innefatta internationell rörlighet i ett EU-program eller ett mångformigt program eller
omfattas av ett avtal mellan två eller fler högskolor.
I detta fall måste du göra en underrättelse om rörlighet till Migrationsverket.
Du får studera i Finland högst 360 dagar när du gör en underrättelse om rörlighet.
Underrättelse om rörlighet i Finlandfinska _ svenska _ engelska
Finsk personbeteckning
Om du får ett uppehållstillstånd i Finland registreras du automatiskt i det finska befolkningsdatasystemet.
Du får samtidigt även en finsk personbeteckning.
När du har flyttat till Finland ska du besöka magistraten på din hemort för att registrera dig som invånare.
Läs mer på InfoFinlands sida Registrering som invånare.
Fortsatt uppehållstillstånd för studerande
Uppehållstillstånd för studerande beviljas högst för två år i taget.
Om dina studier fortsätter men uppehållstillståndet håller på att gå ut ska du ansöka om fortsatt uppehållstillstånd.
Kom ihåg att ansöka om fortsatt uppehållstillstånd för studerande i god tid innan giltighetstiden för det första tillståndet går ut.
Observera att Migrationsverket (Maahanmuuttovirasto) även kontrollerar om grunden för din vistelse i Finland verkligen har varit studier.
Om du till exempel avlägger en grundexamen vid universitet, högskola eller yrkeshögskola bör du avlägga 45 studiepoäng under ett läsår för att uppfylla villkoren för fortsatt uppehållstillstånd.
Du ska bifoga ett studieregisterutdrag till din ansökan om fortsatt uppehållstillstånd.
Fortsatt uppehållstillstånd för studerandefinska _ svenska _ engelska
När du avslutar dina studier
Om du har avlagt en examen i Finland kan du få ett tillfälligt uppehållstillstånd för arbetssökande.
Detta tillstånd kan beviljas endast som ett fortsatt tillstånd till ett uppehållstillstånd för studerande.
Du ska ansöka om tillståndet innan ditt uppehållstillstånd för studerande går ut.
Uppehållstillstånd för arbetssökande kan beviljas för högst ett år.
Om du får ett jobb kan du börja arbeta direkt.
Du måste ansöka om ett nytt uppehållstillstånd på grund av arbete innan ditt uppehållstillstånd för arbetssökande går ut.
Uppehållstillstånd för sökande av arbetefinska _ svenska _ engelska
Till Finland som praktikant
Om du studerar utomlands och vill komma till Finland för arbetspraktik behöver du ett uppehållstillstånd på grund av praktik.
Mer information hittar du på Migrationsverkets webbplats.
Praktik i Finlandfinska _ svenska _ engelska
InfoFinlands sida Utländska studerande i Finland innehåller viktig information om studielivet i Finland.
Information för utländska studerandeengelska
Migrationsverket:
Presentation av e-tjänsten Enter Finland
Arbeta i Finland
Till Finland som företagare
Att studera i Finland
Till familjemedlem i Finland
Kort vistelse i Finland
Om du är medborgare i ett EU-land, Liechtenstein eller Schweiz, behöver du inget uppehållstillstånd eller visum i Finland.
Du kan resa till Finland om du har ett giltigt ID-kort eller pass.
Du har rätt att arbeta, driva ett företag och studera i Finland med lika villkor som finska medborgare.
Du måste själv trygga din försörjning i Finland.
Som EU-medborgare kan du vistas i Finland högst tre månader i sträck utan att registrera din uppehållsrätt.
Om du vill stanna kvar i Finland och registrera dig som invånare, ska du ha ett jobb eller ett aktivt företag, en studieplats, ett långvarigt familjeband eller tillräckliga medel.
Om du avser att bo i Finland i över tre månader, ska du ansöka om Registrering av uppehållsrätten för EU-medborgare hos Migrationsverket.
Ansökan ska ställas senast inom tre månader från datumet för inresa.
Om du flyttar till Finland för att bo här stadigvarande i ett år eller längre, ska du också registrera dig i magistraten på din hemort.
Läs mer på InfoFinlands sida Registrering som invånare.
Om du vistas i Finland tre månader utan avbrott behöver du inte ansöka om registrering av uppehållsrätten.
Vistelsetiden på tre månader räknas alltid från det att du varit utanför Finlands gränser.
linkkiEuropa.eu:
EU-länderfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Rådgivning för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropeiska kommissionen:
Europeiska sjukvårdskortetfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Arbeta i Finland
Som EU-medborgare behöver du inget arbetstillstånd i Finland.
Du kan börja jobba direkt när du har kommit till landet.
Hämta ett skattekort på den närmaste skattebyrån (Verotoimisto) och lämna kortet till din arbetsgivare.
Om du ska jobba i Finland i mer än tre månader ska du ansöka om registrering av uppehållsrätten för EU-medborgare i tjänsten Enter Finland eller på Migrationsverkets (Maahanmuuttovirasto) tjänsteställe.
Om du flyttar till Finland för att bo här stadigvarande i minst ett år ska du också registrera dig som invånare i magistraten (maistraatti).
Personbeteckning
Om du kommer till Finland från utlandet för att arbeta, behöver du en finsk personbeteckning.
Du får personbeteckningen på magistraten (maistraatti) eller skattebyrån (verotoimisto).
Ett giltigt ID-kort eller pass
Ditt anställningsavtal
Du kan även få en finsk personbeteckning hos Migrationsverket i samband med registrering av uppehållsrätten för EU-medborgare.
Skattekort och skattenummer
Alla som arbetar i Finland ska ha ett skattekort.
Din arbetsgivare behöver kortet för utbetalning av lön och för beskattningen.
Om du jobbar inom byggbranschen behöver du också ett skattenummer (veronumero).
Du får skattekort och skattenummer på den närmaste skattebyrån.
På InfoFinlands sida Arbetstagare eller företagare finns mer information för arbetstagare som flyttar till Finland.
Jobbsökning i Finland
Om du är medborgare i ett EU-land kan du komma till Finland för att söka jobb för en rimlig tid.
Du kan inte registrera dig som invånare i Finland eller ansöka om registrering av uppehållsrätten när du är i landet som jobbsökande.
För att kunna bo kvar i Finland ska du ha ett jobb eller någon av de ovan nämnda anledningarna samt tillräckliga medel för din försörjning i Finland.
På InfoFinlands sida Var hittar jag jobb?
finns information om hur du kan hitta ett jobb i Finland.
Om du har rätt till arbetslöshetsersättning i ditt hemland, kan du även få den tillfälligt utbetald till Finland.
Du kan ansöka om utbetalning av arbetslöshetsersättning till Finland med blankett E303 eller U2.
Du får blanketten hos arbetskraftsmyndigheten i ditt hemland.
Om du kommer till Finland för att söka jobb kan du vanligtvis inte få arbetslöshetsersättning från Finland.
linkkiEuropa.eu:
Ta med dig dina arbetslöshetsförmånerfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Till Finland som företagare
Som EU-medborgare kan du starta ett företag i Finland om du är stadigvarande bosatt i ett land som hör till Europeiska ekonomiska samarbetsområdet (EES).
Också ett utländskt företag kan starta verksamhet i Finland.
Om din vistelse i Finland varar mer än tre månader ska du ansöka om registrering av uppehållsrätten för EU-medborgare i tjänsten Enter Finland eller på Migrationsverkets (maahanmuuttovirasto) tjänsteställe.
Om du flyttar till Finland för att bo här stadigvarande i minst ett år ska du också registrera dig som invånare i magistraten.
Etableringsanmälan
När du registrerar ditt företag för första gången ska du fylla i en etableringsanmälan och skicka in erforderliga bilagor.
Du behöver eventuellt bifoga till etableringsanmälan också ett utdrag som motsvarar handelsregisterutdraget i Finland, som en myndighet i ditt hemland utfärdar.
I InfoFinlands avsnitt Arbete och entreprenörskap hittar du mycket information om arbetslivet och företagande i Finland.
Som företagare till Finland:
Vilka tillstånd behöver du?(pdf, 384 kt)finska _ engelska
linkkiPatent- och registerstyrelsen:
Anmälan om grundande av ett företagfinska _ svenska _ engelska
Att studera i Finland
Som EU-medborgare kan du ansöka om studieplats vid en läroanstalt som är godkänd i Finland.
Om din vistelse i Finland varar mer än tre månader utan avbrott ska du ansöka om registrering av uppehållsrätten för EU-medborgare i tjänsten Enter Finland eller på Migrationsverkets (Maahanmuuttovirasto) tjänsteställe.
Om du flyttar till Finland för att bo här stadigvarande i minst ett år ska du också registrera dig som invånare i magistraten (maistraatti).
Om du vistas i Finland tre månader utan avbrott behöver du inte ansöka om registrering av uppehållsrätten.
Vistelsetiden på tre månader räknas alltid från det att du varit utanför Finlands gränser.
Denna regel gäller till exempel utbytesstudenter som endast studerar en kort period i Finland (t.ex. fyra månader). Om du lämnar
Finland under vistelsen och inte stannar i landet tre månader utan avbrott, behöver du inte ansöka om registrering av uppehållsrätten.
I detta fall ska du ansöka om en finsk personbeteckning och meddela din adress till magistraten (maistraatti).
På InfoFinlands sida Studerande finns mer information för studerande som flyttar till Finland.
Om du är EU-medborgare och flyttar till
Finland för att bo hos en familjemedlem ska du ansöka om registrering av uppehållsrätten för EU-medborgare på grund av familjeband i tjänsten Enter Finland eller på Migrationsverkets (Maahanmuuttovirasto) tjänsteställe.
Om du inte är EU-medborgare men din familjemedlem som bor i Finland är EU-medborgare, behöver du ett uppehållskort för en familjemedlem till en EU-medborgare.
Du ansöker om kortet i tjänsten Enter Finland eller vid Migrationsverkets (Maahanmuuttovirasto) tjänsteställe.
Om du flyttar till Finland för att bo här stadigvarande ska du också registrera dig som invånare i magistraten (maistraatti).
För registrering av en familjemedlem till en EU-medborgare krävs också att den person som är bosatt i Finland har tillräckliga medel för att försörja sig själv och sin familjemedlem som ska flytta till Finland.
Familjemedlemmar och andra anhöriga kan vara:
Din sambo som du har bott tillsammans med i minst två år eller med vilken du har gemensam vårdnad om ett barn
Ett barn eller barnbarn under 21 år som är beroende av dig för sin försörjning
Ett barn eller barnbarn under 21 år som är beroende av din sambo för sin försörjning
Din förälder eller mor- eller farförälder som är beroende av dig för sin försörjning
Din förälder eller mor- eller farförälder som är beroende av din sambo för sin försörjning
En förälder till ett barn under 21 år
Också ett barn som föds i Finland och blir medborgare i ett EU-land, Liechtenstein eller Schweiz måste ansöka om registrering av uppehållsrätten.
Registrering ska ansökas inom tre månader efter att barnet föddes.
Läs mer om detta på InfoFinlands sida När ett barn föds i Finland.
När du flyttar till Finland på grund av familjeband, har du obegränsad rätt att arbeta och studera i Finland.
På InfoFinlands sida Familjemedlem finns mer information för dem som flyttar till Finland på grund av familjeskäl.
Kort vistelse i Finland
Som EU-medborgare kan du komma till Finland om du har ett pass eller ett ID-kort förutsatt att du inte har utfärdats ett inreseförbud.
Om du vistas i Finland tillfälligt, kan du få en finsk personbeteckning om det behövs till exempel på grund av ditt arbete.
Du kan hämta en personbeteckning och samtidigt registrera ditt tillfälliga boende i den närmaste magistraten (maistraatti) eller skattebyrån (verotoimisto).
Ta med dig ett giltigt ID-kort eller pass.
Om din tillfälliga vistelse varar i över tre månader, behöver du också ett intyg över registrering av uppehållsrätten för medborgare i Europeiska unionen.
Läs mer om ämnet: Registrering av uppehållsrätten för EU-medborgare.
Om du bor i Finland tillfälligt, registreras ingen hemkommun för dig i Finland och du har inte samma rättigheter som de personer som bor i Finland stadigvarande.
Resor i Finland
Om du är medborgare i ett EU-land, Liechtenstein eller Schweiz och vill resa till Finland för en kort period, till exempel på semester, på affärsresa eller för att besöka släktingar, behöver du inget visum.
Du kan resa till Finland om du har ett giltigt ID-kort eller pass.
Om du är i Finland som turist och råkar ut för någon besvärlig situation, kontakta ditt hemlands beskickning.
Beskickningen kan hjälpa dig om du har råkat ut för en olycka, blivit sjuk eller blivit utsatt för ett brott.
Beskickningen kan också utförda dig ett nytt pass om du har tappat bort eller blivit bestulen på ditt pass.
linkkiVisitFinland.com:
Information om Finland till turistersvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ japanska _ italienska
Andra länders beskickningar i Finlandfinska _ svenska _ engelska
Om du är av finländsk härkomst eller har en nära kontakt med Finland kan du beviljas uppehållstillstånd i Finland på grund av detta.
Då är du återflyttare (paluumuuttaja).
Huruvida du beviljas uppehållstillstånd beror på hur starka och nära släktband du har till Finland.
För att få tillståndet krävs inga andra skäl, som till exempel arbete eller studier.
Personer som aldrig själv har varit finska medborgare men vars ena förälder eller mor- eller farförälder är eller har varit infödd finsk medborgare betraktas som återflyttare (paluumuuttaja) av finsk härkomst.
Också före detta finska medborgare räknas som återflyttare.
Uppehållstillstånd för återflyttarefinska _ svenska _ engelska
Avkomlingar till infödda finska medborgare
Du kan beviljas uppehållstillstånd i Finland om minst en av dina föräldrar eller mor- eller farföräldrar är eller har varit infödd finsk medborgare.
Med infödd finsk medborgare avses en person som har fått finskt medborgarskap vid födseln.
När du ansöker om tillstånd måste du ge en tillförlitlig bild av din härkomst, som till exempel uppvisa den ursprungliga födelseattesten av en förälder eller en mor- eller farförälder samt ett intyg över ert släktskap.
Du krävs inte på redogörelse över din utkomst.
Före detta finska medborgare
Om du är en före detta finsk medborgare kan du på denna grund få uppehållstillstånd i Finland.
Förutsättningen är inte att du är en infödd finsk medborgare, utan du kan också ha fått det finska medborgarskapet på ansökan.
Du krävs inte på redogörelse över din utkomst.
Om du är en före detta finsk medborgare kan du återfå ditt finska medborgarskap genom att göra en medborgarskapsanmälan (kansalaisuusilmoitus).
Läs mer på InfoFinlands sida Finskt medborgarskap.
Ansökan om uppehållstillstånd
Du kan ansöka om uppehållstillstånd antingen utomlands innan du kommer till Finland eller i Finland.
Utomlands kan du ansöka om tillstånd vid den närmaste av Finlands ambassader, i Finland vid Migrationsverkets tjänsteställe.
Du måste personligen gå och lämna in ansökan om uppehållstillstånd.
Ta med dig originalexemplaren av de bilagor som krävs för ansökan när du lämnar in din ansökan vid ambassaden eller Migrationsverkets tjänsteställe.
När du ansöker om uppehållstillstånd måste du ha med dig ett pass för att kunna styrka din identitet.
När du ansöker om tillstånd tas dina fingeravtryck för det biometriska uppehållstillståndskortet.
Ansökan om uppehållstillstånd är avgiftsbelagd.
Avgiften måste betalas i samband med att man lämnar in sin tillståndsansökan.
Finsk personbeteckning
När du ansöker om ditt första uppehållstillstånd i Finland kan du även be om att bli registrerad i Finlands befolkningsdatasystem.
Då får du en finsk personbeteckning på samma gång som du får uppehållstillståndet.
Mer information om personbeteckningen hittar du på InfoFinlands sida Registrering som invånare.
Uppehållstillstånd för avkomlingar till infödda finländarefinska _ svenska _ engelska
Uppehållstillstånd för före detta finska medborgarefinska _ svenska _ engelska
linkkiFinland-Samfundet:
Utlandsfinländarnas intresseorganisationfinska _ svenska _ engelska
Uppehållstillstånd för företagare
Uppehållstillstånd för uppstartsföretagare
Att ansöka om uppehållstillstånd
Företagare i Finland
I Finland kan vem som helst med hemvist i ett land som hör till Europeiska ekonomiska samarbetsområdet (EES) starta ett företag.
Behovet av tillstånd är inte beroende av din nationalitet utan din bosättningsort.
Om du är medborgare i ett EU-land, EES-land, nordiskt land eller Schweiz och vill flytta till Finland för att starta ett företag, behöver du inget uppehållstillstånd.
Läs mer på InfoFinlands sida EU-medborgare.
Om du inte har hemvist inom EES och är medborgare i något annat land än ett medlemsland i den Europeiska unionen, ett EES-land eller Schweiz, behöver du ett uppehållstillstånd för att driva ett företag i Finland.
Din företagsverksamhet ska vara lönsam och dina inkomster från företagsverksamheten måste ge dig en tryggad försörjning.
Du måste ansöka om ditt första uppehållstillstånd innan du kommer till Finland.
Uppehållstillstånd för företagare
Om du vill arbeta som företagare i Finland behöver du ett uppehållstillstånd för företagare.
Som företagare betraktas:
Uppstartsföretagare
Privat näringsidkare, som driver en så kallad firma
Bolagsman i ett öppet bolag
Ansvarig bolagsman i kommanditbolag
Medlem i andelslag med obegränsad tillskottsplikt
Delägare som innehar en ledande ställning i ett aktiebolag (verkställande direktör eller styrelsemedlem) eller person som innehar en ledande ställning i någon annan sammanslutning
För att få uppehållstillstånd för företagare måste du själv arbeta i ditt företag i Finland.
Om du inte har hemvist i Finland eller något annat land inom EES, måste du registrera din företagsverksamhet i Patent- och registerstyrelsens handelsregister innan du ansöker om uppehållstillstånd för företagare.
Om du flyttar stadigvarande till Finland eller EES-området behöver du inte Patent- och registerstyrelsens tillstånd för att grunda företaget.
Tillståndet är alltså inte kopplat till din nationalitet utan till var du har din hemvist.
Ansökan om uppehållstillstånd behandlas i två steg.
Först bedömer NTM-centralen (Närings-, trafik- och miljöcentralen) ditt företags lönsamhet bland annat utifrån affärsverksamhetsplanen och finansieringen.
Därefter fattar Migrationsverket beslut om uppehållstillstånd.
På Migrationsverkets webbplats hittar du mer information om villkoren för att ansöka om uppehållstillstånd.
linkkiPatent- och registerstyrelsen:
Tillstånd för företagare som är bosatta utanför EES-områdetfinska _ svenska _ engelska
Uppehållstillstånd för företagarefinska _ svenska _ engelska
Chatbot-tjänst för utländska företagarefinska _ engelska
Uppehållstillstånd för uppstartsföretagare
Om du vill grunda ett uppstartsföretag i Finland kan du ansöka om uppehållstillstånd för uppstartsföretagare som är avsett för tillväxtföretagare.
För att få uppehållstillstånd för uppstartsföretagare måste du ha en konkret affärsverksamhetsplan.
Ansökan om uppehållstillstånd för uppstartsföretagare är indelat i två steg:
Du behöver ett utlåtande från Business Finland som bifaller verksamheten som tillväxtföretagare.
Ansök om uppehållstillstånd för uppstartsföretagare och besök Finlands beskickning eller Migrationsverkets serviceställe för att styrka din identitet.
Processen är mycket snabb och smidig.
Finland som stöder företag bedömer ditt företags affärsmodell, kunnande och förmåga att få verksamheten att växa.
Du kan skicka uppgifterna om din affärsverksamhetsplan och erforderliga handlingar till Business Finland på elektronisk väg.
När du har fått ett positivt utlåtande från Business Finland kan du ansöka om uppehållstillstånd för uppstartsföretagare hos Migrationsverket.
Bifoga utlåtandet till din ansökan om uppehållstillstånd för uppstartsföretagare som du skickar till Migrationsverket.
Du kan inte få uppehållstillstånd för uppstartsföretagare i Finland utan ett positivt utlåtande från Business Finland.
Du hittar anvisningar och mer information om ansökan om uppehållstillstånd för uppstartsföretagare på Migrationsverkets och Business Finlands webbplatser.
Uppehållstillstånd för uppstartsföretagarefinska _ svenska _ engelska
Uppehållstillstånd för uppstartsföretagareengelska
Att ansöka om uppehållstillstånd
Du kan ansöka om uppehållstillstånd för företagare eller uppehållstillstånd för uppstartsföretagare på internet via tjänsten Enter Finland.
När du ställt ansökan ska du besöka Finlands beskickning närmast dig för att styrka din identitet och visa upp originalexemplaren av ansökningsbilagorna.
Du ska besöka beskickningen inom tre månader efter att ha gjort ansökan på internet.
Ansökningen kan tas för behandling först när du har besökt beskickningen.
Vanligtvis måste du boka en tid hos beskickningen i förväg.
Kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan kommer detta att meddelas via ditt konto.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du också lämna in en pappersansökan jämte bilagor vid Finlands beskickning närmast dig.
Du kan skriva ut ansökningsblanketten på Migrationsverkets webbplats.
Handläggning av tillståndsansökan är avgiftsbelagd.
Du betalar avgiften när du lämnar in din tillståndsansökan.
Läs mer om att grunda ett företag på InfoFinlands sida Att grunda ett företag i Finland.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Finsk personbeteckning
Om du får ett uppehållstillstånd i Finland registreras du automatiskt i det finska befolkningsdatasystemet.
Du får samtidigt även en finsk personbeteckning.
När du har flyttat till Finland ska du besöka magistraten på din hemort för att registrera dig som invånare.
Läs mer på InfoFinlands sida Registrering som invånare.
Företagare i Finland
På InfoFinlands sida Arbete och entreprenörskap hittar du mer information avsedd för företagare och arbetstagare.
Guide om att grunda ett företagfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ turkiska _ kinesiska _ arabiska
Tjänster för företagare-Startup Kitengelska
Migrationsverket:Presentation av e-tjänsten Enter Finland
Visste du..?
Lokal information
På Infobankens sidor hittar du mycket information om tjänsterna på olika orter.
lokal-information
På denna sida finns information riktad till kvotflyktingar.
Information om att ansöka om asyl hittar du på InfoFinlands sida Till Finland som asylsökande.
Kvotflyktingar
Man kan inte ansöka om att bli kvotflykting via myndigheterna i Finland.
Man kan inte heller föreslå en annan person, till exempel en släkting eller vän, som kvotflykting.
Finland tar som kvotflyktingar emot personer som har flyktingstatus enligt Förenta nationernas flyktingorganisation UNHCR.
Kvotflyktingarna väljs bland de personer som UNHCR föreslår till Finland.
De finländska myndigheterna intervjuar dessa flyktingar. Utgående från intervjuerna väljer man de flyktingar som tas emot till Finland.
Intervjuerna görs i de länder där flyktingarna vistas, vanligen i flyktingläger eller i UNHCR:s lokaler.
Information om val av kvotflyktingarfinska _ svenska _ engelska
Flytta till Finland
På webbsidan Movingtofinland.fi finns mycket information avsedd för kvotflyktingar om att flytta till Finland och om livet i Finland.
Information för flyktingarfinska _ engelska _ franska _ persiska _ arabiska _ kurdiska
Stöd till flyktingar
Finlands röda kors (FRK) hjälper kvotflyktingar när de flyttar till Finland.
När flyktingarna anländer till Finland kommer en anställd från röda korset till flygplatsen och tar emot dem.
Röda korsets frivilligarbetare hjälper även flyktingar att bosätta sig och integreras i Finland.
Flyktingar kan be om hjälp och rådgivning i rättsliga frågor bland annat från flyktingrådgivningen r.f. eller från rättshjälpsbyråer.
Finlands flyktinghjälp r.f. är en organisation som strävar efter att främja de grundläggande rättigheterna för flyktingar.
Organisationen utför informations-, utbildnings och socialarbete i Finland.
Flyktinghjälpen hjälper flyktingar och invandrare till exempel med ärenden som gäller integrering, boende och grundande av egna organisationer.
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
linkkiFinlands flyktinghjälp r.f.:
Stöd till flyktingarfinska _ svenska _ engelska
linkkiFinlands röda kors:
Stöd till flyktingarfinska _ svenska _ engelska
Rehabiliteringscentret för tortyrofferfinska _ engelska
Som flykting i Finland
På InfoFinlands sida Flykting hittar du mer information avsedd för flyktingar.
Uppehållstillstånd för arbetstagare
Andra uppehållstillstånd för förvärvsarbete
Uppehållstillstånd för säsongsarbete
Arbete med ett annat uppehållstillstånd
Ansökan om uppehållstillstånd
Arbete utan uppehållstillstånd
Arbetstagare i Finland
Den här sidan är avsedd för dig som är medborgare i något annat land är ett EU-land, Norge, Island, Schweiz eller Liechtenstein.
Om du kommer till Finland för att arbeta behöver du ett uppehållstillstånd.
Innan du kan få ett uppehållstillstånd måste du hitta ett jobb i Finland.
När du har hittat ett jobb kan du ansöka om uppehållstillstånd.
Du måste ansöka om uppehållstillstånd innan du kommer till Finland.
För att kunna arbeta i Finland behöver du vanligen antingen ett uppehållstillstånd för arbetstagare eller någon annan typ av uppehållstillstånd för förvärvsarbete.
Arten av det arbete du ska utföra påverkar typen av tillstånd.
Uppehållstillstånd för arbetstagare
Om du inte kan arbeta med stöd av ett annat uppehållstillstånd eller utan uppehållstillstånd behöver du ett uppehållstillstånd för arbetstagare (työntekijän oleskelulupa).
Uppehållstillstånd för arbetstagare är inte nödvändigt för alla arbetsuppgifter.
Du kan granska hurudant uppehållstillstånd du behöver från Migrationsverkets webbplats.
Du behöver uppehållstillstånd för arbetstagare om du arbetar till exempel som:
städare
hemvårdare eller barnskötare.
Migrationsverket beslutar om du ska beviljas uppehållstillstånd eller inte.
Ett delbeslut av arbets- och näringsbyrån behövs också för tillståndet.
Uppehållstillstånd för arbetstagarefinska _ svenska _ engelska
Andra uppehållstillstånd för förvärvsarbete
För vissa arbetsuppgifter behöver du inte ett uppehållstillstånd för arbetstagare, men du behöver dock ett uppehållstillstånd som beviljas för vissa uppdrag.
Dessa uppdrag kan vara till exempel:
uppdrag inom företagsledning
uppdrag som sakkunnig
forskaruppdrag
uppdrag inom vetenskap, kultur och konst
arbetspraktik.
Migrationsverket beslutar om du får uppehållstillstånd eller inte.
Ett delbeslut av arbets- och näringsbyrån behövs inte för tillståndet.
Arbete i Finlandfinska _ svenska _ engelska
Uppehållstillstånd för säsongsarbete
Om du ska utföra säsongsarbete i Finland behöver du ett säsongsarbetstillstånd.
Säsongsarbetet kan pågå högst nio månader.
Säsongsarbete är till exempel:
växtodling
skogsvårdsarbete
festivalarbete
Om du kommer från ett viseringspliktigt land och ska arbeta i under tre månader, måste du ansöka om ett säsongsarbetsvisum hos den finländska beskickningen.
Om ditt arbete pågår över tre månader ska du ansöka om ett säsongsarbetstillstånd hos Migrationsverket.
Tillstånd för säsongsarbetefinska _ svenska _ engelska
Arbete med ett annat uppehållstillstånd
Om du redan har uppehållstillstånd i Finland utifrån en annan grund, till exempel familjeband, kan du ha rätt att arbeta i Finland.
Då behöver du inte ett separat uppehållstillstånd för att arbeta.
Du kan kontrollera om du har rätt att arbeta i Finland från ditt uppehållstillståndskort eller beslut om uppehållstillstånd.
Rätt att arbetafinska _ svenska _ engelska
Om du har avlagt examen i Finland kan du få ett tillfälligt uppehållstillstånd för att söka arbete.
Detta tillstånd kan beviljas endast som ett fortsatt tillstånd till ett uppehållstillstånd för studerande.
Ansök om tillståndet innan ditt uppehållstillstånd för studerande löper ut.
Du kan få ett tillstånd för högst ett år.
Detta tillstånd kan man endast få en gång.
Om du hittar en arbetsplats, kan du börja arbeta genast.
Du måste ansöka om ett nytt uppehållstillstånd på grund av arbete innan ditt uppehållstillstånd för att söka arbete går ut.
Om du har avlagt examen i Finland, behövs inte ett delbeslut av arbets- och näringsbyrån för ditt tillstånd.
Uppehållstillstånd för sökande av arbetefinska _ svenska _ engelska
Ansökan om uppehållstillstånd
Du måste ansöka om ditt första uppehållstillstånd innan du kommer till Finland.
Du kan ansöka om tillståndet på internet via tjänsten Enter Finland.
När du ställt ansökan ska du besöka Finlands beskickning närmast dig för att styrka din identitet och visa upp originalexemplaren av ansökningsbilagorna.
Du ska besöka beskickningen inom tre månader efter att ha gjort ansökan på internet.
Ansökningen kan tas för behandling först när du besökt beskickningen.
Vanligtvis måste du boka en tid hos beskickningen i förväg.
Kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan kommer detta att meddelas via ditt konto.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du också lämna in en pappersansökan jämte bilagor vid Finlands beskickning närmast dig.
Du kan skriva ut ansökningsblanketten på Migrationsverkets webbplats.
Handläggningen av din ansökan om tillstånd är avgiftsbelagd.
Du måste betala avgiften när du lämnar in ansökan om uppehållstillstånd.
Till ansökan om uppehållstillstånd för arbetstagare ska du bifoga blanketten TEM054 som din arbetsgivare fyller i och undertecknar.
Arbetsgivaren kan lämna uppgifterna om arbetet och sitt företag själv samt följa handläggning av ansökan direkt via tjänsten Enter Finland.
Arbetsgivaren kan även betala handläggningsavgiften för arbetstagaren.
Fråga din arbetsgivare som hen använder tjänsten Enter Finland för arbetsgivare.
Kom ändå ihåg att arbetsgivaren inte kan ansöka om uppehållstillstånd för dig, utan hen kompletterar din ansökan för egen del i tjänsten Enter Finland.
Så länge handläggningen av din första ansökan om uppehållstillstånd pågår har du inte rätt att arbeta.
Om du har ansökt om uppehållstillstånd utomlands, kan du inte komma till Finland innan tillstånd har beviljats.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Handläggningstider för tillståndsansökningarfinska _ svenska _ engelska
Ansökan om uppehållstillstånd för specialist
Om du ska arbeta i Finland som specialist kan du även komma till Finland utan uppehållstillstånd.
Du måste dock ha visum eller rätt att vistas i Finland tre månader utan visum.
Du ska också ha en arbetsplats som uppfyller kraven.
Om du arbetar i Finland längre än tre månader måste du ansöka om uppehållstillstånd.
Du kan ansöka om tillståndet elektroniskt via tjänsten Enter Finland eller på Migrationsverkets tjänsteställe.
Finsk personbeteckning
Om du får ett uppehållstillstånd i Finland registreras du automatiskt i det finska befolkningsdatasystemet.
Du får samtidigt även en finsk personbeteckning.
När du har flyttat till Finland ska du besöka magistraten på din hemort för att registrera dig som invånare.
Läs mer på InfoFinlands sida Registrering som invånare.
Arbete utan uppehållstillstånd
Oberoende av vilket land du är medborgare i kan du i vissa fall arbeta i Finland utan uppehållstillstånd.
Du måste dock ha ett visum, om du behöver visum till Finland.
Du kan arbeta i Finland utan uppehållstillstånd till exempel om:
du kommer till Finland för att arbeta som tolk, lärare, sakkunnig eller idrottsdomare i högst tre månader utifrån en inbjudan eller ett avtal;
du är fast anställd vid ett företag som bedriver verksamhet i ett annat EU/EES-land och ska komma till Finland för att utföra tillfälligt leverans- eller underleveransarbete och ditt arbete pågår högst tre månader;
du är asylsökande i Finland och har ett giltigt resedokument som berättigar till gränsövergång.
Trots att du inte har uppehållstillstånd kan du börja arbeta tre månader efter att du har lämnat in din asylansökan;
du är asylsökande i Finland och har inte ett giltigt resedokument som berättigar till gränsövergång.
Trots att du inte har uppehållstillstånd kan du börja arbeta när du vistats i sex månader i landet.
Du kan granska om du har rätt att arbeta i Finland utan uppehållstillstånd från Migrationsverkets webbplats.
Arbete utan uppehållstillståndfinska _ svenska _ engelska
Arbetstagare i Finland
På InfoFinlands sida Var hittar jag jobb? finns information om hur du kan hitta ett jobb i Finland.
InfoFinlands sidor Arbete och entreprenörskap innehåller mer information för arbetstagare och företagare.
linkkiArbets- och näringsministeriet:
Arbeta i Finlandfinska _ svenska _ engelska
linkkiArbets- och näringsbyrån:
Broschyren Jobba i Finland(pdf, 5,51 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ polska
linkkiArbetshälsoinstitutet:
Handboken Jobba i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ kurdiska _ tyska _ thai _ vietnamesiska
Migrationsverket:
Presentation av e-tjänsten Enter Finland
Söka asyl
Asylsökande från Europeiska unionens område
Minderåriga asylsökande
Handläggning av asylansökan
Asylsamtal
Positivt beslut
Negativt beslut
Rättshjälp för asylsökande
Asylsökandes rätt att arbeta
Du kan söka asyl i Finland om du har välgrundad fruktan för förföljelse i ditt hemland.
Orsaker till förföljelse kan vara etniskt ursprung, religion, medborgarskap, tillhörighet till en viss grupp i samhället eller politiska åsikter.
Migrationsverket utreder om det finns asylskäl och fattar ett beslut.
Du kan endast söka asyl för dig själv.
Broschyren Information till asylsökandefinska _ svenska _ engelska _ ryska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
Söka asyl
Du kan endast söka asyl i Finland på det finska territoriet.
Det finns ingen särskild asylansökningsblankett som du skulle kunna fylla i förväg.
När du kommer till Finland, meddela gränskontrollmyndigheten eller polisen genast att du vill söka asyl.
Gränskontrollmyndigheten eller polisen registrerar dig som asylsökande, antecknar uppgifter om dig och tar dina fingeravtryck.
När myndigheten har mottagit din asylansökan, hänvisas du till ett mottagningscenter.
Där kan du bo under tiden då Migrationsverket behandlar din ansökan.
Du kan även bo någon annanstans, men då måste du själv bekosta boendet.
Att söka asyl i Finlandfinska _ svenska _ engelska
Asylsökande från Europeiska unionens område
Inom EU (och i Schweiz, Norge, Island och Liechtenstein) måste man söka asyl i det land, till vars territorium man kommer först.
Om du har sökt asyl eller vistats i något annat EU-land (eller i Schweiz, Norge, Island eller Liechtenstein) innan du kom till Finland, behandlas din ansökan inte i Finland.
I detta fall avvisas du tillbaka till det land där du var innan du kom till Finland.
Detta kallas för Dublinprocessen.
Om du är medborgare i ett EU-land, får du sannolikt inte asyl i Finland.
Finland anser att alla EU-länder är trygga för medborgarna.
Likväl utreds alla ansökningar som EU-medborgare skickar in.
På InfoFinlands sida EU-medborgare hittar du information om flytt till Finland av andra skäl än som asylsökande.
Att lämna asylansökan utan prövningfinska _ svenska _ engelska
Minderåriga asylsökande
Om du är under 18 år gammal och kommer till Finland som asylsökande utan vårdnadshavare, förordnas du ett ombud.
Ombudet är en pålitlig vuxen person som hjälper dig med olika ärenden under tiden då Migrationsverket behandlar din ansökan.
Ombudet följer med dig när du ska prata med myndigheter.
Dessutom utreder ditt ombud om du kan återförenas med din familj.
Du har rätt till boende, mat och hälsovård.
Du har även rätt att gå i skola.
Ensamkommande barn(pdf, 674)finska _ svenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ persiska _ arabiska _ kurdiska
Handläggning av asylansökan
Migrationsverket handlägger din ansökan och fattar ett beslut.
Migrationsverket utreder din identitet och resväg till Finland och bedömer om du kan beviljas asyl i Finland.
Det är vanligt att behandlingen av ansökan tar flera månader.
När du har sökt asyl har du rätt att vistas i Finland medan din ansökan behandlas.
Under denna tid kan du inte resa utomlands.
Om du reser kan myndigheterna besluta att din ansökan inte längre gäller.
Migrationsverket skickar dig en kallelse till asylsamtal.
I kallelsen anges tolkningsspråket, den exakta adressen till verksamhetsstället där samtalet hålls och klockslaget.
Handläggning av asylansökanfinska _ svenska _ engelska
Asylsamtal
Asylsamtalet (turvapaikkapuhuttelu) är den viktigaste händelsen under behandlingen av din ansökan.
Under samtalet ställs frågor om de händelser och orsaker som tvingade dig att lämna ditt hemland.
Det är viktigt att du beskriver allt som hänt så exakt som möjligt.
Migrationsverket beslutar baserat på din berättelse om du beviljas asyl i Finland.
Som asylsökande har du rätt att använda ett rättsbiträde under samtalet.
Biträdet deltar i asylsamtalet efter sitt eget omdöme.
Om du behöver en tolk, skaffar Migrationsverket tolken.
Positivt beslut
Du får stanna i Finland om du beviljas asyl eller uppehållstillstånd på andra grunder.
Du kan beviljas asyl i Finland om myndigheterna anser att du blir förföljd i ditt hemland på grund av
etniskt ursprung,
religion,
medborgarskap,
tillhörighet till en viss grupp i samhället eller
politiska åsikter.
Om du inte får asyl kan du i vissa fall beviljas uppehållstillstånd på grund av alternativt skydd.
Du kan beviljas uppehållstillstånd på grund av alternativt skydd om du hotas av:
dödsstraff eller avrättning,
tortyr eller någon annan behandling eller bestraffning som är omänsklig eller kränker människovärdet eller
om du utsätts för allvarlig personlig fara på grund av en väpnad konflikt.
När du söker asyl utreder Migrationsverket samtidigt om du kan få uppehållstillstånd på någon annan grund.
Asylfinska _ svenska _ engelska
Negativt beslut
Om du inte beviljas asyl eller uppehållstillstånd på någon annan grund blir du avvisad från Finland.
Du har även möjlighet att överklaga ett negativt beslut till förvaltningsdomstolen.
Bifogat till beslutet finns en anvisning om hur du överklagar.
På InfoFinlands sida Negativt beslut om uppehållstillstånd hittar du information om vad du kan göra om du får ett negativt beslut.
Ändringssökande i asylbeslutfinska _ svenska _ engelska
Avvisning av en asylsökandefinska _ svenska _ engelska
Rättshjälp för asylsökande
Under tiden då din ansökan behandlas kan du få rådgivning och rättshjälp vid den offentliga rättshjälpsbyrån.
Kontakta rättshjälpsbyrån om du vill ha ett rättsbiträde.
Vid behov hjälper mottagningscentret dig.
Rättshjälpsbyrån (oikeusaputoimisto) kan även hänvisa dig till en privat jurist eller en privat juristbyrå.
Du kan även få rådgivning hos Flyktingrådgivningen rf (Pakolaisneuvonta ry).
Flyktingrådgivningen ger rådgivning även till personer som vistas i Finland utan uppehållstillstånd.
linkkiRättsväsendet:
Rättshjälpsbyråerfinska _ svenska _ engelska
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Asylsökandes rätt att arbeta
Du får förvärvsarbeta i Finland om det har gått tre månader sedan du lämnade in din asylansökan och du har ett giltigt pass eller någon annan resehandling som du har företett till myndigheten när du sökte asyl.
Om du inte företedde en giltig resehandling till myndigheten i samband med din asylansökan får du förvärvsarbeta i Finland när det har gått sex månader sedan du lämnade in din asylansökan.
Du har rätt att arbeta tills du har fått ett lagakraftvunnet beslut på din asylansökan.
Om Migrationsverket ger dig ett positivt beslut på din asylansökan, får du uppehållstillstånd.
I det ingår nästan alltid rätt att arbeta.
Om Migrationsverket fattar ett negativt beslut på din asylansökan, har du rätt att arbeta under tiden då en eventuell överklagan behandlas.
För att arbeta måste du ha ett finländskt skattekort.
Hämta ett skattekort på den närmaste skattebyrån och lämna kortet till din arbetsgivare.
Läs mer på InfoFinlands sida Skattekort.
Om du arbetar permanent kan du även ansöka om uppehållstillstånd i Finland på grund av arbete.
På InfoFinlands sida Arbeta i Finland hittar du mer information om uppehållstillstånd för arbetstagare.
Asylsökandes rätt att arbetafinska _ svenska _ engelska
Uppehållstillstånd på andra grunderfinska _ svenska _ engelska
Hur ansöker jag?
Vad behövs för registreringen?
Kan jag bli av med uppehållsrätten?
Registrering av uppehållsrätten för EU-medborgare sker inte per automatik.
Du kan ansöka om registrering av uppehållsrätten om din försörjning i Finland är tryggad.
Den kan vara baserad på ett jobb, studier, företagsverksamhet, familjeband eller tillräckliga medel.
Om du avser att bo i Finland längre än tre månader, måste du registrera din uppehållsrätt hos Migrationsverket (Maahanmuuttovirasto).
Ansökan ska lämnas in senast inom tre månader från datumet för inresa.
Registreringen hos Migrationsverket är inte samma sak som registreringen av din bosättningsort i befolkningsdatasystemet (väestötietojärjestelmä) vid magistraten (maistraatti).
Om din sammanhängande vistelse i Finland är kortare än tre månader behöver du inte registrera vistelsen vid Migrationsverket.
Vistelsetiden på tre månader räknas alltid från det att du varit utanför Finlands gränser.
Läs mer om förutsättningarna på sidan EU-medborgare.
Hur ansöker jag?
Handläggning av ansökan om registrering av uppehållsrätt är avgiftsbelagd.
Du betalar avgiften när du lämnar in din ansökan.
Ansök om registrering av uppehållsrätten för EU-medborgare i tjänsten Enter Finland:
Fyll i ansökningsblanketten och bifoga erforderliga bilagor.
Du hittar information om vilka bilagor som behövs till ansökningen i avsnittet
Vad behövs för registreringen?
Besök Migrationsverkets tjänsteställe; du måste styrka din identitet och visa upp originalexemplaren av ansökningsbilagorna.
Ta med dig ett giltigt ID-kort eller pass.
Du ska besöka tjänstestället inom tre månader efter att ha gjort ansökan.
Det är bra att boka en tid på tjänstestället i förväg.
Boka tiden via Migrationsverkets elektroniska tidsbokningssystem.
Kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan, kommer detta att meddelas via ditt Enter Finland-konto.
Du får också ett meddelande när beslutet är klart.
Om du inte kan eller inte vet hur du ska göra ansökan på internet:
Gör registreringsansökan på en pappersblankett.
Du kan även göra det personligen på Migrationsverkets tjänsteställe.
Gör ansökan inom tre månader efter datumet för inresa.
Skriv ut registreringsblanketten på Migrationsverkets webbplats och fyll i den färdigt.
Var noga när du fyller i ansökan.
Felaktigt ifyllda ansökningar tas inte emot.
Boka en tid på Migrationsverkets tjänsteställe i det elektroniska tidsbokningssystemet.
Det är bra att boka en tid på tjänstestället i förväg.
Ta med dig den ifyllda registreringsblanketten, ett giltigt ID-kort eller pass och erforderliga bilagor.
Du hittar information om vilka bilagor som behövs till ansökningen i avsnittet
Vad behövs för registreringen?
Om kraven på grund och förutsättningar för vistelsen Finland uppfylls, kan du få ett intyg över registrering av uppehållsrätten för medborgare i Europeiska unionen från Migrationsverket.
Registreringen av uppehållsrätten gäller tillsvidare.
När du har bott lagligt och utan avbrott i Finland i fem år, har du permanent uppehållsrätt.
Permanent uppehållsrätt för EU-medborgare ansöks separat från Migrationsverket.
Registrering av uppehållsrätt för EU-medborgarefinska _ svenska _ engelska
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Permanent uppehållstillståndfinska _ svenska _ engelska
Om magistraten registrerar din uppehållsrätt, registreras dina personuppgifter automatiskt även i befolkningsdatasystemet.
Du får samtidigt även en finsk personbeteckning.
Du kan få en finsk personbeteckning även vid magistraten eller skattebyrån på din hemort.
Om du flyttar till Finland för att bo här stadigvarande i ett år eller längre, ska du också registrera dig i magistraten på din hemort.
Läs mer på InfoFinlands sida Registrering som invånare.
På InfoFinlands sida Komihåglista för dig som flyttar till Finland hittar du nyttig information om allt som du ska ta hand om när du flyttar till Finland.
Vad behövs för registreringen?
Arbetstagare eller företagare
Din uppehållsrätt kan registreras om du är anställd eller har ett eget företag i Finland.
Du behöver följande handlingar:
EU-registreringsblankett
Giltigt ID-kort eller pass
Anställningsavtal (om du är anställd)
En utredning över företagsverksamheten (om du är egenföretagare)
Studerande
Din uppehållsrätt kan registreras om du studerar vid en läroanstalt som är godkänd i Finland.
Du behöver följande handlingar:
EU-registreringsblankett
Giltigt ID-kort eller pass
Närvarointyg (intyg över att du är studerande vid en läroanstalt som är godkänd i Finland)
Du har en sjukförsäkring (t.ex. det europeiska sjukvårdskortet)
En utredning över din försörjning i Finland
Familjemedlem till en person bosatt i Finland
Din uppehållsrätt kan registreras om du har en familjemedlem som är stadigvarande bosatt i Finland.
Du behöver följande handlingar:
EU-registreringsblankett
Giltigt ID-kort eller pass
Intyg över äktenskap eller registrerat parförhållande
En utredning över att ni har bott tillsammans i två år eller har gemensam vårdnad om ett barn, om du är i ett samboförhållande
Barnets födelseattest om du har vårdnaden om ett barn
En utredning över grunden för att den person som ansöker om familjeförening vistas i Finland.
Uppehållskort för en familjemedlem till en EU-medborgare
Om du inte själv är medborgare i ett EU-land, Liechtenstein eller Schweiz men avser att flytta till Finland till en familjemedlem som är EU-medborgare, måste du ansöka om uppehållskort för en familjemedlem till en EU-medborgare.
Du kan ansöka om uppehållskortet elektroniskt via tjänsten Enter Finland eller på Migrationsverkets (Maahanmuuttovirasto) tjänsteställe.
Handläggning av ansökan om uppehållskort är avgiftsbelagd.
Du betalar avgiften när du lämnar in din ansökan.
Du behöver följande handlingar:
Ansökan om uppehållskort
Giltigt pass
Intyg över äktenskap eller registrerat parförhållande
Registreringsintyget för den EU-medborgare, med vem du kommer till Finland
Utredning över släktskapsförhållandet (barn till EU-medborgaren eller andra släktingar som står under dennes vårdnad)
Utredning över samboskap (om du är sambo med EU-medborgaren och ni inte har gemensam vårdnad om barn)
Uppehållskortet för en familjemedlem till en EU-medborgare beviljas för fem år eller en kortare tid om boendet i Finland varar mindre än fem år.
Uppehållskort för EU-medborgares familjemedlemfinska _ svenska _ engelska
Tillräckliga medel
Om din uppehållsrätt inte kan registreras på någon av de ovan nämnda grunderna kan du ansöka om registrering om du har tillräckliga medel för din försörjning i Finland.
Också tillräckliga medel är en grund.
Du behöver följande handlingar:
EU-registreringsblankett
Giltigt ID-kort eller pass
En utredning över att du har tillräckliga medel för din försörjning i Finland.
Kan jag bli av med uppehållsrätten?
Registreringen av uppehållsrätten för en EU-medborgare och uppehållskortet för en familjemedlem till en EU-medborgare kan återkallas eller bli ogiltigt om:
du flyttar permanent från Finland
du har vistats utomlands utan avbrott i två år
du lämnade felaktiga uppgifter när du ansökte om registreringen eller om uppehållskortet för en familjemedlem till en EU-medborgare
du har undanhållit sådan information som skulle kunna ha hindrat dig från att få registreringen eller uppehållskortet
du utvisas från Finland
du får finskt medborgarskap.
Tänk på att ändringar i din livssituation kan påverka din uppehållsrätt.
Om din uppehållsrätt registrerades på basis av arbete, ett aktivt företag, en studieplats, familjeband eller tillräckliga medel, och detta skäl inte längre existerar, kan registreringen återkallas.
Beslut om återkallande eller upphörande av uppehållsrätten fattas av Migrationsverket.
Om du flyttar utomlands
Om du inte vill att ditt uppehållstillstånd eller uppehållskort ska återkallas ska du lämna in en ansökan om detta hos Migrationsverket senast inom två år efter att du har flyttat utomlands.
Återkallande av uppehållsrättfinska _ svenska _ engelska
Också andra anhöriga till finska medborgare än en make/maka, en sambo, föräldrar till minderåriga barn eller minderåriga barn kan i vissa fall få uppehållstillstånd i Finland på grund av familjeband.
Även andra anhöriga till en person som har ett uppehållstillstånd på grund av internationellt skydd kan beviljas uppehållstillstånd.
Om uppehållstillståndet beviljats på någon annan grund än internationellt skydd, kan andra anhöriga inte få uppehållstillstånd.
En annan anhörig kan få uppehållstillstånd om han eller hon är helt beroende av den anhöriga som bor i Finland.
På denna grund kan uppehållstillstånd beviljas till exempel för en förälder till en myndig (18 år gammal) person.
Enbart ekonomiskt beroende eller svag hälsa räcker ändå inte för att beviljas uppehållstillstånd.
En annan anhörig kan få uppehållstillstånd också om han eller hon levt tillsammans som en familjemedlem till den anhöriga som är bosatt i Finland, innan denna person kom till Finland.
Dessutom krävs det att familjelivet upphört på grund av ett tvingande skäl, till exempel för att man blivit flyktingar.
Annan anhörig till en finsk medborgarefinska _ svenska _ engelska
Annan anhörig till en person som fått internationellt skyddfinska _ svenska _ engelska
Att ansöka om uppehållstillstånd
Vanligtvis måste du ansöka om ditt första uppehållstillstånd innan du kommer till Finland.
Ansök om tillståndet i ditt hemland eller i ett annat land där du vistas lagligt.
Du kan ansöka om tillståndet på internet via tjänsten Enter Finland.
När du ställt ansökan ska du besöka Finlands beskickning närmast dig eller Migrationsverkets tjänsteställe för att styrka din identitet och visa upp originalexemplaren av ansökningsbilagorna.
Du ska besöka beskickningen eller tjänstestället inom tre månader efter att ha gjort ansökan på internet.
Ansökningen kan tas för behandling först när du besökt beskickningen eller tjänstestället.
Vanligtvis måste du boka en tid hos beskickningen eller tjänstestället i förväg.
Kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan, kommer detta att meddelas via ditt Enter Finland-konto.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du också lämna in en pappersansökan jämte bilagor vid Finlands beskickning närmast dig eller på Migrationsverkets tjänsteställe i Finland.
Du kan skriva ut ansökningsblanketten på Migrationsverkets webbplats.
Ansökan om uppehållstillstånd är avgiftsbelagd.
Avgiften ska betalas då ansökan ställs.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Finlands beskickningar utomlandsfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Finsk personbeteckning
När du ansöker om det första uppehållstillståndet i Finland kan du även be om registrering i det finska befolkningsdatasystemet.
Då får du en finsk personbeteckning samtidigt som du får ditt uppehållstillstånd.
Mer information om personbeteckningen hittar du på InfoFinlands sida Registrering som invånare.
Arbeta i Finland
Till Finland som företagare
Att studera i Finland
Till familjemedlem i Finland
Kort vistelse i Finland
Om du är medborgare i ett EU-land, Liechtenstein eller Schweiz, behöver du inget uppehållstillstånd eller visum i Finland.
Du kan resa till Finland om du har ett giltigt ID-kort eller pass.
Du har rätt att arbeta, driva ett företag och studera i Finland med lika villkor som finska medborgare.
Du måste själv trygga din försörjning i Finland.
Som EU-medborgare kan du vistas i Finland högst tre månader i sträck utan att registrera din uppehållsrätt.
Om du vill stanna kvar i Finland och registrera dig som invånare, ska du ha ett jobb eller ett aktivt företag, en studieplats, ett långvarigt familjeband eller tillräckliga medel.
Om du avser att bo i Finland i över tre månader, ska du ansöka om Registrering av uppehållsrätten för EU-medborgare hos Migrationsverket.
Ansökan ska ställas senast inom tre månader från datumet för inresa.
Om du flyttar till Finland för att bo här stadigvarande i ett år eller längre, ska du också registrera dig i magistraten på din hemort.
Läs mer på InfoFinlands sida Registrering som invånare.
Om du vistas i Finland tre månader utan avbrott behöver du inte ansöka om registrering av uppehållsrätten.
Vistelsetiden på tre månader räknas alltid från det att du varit utanför Finlands gränser.
linkkiEuropa.eu:
EU-länderfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Rådgivning för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropeiska kommissionen:
Europeiska sjukvårdskortetfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Arbeta i Finland
Som EU-medborgare behöver du inget arbetstillstånd i Finland.
Du kan börja jobba direkt när du har kommit till landet.
Hämta ett skattekort på den närmaste skattebyrån (Verotoimisto) och lämna kortet till din arbetsgivare.
Om du ska jobba i Finland i mer än tre månader ska du ansöka om registrering av uppehållsrätten för EU-medborgare i tjänsten Enter Finland eller på Migrationsverkets (Maahanmuuttovirasto) tjänsteställe.
Om du flyttar till Finland för att bo här stadigvarande i minst ett år ska du också registrera dig som invånare i magistraten (maistraatti).
Personbeteckning
Om du kommer till Finland från utlandet för att arbeta, behöver du en finsk personbeteckning.
Du får personbeteckningen på magistraten (maistraatti) eller skattebyrån (verotoimisto).
Ett giltigt ID-kort eller pass
Ditt anställningsavtal
Du kan även få en finsk personbeteckning hos Migrationsverket i samband med registrering av uppehållsrätten för EU-medborgare.
Skattekort och skattenummer
Alla som arbetar i Finland ska ha ett skattekort.
Din arbetsgivare behöver kortet för utbetalning av lön och för beskattningen.
Om du jobbar inom byggbranschen behöver du också ett skattenummer (veronumero).
Du får skattekort och skattenummer på den närmaste skattebyrån.
På InfoFinlands sida Arbetstagare eller företagare finns mer information för arbetstagare som flyttar till Finland.
Jobbsökning i Finland
Om du är medborgare i ett EU-land kan du komma till Finland för att söka jobb för en rimlig tid.
Du kan inte registrera dig som invånare i Finland eller ansöka om registrering av uppehållsrätten när du är i landet som jobbsökande.
För att kunna bo kvar i Finland ska du ha ett jobb eller någon av de ovan nämnda anledningarna samt tillräckliga medel för din försörjning i Finland.
På InfoFinlands sida Var hittar jag jobb?
finns information om hur du kan hitta ett jobb i Finland.
Om du har rätt till arbetslöshetsersättning i ditt hemland, kan du även få den tillfälligt utbetald till Finland.
Du kan ansöka om utbetalning av arbetslöshetsersättning till Finland med blankett E303 eller U2.
Du får blanketten hos arbetskraftsmyndigheten i ditt hemland.
Om du kommer till Finland för att söka jobb kan du vanligtvis inte få arbetslöshetsersättning från Finland.
linkkiEuropa.eu:
Ta med dig dina arbetslöshetsförmånerfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Till Finland som företagare
Som EU-medborgare kan du starta ett företag i Finland om du är stadigvarande bosatt i ett land som hör till Europeiska ekonomiska samarbetsområdet (EES).
Också ett utländskt företag kan starta verksamhet i Finland.
Om din vistelse i Finland varar mer än tre månader ska du ansöka om registrering av uppehållsrätten för EU-medborgare i tjänsten Enter Finland eller på Migrationsverkets (maahanmuuttovirasto) tjänsteställe.
Om du flyttar till Finland för att bo här stadigvarande i minst ett år ska du också registrera dig som invånare i magistraten.
Etableringsanmälan
När du registrerar ditt företag för första gången ska du fylla i en etableringsanmälan och skicka in erforderliga bilagor.
Du behöver eventuellt bifoga till etableringsanmälan också ett utdrag som motsvarar handelsregisterutdraget i Finland, som en myndighet i ditt hemland utfärdar.
I InfoFinlands avsnitt Arbete och entreprenörskap hittar du mycket information om arbetslivet och företagande i Finland.
Som företagare till Finland:
Vilka tillstånd behöver du?(pdf, 384 kt)finska _ engelska
linkkiPatent- och registerstyrelsen:
Anmälan om grundande av ett företagfinska _ svenska _ engelska
Att studera i Finland
Som EU-medborgare kan du ansöka om studieplats vid en läroanstalt som är godkänd i Finland.
Om din vistelse i Finland varar mer än tre månader utan avbrott ska du ansöka om registrering av uppehållsrätten för EU-medborgare i tjänsten Enter Finland eller på Migrationsverkets (Maahanmuuttovirasto) tjänsteställe.
Om du flyttar till Finland för att bo här stadigvarande i minst ett år ska du också registrera dig som invånare i magistraten (maistraatti).
Om du vistas i Finland tre månader utan avbrott behöver du inte ansöka om registrering av uppehållsrätten.
Vistelsetiden på tre månader räknas alltid från det att du varit utanför Finlands gränser.
Denna regel gäller till exempel utbytesstudenter som endast studerar en kort period i Finland (t.ex. fyra månader).
Om du lämnar Finland under vistelsen och inte stannar i landet tre månader utan avbrott, behöver du inte ansöka om registrering av uppehållsrätten.
I detta fall ska du ansöka om en finsk personbeteckning och meddela din adress till magistraten (maistraatti).
På InfoFinlands sida Studerande finns mer information för studerande som flyttar till Finland.
Till familjemedlem i Finland
Om du är EU-medborgare och flyttar till Finland för att bo hos en familjemedlem ska du ansöka om registrering av uppehållsrätten för EU-medborgare på grund av familjeband i tjänsten Enter Finland eller på Migrationsverkets (Maahanmuuttovirasto) tjänsteställe.
Om du inte är EU-medborgare men din familjemedlem som bor i Finland är EU-medborgare, behöver du ett uppehållskort för en familjemedlem till en EU-medborgare.
Du ansöker om kortet i tjänsten Enter Finland eller vid Migrationsverkets (Maahanmuuttovirasto) tjänsteställe.
Om du flyttar till Finland för att bo här stadigvarande ska du också registrera dig som invånare i magistraten (maistraatti).
För registrering av en familjemedlem till en EU-medborgare krävs också att den person som är bosatt i Finland har tillräckliga medel för att försörja sig själv och sin familjemedlem som ska flytta till Finland.
Familjemedlemmar och andra anhöriga kan vara:
Din sambo som du har bott tillsammans med i minst två år eller med vilken du har gemensam vårdnad om ett barn
Ett barn eller barnbarn under 21 år som är beroende av dig för sin försörjning
Ett barn eller barnbarn under 21 år som är beroende av din sambo för sin försörjning
Din förälder eller mor- eller farförälder som är beroende av dig för sin försörjning
Din förälder eller mor- eller farförälder som är beroende av din sambo för sin försörjning
En förälder till ett barn under 21 år
Också ett barn som föds i Finland och blir medborgare i ett EU-land, Liechtenstein eller Schweiz måste ansöka om registrering av uppehållsrätten.
Registrering ska ansökas inom tre månader efter att barnet föddes.
Läs mer om detta på InfoFinlands sida När ett barn föds i Finland.
När du flyttar till Finland på grund av familjeband, har du obegränsad rätt att arbeta och studera i Finland.
På InfoFinlands sida Familjemedlem finns mer information för dem som flyttar till Finland på grund av familjeskäl.
Kort vistelse i Finland
Som EU-medborgare kan du komma till Finland om du har ett pass eller ett ID-kort förutsatt att du inte har utfärdats ett inreseförbud.
Om du vistas i Finland tillfälligt, kan du få en finsk personbeteckning om det behövs till exempel på grund av ditt arbete.
Du kan hämta en personbeteckning och samtidigt registrera ditt tillfälliga boende i den närmaste magistraten (maistraatti) eller skattebyrån (verotoimisto).
Ta med dig ett giltigt ID-kort eller pass.
Om din tillfälliga vistelse varar i över tre månader, behöver du också ett intyg över registrering av uppehållsrätten för medborgare i Europeiska unionen.
Läs mer om ämnet: Registrering av uppehållsrätten för EU-medborgare.
Om du bor i Finland tillfälligt, registreras ingen hemkommun för dig i Finland och du har inte samma rättigheter som de personer som bor i Finland stadigvarande.
Resor i Finland
Om du är medborgare i ett EU-land, Liechtenstein eller Schweiz och vill resa till Finland för en kort period, till exempel på semester, på affärsresa eller för att besöka släktingar, behöver du inget visum.
Du kan resa till Finland om du har ett giltigt ID-kort eller pass.
Om du är i Finland som turist och råkar ut för någon besvärlig situation, kontakta ditt hemlands beskickning.
Beskickningen kan hjälpa dig om du har råkat ut för en olycka, blivit sjuk eller blivit utsatt för ett brott.
Beskickningen kan också utförda dig ett nytt pass om du har tappat bort eller blivit bestulen på ditt pass.
linkkiVisitFinland.com:
Information om Finland till turistersvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ japanska _ italienska
Andra länders beskickningar i Finlandfinska _ svenska _ engelska
Barn till en finsk medborgare
Barnet kan få uppehållstillstånd på grund av familjeband om hans/hennes förälder är finsk medborgare eller gift med en finsk medborgare och bor i Finland.
Barnet måste vara under 18 år gammalt och ogift den dag då beslutet om uppehållstillstånd fattas.
Den förälder till barnet som är bosatt i Finland måste vara barnets vårdnadshavare för att barnet ska kunna få uppehållstillstånd.
Om båda föräldrarna är vårdnadshavare måste även den andra föräldern ge sitt samtycke till att barnet flyttar till Finland.
En myndighet, till exempel en notaries publicus, måste verifiera överenskommelsen.
Familjebandet mellan föräldern och barnet måste bevisas, till exempel med en födelseattest med föräldrarnas namn.
Barnets vårdnadshavare gör ansökan för det minderåriga barnets del.
Även barnet måste vara närvarande när tillståndsansökan lämnas in.
Barn till en finsk medborgarefinska _ svenska _ engelska
Barn till en utländsk medborgare
Barnet kan få uppehållstillstånd på grund av familjeband om hans/hennes föräldrar har uppehållstillstånd i Finland och en förälder bor i Finland.
Barnet måste vara under 18 år gammalt och ogift den dag då beslutet om uppehållstillstånd fattas.
Även ett barn som föds i Finland behöver ett uppehållstillstånd i Finland.
Tillståndet måste sökas inom tre månader från barnets födelse.
Den förälder till barnet som är bosatt i Finland måste vara barnets vårdnadshavare för att barnet ska kunna få uppehållstillstånd.
Om båda föräldrarna är vårdnadshavare måste även den andra föräldern ge sitt samtycke till att barnet flyttar till Finland.
En myndighet, till exempel en notaries publicus, måste verifiera överenskommelsen.
Familjebandet mellan föräldern och barnet måste bevisas till exempel med en födelseattest med föräldrarnas namn.
För att barnet ska kunna få uppehållstillstånd måste hans/hennes uppehälle i Finland vara tryggat, till exempel genom förälderns löneinkomster.
Kravet på tillräcklig inkomst tillämpas dock inte på föräldern om barnet fötts innan föräldern anlänt till Finland och föräldern har flyktingstatus i Finland.
Om föräldern har fått flyktingstatus den 1.7.2016 eller senare, ska man ansöka om uppehållstillstånd för barnet inom tre månader från att föräldern fått flyktingstatus.
Ansökan kan även göras senare, men då tillämpas kravet på tillräcklig inkomst.
Om barnets förälder har uppehållstillstånd på grund av internetionellt skydd, men inte flyktingstatus, krävs att föräldern har en tillräcklig inkomst för att barnet ska kunna få uppehållstillstånd.
Barnets vårdnadshavare gör ansökan för det minderåriga barnets del.
Även barnet måste vara närvarande när tillståndsansökan lämnas in.
Barn till en utländsk medborgarefinska _ svenska _ engelska
Utkomstförutsättningfinska _ svenska _ engelska
Barn till en person som fått internationellt skyddfinska _ svenska _ engelska
Förälder eller annan vårdnadshavare
Du kan få uppehållstillstånd på grund av familjeband om ditt barn bor i Finland.
Barnet måste vara under 18 år gammalt och ogift den dag då beslutet om uppehållstillstånd fattas.
För att få uppehållstillstånd på grund av familjeband måste du vara barnets vårdnadshavare.
Vanligtvis är barnets mor eller far vårdnadshavare.
Vårdnadshavaren kan dock även vara någon annan, till exempel en mor- eller farförälder.
Familjebandet mellan barnet och föräldern måste bevisas till exempel med en födelseattest med föräldrarnas namn.
Om en annan vårdnadshavare än barnets mor eller far ansöker om uppehållstillstånd måste vårdnaden bevisas till exempel genom uppvisande av ett domstolsbeslut.
För att du ska kunna få uppehållstillstånd måste du ha tillräckliga medel för att leva i Finland.
Kravet på tillräcklig inkomst tillämpas dock inte på dig om ditt barn är en finsk medborgare.
Kravet på tillräcklig inkomst tillämpas inte heller om du varit barnets vårdnadshavare redan innan barnet anlänt till Finland och barnet har flyktingstatus i Finland.
Om barnet fått flyktingstatus den 1.7.2016 eller senare, ska du ansöka om uppehållstillstånd inom tre månader från att barnet fått flyktingstatus i Finland.
Ansökan kan även göras senare, men då tillämpas kravet på tillräcklig inkomst.
Vårdnadshavare till en finsk medborgarefinska _ svenska _ engelska
Vårdnadshavare till en utländsk medborgarefinska _ svenska _ engelska
Utkomstförutsättningfinska _ svenska _ engelska
Vårdnadshavare till en person som fått internationellt skyddfinska _ svenska _ engelska
Att ansöka om uppehållstillstånd
Vanligtvis måste du ansöka om ditt första uppehållstillstånd innan du kommer till Finland.
Ansök om tillståndet i ditt hemland eller i ett annat land där du vistas lagligt.
Du kan också ansöka om ditt första visum i Finland, om din familjemedlem är finsk medborgare och du själv är medborgare i ett visumfritt land, det vill säga du inte behöver visum för att komma till Finland.
Du kan ansöka om tillståndet på internet via tjänsten Enter Finland.
När du ställt ansökan ska du besöka Finlands beskickning närmast dig eller Migrationsverkets tjänsteställe för att styrka din identitet och visa upp originalexemplaren av ansökningsbilagorna.
Du ska besöka beskickningen eller tjänstestället inom tre månader efter att ha gjort ansökan på internet.
Ansökningen kan tas för behandling först när du besökt beskickningen eller tjänstestället.
Det är bra att boka en tid hos beskickningen eller tjänstestället i förväg.
Kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan, kommer detta att meddelas via ditt Enter Finland-konto.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du också lämna in en pappersansökan jämte bilagor vid Finlands beskickning närmast dig eller på Migrationsverkets tjänsteställe i Finland.
Du kan skriva ut ansökningsblanketten på Migrationsverkets webbplats.
Ansökan om uppehållstillstånd är avgiftsbelagd.
Avgiften ska betalas då ansökan ställs.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Finlands beskickningar utomlandsfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Finsk personbeteckning
När du ansöker om det första uppehållstillståndet i Finland kan du även be om registrering i det finska befolkningsdatasystemet.
Då får du en finsk personbeteckning samtidigt som du får ditt uppehållstillstånd.
Mer information om personbeteckningen hittar du på InfoFinlands sida Registrering som invånare.
Visste du..?
Lokal information
På Infobankens sidor hittar du mycket information om tjänsterna på olika orter.
lokal-information
Make/maka till en finsk medborgare
Make/maka till en utländsk medborgare
Make/maka till en flykting
Partner
Att ansöka om uppehållstillstånd
Om maken/makan/sambon/partnern inte får uppehållstillstånd
Make/maka till en finsk medborgare
Om du har ingått äktenskap med en finländsk medborgare som är bosatt i Finland kan du få uppehållstillstånd i Finland på grund av familjeband.
Även en maka/make av samma kön kan få uppehållstillstånd, om ni är gifta eller i ett registrerat parförhållande.
Sambo med en finsk medborgare
Om du är sambo med en finsk medborgare som bor i Finland kan du få uppehållstillstånd på grund av familjeband.
Tillståndet kan beviljas om:
du har bott tillsammans med din sambo minst två år eller
du har ett gemensamt barn med din sambo (då uteblir kravet på gemensamt boende under två års tid) eller
det finns något annat vägande skäl för att bevilja tillståndet
Ifall du ansöker om tillstånd på dessa grunder måste du och din sambo bevisa att ni har bott tillsammans två år.
Som bevis godtas till exempel ett utdrag ur boenderegistret eller ett hyreskontrakt med bådas namn.
Om du och din sambo är bosatta i olika stater anses gemensamt boende till exempel under semesterresor inte som en tillräcklig grund för beviljande av uppehållstillstånd.
Varken du eller din sambo får vara gift med någon annan.
Försörjningsförutsättning för make/maka till en finsk medborgare
Om du är familjemedlem till en finsk medborgare, behöver din försörjning inte vara tryggad.
Du har obegränsad rätt att arbeta.
Du får börja arbeta först när du har fått ett uppehållstillstånd.
Information om hur du ansöker om tillståndet finns under rubriken Att ansöka om uppehållstillstånd.
Make eller maka till en finsk medborgarefinska _ svenska _ engelska
Sambo till en finsk medborgarefinska _ svenska _ engelska
Make/maka till en utländsk medborgare
Om din make/maka har uppehållstillstånd i Finland och bor i Finland kan du få uppehållstillstånd
Sambo med en utländsk medborgare
Om din sambo har uppehållstillstånd i Finland och bor i Finland kan du få uppehållstillstånd i Finland på grund av familjeband.
Du kan få tillståndet om:
du har bott tillsammans med din sambo minst två år eller
du har ett gemensamt barn tillsammans med din sambo (då uteblir kravet på gemensamt boende under två års tid)
Ifall du ansöker om tillstånd på dessa grunder måste du och din sambo bevisa att ni har bott tillsammans två år.
Som bevis duger till exempel ett utdrag ur boenderegistret eller ett hyreskontrakt med bådas namn.
Om du och din sambo är bosatta i olika stater anses gemensamt boende till exempel under semesterresor inte som en tillräcklig grund för beviljande av uppehållstillstånd.
Varken du eller din sambo får vara gift med någon annan.
Försörjningsförutsättning för make/maka till en utländsk medborgare
För att du ska få uppehållstillstånd i Finland måste du eller din make/maka ha tillräcklig inkomst även för din försörjning.
På Migrationsverkets sidor kan du kontrollera hur stor inkomst ni måste ha.
Om din maka/make fått uppehållstillstånd på grund av internationellt skydd, tillämpas kravet på tillräcklig inkomst på er.
Det är möjligt att i enskilda fall avvika från försörjningsförutsättningen, om det finns exceptionellt vägande skäl eller om barnets bästa kräver detta.
Information om hur du ansöker om tillståndet finns under rubriken Att ansöka om uppehållstillstånd.
Make eller maka till en utländsk medborgarefinska _ svenska _ engelska
Sambo till en utländsk medborgarefinska _ svenska _ engelska
Utkomstförutsättningfinska _ svenska _ engelska
Make/maka till en flykting
Om din maka/make har uppehållstillstånd i Finland på grund av internationellt skydd och flyktingstatus, kan du få uppehållstillstånd i Finland på grund av familjeband.
Sambo med flykting
Om din sambo har uppehållstillstånd i Finland på grund av internationellt skydd och flyktingstatus, kan du få uppehållstillstånd i Finland på grund av familjeband.
Du kan få tillståndet om:
du har bott tillsammans med din sambo minst två år eller
du har ett gemensamt barn tillsammans med din sambo (då uteblir kravet på gemensamt boende under två års tid)
Ifall du ansöker om tillstånd på dessa grunder måste du och din sambo bevisa att ni har bott tillsammans två år.
Som bevis duger till exempel ett utdrag ur boenderegistret eller ett hyreskontrakt med bådas namn.
Om du och din sambo är bosatta i olika stater anses gemensamt boende till exempel under semesterresor inte som en tillräcklig grund för beviljande av uppehållstillstånd.
Varken du eller din sambo får vara gift med någon annan.
Försörjningsförutsättning för make/maka/sambo/partner till en flykting
Försörjningsförutsättningen tillämpas på er på olika sätt, om din make/maka/sambo/partner har fått uppehållstillstånd på grund av internationellt skydd och har flyktingstatus i Finland.
Din försörjning behöver inte vara tryggad i följande fall:
Om din make/maka/sambo/partner har beviljats asyl eller godkänts som kvotflykting före den 1 juli 2016 och familjen har bildats före hen kom till Finland.
Om din make/maka/sambo/partner har fått flyktingstatus den 1 juli 2016 eller efter detta ska ansökan om uppehållstillstånd lämnas in inom tre månader efter att hen fått beslut på sin ansökan.
De tre månaderna räknas från den dag då din maka/make/sambo/partner delgivits beslutet.
Om du, av anledningar som du inte själv kan påverka, inte hinner ansöka om uppehållstillstånd inom tre månader, kan du ändå ansöka om familjeåterförening.
I din ansökan ska du ange varför tidsfristen på tre månader överskreds.
Du kan ansöka om familjeåterförening även senare, men då tillämpas kravet på tillräcklig inkomst på er.
Försörjningsförutsättningen gäller er även i det fall att ni gifte er efter att din make/maka kom till Finland.
I vissa enskilda fall kan man avvika från försörjningsförutsättningen om det finns exceptionellt vägande skäl eller om barnets bästa kräver detta.
Information om hur du ansöker om tillståndet finns under rubriken Att ansöka om uppehållstillstånd.
Maka eller make till en person som fått internationellt skyddfinska _ svenska _ engelska
Sambo till en person som fått internationellt skyddfinska _ svenska _ engelska
Försörjningsförutsättning för familjemedlemmar till personer som får internationellt skyddfinska _ svenska _ engelska
Partner
Man kan vanligen inte få uppehållstillstånd på grund av sällskapande.
I Finland är en person man sällskapar med inte en familjemedlem enligt lagen.
I vissa fall kan du ändå få ett tillfälligt (B) uppehållstillstånd i Finland på grund av sällskapande.
För att du ska kunna beviljas uppehållstillstånd i Finland måste ditt och din partners förhållande vara stadigt.
Ett bevis på stadigt sällskapande kan till exempel vara att er avsikt är att ingå äktenskap i Finland.
Varken du eller din partner får vara gift med någon annan.
För att du ska kunna få uppehållstillstånd måste du ha tillräckliga medel för ditt uppehälle.
Dessa medel bör vara fritt tillgängliga för dig till exempel på ditt eget bankkonto.
Inkomsterna för din partner som är bosatt i Finland beaktas inte.
Flick- eller pojkvän till en finsk medborgarefinska _ svenska _ engelska
Att ansöka om uppehållstillstånd
Vanligtvis måste du ansöka om ditt första uppehållstillstånd innan du kommer till Finland.
Ansök om tillståndet i ditt hemland eller i ett annat land där du vistas lagligt. Du kan också ansöka om ditt första uppehållstillstånd i Finland om din make eller maka är finsk medborgare och du själv är medborgare i ett visumfritt land, det vill säga du inte behöver visum för att komma till Finland.
Du kan ansöka om tillståndet på internet via tjänsten Enter Finland.
När du ställt ansökan ska du besöka Finlands beskickning närmast dig eller Migrationsverkets tjänsteställe för att styrka din identitet och visa upp originalexemplaren av ansökningsbilagorna.
Du ska besöka beskickningen eller tjänstestället inom tre månader efter att ha gjort ansökan på internet.
Ansökningen kan tas för behandling först när du besökt beskickningen eller tjänstestället.
Vanligtvis måste du boka en tid hos beskickningen eller tjänstestället i förväg.
Kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan, kommer detta att meddelas via ditt Enter Finland-konto.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du också lämna in en pappersansökan jämte bilagor vid Finlands beskickning närmast dig eller på Migrationsverkets tjänsteställe i Finland.
Du kan skriva ut ansökningsblanketten på Migrationsverkets webbplats.
Ansökan om uppehållstillstånd är avgiftsbelagd.
Avgiften ska betalas då ansökan ställs.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Finlands beskickningar utomlandsfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Handläggningstider för tillståndsansökningarfinska _ svenska _ engelska
Finsk personbeteckning
När du ansöker om det första uppehållstillståndet i Finland kan du även be om registrering i det finska befolkningsdatasystemet.
Då får du en finsk personbeteckning samtidigt som du får ditt uppehållstillstånd.
Mer information om personbeteckningen hittar du på InfoFinlands sida Registrering som invånare.
Om maken/makan/sambon/partnern inte får uppehållstillstånd
En make/maka/sambo/partner beviljas inte uppehållstillstånd om förutsättningarna för uppehållstillstånd inte uppfylls.
Man kan låta bli att bevilja tillståndet även då de finländska myndigheterna anser att parterna har ingått äktenskap endast för uppehållstillståndets skull och att makarna inte avser att leva tillsammans som en familj.
Myndigheterna kan misstänka att parterna ingått äktenskap endast för uppehållstillståndets skull till exempel om ni har ingått äktenskap efter endast en kort bekantskap, om det är stor åldersskillnad mellan er eller om den ena av er har haft flera korta äktenskap.
Om du får ett nekande beslut på din tillståndsansökan kan du överklaga den till förvaltningsdomstolen.
Du får instruktioner för detta bifogade till tillståndsbeslutet.
Läs mer om problem med uppehållstillståndet på InfoFinlands sida Problem med uppehållstillståndet.
Om du vill flytta till en familjemedlem som bor i Finland behöver du ett uppehållstillstånd.
Om du bara vill hälsa på hos din familjemedlem i Finland hittar du mer information på InfoFinlands sida Kort vistelse i Finland.
Alla familjemedlemmar kan inte få uppehållstillstånd.
Vanligen kan man få tillstånd om man är make/maka, sambo, minderårigt barn eller förälder till minderårigt barn till personen bosatt i Finland.
Ofta krävs det även att personen bosatt i Finland ska ha tillräckliga medel för att försörja en familjemedlem som flyttar till Finland.
Notera att separata regler gäller för familjemedlemmar till EU-medborgare (inte finländska medborgare).
Om du är familjemedlem till en EU-medborgare bosatt i Finland hittar du mer information om tillståndsärenden på InfoFinlands sidan EU-medborgare.
Mer information om hur familjemedlemmar kan få uppehållstillstånd finns på InfoFinlands sidor Uppehållstillstånd för make eller maka, Uppehållstillstånd för barn eller förälder, Uppehållstillstånd för övriga anhöriga.
På InfoFinlands sida Familjemedlem hittar du mer information avsedd för personer som flyttar av familjeskäl.
Till Finland på grund av familjebandfinska _ svenska _ engelska
Ansök om studieplats
Teckna en tillräckligt omfattande sjukförsäkring i ditt hemland
Reservera tillräckliga medel för din försörjning
Ansök om uppehållstillstånd för studerande
Uppehållstillstånd för studerande från andra EU-länder
Fortsatt uppehållstillstånd för studerande
När du avslutar dina studier
För praktik till Finland
Studier i Finland
Den här sidan är avsedd för dig som är medborgare i något annat land än ett EU-land, Norge, Island, Schweiz eller Liechtenstein.
Om du ska studera i Finland längre än 90 dagar behöver du ett uppehållstillstånd på grund av studier.
Du kan studera mindre än 90 dagar i Finland utan uppehållstillstånd.
Om du ska flytta till Finland för studier måste du ta hand om följande:
Ansök om studieplats
Innan du kan ansöka om uppehållstillstånd måste du skaffa dig en studieplats i Finland.
Godkända läroanstalter är läroanstalter efter grundskolan, till exempel universitet, högskolor och yrkesläroanstalter.
Studieplatsen ska uppfylla ett av följande villkor:
studierna leder till yrke eller examen
du deltar i ett utbytesprogram mellan läroanstalter eller något annat utbytesprogram
du avlägger en kompletterande utbildning eller en specialutbildning som hör till din examen.
Du kan ansöka om studieplats i skolornas gemensamma ansökan på våren eller hösten.
Till vissa utbildningar är den gemensamma ansökan (yhteishaku) redan i januari.
Ta i god tid reda på när du kan ansöka om en studieplats.
Fyll i ansökan i tjänsten Opintopolku.fi.
På InfoFinlands sida Ansökan till utbildning hittar du mer information om hur du ansöker om en studieplats i Finland.
Teckna en tillräckligt omfattande sjukförsäkring i ditt hemland
Som studerande betalar du själv vårdkostnaderna om du insjuknar i Finland.
För ditt uppehållstillstånd behöver du en privat försäkring som täcker kostnaderna för sjukdom och läkemedel.
Du kan teckna en försäkring hos ett försäkringsbolag i ditt hemland eller fråga om en lämplig försäkring hos internationella försäkringsbolag.
Alla försäkringar ska uppfylla följande villkor:
Försäkringens självrisk får inte överstiga 300 euro.
Försäkringen ska gälla under hela din vistelse i Finland.
Försäkringen ska gälla när du kommer till Finland.
Försäkringen får inte vara en vanlig reseförsäkring.
Säg inte upp din försäkring.
Om du insjuknar måste du själv betala läkar- och sjukhuskostnaderna.
Hur stora vårdkostnader som försäkringen måste täcka beror på hur länge dina studier varar.
Om dina studier i Finland till exempel varar mindre än två år, ska försäkringen täcka sjukvårdskostnader upp till minst 100 000 euro.
Om du har det europeiska sjukvårdskortet (European Health Insurance Card, EHIC), behöver du ingen separat försäkring.
Sjukvårdskortet ska vara giltigt under hela din vistelse i Finland.
Försäkring för studerandefinska _ svenska _ engelska
Reservera tillräckliga medel för din försörjning
Du måste också själv ansvara för levnadskostnaderna i Finland.
Du behöver ha minst 560 euro disponibla medel i månaden för att kunna betala för boende, mat och andra utgifter.
För en vistelse som varar ett år ska du alltså ha 6 720 euro i disponibla medel.
Försörjningsförutsättningen kan i vissa fall undgås.
Om till exempel läroanstalten ordnar dig en gratis bostad och även gratis måltider behöver du ha en mindre summa i disponibla medel.
Om studierna är avgiftsbelagda måste du även se till att du har tillräckliga medel för din försörjning efter att du har betalat läsårsavgiften.
Beloppet som krävs ska finnas på ditt bankkonto eller också ska du ha ett intyg över ett stipendium som beviljats av en officiell instans.
Sådana stipendier är till exempel de som beviljats av staten, läroanstalter eller organisationer.
Sponsringslöften eller kontoutdrag från privatpersoner, såsom släktingar, bekanta eller arbetsgivare, godkänns inte.
Försörjningsförutsättning för studerandefinska _ svenska _ engelska
Ansök om uppehållstillstånd för studerande
Du måste ansöka om ditt första uppehållstillstånd innan du kommer till Finland.
Du kan ansöka om tillståndet på internet via tjänsten Enter Finland.
När du ställt ansökan ska du besöka Finlands beskickning närmast dig för att styrka din identitet och visa upp originalexemplaren av ansökningsbilagorna.
Du ska besöka beskickningen inom tre månader efter att ha gjort ansökan på internet.
Ansökningen kan tas för behandling först när du besökt beskickningen.
Vanligtvis måste du boka en tid hos beskickningen i förväg.
Kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan kommer detta att meddelas via ditt konto.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du också lämna in en pappersansökan jämte bilagor vid Finlands beskickning närmast dig.
Du kan skriva ut ansökningsblanketten på Migrationsverkets webbplats.
Handläggningen av ansökan är avgiftsbelagd.
Du måste betala avgiften när du lämnar in ansökan om uppehållstillstånd.
Du ska bifoga följande handlingar till din ansökan om uppehållstillstånd för studerande:
Giltigt pass
Passfoto (anvisningar för fotot finns på Migrationsverkets webbplats)
Närvarointyg (intyg över att du är studerande vid en läroanstalt som är godkänd i Finland)
En utredning över att du har tillräckliga medel för din försörjning
Ett försäkringsintyg eller en kopia av det europeiska sjukvårdskortet
En utredning över att du har betalat läsårsavgiften eller har ett stipendium
Tidigare examensbetyg (om du inte ska avlägga examen eller är en utbytesstudent)
Eventuella arbetsintyg (om du inte ska avlägga examen eller är en utbytesstudent)
Information om uppehållstillstånd för studierfinska _ svenska _ engelska
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Finlands beskickningar utomlandsfinska _ svenska _ engelska
Uppehållstillstånd för studerande från andra EU-länder
Du behöver inget uppehållstillstånd i Finland om du har ett uppehållstillstånd som beviljats i ett annat EU-land och om du studerar vid en högskola.
Dessutom måste dina studier:
innefatta internationell rörlighet i ett EU-program eller ett mångformigt program eller
omfattas av ett avtal mellan två eller fler högskolor.
I detta fall måste du göra en underrättelse om rörlighet till Migrationsverket.
Du får studera i Finland högst 360 dagar när du gör en underrättelse om rörlighet.
Underrättelse om rörlighet i Finlandfinska _ svenska _ engelska
Fortsatt uppehållstillstånd för studerande
Uppehållstillstånd för studerande beviljas högst för två år i taget.
Om dina studier fortsätter men uppehållstillståndet håller på att gå ut ska du ansöka om fortsatt uppehållstillstånd.
Kom ihåg att ansöka om fortsatt uppehållstillstånd för studerande i god tid innan giltighetstiden för det första tillståndet går ut.
Observera att Migrationsverket (Maahanmuuttovirasto) även kontrollerar om grunden för din vistelse i Finland verkligen har varit studier.
Om du till exempel avlägger en grundexamen vid universitet, högskola eller yrkeshögskola bör du avlägga 45 studiepoäng under ett läsår för att uppfylla villkoren för fortsatt uppehållstillstånd.
Du ska bifoga ett studieregisterutdrag till din ansökan om fortsatt uppehållstillstånd.
Fortsatt uppehållstillstånd för studerandefinska _ svenska _ engelska
När du avslutar dina studier
Om du har avlagt en examen i Finland kan du få ett tillfälligt uppehållstillstånd för arbetssökande.
Detta tillstånd kan beviljas endast som ett fortsatt tillstånd till ett uppehållstillstånd för studerande.
Du ska ansöka om tillståndet innan ditt uppehållstillstånd för studerande går ut.
Uppehållstillstånd för arbetssökande kan beviljas för högst ett år.
Om du får ett jobb kan du börja arbeta direkt.
Du måste ansöka om ett nytt uppehållstillstånd på grund av arbete innan ditt uppehållstillstånd för arbetssökande går ut.
Uppehållstillstånd för sökande av arbetefinska _ svenska _ engelska
Till Finland som praktikant
Om du studerar utomlands och vill komma till Finland för arbetspraktik behöver du ett uppehållstillstånd på grund av praktik.
Mer information hittar du på Migrationsverkets webbplats.
Praktik i Finlandfinska _ svenska _ engelska
Att studera i Finland
Om du flyttar till Finland för att bo här stadigvarande i ett år eller längre, ska du också registrera dig i magistraten på din hemort.
Läs mer på InfoFinlands sida Registrering som invånare.
InfoFinlands sida Utländska studerande i Finland innehåller viktig information om studielivet i Finland.
Information för utländska studerandeengelska
Migrationsverket:
Presentation av e-tjänsten Enter Finland
Uppehållstillstånd för företagare
Uppehållstillstånd för uppstartsföretagare
Att ansöka om uppehållstillstånd
Företagare i Finland
I Finland kan vem som helst med hemvist i ett land som hör till Europeiska ekonomiska samarbetsområdet (EES) starta ett företag.
Behovet av tillstånd är inte beroende av din nationalitet utan din bosättningsort.
Om du är medborgare i ett EU-land, EES-land, nordiskt land eller Schweiz och vill flytta till Finland för att starta ett företag, behöver du inget uppehållstillstånd.
Läs mer på InfoFinlands sida EU-medborgare.
Om du inte har hemvist inom EES och är medborgare i något annat land än ett medlemsland i den Europeiska unionen, ett EES-land eller Schweiz, behöver du ett uppehållstillstånd för att driva ett företag i Finland.
Din företagsverksamhet ska vara lönsam och dina inkomster från företagsverksamheten måste ge dig en tryggad försörjning.
Du måste ansöka om ditt första uppehållstillstånd innan du kommer till Finland.
Uppehållstillstånd för företagare
Om du vill arbeta som företagare i Finland behöver du ett uppehållstillstånd för företagare.
Som företagare betraktas:
Uppstartsföretagare
Privat näringsidkare, som driver en så kallad firma
Bolagsman i ett öppet bolag
Ansvarig bolagsman i kommanditbolag
Medlem i andelslag med obegränsad tillskottsplikt
Delägare som innehar en ledande ställning i ett aktiebolag (verkställande direktör eller styrelsemedlem) eller person som innehar en ledande ställning i någon annan sammanslutning
För att få uppehållstillstånd för företagare måste du själv arbeta i ditt företag i Finland.
Om du inte har hemvist i Finland eller något annat land inom EES, måste du registrera din företagsverksamhet i Patent- och registerstyrelsens handelsregister innan du ansöker om uppehållstillstånd för företagare.
Om du flyttar stadigvarande till Finland eller EES-området behöver du inte Patent- och registerstyrelsens tillstånd för att grunda företaget.
Tillståndet är alltså inte kopplat till din nationalitet utan till var du har din hemvist.
Ansökan om uppehållstillstånd behandlas i två steg.
Först bedömer NTM-centralen (Närings-, trafik- och miljöcentralen) ditt företags lönsamhet bland annat utifrån affärsverksamhetsplanen och finansieringen.
Därefter fattar Migrationsverket beslut om uppehållstillstånd.
På Migrationsverkets webbplats hittar du mer information om villkoren för att ansöka om uppehållstillstånd.
linkkiPatent- och registerstyrelsen:
Tillstånd för företagare som är bosatta utanför EES-områdetfinska _ svenska _ engelska
Uppehållstillstånd för företagarefinska _ svenska _ engelska
Chatbot-tjänst för utländska företagarefinska _ engelska
Uppehållstillstånd för uppstartsföretagare
Om du vill grunda ett uppstartsföretag i Finland kan du ansöka om uppehållstillstånd för uppstartsföretagare som är avsett för tillväxtföretagare.
För att få uppehållstillstånd för uppstartsföretagare måste du ha en konkret affärsverksamhetsplan.
Ansökan om uppehållstillstånd för uppstartsföretagare är indelat i två steg:
Du behöver ett utlåtande från Business Finland som bifaller verksamheten som tillväxtföretagare.
Ansök om uppehållstillstånd för uppstartsföretagare och besök Finlands beskickning eller Migrationsverkets serviceställe för att styrka din identitet.
Processen är mycket snabb och smidig.
Finland som stöder företag bedömer ditt företags affärsmodell, kunnande och förmåga att få verksamheten att växa.
Du kan skicka uppgifterna om din affärsverksamhetsplan och erforderliga handlingar till Business Finland på elektronisk väg.
När du har fått ett positivt utlåtande från Business Finland kan du ansöka om uppehållstillstånd för uppstartsföretagare hos Migrationsverket.
Bifoga utlåtandet till din ansökan om uppehållstillstånd för uppstartsföretagare som du skickar till Migrationsverket.
Du kan inte få uppehållstillstånd för uppstartsföretagare i Finland utan ett positivt utlåtande från Business Finland.
Du hittar anvisningar och mer information om ansökan om uppehållstillstånd för uppstartsföretagare på Migrationsverkets och Business Finlands webbplatser.
Uppehållstillstånd för uppstartsföretagarefinska _ svenska _ engelska
Uppehållstillstånd för uppstartsföretagareengelska
Att ansöka om uppehållstillstånd
Du kan ansöka om uppehållstillstånd för företagare eller uppehållstillstånd för uppstartsföretagare på internet via tjänsten Enter Finland.
När du ställt ansökan ska du besöka Finlands beskickning närmast dig för att styrka din identitet och visa upp originalexemplaren av ansökningsbilagorna.
Du ska besöka beskickningen inom tre månader efter att ha gjort ansökan på internet.
Ansökningen kan tas för behandling först när du har besökt beskickningen.
Vanligtvis måste du boka en tid hos beskickningen i förväg.
Kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan kommer detta att meddelas via ditt konto.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du också lämna in en pappersansökan jämte bilagor vid Finlands beskickning närmast dig.
Du kan skriva ut ansökningsblanketten på Migrationsverkets webbplats.
Handläggning av tillståndsansökan är avgiftsbelagd.
Du betalar avgiften när du lämnar in din tillståndsansökan.
Läs mer om att grunda ett företag på InfoFinlands sida Att grunda ett företag.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Finsk personbeteckning
När du ansöker om ditt första uppehållstillstånd i Finland kan du även be om att bli registrerad i Finlands befolkningsdatasystem.
Då får du en finsk personbeteckning på samma gång som du får uppehållstillståndet.
Mer information om personbeteckningen hittar du på InfoFinlands sida Registrering som invånare.
Företagare i Finland
På InfoFinlands sida Arbete och entreprenörskap hittar du mer information avsedd för företagare och arbetstagare.
Guide om att grunda ett företagfinska _ engelska _ kinesiska
Tjänster för företagare-Startup Kitfinska
Migrationsverket:Presentation av e-tjänsten Enter Finland
Uppehållstillstånd för arbetstagare
Andra uppehållstillstånd för förvärvsarbete
Uppehållstillstånd för säsongsarbete
Arbete med ett annat uppehållstillstånd
Ansökan om uppehållstillstånd
Arbete utan uppehållstillstånd
Arbetstagare i Finland
Den här sidan är avsedd för dig som är medborgare i något annat land är ett EU-land, Norge, Island, Schweiz eller Liechtenstein.
Om du kommer till Finland för att arbeta behöver du ett uppehållstillstånd.
Innan du kan få ett uppehållstillstånd måste du hitta ett jobb i Finland.
När du har hittat ett jobb kan du ansöka om uppehållstillstånd.
Du måste ansöka om uppehållstillstånd innan du kommer till Finland.
För att kunna arbeta i Finland behöver du vanligen antingen ett uppehållstillstånd för arbetstagare eller någon annan typ av uppehållstillstånd för förvärvsarbete.
Arten av det arbete du ska utföra påverkar typen av tillstånd.
Uppehållstillstånd för arbetstagare
Om du inte kan arbeta med stöd av ett annat uppehållstillstånd eller utan uppehållstillstånd behöver du ett uppehållstillstånd för arbetstagare (työntekijän oleskelulupa).
Uppehållstillstånd för arbetstagare är inte nödvändigt för alla arbetsuppgifter.
Du kan granska hurudant uppehållstillstånd du behöver från Migrationsverkets webbplats.
Du behöver uppehållstillstånd för arbetstagare om du arbetar till exempel som:
städare
hemvårdare eller barnskötare.
Migrationsverket beslutar om du ska beviljas uppehållstillstånd eller inte.
Ett delbeslut av arbets- och näringsbyrån behövs också för tillståndet.
Uppehållstillstånd för arbetstagarefinska _ svenska _ engelska
Andra uppehållstillstånd för förvärvsarbete
För vissa arbetsuppgifter behöver du inte ett uppehållstillstånd för arbetstagare, men du behöver dock ett uppehållstillstånd som beviljas för vissa uppdrag.
Dessa uppdrag kan vara till exempel:
uppdrag inom företagsledning
uppdrag som sakkunnig
forskaruppdrag
uppdrag inom vetenskap, kultur och konst
arbetspraktik.
Migrationsverket beslutar om du får uppehållstillstånd eller inte.
Ett delbeslut av arbets- och näringsbyrån behövs inte för tillståndet.
Arbete i Finlandfinska _ svenska _ engelska
Uppehållstillstånd för säsongsarbete
Om du ska utföra säsongsarbete i Finland behöver du ett säsongsarbetstillstånd.
Säsongsarbetet kan pågå högst nio månader.
Säsongsarbete är till exempel:
växtodling
skogsvårdsarbete
festivalarbete
Om du kommer från ett viseringspliktigt land och ska arbeta i under tre månader, måste du ansöka om ett säsongsarbetsvisum hos den finländska beskickningen.
Om ditt arbete pågår över tre månader ska du ansöka om ett säsongsarbetstillstånd hos Migrationsverket.
Tillstånd för säsongsarbetefinska _ svenska _ engelska
Arbete med ett annat uppehållstillstånd
Om du redan har uppehållstillstånd i Finland utifrån en annan grund, till exempel familjeband, kan du ha rätt att arbeta i Finland.
Då behöver du inte ett separat uppehållstillstånd för att arbeta.
Du kan kontrollera om du har rätt att arbeta i Finland från ditt uppehållstillståndskort eller beslut om uppehållstillstånd.
Rätt att arbetafinska _ svenska _ engelska
Om du har avlagt examen i Finland kan du få ett tillfälligt uppehållstillstånd för att söka arbete.
Detta tillstånd kan beviljas endast som ett fortsatt tillstånd till ett uppehållstillstånd för studerande.
Ansök om tillståndet innan ditt uppehållstillstånd för studerande löper ut.
Du kan få ett tillstånd för högst ett år.
Detta tillstånd kan man endast få en gång.
Om du hittar en arbetsplats, kan du börja arbeta genast.
Du måste ansöka om ett nytt uppehållstillstånd på grund av arbete innan ditt uppehållstillstånd för att söka arbete går ut.
Om du har avlagt examen i Finland, behövs inte ett delbeslut av arbets- och näringsbyrån för ditt tillstånd.
Uppehållstillstånd för sökande av arbetefinska _ svenska _ engelska
Ansökan om uppehållstillstånd
Du måste ansöka om ditt första uppehållstillstånd innan du kommer till Finland.
Du kan ansöka om tillståndet på internet via tjänsten Enter Finland.
När du ställt ansökan ska du besöka Finlands beskickning närmast dig för att styrka din identitet och visa upp originalexemplaren av ansökningsbilagorna.
Du ska besöka beskickningen inom tre månader efter att ha gjort ansökan på internet.
Ansökningen kan tas för behandling först när du besökt beskickningen.
Vanligtvis måste du boka en tid hos beskickningen i förväg.
Kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan kommer detta att meddelas via ditt konto.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du också lämna in en pappersansökan jämte bilagor vid Finlands beskickning närmast dig.
Du kan skriva ut ansökningsblanketten på Migrationsverkets webbplats.
Handläggningen av din ansökan om tillstånd är avgiftsbelagd.
Du måste betala avgiften när du lämnar in ansökan om uppehållstillstånd.
Till ansökan om uppehållstillstånd för arbetstagare ska du bifoga blanketten TEM054 som din arbetsgivare fyller i och undertecknar.
Arbetsgivaren kan lämna uppgifterna om arbetet och sitt företag själv samt följa handläggning av ansökan direkt via tjänsten Enter Finland.
Arbetsgivaren kan även betala handläggningsavgiften för arbetstagaren.
Fråga din arbetsgivare som hen använder tjänsten Enter Finland för arbetsgivare.
Kom ändå ihåg att arbetsgivaren inte kan ansöka om uppehållstillstånd för dig, utan hen kompletterar din ansökan för egen del i tjänsten Enter Finland.
Så länge handläggningen av din första ansökan om uppehållstillstånd pågår har du inte rätt att arbeta.
Om du har ansökt om uppehållstillstånd utomlands, kan du inte komma till Finland innan tillstånd har beviljats.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Handläggningstider för tillståndsansökningarfinska _ svenska _ engelska
Ansökan om uppehållstillstånd för specialist
Om du ska arbeta i Finland som specialist kan du även komma till Finland utan uppehållstillstånd.
Du måste dock ha visum eller rätt att vistas i Finland tre månader utan visum.
Du ska också ha en arbetsplats som uppfyller kraven.
Om du arbetar i Finland längre än tre månader måste du ansöka om uppehållstillstånd.
Du kan ansöka om tillståndet elektroniskt via tjänsten Enter Finland eller på Migrationsverkets tjänsteställe.
Finsk personbeteckning
När du ansöker om ditt första uppehållstillstånd i Finland kan du även be om att bli registrerad i Finlands befolkningsdatasystem.
Då får du en finsk personbeteckning på samma gång som du får uppehållstillståndet.
Mer information om personbeteckningen hittar du på InfoFinlands sida Registrering som invånare.
Arbete utan uppehållstillstånd
Oberoende av vilket land du är medborgare i kan du i vissa fall arbeta i Finland utan uppehållstillstånd.
Du måste dock ha ett visum, om du behöver visum till Finland.
Du kan arbeta i Finland utan uppehållstillstånd till exempel om:
du kommer till Finland för att arbeta som tolk, lärare, sakkunnig eller idrottsdomare i högst tre månader utifrån en inbjudan eller ett avtal;
du är fast anställd vid ett företag som bedriver verksamhet i ett annat EU/EES-land och ska komma till Finland för att utföra tillfälligt leverans- eller underleveransarbete och ditt arbete pågår högst tre månader;
du är asylsökande i Finland och har ett giltigt resedokument som berättigar till gränsövergång.
Trots att du inte har uppehållstillstånd kan du börja arbeta tre månader efter att du har lämnat in din asylansökan;
du är asylsökande i Finland och har inte ett giltigt resedokument som berättigar till gränsövergång.
Trots att du inte har uppehållstillstånd kan du börja arbeta när du vistats i sex månader i landet.
Du kan granska om du har rätt att arbeta i Finland utan uppehållstillstånd från Migrationsverkets webbplats.
Arbete utan uppehållstillståndfinska _ svenska _ engelska
Arbetstagare i Finland
På InfoFinlands sida Var hittar jag jobb? finns information om hur du kan hitta ett jobb i Finland.
InfoFinlands sidor Arbete och entreprenörskap innehåller mer information för arbetstagare och företagare.
linkkiArbets- och näringsministeriet:
Arbeta i Finlandfinska _ svenska _ engelska
linkkiArbets- och näringsbyrån:
Broschyren Jobba i Finland(pdf, 5,51 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ polska
linkkiArbetshälsoinstitutet:
Handboken Jobba i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ kurdiska _ tyska _ thai _ vietnamesiska
Migrationsverket:
Presentation av e-tjänsten Enter Finland
Hur ansöker jag?
Vad behövs för registreringen?
Kan jag bli av med uppehållsrätten?
Registrering av uppehållsrätten för EU-medborgare sker inte per automatik.
Du kan ansöka om registrering av uppehållsrätten om din försörjning i Finland är tryggad.
Den kan vara baserad på ett jobb, studier, företagsverksamhet, familjeband eller tillräckliga medel.
Om du avser att bo i Finland längre än tre månader, måste du registrera din uppehållsrätt hos Migrationsverket (Maahanmuuttovirasto).
Ansökan ska lämnas in senast inom tre månader från datumet för inresa.
Registreringen hos Migrationsverket är inte samma sak som registreringen av din bosättningsort i befolkningsdatasystemet (väestötietojärjestelmä) vid magistraten (maistraatti).
Om din sammanhängande vistelse i Finland är kortare än tre månader behöver du inte registrera vistelsen vid Migrationsverket.
Vistelsetiden på tre månader räknas alltid från det att du varit utanför Finlands gränser.
Läs mer om förutsättningarna på sidan EU-medborgare.
Hur ansöker jag?
Handläggning av ansökan om registrering av uppehållsrätt är avgiftsbelagd.
Du betalar avgiften när du lämnar in din ansökan.
Ansök om registrering av uppehållsrätten för EU-medborgare i tjänsten Enter Finland:
Fyll i ansökningsblanketten och bifoga erforderliga bilagor.
Du hittar information om vilka bilagor som behövs till ansökningen i avsnittet
Vad behövs för registreringen?
Besök Migrationsverkets tjänsteställe; du måste styrka din identitet och visa upp originalexemplaren av ansökningsbilagorna.
Ta med dig ett giltigt ID-kort eller pass.
Du ska besöka tjänstestället inom tre månader efter att ha gjort ansökan.
Det är bra att boka en tid på tjänstestället i förväg.
Boka tiden via Migrationsverkets elektroniska tidsbokningssystem.
Kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Om det behövs ytterligare utredningar för din ansökan, kommer detta att meddelas via ditt Enter Finland-konto.
Du får också ett meddelande när beslutet är klart.
Om du inte kan eller inte vet hur du ska göra ansökan på internet:
Gör registreringsansökan på en pappersblankett.
Du kan även göra det personligen på Migrationsverkets tjänsteställe.
Gör ansökan inom tre månader efter datumet för inresa.
Skriv ut registreringsblanketten på Migrationsverkets webbplats och fyll i den färdigt.
Var noga när du fyller i ansökan.
Felaktigt ifyllda ansökningar tas inte emot.
Boka en tid på Migrationsverkets tjänsteställe i det elektroniska tidsbokningssystemet.
Det är bra att boka en tid på tjänstestället i förväg.
Ta med dig den ifyllda registreringsblanketten, ett giltigt ID-kort eller pass och erforderliga bilagor.
Du hittar information om vilka bilagor som behövs till ansökningen i avsnittet
Vad behövs för registreringen?
Om kraven på grund och förutsättningar för vistelsen Finland uppfylls, kan du få ett intyg över registrering av uppehållsrätten för medborgare i Europeiska unionen från Migrationsverket.
Registreringen av uppehållsrätten gäller tillsvidare.
När du har bott lagligt och utan avbrott i Finland i fem år, har du permanent uppehållsrätt.
Permanent uppehållsrätt för EU-medborgare ansöks separat från Migrationsverket.
Registrering av uppehållsrätt för EU-medborgarefinska _ svenska _ engelska
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Permanent uppehållstillståndfinska _ svenska _ engelska
När du ansöker om registrering av uppehållsrätt, kan du på samma blankett också begära att få en finsk personbeteckning.
Då sparas dina personuppgifter, din adress, ditt modersmål och ditt yrke i det finländska befolkningsdatasystemet.
Du behöver ha en personbeteckning när du sköter ärenden med myndigheter.
Det underlättar dessutom skötseln av ärenden i banken och med arbetsgivaren.
Du kan också ansöka om personbeteckning i magistraten (maistraatti) eller skattebyrån (verotoimisto) på din hemort.
Om du flyttar till Finland för att bo här stadigvarande i ett år eller längre, ska du också registrera dig i magistraten på din hemort.
Läs mer på InfoFinlands sida Registrering som invånare.
På InfoFinlands sida Komihåglista för dig som flyttar till Finland hittar du nyttig information om allt som du ska ta hand om när du flyttar till Finland.
Vad behövs för registreringen?
Arbetstagare eller företagare
Din uppehållsrätt kan registreras om du är anställd eller har ett eget företag i Finland.
Du behöver följande handlingar:
EU-registreringsblankett
Giltigt ID-kort eller pass
Anställningsavtal (om du är anställd)
En utredning över företagsverksamheten (om du är egenföretagare)
Studerande
Din uppehållsrätt kan registreras om du studerar vid en läroanstalt som är godkänd i Finland.
Du behöver följande handlingar:
EU-registreringsblankett
Giltigt ID-kort eller pass
Närvarointyg (intyg över att du är studerande vid en läroanstalt som är godkänd i Finland)
Du har en sjukförsäkring (t.ex. det europeiska sjukvårdskortet)
En utredning över din försörjning i Finland
Familjemedlem till en person bosatt i Finland
Din uppehållsrätt kan registreras om du har en familjemedlem som är stadigvarande bosatt i Finland.
Du behöver följande handlingar:
EU-registreringsblankett
Giltigt ID-kort eller pass
Intyg över äktenskap eller registrerat parförhållande
En utredning över att ni har bott tillsammans i två år eller har gemensam vårdnad om ett barn, om du är i ett samboförhållande
Barnets födelseattest om du har vårdnaden om ett barn
En utredning över grunden för att den person som ansöker om familjeförening vistas i Finland.
Uppehållskort för en familjemedlem till en EU-medborgare
Om du inte själv är medborgare i ett EU-land, Liechtenstein eller Schweiz men avser att flytta till Finland till en familjemedlem som är EU-medborgare, måste du ansöka om uppehållskort för en familjemedlem till en EU-medborgare.
Du kan ansöka om uppehållskortet elektroniskt via tjänsten Enter Finland eller på Migrationsverkets (Maahanmuuttovirasto) tjänsteställe.
Handläggning av ansökan om uppehållskort är avgiftsbelagd.
Du betalar avgiften när du lämnar in din ansökan.
Du behöver följande handlingar:
Ansökan om uppehållskort
Giltigt pass
Intyg över äktenskap eller registrerat parförhållande
Registreringsintyget för den EU-medborgare, med vem du kommer till Finland
Utredning över släktskapsförhållandet (barn till EU-medborgaren eller andra släktingar som står under dennes vårdnad)
Utredning över samboskap (om du är sambo med EU-medborgaren och ni inte har gemensam vårdnad om barn)
Uppehållskortet för en familjemedlem till en EU-medborgare beviljas för fem år eller en kortare tid om boendet i Finland varar mindre än fem år.
Uppehållskort för EU-medborgares familjemedlemfinska _ svenska _ engelska
Tillräckliga medel
Om din uppehållsrätt inte kan registreras på någon av de ovan nämnda grunderna kan du ansöka om registrering om du har tillräckliga medel för din försörjning i Finland.
Också tillräckliga medel är en grund.
Du behöver följande handlingar:
EU-registreringsblankett
Giltigt ID-kort eller pass
En utredning över att du har tillräckliga medel för din försörjning i Finland.
Kan jag bli av med uppehållsrätten?
Registreringen av uppehållsrätten för en EU-medborgare och uppehållskortet för en familjemedlem till en EU-medborgare kan återkallas eller bli ogiltigt om:
du flyttar permanent från Finland
du har vistats utomlands utan avbrott i två år
du lämnade felaktiga uppgifter när du ansökte om registreringen eller om uppehållskortet för en familjemedlem till en EU-medborgare
du har undanhållit sådan information som skulle kunna ha hindrat dig från att få registreringen eller uppehållskortet
du utvisas från Finland
du får finskt medborgarskap.
Tänk på att ändringar i din livssituation kan påverka din uppehållsrätt.
Om din uppehållsrätt registrerades på basis av arbete, ett aktivt företag, en studieplats, familjeband eller tillräckliga medel, och detta skäl inte längre existerar, kan registreringen återkallas.
Beslut om återkallande eller upphörande av uppehållsrätten fattas av Migrationsverket.
Om du flyttar utomlands
Om du inte vill att ditt uppehållstillstånd eller uppehållskort ska återkallas ska du lämna in en ansökan om detta hos Migrationsverket senast inom två år efter att du har flyttat utomlands.
Återkallande av uppehållsrättfinska _ svenska _ engelska
Arbeta i Finland
Till Finland som företagare
Att studera i Finland
Till familjemedlem i Finland
Kort vistelse i Finland
Om du är medborgare i ett EU-land, Liechtenstein eller Schweiz, behöver du inget uppehållstillstånd eller visum i Finland.
Du kan resa till Finland om du har ett giltigt ID-kort eller pass.
Du har rätt att arbeta, driva ett företag och studera i Finland med lika villkor som finska medborgare.
Du måste själv trygga din försörjning i Finland.
Som EU-medborgare kan du vistas i Finland högst tre månader i sträck utan att registrera din uppehållsrätt.
Om du vill stanna kvar i Finland och registrera dig som invånare, ska du ha ett jobb eller ett aktivt företag, en studieplats, ett långvarigt familjeband eller tillräckliga medel.
Om du avser att bo i Finland i över tre månader, ska du ansöka om Registrering av uppehållsrätten för EU-medborgare hos Migrationsverket.
Ansökan ska ställas senast inom tre månader från datumet för inresa.
Om du flyttar till Finland för att bo här stadigvarande i ett år eller längre, ska du också registrera dig i magistraten på din hemort.
Läs mer på InfoFinlands sida Registrering som invånare.
Om du vistas i Finland tre månader utan avbrott behöver du inte ansöka om registrering av uppehållsrätten.
Vistelsetiden på tre månader räknas alltid från det att du varit utanför Finlands gränser.
linkkiEuropa.eu:
EU-länderfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
linkkiEuropa.eu:
Rådgivning för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
_ skotsk gäliska
linkkiEuropeiska kommissionen:
Europeiska sjukvårdskortetfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Arbeta i Finland
Som EU-medborgare behöver du inget arbetstillstånd i Finland.
Du kan börja jobba direkt när du har kommit till landet.
Hämta ett skattekort på den närmaste skattebyrån (Verotoimisto) och lämna kortet till din arbetsgivare.
Om du ska jobba i Finland i mer än tre månader ska du ansöka om registrering av uppehållsrätten för EU-medborgare i tjänsten Enter Finland eller på Migrationsverkets (Maahanmuuttovirasto) tjänsteställe.
Om du flyttar till Finland för att bo här stadigvarande i minst ett år ska du också registrera dig som invånare i magistraten (maistraatti).
Personbeteckning
Om du kommer till Finland från utlandet för att arbeta, behöver du en finsk personbeteckning.
Du får personbeteckningen på magistraten (maistraatti) eller skattebyrån (verotoimisto).
Ett giltigt ID-kort eller pass
Ditt anställningsavtal
Du kan lämna in begäran om personbeteckning också hos Migrationsverket samtidigt som du ansöker om registrering av uppehållsrätten för EU-medborgare.
Skattekort och skattenummer
Alla som arbetar i Finland ska ha ett skattekort.
Din arbetsgivare behöver kortet för utbetalning av lön och för beskattningen.
Om du jobbar inom byggbranschen behöver du också ett skattenummer (veronumero).
Du får skattekort och skattenummer på den närmaste skattebyrån.
På InfoFinlands sida Arbetstagare eller företagare finns mer information för arbetstagare som flyttar till Finland.
Jobbsökning i Finland
Om du är medborgare i ett EU-land kan du komma till Finland för att söka jobb för en rimlig tid.
Du kan inte registrera dig som invånare i Finland eller ansöka om registrering av uppehållsrätten när du är i landet som jobbsökande.
För att kunna bo kvar i Finland ska du ha ett jobb eller någon av de ovan nämnda anledningarna samt tillräckliga medel för din försörjning i Finland.
På InfoFinlands sida Var hittar jag jobb?
finns information om hur du kan hitta ett jobb i Finland.
Om du har rätt till arbetslöshetsersättning i ditt hemland, kan du även få den tillfälligt utbetald till Finland.
Du kan ansöka om utbetalning av arbetslöshetsersättning till Finland med blankett E303 eller U2.
Du får blanketten hos arbetskraftsmyndigheten i ditt hemland.
Om du kommer till Finland för att söka jobb kan du vanligtvis inte få arbetslöshetsersättning från Finland.
linkkiEuropa.eu:
Ta med dig dina arbetslöshetsförmånerfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
_ lettiska
_ litauiska
_ danska
_ bulgariska
_ slovakiska
_ grekiska
_ tjeckiska
Till Finland som företagare
Som EU-medborgare kan du starta ett företag i Finland om du är stadigvarande bosatt i ett land som hör till Europeiska ekonomiska samarbetsområdet (EES).
Också ett utländskt företag kan starta verksamhet i Finland.
Om din vistelse i Finland varar mer än tre månader ska du ansöka om registrering av uppehållsrätten för EU-medborgare i tjänsten Enter Finland eller på Migrationsverkets (maahanmuuttovirasto) tjänsteställe.
Om du flyttar till Finland för att bo här stadigvarande i minst ett år ska du också registrera dig som invånare i magistraten.
Etableringsanmälan
När du registrerar ditt företag för första gången ska du fylla i en etableringsanmälan och skicka in erforderliga bilagor.
Du behöver eventuellt bifoga till etableringsanmälan också ett utdrag som motsvarar handelsregisterutdraget i Finland, som en myndighet i ditt hemland utfärdar.
I InfoFinlands avsnitt Arbete och entreprenörskap hittar du mycket information om arbetslivet och företagande i Finland.
Som företagare till Finland:
Vilka tillstånd behöver du?(pdf, 384 kt)finska _ engelska
linkkiPatent- och registerstyrelsen:
Anmälan om grundande av ett företagfinska _ svenska _ engelska
Att studera i Finland
Som EU-medborgare kan du ansöka om studieplats vid en läroanstalt som är godkänd i Finland.
Om din vistelse i Finland varar mer än tre månader utan avbrott ska du ansöka om registrering av uppehållsrätten för EU-medborgare i tjänsten Enter Finland eller på Migrationsverkets (Maahanmuuttovirasto) tjänsteställe.
Om du flyttar till Finland för att bo här stadigvarande i minst ett år ska du också registrera dig som invånare i magistraten (maistraatti).
Om du vistas i Finland tre månader utan avbrott behöver du inte ansöka om registrering av uppehållsrätten.
Vistelsetiden på tre månader räknas alltid från det att du varit utanför Finlands gränser.
Denna regel gäller till exempel utbytesstudenter som endast studerar en kort period i Finland (t.ex. fyra månader).
Om du lämnar Finland under vistelsen och inte stannar i landet tre månader utan avbrott, behöver du inte ansöka om registrering av uppehållsrätten.
I detta fall ska du ansöka om en finsk personbeteckning och meddela din adress till magistraten (maistraatti).
På InfoFinlands sida Studerande finns mer information för studerande som flyttar till Finland.
Till familjemedlem i Finland
Om du är EU-medborgare och flyttar till Finland för att bo hos en familjemedlem ska du ansöka om registrering av uppehållsrätten för EU-medborgare på grund av familjeband i tjänsten Enter Finland eller på Migrationsverkets (Maahanmuuttovirasto) tjänsteställe.
Om du inte är EU-medborgare men din familjemedlem som bor i Finland är EU-medborgare, behöver du ett uppehållskort för en familjemedlem till en EU-medborgare.
Du ansöker om kortet i tjänsten Enter Finland eller vid Migrationsverkets (Maahanmuuttovirasto) tjänsteställe.
Om du flyttar till Finland för att bo här stadigvarande ska du också registrera dig som invånare i magistraten (maistraatti).
För registrering av en familjemedlem till en EU-medborgare krävs också att den person som är bosatt i Finland har tillräckliga medel för att försörja sig själv och sin familjemedlem som ska flytta till Finland.
Familjemedlemmar och andra anhöriga kan vara:
Din sambo som du har bott tillsammans med i minst två år eller med vilken du har gemensam vårdnad om ett barn
Ett barn eller barnbarn under 21 år som är beroende av dig för sin försörjning
Ett barn eller barnbarn under 21 år som är beroende av din sambo för sin försörjning
Din förälder eller mor- eller farförälder som är beroende av dig för sin försörjning
Din förälder eller mor- eller farförälder som är beroende av din sambo för sin försörjning
En förälder till ett barn under 21 år
Också ett barn som föds i Finland och blir medborgare i ett EU-land, Liechtenstein eller Schweiz måste ansöka om registrering av uppehållsrätten.
Registrering ska ansökas inom tre månader efter att barnet föddes.
Läs mer om detta på InfoFinlands sida När ett barn föds i Finland.
När du flyttar till Finland på grund av familjeband, har du obegränsad rätt att arbeta och studera i Finland.
På InfoFinlands sida Familjemedlem finns mer information för dem som flyttar till Finland på grund av familjeskäl.
Kort vistelse i Finland
Som EU-medborgare kan du komma till Finland om du har ett pass eller ett ID-kort förutsatt att du inte har utfärdats ett inreseförbud.
Om du vistas i Finland tillfälligt, kan du få en finsk personbeteckning om det behövs till exempel på grund av ditt arbete.
Du kan hämta en personbeteckning och samtidigt registrera ditt tillfälliga boende i den närmaste magistraten (maistraatti) eller skattebyrån (verotoimisto).
Ta med dig ett giltigt ID-kort eller pass.
Om din tillfälliga vistelse varar i över tre månader, behöver du också ett intyg över registrering av uppehållsrätten för medborgare i Europeiska unionen.
Läs mer om ämnet: Registrering av uppehållsrätten för EU-medborgare.
Om du bor i Finland tillfälligt, registreras ingen hemkommun för dig i Finland och du har inte samma rättigheter som de personer som bor i Finland stadigvarande.
Resor i Finland
Om du är medborgare i ett EU-land, Liechtenstein eller Schweiz och vill resa till Finland för en kort period, till exempel på semester, på affärsresa eller för att besöka släktingar, behöver du inget visum.
Du kan resa till Finland om du har ett giltigt ID-kort eller pass.
Om du är i Finland som turist och råkar ut för någon besvärlig situation, kontakta ditt hemlands beskickning.
Beskickningen kan hjälpa dig om du har råkat ut för en olycka, blivit sjuk eller blivit utsatt för ett brott.
Beskickningen kan också utförda dig ett nytt pass om du har tappat bort eller blivit bestulen på ditt pass.
linkkiVisitFinland.com:
Information om Finland till turistersvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ japanska _ italienska
Andra länders beskickningar i Finlandfinska _ svenska _ engelska
Visste du..?
Lokal information
På Infobankens sidor hittar du mycket information om tjänsterna på olika orter.
lokal-information
Kom med och bygg framtidens InfoFinland!
Som medlem i InfoFinlands användarpanel kan du påverka utvecklingen av webbtjänsten InfoFinland, som finns översatt till flera språk.
Användarpanelen är öppen för alla som är intresserade av InfoFinland.
Vi hoppas på att hitta medlemmar med olika modersmål och i olika åldrar i Finland och andra länder.
Gå med i InfoFinlands användarpanel här:
Hur fungerar användarpanelen?
För användarpanelen behöver vi din e-postadress.
Vi skickar ut korta webbenkäter högst varannan månad som rör innehållet i InfoFinland, webbplatsen eller kommunikation.
Din e-post används inte för några andra syften.
Enkäterna är oftast på engelska, ibland även på andra språk.
Några gånger per år lottar vi ut priser bland alla som svarat.
Medlemskapet i panelen binder dig inte till någonting.
Du kan även lämna panelen när som helst.
Registerbeskrivning
Registerbeskrivning för InfoFinland finns på Helsingfors stads webbplats.
Registerbeskrivning:
Kom med och bygg framtidens InfoFinland!
Som medlem i InfoFinlands användarpanel kan du påverka utvecklingen av webbtjänsten InfoFinland, som finns översatt till flera språk.
Användarpanelen är öppen för alla som är intresserade av InfoFinland.
Vi hoppas på att hitta medlemmar med olika modersmål och i olika åldrar i Finland och andra länder.
Gå med i InfoFinlands användarpanel här:
Hur fungerar användarpanelen?
För användarpanelen behöver vi din e-postadress.
Vi skickar ut korta webbenkäter högst varannan månad som rör innehållet i InfoFinland, webbplatsen eller kommunikation.
Din e-post används inte för några andra syften.
Enkäterna är oftast på engelska, ibland även på andra språk.
Några gånger per år lottar vi ut priser bland alla som svarat.
Medlemskapet i panelen binder dig inte till någonting.
Du kan även lämna panelen när som helst.
Registerbeskrivning
Registerbeskrivning för InfoFinland finns på Helsingfors stads webbplats.
Registerbeskrivning:
Kom med och bygg framtidens InfoFinland!
Som medlem i InfoFinlands användarpanel kan du påverka utvecklingen av webbtjänsten InfoFinland, som finns översatt till flera språk.
Användarpanelen är öppen för alla som är intresserade av InfoFinland.
Vi hoppas på att hitta medlemmar med olika modersmål och i olika åldrar i Finland och andra länder.
Gå med i InfoFinlands användarpanel här:
Hur fungerar användarpanelen?
För användarpanelen behöver vi din e-postadress.
Vi skickar ut korta webbenkäter högst varannan månad som rör innehållet i InfoFinland, webbplatsen eller kommunikation.
Din e-post används inte för några andra syften.
Enkäterna är oftast på engelska, ibland även på andra språk.
Några gånger per år lottar vi ut priser bland alla som svarat.
Medlemskapet i panelen binder dig inte till någonting.
Du kan även lämna panelen när som helst.
Registerbeskrivning
Registerbeskrivning för InfoFinland finns på Helsingfors stads webbplats.
Registerbeskrivning:
Register över stadskansliets kundkommunikation, marknadsföring och evenemangshanteringfinska _ svenska _ engelska
Tjänsten InfoFinland.fi upprätthålls av Helsingfors stad.
Staden har åtagit sig att sörja för integritetsskyddet för användarna av stadens webbtjänster.
Vi följer automatiskt besökarna i tjänsten och använder informationen till att utveckla tjänsten.
Med hjälp av uppföljningen vet vi till exempel följande:
Hur många besökare webbplatsen har
Hur mycket de olika sidorna används
På vilka språk webbplatsen används
Hur länge användarna stannar kvar på sidorna
Hur användarna rör sig på webbplatsen
I vilket land användarna befinner sig
Med vilka apparater och webbläsare sidorna används
Vi använder cookies
På webbplatsen används cookies.
Vi följer användningen av sidorna, men samlar inte in några sådana uppgifter som kan kopplas till en person.
Användaren kan förhindra användningen av cookies i sina webbläsarinställningar.
Förändringen kan påverka webbplatsens funktionalitet.
På sidorna finns inbäddat innehåll som producerats av andra.
Integritetsskyddet för till exempel sociala mediers och videokanalers innehåll åligger producentorganisationen.
Tjänsten InfoFinland.fi upprätthålls av Helsingfors stad.
Staden har åtagit sig att sörja för integritetsskyddet för användarna av stadens webbtjänster.
Vi följer automatiskt besökarna i tjänsten och använder informationen till att utveckla tjänsten.
Med hjälp av uppföljningen vet vi till exempel följande:
Hur många besökare webbplatsen har
Hur mycket de olika sidorna används
På vilka språk webbplatsen används
Hur länge användarna stannar kvar på sidorna
Hur användarna rör sig på webbplatsen
I vilket land användarna befinner sig
Med vilka apparater och webbläsare sidorna används
Vi använder cookies
På webbplatsen används cookies.
Vi följer användningen av sidorna, men samlar inte in några sådana uppgifter som kan kopplas till en person.
Användaren kan förhindra användningen av cookies i sina webbläsarinställningar.
Förändringen kan påverka webbplatsens funktionalitet.
På sidorna finns inbäddat innehåll som producerats av andra.
Integritetsskyddet för till exempel sociala mediers och videokanalers innehåll åligger producentorganisationen.
Tjänsten InfoFinland.fi upprätthålls av Helsingfors stad.
Staden har åtagit sig att sörja för integritetsskyddet för användarna av stadens webbtjänster.
Vi följer automatiskt besökarna i tjänsten och använder informationen till att utveckla tjänsten.
Med hjälp av uppföljningen vet vi till exempel följande:
Hur många besökare webbplatsen har
Hur mycket de olika sidorna används
På vilka språk webbplatsen används
Hur länge användarna stannar kvar på sidorna
Hur användarna rör sig på webbplatsen
I vilket land användarna befinner sig
Med vilka apparater och webbläsare sidorna används
Vi använder cookies
På webbplatsen används cookies.
Vi följer användningen av sidorna, men samlar inte in några sådana uppgifter som kan kopplas till en person.
Användaren kan förhindra användningen av cookies i sina webbläsarinställningar.
Förändringen kan påverka webbplatsens funktionalitet.
På sidorna finns inbäddat innehåll som producerats av andra.
Integritetsskyddet för till exempel sociala mediers och videokanalers innehåll åligger producentorganisationen.
Skicka oss respons på InfoFinlands webbplats via länken ”Ge respons på denna sida” nedan!
Längst ner på varje undersida i InfoFinland hittar du en responslänk, via vilken du kan skicka respons som direkt berör innehållet på sidan.
Vi svarar på responsen på följande språk: finska, svenska och engelska.
Skicka oss respons på InfoFinlands webbplats via länken ”Ge respons på denna sida” nedan!
Längst ner på varje undersida i InfoFinland hittar du en responslänk, via vilken du kan skicka respons som direkt berör innehållet på sidan.
Vi svarar på responsen på följande språk: finska, svenska och engelska.
Skicka oss respons på InfoFinlands webbplats via länken ”Ge respons på denna sida” nedan!
Längst ner på varje undersida i InfoFinland hittar du en responslänk, via vilken du kan skicka respons som direkt berör innehållet på sidan.
Vi svarar på responsen på följande språk: finska, svenska och engelska.
Infobankens videotävling är avslutad.
Min Infobank – fem tips för dig som flyttar till Finland
Infobanken bjuder in alla som flyttat till Finland till videotävlingen ”Min Infobank – fem tips för dig som flyttar till Finland”.
Delta i tävlingen med ditt eget videoklipp!
Instruktioner
Gå in på sidan www.infopankki.fi och bekanta dig med Infobankens webbplats.
Gör ditt eget videoklipp med rubriken ”Min Infobank – fem tips för dig som flyttar till Finland”.
Berätta på ditt sätt vad som är bra att veta när man ska flytta till Finland.
Det kan till exempel vara vardagliga tips om arbete, studier, tillståndsärenden, boende eller språkinlärning.
Filmklippet ska vara 1–3 minuter långt.
Gör videoklippet på något av de språk som används i Infobanken.
Språken i Infobanken är finska, svenska, engelska, ryska, estniska, franska, serbokroatiska, somaliska, spanska, turkiska, albanska, kinesiska, kurdiska (sorani), persiska och arabiska.
Använd inte material, såsom bakgrundsmusik eller bilder, som en tredje part har upphovsrätt till.
Skapa dig ett YouTube-konto och ladda upp videoklippet på YouTube.
Skicka länken till ditt videoklipp och dina kontaktuppgifter till Infobanken till adressen infopankki@hel.fi.
Vi hoppas att få se videoklipp från personer i olika livssituationer, med olika yrken och av studerande.
Vi hoppas att få se känslofyllda, intelligenta, smarta och roliga videoklipp.
Du kan delta i tävlingen fram till den 1 december 2013.
Regler
Uppgifter om medverkande:
Ange i slutet av videoklippet namnen på samtliga personer som medverkat i skapandet av videoklippet.
Om flera personer har medverkat ska man i sluttexterna ange en ansvarig person som fyllt 15 år.
Denna person ansvarar i sista hand för att de tillstånd som krävs för att göra videoklippet skaffas, att tillstånden är vederbörliga, att eventuellt material i videoklippet som en tredje part har upphovsrätt till används vederbörligt samt för eventuella upphovsrättsavgifter och upphovsrättsliga krav.
Upphovsrätt:
Använd inte material, såsom bakgrundsmusik eller bilder, som en tredje part har upphovsrätt till.
Observera att tävlingsdeltagaren ansvarar för att verket eller en del av verket, till exempel musik eller bilder, som skickas till tävlingen inte gör intrång på en tredje parts upphovsrätt, varumärkesrätt eller immateriella rättighet.
Tävlingsarrangören ansvarar inte för krav som tredje parter ställer, och som hänför sig till avtalsvidrig användning, kopiering, modifiering eller spridning av material, som utgör en del av verket, eller till någon annan motsvarande orsak.
Sändaren (upphovsmannen) ansvarar för att han eller hon har rätt att överlåta upphovsrätten till verket som skickas till tävlingen.
Mer information om upphovsrätt finns på adresserna www.teosto.fi, www.kopiosto.fi, www.gramex.fi, www.tuotos.fi.
Om videoklippet/verket innehåller material, vars upphovsrätt innehas av en tredje part, ska upphovsmannen säkerställa att han eller hon har vederbörliga tillstånd till att använda materialet.
Upphovsmannen/den ansvariga personen ansvarar för alla eventuella upphovsrätts- och lagringsavgifter och rättsliga krav från tredje parter.
Upphovsrätten till verket förblir i upphovsmannens ägo.
Kränkande eller osakligt innehåll
Videoklipp som inte anknyter till tävlingens tema eller är osakliga på andra sätt godkänns inte.
Videoklippet får inte vara kränkande, nedsättande eller diskriminerande mot kön, etniskt ursprung eller religiös övertygelse.
Videoklippet ska vara i enlighet med Finlands lag och följa god sed.
Personer som uppträder i videoklippet och tillstånd
Sändaren ska inhämta ett skriftligt tillstånd för offentlig visning av videoklippet av samtliga personer som uppträder i videoklippet och kan identifieras, samt av de personer som medverkat i framställningen av videoklippet.
För minderåriga barn krävs tillstånd av deras vårdnadshavare.
Sändaren ska inhämta skriftliga tillstånd för framställning av videoklippet och för tillverkning av kopior av samtliga personer som medverkat i framställningen av videoklippet.
Det är tillåtet att spela in material på offentliga platser, för inspelning i privata lokaler ska tillstånd inhämtas.
Rättigheter
Upphovsmannen som deltar i tävlingen överlåter till tävlingsarrangören, Helsingfors stad, obegränsad rätt att kostnadsfritt visa verket offentligt och att utnyttja verket eller delar av verket i sin marknadsföring av Infobanken på Internet och i andra motsvarande medier samt internationella evenemang.
Videoklippen kan publiceras bland annat på Infobankens webbplats och på Infobankens YouTube-kanal.
Upphovsmannen som deltar i tävlingen överlåter rätten att kopiera verket och ändra verkets format och storlek i den omfattning som krävs för att visa verket.
Val av tävlingens vinnare och pris
Infobankens redaktion utser tävlingens vinnare i samråd med Infobankens användarråd.
Vinnaren belönas med en tabletdator.
Godkännande av reglerna
Sändaren/upphovsmannen till verket godkänner dessa regler genom att skicka in videoklippet till tävlingen.
Infobankens videotävling är avslutad.
Min Infobank – fem tips för dig som flyttar till Finland
Infobanken bjuder in alla som flyttat till Finland till videotävlingen ”Min Infobank – fem tips för dig som flyttar till Finland”.
Delta i tävlingen med ditt eget videoklipp!
Instruktioner
Gå in på sidan www.infopankki.fi och bekanta dig med Infobankens webbplats.
Gör ditt eget videoklipp med rubriken ”Min Infobank – fem tips för dig som flyttar till Finland”.
Berätta på ditt sätt vad som är bra att veta när man ska flytta till Finland.
Det kan till exempel vara vardagliga tips om arbete, studier, tillståndsärenden, boende eller språkinlärning.
Filmklippet ska vara 1–3 minuter långt.
Gör videoklippet på något av de språk som används i Infobanken.
Språken i Infobanken är finska, svenska, engelska, ryska, estniska, franska, serbokroatiska, somaliska, spanska, turkiska, albanska, kinesiska, kurdiska (sorani), persiska och arabiska.
Använd inte material, såsom bakgrundsmusik eller bilder, som en tredje part har upphovsrätt till.
Skapa dig ett YouTube-konto och ladda upp videoklippet på YouTube.
Skicka länken till ditt videoklipp och dina kontaktuppgifter till Infobanken till adressen infopankki@hel.fi.
Vi hoppas att få se videoklipp från personer i olika livssituationer, med olika yrken och av studerande.
Vi hoppas att få se känslofyllda, intelligenta, smarta och roliga videoklipp.
Du kan delta i tävlingen fram till den 1 december 2013.
Regler
Uppgifter om medverkande:
Ange i slutet av videoklippet namnen på samtliga personer som medverkat i skapandet av videoklippet.
Om flera personer har medverkat ska man i sluttexterna ange en ansvarig person som fyllt 15 år.
Denna person ansvarar i sista hand för att de tillstånd som krävs för att göra videoklippet skaffas, att tillstånden är vederbörliga, att eventuellt material i videoklippet som en tredje part har upphovsrätt till används vederbörligt samt för eventuella upphovsrättsavgifter och upphovsrättsliga krav.
Upphovsrätt:
Använd inte material, såsom bakgrundsmusik eller bilder, som en tredje part har upphovsrätt till.
Observera att tävlingsdeltagaren ansvarar för att verket eller en del av verket, till exempel musik eller bilder, som skickas till tävlingen inte gör intrång på en tredje parts upphovsrätt, varumärkesrätt eller immateriella rättighet.
Tävlingsarrangören ansvarar inte för krav som tredje parter ställer, och som hänför sig till avtalsvidrig användning, kopiering, modifiering eller spridning av material, som utgör en del av verket, eller till någon annan motsvarande orsak.
Sändaren (upphovsmannen) ansvarar för att han eller hon har rätt att överlåta upphovsrätten till verket som skickas till tävlingen.
Mer information om upphovsrätt finns på adresserna www.teosto.fi, www.kopiosto.fi, www.gramex.fi, www.tuotos.fi.
Om videoklippet/verket innehåller material, vars upphovsrätt innehas av en tredje part, ska upphovsmannen säkerställa att han eller hon har vederbörliga tillstånd till att använda materialet.
Upphovsmannen/den ansvariga personen ansvarar för alla eventuella upphovsrätts- och lagringsavgifter och rättsliga krav från tredje parter.
Upphovsrätten till verket förblir i upphovsmannens ägo.
Kränkande eller osakligt innehåll
Videoklipp som inte anknyter till tävlingens tema eller är osakliga på andra sätt godkänns inte.
Videoklippet får inte vara kränkande, nedsättande eller diskriminerande mot kön, etniskt ursprung eller religiös övertygelse.
Videoklippet ska vara i enlighet med Finlands lag och följa god sed.
Personer som uppträder i videoklippet och tillstånd
Sändaren ska inhämta ett skriftligt tillstånd för offentlig visning av videoklippet av samtliga personer som uppträder i videoklippet och kan identifieras, samt av de personer som medverkat i framställningen av videoklippet.
För minderåriga barn krävs tillstånd av deras vårdnadshavare.
Sändaren ska inhämta skriftliga tillstånd för framställning av videoklippet och för tillverkning av kopior av samtliga personer som medverkat i framställningen av videoklippet.
Det är tillåtet att spela in material på offentliga platser, för inspelning i privata lokaler ska tillstånd inhämtas.
Rättigheter
Upphovsmannen som deltar i tävlingen överlåter till tävlingsarrangören, Helsingfors stad, obegränsad rätt att kostnadsfritt visa verket offentligt och att utnyttja verket eller delar av verket i sin marknadsföring av Infobanken på Internet och i andra motsvarande medier samt internationella evenemang.
Videoklippen kan publiceras bland annat på Infobankens webbplats och på Infobankens YouTube-kanal.
Upphovsmannen som deltar i tävlingen överlåter rätten att kopiera verket och ändra verkets format och storlek i den omfattning som krävs för att visa verket.
Val av tävlingens vinnare och pris
Infobankens redaktion utser tävlingens vinnare i samråd med Infobankens användarråd.
Vinnaren belönas med en tabletdator.
Godkännande av reglerna
Sändaren/upphovsmannen till verket godkänner dessa regler genom att skicka in videoklippet till tävlingen.
Infobankens videotävling är avslutad.
Min Infobank – fem tips för dig som flyttar till Finland
Infobanken bjuder in alla som flyttat till Finland till videotävlingen ”Min Infobank – fem tips för dig som flyttar till Finland”.
Delta i tävlingen med ditt eget videoklipp!
Instruktioner
Gå in på sidan www.infopankki.fi och bekanta dig med Infobankens webbplats.
Gör ditt eget videoklipp med rubriken ”Min Infobank – fem tips för dig som flyttar till Finland”.
Berätta på ditt sätt vad som är bra att veta när man ska flytta till Finland.
Det kan till exempel vara vardagliga tips om arbete, studier, tillståndsärenden, boende eller språkinlärning.
Filmklippet ska vara 1–3 minuter långt.
Gör videoklippet på något av de språk som används i Infobanken.
Språken i Infobanken är finska, svenska, engelska, ryska, estniska, franska, serbokroatiska, somaliska, spanska, turkiska, albanska, kinesiska, kurdiska (sorani), persiska och arabiska.
Använd inte material, såsom bakgrundsmusik eller bilder, som en tredje part har upphovsrätt till.
Skapa dig ett YouTube-konto och ladda upp videoklippet på YouTube.
Skicka länken till ditt videoklipp och dina kontaktuppgifter till Infobanken till adressen infopankki@hel.fi.
Vi hoppas att få se videoklipp från personer i olika livssituationer, med olika yrken och av studerande.
Vi hoppas att få se känslofyllda, intelligenta, smarta och roliga videoklipp.
Du kan delta i tävlingen fram till den 1 december 2013.
Regler
Uppgifter om medverkande:
Ange i slutet av videoklippet namnen på samtliga personer som medverkat i skapandet av videoklippet.
Om flera personer har medverkat ska man i sluttexterna ange en ansvarig person som fyllt 15 år.
Denna person ansvarar i sista hand för att de tillstånd som krävs för att göra videoklippet skaffas, att tillstånden är vederbörliga, att eventuellt material i videoklippet som en tredje part har upphovsrätt till används vederbörligt samt för eventuella upphovsrättsavgifter och upphovsrättsliga krav.
Upphovsrätt:
Använd inte material, såsom bakgrundsmusik eller bilder, som en tredje part har upphovsrätt till.
Observera att tävlingsdeltagaren ansvarar för att verket eller en del av verket, till exempel musik eller bilder, som skickas till tävlingen inte gör intrång på en tredje parts upphovsrätt, varumärkesrätt eller immateriella rättighet.
Tävlingsarrangören ansvarar inte för krav som tredje parter ställer, och som hänför sig till avtalsvidrig användning, kopiering, modifiering eller spridning av material, som utgör en del av verket, eller till någon annan motsvarande orsak.
Sändaren (upphovsmannen) ansvarar för att han eller hon har rätt att överlåta upphovsrätten till verket som skickas till tävlingen.
Mer information om upphovsrätt finns på adresserna www.teosto.fi, www.kopiosto.fi, www.gramex.fi, www.tuotos.fi.
Om videoklippet/verket innehåller material, vars upphovsrätt innehas av en tredje part, ska upphovsmannen säkerställa att han eller hon har vederbörliga tillstånd till att använda materialet.
Upphovsmannen/den ansvariga personen ansvarar för alla eventuella upphovsrätts- och lagringsavgifter och rättsliga krav från tredje parter.
Upphovsrätten till verket förblir i upphovsmannens ägo.
Kränkande eller osakligt innehåll
Videoklipp som inte anknyter till tävlingens tema eller är osakliga på andra sätt godkänns inte.
Videoklippet får inte vara kränkande, nedsättande eller diskriminerande mot kön, etniskt ursprung eller religiös övertygelse.
Videoklippet ska vara i enlighet med Finlands lag och följa god sed.
Personer som uppträder i videoklippet och tillstånd
Sändaren ska inhämta ett skriftligt tillstånd för offentlig visning av videoklippet av samtliga personer som uppträder i videoklippet och kan identifieras, samt av de personer som medverkat i framställningen av videoklippet.
För minderåriga barn krävs tillstånd av deras vårdnadshavare.
Sändaren ska inhämta skriftliga tillstånd för framställning av videoklippet och för tillverkning av kopior av samtliga personer som medverkat i framställningen av videoklippet.
Det är tillåtet att spela in material på offentliga platser, för inspelning i privata lokaler ska tillstånd inhämtas.
Rättigheter
Upphovsmannen som deltar i tävlingen överlåter till tävlingsarrangören, Helsingfors stad, obegränsad rätt att kostnadsfritt visa verket offentligt och att utnyttja verket eller delar av verket i sin marknadsföring av Infobanken på Internet och i andra motsvarande medier samt internationella evenemang.
Videoklippen kan publiceras bland annat på Infobankens webbplats och på Infobankens YouTube-kanal.
Upphovsmannen som deltar i tävlingen överlåter rätten att kopiera verket och ändra verkets format och storlek i den omfattning som krävs för att visa verket.
Val av tävlingens vinnare och pris
Infobankens redaktion utser tävlingens vinnare i samråd med Infobankens användarråd.
Vinnaren belönas med en tabletdator.
Godkännande av reglerna
Sändaren/upphovsmannen till verket godkänner dessa regler genom att skicka in videoklippet till tävlingen.
Kontaktuppgifter till InfoFinlands redaktion:
Vi tar gärna emot respons på och utvecklingsidéer med koppling till InfoFinlands verksamhet, översättningarna och samarbetsmöjligheter.
Om du behöver hjälp eller råd i skötseln av dina personliga ärenden, ta då direkt kontakt med myndigheterna.
Vi har samlat kontaktuppgifter till myndigheterna på InfoFinlands sida Ring och fråga om råd.
PB 1
Kontaktuppgifter till InfoFinlands redaktion:
Vi tar gärna emot respons på och utvecklingsidéer med koppling till InfoFinlands verksamhet, översättningarna och samarbetsmöjligheter.
Om du behöver hjälp eller råd i skötseln av dina personliga ärenden, ta då direkt kontakt med myndigheterna.
Vi har samlat kontaktuppgifter till myndigheterna på InfoFinlands sida Ring och fråga om råd.
PB 1
Kontaktuppgifter till InfoFinlands redaktion:
Vi tar gärna emot respons på och utvecklingsidéer med koppling till InfoFinlands verksamhet, översättningarna och samarbetsmöjligheter.
Om du behöver hjälp eller råd i skötseln av dina personliga ärenden, ta då direkt kontakt med myndigheterna.
Vi har samlat kontaktuppgifter till myndigheterna på InfoFinlands sida Ring och fråga om råd.
PB 1
