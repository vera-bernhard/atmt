��R�      ]�(�numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i4�����R�(K�<�NNNJ����J����K t�b�CX  �      �t�bhhK ��h��R�(KK��h�C8      �   :   �     
      "   S     *         �t�bhhK ��h��R�(KK��h�C@   �        �   �  ;   -   
   *   4      J   S        �t�bhhK ��h��R�(KK��h�C8      �   }   d      �     *      �  �        �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C(      <            �t�bhhK ��h��R�(KK��h�C       �   �     \        �t�bhhK ��h��R�(KK��h�CD
      5   �      s  	   w   �      0      �               �t�bhhK ��h��R�(KK��h�C0      �            �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C(      <            �t�bhhK ��h��R�(KK��h�C      \        �t�bhhK ��h��R�(KK��h�CL
      5        �     ?   B  	         =   W       9         �t�bhhK ��h��R�(KK��h�C\�      W    "   �   \  y      p     F              y      �     F        �t�bhhK ��h��R�(KK��h�C(      <      �        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C    *      D   �   �        �t�bhhK ��h��R�(KK��h�CT              �   �  -   
      4   "   �       �   &   �   �  ;         �t�bhhK ��h��R�(KK	��h�C$�   �      �  B  X  �         �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�  Y     �t�bhhK ��h��R�(KK��h�C�   G      �t�bhhK ��h��R�(KK��h�CP
      5   +      V      �     �        	   �   }                  �t�bhhK ��h��R�(KK��h�C<      �   }   \  y      �     /     �  �        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C    
   4                 �t�bhhK ��h��R�(KK��h�C   "        �        �t�bhhK ��h��R�(KK��h�C      L         -        �t�bhhK ��h��R�(KK&��h�C�      -   �   �          �     �           �     �   b  �     �  y                  �   �        y      r              �t�bhhK ��h��R�(KK
��h�C(�         C  	   }  �           �t�bhhK ��h��R�(KK��h�CT
      5   �  s  	   w   �      *   0           D  )  }  *           �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C(      <      D     �t�bhhK ��h��R�(KK��h�C�         �   �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C 0                       �t�bhhK ��h��R�(KK��h�C         �   G         �t�bhhK ��h��R�(KK��h�C 9     �   G      1         �t�bhhK ��h��R�(KK��h�C@�     �                  E      �      �      �     �t�bhhK ��h��R�(KK��h�C    
   4                 �t�bhhK ��h��R�(KK��h�C4  G      �t�bhhK ��h��R�(KK��h�C<                  O      +      �     �        �t�bhhK ��h��R�(KK��h�C<�      �  �   :  4  G      ?     �  �           �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�C4
      5      �	  �  	   w   �      �         �t�bhhK ��h��R�(KK��h�CT      D   �   }      �   
      5   '         
     
      �  �        �t�bhhK ��h��R�(KK	��h�C$   �         *   Q   2         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Ct                 �t�bhhK ��h��R�(KK��h�C0�  Z     �      t     �     9         �t�bhhK ��h��R�(KK��h�C�      ~   q  �        �t�bhhK ��h��R�(KK��h�C t     [                 �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�C8=   L     �     N      _            �        �t�bhhK ��h��R�(KK��h�C8   L  6  �  	   ]     �  A  ^  ?   �        �t�bhhK ��h��R�(KK��h�C0   *      ^   Q     >   �     �         �t�bhhK ��h��R�(KK��h�C0      �   }         Q       �        �t�bhhK ��h��R�(KK��h�Cc            �     �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK	��h�C$         N      u  $         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cj  �                  �t�bhhK ��h��R�(KK��h�CT     �t�bhhK ��h��R�(KK��h�C0   *      W  �   v   B      �  $         �t�bhhK ��h��R�(KK��h�C\
      �         -   �  z      �   e   �   �   �  9      ~   q     �           �t�bhhK ��h��R�(KK	��h�C$      7         �  2         �t�bhhK ��h��R�(KK��h�C         T        �t�bhhK ��h��R�(KK��h�C�      ~   q  �        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�      ~   q        �t�bhhK ��h��R�(KK��h�C`  a                 �t�bhhK ��h��R�(KK��h�C�   Y      �t�bhhK ��h��R�(KK��h�C<*      �   >   ;      �   	      F   �              �t�bhhK ��h��R�(KK��h�C8Y      "   �  S     *   "   �      �  ;         �t�bhhK ��h��R�(KK��h�C0      i   
   ;      �	  d   H   %        �t�bhhK ��h��R�(KK��h�C8      
   �      �   7         *   Q            �t�bhhK ��h��R�(KK��h�C*         �t�bhhK ��h��R�(KK��h�C �    �  	   �     1     �t�bhhK ��h��R�(KK��h�C(      <            �t�bhhK ��h��R�(KK��h�C         �   Y      �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C �                        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C      �                 �t�bhhK ��h��R�(KK��h�C'   �  $      �t�bhhK ��h��R�(KK��h�C\
      "   '   �  $         =   �           r   �   �  �     �              �t�bhhK ��h��R�(KK��h�Cl�      �        '   �  $         &                 \                                 �t�bhhK ��h��R�(KK��h�C         '   �  $      �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                  �t�bhhK ��h��R�(KK��h�C�     *      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�   G      �t�bhhK ��h��R�(KK��h�C4  G      �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�C�   Y      �t�bhhK ��h��R�(KK��h�C4�   �   �   
   .      �   
      �   M        �t�bhhK ��h��R�(KK��h�CD�   �      F         �  �     N     �        L        �t�bhhK ��h��R�(KK��h�C,�   4   �   
   .   4         M        �t�bhhK ��h��R�(KK��h�C<
      "   J   S     *         �  :   �   �        �t�bhhK ��h��R�(KK��h�C4�   �   8     5  	   �  	   Q     �         �t�bhhK ��h��R�(KK��h�CP
      4   "   �      :   �   �  	         g   +         �   �        �t�bhhK ��h��R�(KK��h�C0      �   �  �      �  3  ~  %        �t�bhhK ��h��R�(KK��h�C         G         �t�bhhK ��h��R�(KK��h�C�     *      �t�bhhK ��h��R�(KK
��h�C(�   �   8     �     )           �t�bhhK ��h��R�(KK
��h�C(�  "   �   \     �     /        �t�bhhK ��h��R�(KK��h�C0   �     �  N  	   O     P  Q        �t�bhhK ��h��R�(KK
��h�C(      �   }      �   �   ]         �t�bhhK ��h��R�(KK��h�C0   *   Q   2      P     �     �        �t�bhhK ��h��R�(KK��h�C4N      �  �   	   �  r   �  4               �t�bhhK ��h��R�(KK��h�C4r   �     �        �                   �t�bhhK ��h��R�(KK��h�C      }      �        �t�bhhK ��h��R�(KK��h�CX
      4      �     �  	             �  J   }            �     p        �t�bhhK ��h��R�(KK��h�C@
      5   �  �  s  	         �     �   �            �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Ct                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C,      a             �   �         �t�bhhK ��h��R�(KK��h�CLD   :   Y      4   "   �      &   �   �     1      �   �   5        �t�bhhK ��h��R�(KK��h�C0      �   �   �      %  �  3  ~        �t�bhhK ��h��R�(KK��h�C    *      ^   �   *        �t�bhhK ��h��R�(KK��h�C0�      �   @  7         F      �        �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C�   �                 �t�bhhK ��h��R�(KK��h�C�   �                 �t�bhhK ��h��R�(KK��h�C-     �t�bhhK ��h��R�(KK��h�C4   
   �     -  7         j   �   �        �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�CL   9      3  X  	   v   Y      �     1   �   >     @   �        �t�bhhK ��h��R�(KK
��h�C(�      3  X     v     Q        �t�bhhK ��h��R�(KK��h�C03  X  �  4   Q     �     W   {        �t�bhhK ��h��R�(KK��h�C4       �  Q  �  4   �  �      �  �        �t�bhhK ��h��R�(KK
��h�C(l     3  X     9      �        �t�bhhK ��h��R�(KK
��h�C(�  �        �        @        �t�bhhK ��h��R�(KK��h�C@�     �           E      �      �      �     �     �t�bhhK ��h��R�(KK��h�C         �      1      �t�bhhK ��h��R�(KK	��h�C$�     ?   B  "   �   �        �t�bhhK ��h��R�(KK��h�C4�     z        �     �      �           �t�bhhK ��h��R�(KK��h�C,&   |  �      �         W  �         �t�bhhK ��h��R�(KK��h�C8�   &   R  �     (          U     �         �t�bhhK ��h��R�(KK��h�C�      W  �      �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C@      $   ?   /  I         W        �     9         �t�bhhK ��h��R�(KK	��h�C$   5   4   �   }      �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C         �      1      �t�bhhK ��h��R�(KK��h�Cn   G      �t�bhhK ��h��R�(KK��h�CX   �     C     �     H  $   O   B   +            �     0     @        �t�bhhK ��h��R�(KK��h�C<#        �   
   f      @   +      �     $         �t�bhhK ��h��R�(KK��h�C8   �  6      z                  .   6         �t�bhhK ��h��R�(KK��h�C0   *      ^   Q     >   �     �         �t�bhhK ��h��R�(KK	��h�C$j  �         *   Q   2         �t�bhhK ��h��R�(KK��h�C0      �   }         Q       �        �t�bhhK ��h��R�(KK��h�CL
   '   $     �     5   s  o   	   w   �      �      )           �t�bhhK ��h��R�(KK��h�C �  "   �   
   �  G         �t�bhhK ��h��R�(KK��h�CT?   �     B     �      $   ?   /  I      W  �         �     9         �t�bhhK ��h��R�(KK��h�C0      D   w   r   $         �   �        �t�bhhK ��h��R�(KK��h�C         n   G         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C   �                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cj  �                  �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Ct                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK
��h�C(   
   �     �                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CX  �      �t�bhhK ��h��R�(KK��h�C8      �   :   �     
      "   S     *         �t�bhhK ��h��R�(KK��h�C@   �        �   �  ;   -   
   *   4      J   S        �t�bhhK ��h��R�(KK��h�C8      �   }   d      �     *      �  �        �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C(      <            �t�bhhK ��h��R�(KK��h�C       �   �     \        �t�bhhK ��h��R�(KK��h�CD
      5   �      s  	   w   �      0      �               �t�bhhK ��h��R�(KK��h�C0      �            �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C(      <            �t�bhhK ��h��R�(KK��h�C      \        �t�bhhK ��h��R�(KK��h�CL
      5        �     ?   B  	         =   W       9         �t�bhhK ��h��R�(KK��h�C\�      W    "   �   \  y      p     F              y      �     F        �t�bhhK ��h��R�(KK��h�C(      <      �        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C    *      D   �   �        �t�bhhK ��h��R�(KK��h�CT              �   �  -   
      4   "   �       �   &   �   �  ;         �t�bhhK ��h��R�(KK	��h�C$�   �      �  B  X  �         �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�  Y     �t�bhhK ��h��R�(KK��h�C�   G      �t�bhhK ��h��R�(KK��h�CP
      5   +      V      �     �        	   �   }                  �t�bhhK ��h��R�(KK��h�C<      �   }   \  y      �     /     �  �        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C    
   4                 �t�bhhK ��h��R�(KK��h�C   "        �        �t�bhhK ��h��R�(KK��h�C      L         -        �t�bhhK ��h��R�(KK&��h�C�      -   �   �          �     �           �     �   b  �     �  y                  �   �        y      r              �t�bhhK ��h��R�(KK
��h�C(�         C  	   }  �           �t�bhhK ��h��R�(KK��h�CT
      5   �  s  	   w   �      *   0           D  )  }  *           �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C(      <      D     �t�bhhK ��h��R�(KK��h�C�         �   �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C 0                       �t�bhhK ��h��R�(KK��h�C         �   G         �t�bhhK ��h��R�(KK��h�C 9     �   G      1         �t�bhhK ��h��R�(KK��h�C@�     �                  E      �      �      �     �t�bhhK ��h��R�(KK��h�C    
   4                 �t�bhhK ��h��R�(KK��h�C4  G      �t�bhhK ��h��R�(KK��h�C<                  O      +      �     �        �t�bhhK ��h��R�(KK��h�C<�      �  �   :  4  G      ?     �  �           �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�C4
      5      �	  �  	   w   �      �         �t�bhhK ��h��R�(KK��h�CT      D   �   }      �   
      5   '         
     
      �  �        �t�bhhK ��h��R�(KK	��h�C$   �         *   Q   2         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Ct                 �t�bhhK ��h��R�(KK��h�C0�  Z     �      t     �     9         �t�bhhK ��h��R�(KK��h�C�      ~   q  �        �t�bhhK ��h��R�(KK��h�C t     [                 �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�C8=   L     �     N      _            �        �t�bhhK ��h��R�(KK��h�C8   L  6  �  	   ]     �  A  ^  ?   �        �t�bhhK ��h��R�(KK��h�C0   *      ^   Q     >   �     �         �t�bhhK ��h��R�(KK��h�C0      �   }         Q       �        �t�bhhK ��h��R�(KK��h�Cc            �     �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK	��h�C$         N      u  $         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cj  �                  �t�bhhK ��h��R�(KK��h�CT     �t�bhhK ��h��R�(KK��h�C0   *      W  �   v   B      �  $         �t�bhhK ��h��R�(KK��h�C\
      �         -   �  z      �   e   �   �   �  9      ~   q     �           �t�bhhK ��h��R�(KK	��h�C$      7         �  2         �t�bhhK ��h��R�(KK��h�C         T        �t�bhhK ��h��R�(KK��h�C�      ~   q  �        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�      ~   q        �t�bhhK ��h��R�(KK��h�C`  a                 �t�bhhK ��h��R�(KK��h�C�   Y      �t�bhhK ��h��R�(KK��h�C<*      �   >   ;      �   	      F   �              �t�bhhK ��h��R�(KK��h�C8Y      "   �  S     *   "   �      �  ;         �t�bhhK ��h��R�(KK��h�C0      i   
   ;      �	  d   H   %        �t�bhhK ��h��R�(KK��h�C8      
   �      �   7         *   Q            �t�bhhK ��h��R�(KK��h�C*         �t�bhhK ��h��R�(KK��h�C �    �  	   �     1     �t�bhhK ��h��R�(KK��h�C(      <            �t�bhhK ��h��R�(KK��h�C�               �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C      �                 �t�bhhK ��h��R�(KK��h�C'   �  $      �t�bhhK ��h��R�(KK��h�C\
      "   '   �  $         =   �           r   �   �  �     �              �t�bhhK ��h��R�(KK��h�Cl�      �        '   �  $         &                 \                                 �t�bhhK ��h��R�(KK��h�C         '   �  $      �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                  �t�bhhK ��h��R�(KK��h�C�     *      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�   G      �t�bhhK ��h��R�(KK��h�C4  G      �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�C�   Y      �t�bhhK ��h��R�(KK��h�C4�   �   �   
   .      �   
      �   M        �t�bhhK ��h��R�(KK��h�CD�   �      F         �  �     N     �        L        �t�bhhK ��h��R�(KK��h�C,�   4   �   
   .   4         M        �t�bhhK ��h��R�(KK��h�C<
      "   J   S     *         �  :   �   �        �t�bhhK ��h��R�(KK��h�C4�   �   8     5  	   �  	   Q     �         �t�bhhK ��h��R�(KK��h�CP
      4   "   �      :   �   �  	         g   +         �   �        �t�bhhK ��h��R�(KK��h�C0      �   �  �      �  3  ~  %        �t�bhhK ��h��R�(KK��h�C         G         �t�bhhK ��h��R�(KK��h�C�     *      �t�bhhK ��h��R�(KK
��h�C(�   �   8     �     )           �t�bhhK ��h��R�(KK
��h�C(�  "   �   \     �     /        �t�bhhK ��h��R�(KK��h�C0   �     �  N  	   O     P  Q        �t�bhhK ��h��R�(KK
��h�C(      �   }      �   �   ]         �t�bhhK ��h��R�(KK��h�C0   *   Q   2      P     �     �        �t�bhhK ��h��R�(KK��h�C4N      �  �   	   �  r   �  4               �t�bhhK ��h��R�(KK��h�C4r   �     �        �                   �t�bhhK ��h��R�(KK��h�C      }      �        �t�bhhK ��h��R�(KK��h�CX
      4      �     �  	             �  J   }            �     p        �t�bhhK ��h��R�(KK��h�C@
      5   �  �  s  	         �     �   �            �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Ct                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C,      a             �   �         �t�bhhK ��h��R�(KK��h�CLD   :   Y      4   "   �      &   �   �     1      �   �   5        �t�bhhK ��h��R�(KK��h�C0      �   �   �      %  �  3  ~        �t�bhhK ��h��R�(KK��h�C    *      ^   �   *        �t�bhhK ��h��R�(KK��h�C0�      �   @  7         F      �        �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C�   �                 �t�bhhK ��h��R�(KK��h�C�   �                 �t�bhhK ��h��R�(KK��h�C-     �t�bhhK ��h��R�(KK��h�C4   
   �     -  7         j   �   �        �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�CL   9      3  X  	   v   Y      �     1   �   >     @   �        �t�bhhK ��h��R�(KK
��h�C(�      3  X     v     Q        �t�bhhK ��h��R�(KK��h�C03  X  �  4   Q     �     W   {        �t�bhhK ��h��R�(KK��h�C4       �  Q  �  4   �  �      �  �        �t�bhhK ��h��R�(KK
��h�C(l     3  X     9      �        �t�bhhK ��h��R�(KK
��h�C(�  �        �        @        �t�bhhK ��h��R�(KK��h�C@�     �           E      �      �      �     �     �t�bhhK ��h��R�(KK��h�C         �      1      �t�bhhK ��h��R�(KK	��h�C$�     ?   B  "   �   �        �t�bhhK ��h��R�(KK��h�C4�     z        �     �      �           �t�bhhK ��h��R�(KK��h�C,&   |  �      �         W  �         �t�bhhK ��h��R�(KK��h�C8�   &   R  �     (          U     �         �t�bhhK ��h��R�(KK��h�C�      W  �      �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C@      $   ?   /  I         W        �     9         �t�bhhK ��h��R�(KK	��h�C$   5   4   �   }      �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C         �      1      �t�bhhK ��h��R�(KK��h�Cn   G      �t�bhhK ��h��R�(KK��h�CX   �     C     �     H  $   O   B   +            �     0     @        �t�bhhK ��h��R�(KK��h�C<#        �   
   f      @   +      �     $         �t�bhhK ��h��R�(KK��h�C8   �  6      z                  .   6         �t�bhhK ��h��R�(KK��h�C0   *      ^   Q     >   �     �         �t�bhhK ��h��R�(KK	��h�C$j  �         *   Q   2         �t�bhhK ��h��R�(KK��h�C0      �   }         Q       �        �t�bhhK ��h��R�(KK��h�CL
   '   $     �     5   s  o   	   w   �      �      )           �t�bhhK ��h��R�(KK��h�C �  "   �   
   �  G         �t�bhhK ��h��R�(KK��h�CT?   �     B     �      $   ?   /  I      W  �         �     9         �t�bhhK ��h��R�(KK��h�C0      D   w   r   $         �   �        �t�bhhK ��h��R�(KK��h�C         n   G         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C   �                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cj  �                  �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Ct                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK
��h�C(   
   �     �                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CX  �      �t�bhhK ��h��R�(KK��h�C8      �   :   �     
      "   S     *         �t�bhhK ��h��R�(KK��h�C@   �        �   �  ;   -   
   *   4      J   S        �t�bhhK ��h��R�(KK��h�C8      �   }   d      �     *      �  �        �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C(      <            �t�bhhK ��h��R�(KK��h�C       �   �     \        �t�bhhK ��h��R�(KK��h�CD
      5   �      s  	   w   �      0      �               �t�bhhK ��h��R�(KK��h�C0      �            �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C(      <            �t�bhhK ��h��R�(KK��h�C      \        �t�bhhK ��h��R�(KK��h�CL
      5        �     ?   B  	         =   W       9         �t�bhhK ��h��R�(KK��h�C\�      W    "   �   \  y      p     F              y      �     F        �t�bhhK ��h��R�(KK��h�C(      <      �        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C    *      D   �   �        �t�bhhK ��h��R�(KK��h�CT              �   �  -   
      4   "   �       �   &   �   �  ;         �t�bhhK ��h��R�(KK	��h�C$�   �      �  B  X  �         �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�  Y     �t�bhhK ��h��R�(KK��h�C�   G      �t�bhhK ��h��R�(KK��h�CP
      5   +      V      �     �        	   �   }                  �t�bhhK ��h��R�(KK��h�C<      �   }   \  y      �     /     �  �        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C    
   4                 �t�bhhK ��h��R�(KK��h�C   "        �        �t�bhhK ��h��R�(KK��h�C      L         -        �t�bhhK ��h��R�(KK&��h�C�      -   �   �          �     �           �     �   b  �     �  y                  �   �        y      r              �t�bhhK ��h��R�(KK
��h�C(�         C  	   }  �           �t�bhhK ��h��R�(KK��h�CT
      5   �  s  	   w   �      *   0           D  )  }  *           �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C(      <      D     �t�bhhK ��h��R�(KK��h�C�         �   �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C 0                       �t�bhhK ��h��R�(KK��h�C         �   G         �t�bhhK ��h��R�(KK��h�C 9     �   G      1         �t�bhhK ��h��R�(KK��h�C@�     �                  E      �      �      �     �t�bhhK ��h��R�(KK��h�C    
   4                 �t�bhhK ��h��R�(KK��h�C4  G      �t�bhhK ��h��R�(KK��h�C<                  O      +      �     �        �t�bhhK ��h��R�(KK��h�C<�      �  �   :  4  G      ?     �  �           �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�C4
      5      �	  �  	   w   �      �         �t�bhhK ��h��R�(KK��h�CT      D   �   }      �   
      5   '         
     
      �  �        �t�bhhK ��h��R�(KK	��h�C$   �         *   Q   2         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Ct                 �t�bhhK ��h��R�(KK��h�C0�  Z     �      t     �     9         �t�bhhK ��h��R�(KK��h�C�      ~   q  �        �t�bhhK ��h��R�(KK��h�C t     [                 �t�bhhK ��h��R�(KK��h�C         K     �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�C8=   L     �     N      _            �        �t�bhhK ��h��R�(KK��h�C8   L  6  �  	   ]     �  A  ^  ?   �        �t�bhhK ��h��R�(KK��h�C0   *      ^   Q     >   �     �         �t�bhhK ��h��R�(KK��h�C0      �   }         Q       �        �t�bhhK ��h��R�(KK��h�Cc            �     �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C          �     T        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cj  �                  �t�bhhK ��h��R�(KK��h�CT     �t�bhhK ��h��R�(KK��h�C0   *      W  �   v   B      �  $         �t�bhhK ��h��R�(KK��h�C\
      �         -   �  z      �   e   �   �   �  9      ~   q     �           �t�bhhK ��h��R�(KK	��h�C$      7         �  2         �t�bhhK ��h��R�(KK��h�C�      ~   q  �        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�      ~   q        �t�bhhK ��h��R�(KK��h�C`  a                 �t�bhhK ��h��R�(KK��h�C�   Y      �t�bhhK ��h��R�(KK��h�C<*      �   >   ;      �   	      F   �              �t�bhhK ��h��R�(KK��h�C8Y      "   �  S     *   "   �      �  ;         �t�bhhK ��h��R�(KK��h�C0      i   
   ;      �	  d   H   %        �t�bhhK ��h��R�(KK��h�C8      
   �      �   7         *   Q            �t�bhhK ��h��R�(KK��h�C*         �t�bhhK ��h��R�(KK��h�C �    �  	   �     1     �t�bhhK ��h��R�(KK��h�C(      <            �t�bhhK ��h��R�(KK��h�C         �   Y      �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C      �                 �t�bhhK ��h��R�(KK��h�C'   �  $      �t�bhhK ��h��R�(KK��h�C\
      "   '   �  $         =   �           r   �   �  �     �              �t�bhhK ��h��R�(KK��h�Cl�      �        '   �  $         &                 \                                 �t�bhhK ��h��R�(KK��h�C         '   �  $      �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                  �t�bhhK ��h��R�(KK��h�C4�  �     4      .   k         "           �t�bhhK ��h��R�(KK��h�C  �   e   k         �t�bhhK ��h��R�(KK��h�C)      �t�bhhK ��h��R�(KK��h�C4�  �     4      .   k         "           �t�bhhK ��h��R�(KK��h�C  �   e   k         �t�bhhK ��h��R�(KK��h�C)      �t�bhhK ��h��R�(KK��h�C4�  �     4      .   k         "           �t�bhhK ��h��R�(KK��h�C  �   e   k         �t�bhhK ��h��R�(KK��h�C)      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK��h�C�     C      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CV           L      �t�bhhK ��h��R�(KK��h�Cz     �t�bhhK ��h��R�(KK��h�CW   �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK
��h�C(   *      �  �     �   �         �t�bhhK ��h��R�(KK��h�C   *      �   l        �t�bhhK ��h��R�(KK	��h�C$�   �     )                  �t�bhhK ��h��R�(KK��h�C8�  
   �  w  �   n    z   6   f     &        �t�bhhK ��h��R�(KK��h�CH
         F   D  O   �         �         i   
   l  �        �t�bhhK ��h��R�(KK��h�C4N      �   
   l  6              x        �t�bhhK ��h��R�(KK	��h�C$      D   g   �  M   �        �t�bhhK ��h��R�(KK��h�CP     �     *      D   g   �     v  $      9   	   !      8         �t�bhhK ��h��R�(KK��h�C,   6   c  �   �   J   `      *         �t�bhhK ��h��R�(KK	��h�C$      O      M   q   �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C`   
   d     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C                   �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C,   *   �       �        U        �t�bhhK ��h��R�(KK	��h�C$�   V     )                  �t�bhhK ��h��R�(KK��h�C,     �  B   a   M   *   Q   2         �t�bhhK ��h��R�(KK��h�C               �t�bhhK ��h��R�(KK��h�Cf     �             �t�bhhK ��h��R�(KK��h�CT   �   :        �         D   =         H         i                 �t�bhhK ��h��R�(KK��h�CP        H   2         �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C `                       �t�bhhK ��h��R�(KK��h�C[   X      �t�be.