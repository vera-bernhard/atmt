��      ]�(�numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i4�����R�(K�<�NNNJ����J����K t�b�C[         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK
��h�C(#         t   �  �  �  �        �t�bhhK ��h��R�(KK��h�C,#         �  �     �  �   �        �t�bhhK ��h��R�(KK��h�C �  �   �  H   )   �        �t�bhhK ��h��R�(KK��h�C4   #   I           �  �  �  �  �        �t�bhhK ��h��R�(KK��h�C �     U   �     Z        �t�bhhK ��h��R�(KK��h�C,&   �  J  �     �  �     �        �t�bhhK ��h��R�(KK��h�C,:   �     �     U   �     Z        �t�bhhK ��h��R�(KK��h�C0#         �     [      �     �        �t�bhhK ��h��R�(KK��h�C@#   �  �      �  �              �   �  �  �        �t�bhhK ��h��R�(KK��h�C,�     �     #      &   ~  �        �t�bhhK ��h��R�(KK��h�C@   #      &   �  �     �     �     �  .  K        �t�bhhK ��h��R�(KK��h�C #      -      �  �        �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C8  ?   �  �  .   �  	   �     �     #         �t�bhhK ��h��R�(KK��h�C,�  "   �     �  �     �          �t�bhhK ��h��R�(KK��h�CH&   "   �  �     �  �     �   e   �  �     �     �        �t�bhhK ��h��R�(KK��h�CT�  �  �     �  �  �     �  	   �  	   L     �  u   -   �  �        �t�bhhK ��h��R�(KK��h�CP�     �  	      �   [  K     �    	   �       �     Z        �t�bhhK ��h��R�(KK��h�Ch&   �  �  �  �  �  �  �  �  �     �     �  &   �  �     �     �  �              �t�bhhK ��h��R�(KK��h�C<�  �  u   �      �  �     �  a   �     �        �t�bhhK ��h��R�(KK��h�C8�  5  �  �   #      K        �     �        �t�bhhK ��h��R�(KK��h�C0�  �  �   e      �  	   �     �        �t�bhhK ��h��R�(KK��h�CP�  �  B   x           �  	     #      �     4   �            �t�bhhK ��h��R�(KK��h�C`I       �     	     �          	   �  M  N  &            	  �        �t�bhhK ��h��R�(KK��h�CX#   �   s     
        �          Z  M  N    �     �             �t�bhhK ��h��R�(KK��h�CPH       �            &   	   O                          �t�bhhK ��h��R�(KK	��h�C$#     u   ?     �   P        �t�bhhK ��h��R�(KK��h�Cd&     Q  �                 Z  	   5           �       M  N          �t�bhhK ��h��R�(KK��h�C4#   �      K    �  M  N               �t�bhhK ��h��R�(KK��h�C�                   �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C#   "   R          �t�bhhK ��h��R�(KK	��h�C$M   #      !  �     r        �t�bhhK ��h��R�(KK��h�C"        H   I        �t�bhhK ��h��R�(KK��h�C,#     �     9        �   �        �t�bhhK ��h��R�(KK��h�C8        �     x  �  $  %  U   #   I        �t�bhhK ��h��R�(KK��h�CH&    -   '   '  	   �  	   (     )  �     &   *  	        �t�bhhK ��h��R�(KK��h�C,#   "   +         �  ,     -        �t�bhhK ��h��R�(KK��h�C,.  /  :   >   0     �      \        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C1     
           �t�bhhK ��h��R�(KK��h�C2           �t�bhhK ��h��R�(KK��h�C3        �t�bhhK ��h��R�(KK��h�C 4                 E      �t�bhhK ��h��R�(KK��h�C5                 �t�bhhK ��h��R�(KK��h�C,�  U   #      �  6                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK	��h�C$   #      ^   >     S        �t�bhhK ��h��R�(KK��h�CH   q   �  �     7     1            
     S  6          �t�bhhK ��h��R�(KK��h�CD&   �      �   �  "   �   �  �        �  �     #         �t�bhhK ��h��R�(KK	��h�C$         #   �   �  2         �t�bhhK ��h��R�(KK��h�C    #         �  �        �t�bhhK ��h��R�(KK��h�CD      
   &   �   8  +     #         �  �   �  2         �t�bhhK ��h��R�(KK
��h�C(         T     �     1         �t�bhhK ��h��R�(KK��h�CU  �   �        �t�bhhK ��h��R�(KK��h�C #   �   �                 �t�bhhK ��h��R�(KK��h�C9  �   �        �t�bhhK ��h��R�(KK��h�C �  �   :           E      �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C0&   ;    <     #      =     �        �t�bhhK ��h��R�(KK��h�C0>     �  ?  �     �  �  �  I         �t�bhhK ��h��R�(KK��h�C0   H   2         
   �     �  �        �t�bhhK ��h��R�(KK��h�C,     �  H       �   �  @        �t�bhhK ��h��R�(KK��h�C8   
   >   �      �      �        H   2         �t�bhhK ��h��R�(KK��h�CPt  |   "   6  A  �       �   �   B     ]     �      V  �  +        �t�bhhK ��h��R�(KK��h�C@   #      C  	   D     E  \   '   f      F  G        �t�bhhK ��h��R�(KK��h�C0         �   H  	        I     1      �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK
��h�C(#         t   �  �  �  �        �t�bhhK ��h��R�(KK��h�C,#         �  �     �  �   �        �t�bhhK ��h��R�(KK��h�C �  �   �  H   )   �        �t�bhhK ��h��R�(KK��h�C4   #   I           �  �  �  �  �        �t�bhhK ��h��R�(KK��h�C �     U   �     Z        �t�bhhK ��h��R�(KK��h�C,&   �  J  �     �  �     �        �t�bhhK ��h��R�(KK��h�C,:   �     �     U   �     Z        �t�bhhK ��h��R�(KK��h�C0#         �     [      �     �        �t�bhhK ��h��R�(KK��h�C@#   �  �      �  �              �   �  �  �        �t�bhhK ��h��R�(KK��h�C,�     �     #      &   ~  �        �t�bhhK ��h��R�(KK��h�C@   #      &   �  �     �     �     �  .  K        �t�bhhK ��h��R�(KK��h�C #      -      �  �        �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C8  ?   �  �  .   �  	   �     �     #         �t�bhhK ��h��R�(KK��h�C,�  "   �     �  �     �          �t�bhhK ��h��R�(KK��h�CH&   "   �  �     �  �     �   e   �  �     �     �        �t�bhhK ��h��R�(KK��h�CT�  �  �     �  �  �     �  	   �  	   L     �  u   -   �  �        �t�bhhK ��h��R�(KK��h�CP�     �  	      �   [  K     �    	   �       �     Z        �t�bhhK ��h��R�(KK��h�Ch&   �  �  �  �  �  �  �  �  �     �     �  &   �  �     �     �  �              �t�bhhK ��h��R�(KK��h�C<�  �  u   �      �  �     �  a   �     �        �t�bhhK ��h��R�(KK��h�C8�  5  �  �   #      K        �     �        �t�bhhK ��h��R�(KK��h�C0�  �  �   e      �  	   �     �        �t�bhhK ��h��R�(KK��h�CP�  �  B   x           �  	     #      �     4   �            �t�bhhK ��h��R�(KK��h�C`I       �     	     �          	   �  M  N  &            	  �        �t�bhhK ��h��R�(KK��h�CX#   �   s     
        �          Z  M  N    �     �             �t�bhhK ��h��R�(KK��h�CPH       �            &   	   O                          �t�bhhK ��h��R�(KK	��h�C$#     u   ?     �   P        �t�bhhK ��h��R�(KK��h�Cd&     Q  �                 Z  	   5           �       M  N          �t�bhhK ��h��R�(KK��h�C4#   �      K    �  M  N               �t�bhhK ��h��R�(KK��h�C�                   �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C#   "   R          �t�bhhK ��h��R�(KK	��h�C$M   #      !  �     r        �t�bhhK ��h��R�(KK��h�C"        H   I        �t�bhhK ��h��R�(KK��h�C,#     �     9        �   �        �t�bhhK ��h��R�(KK��h�C8        �     x  �  $  %  U   #   I        �t�bhhK ��h��R�(KK��h�CH&    -   '   '  	   �  	   (     )  �     &   *  	        �t�bhhK ��h��R�(KK��h�C,#   "   +         �  ,     -        �t�bhhK ��h��R�(KK��h�C,.  /  :   >   0     �      \        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C1     
           �t�bhhK ��h��R�(KK��h�C2           �t�bhhK ��h��R�(KK��h�C3        �t�bhhK ��h��R�(KK��h�C 4                 E      �t�bhhK ��h��R�(KK��h�C5                 �t�bhhK ��h��R�(KK��h�C,�  U   #      �  6                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK	��h�C$   #      ^   >     S        �t�bhhK ��h��R�(KK��h�CH   q   �  �     7     1            
     S  6          �t�bhhK ��h��R�(KK��h�CD&   �      �   �  "   �   �  �        �  �     #         �t�bhhK ��h��R�(KK	��h�C$         #   �   �  2         �t�bhhK ��h��R�(KK��h�C    #         �  �        �t�bhhK ��h��R�(KK��h�CD      
   &   �   8  +     #         �  �   �  2         �t�bhhK ��h��R�(KK
��h�C(         T     �     1         �t�bhhK ��h��R�(KK��h�CU  �   �        �t�bhhK ��h��R�(KK��h�C #   �   �                 �t�bhhK ��h��R�(KK��h�C9  �   �        �t�bhhK ��h��R�(KK��h�C �  �   :           E      �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C0&   ;    <     #      =     �        �t�bhhK ��h��R�(KK��h�C0>     �  ?  �     �  �  �  I         �t�bhhK ��h��R�(KK��h�C0   H   2         
   �     �  �        �t�bhhK ��h��R�(KK��h�C,     �  H       �   �  @        �t�bhhK ��h��R�(KK��h�C8   
   >   �      �      �        H   2         �t�bhhK ��h��R�(KK��h�CPt  |   "   6  A  �       �   �   B     ]     �      V  �  +        �t�bhhK ��h��R�(KK��h�C@   #      C  	   D     E  \   '   f      F  G        �t�bhhK ��h��R�(KK��h�C0         �   H  	        I     1      �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK
��h�C(#         t   �  �  �  �        �t�bhhK ��h��R�(KK��h�C,#         �  �     �  �   �        �t�bhhK ��h��R�(KK��h�C �  �   �  H   )   �        �t�bhhK ��h��R�(KK��h�C4   #   I           �  �  �  �  �        �t�bhhK ��h��R�(KK��h�C �     U   �     Z        �t�bhhK ��h��R�(KK��h�C,&   �  J  �     �  �     �        �t�bhhK ��h��R�(KK��h�C,:   �     �     U   �     Z        �t�bhhK ��h��R�(KK��h�C0#         �     [      �     �        �t�bhhK ��h��R�(KK��h�C@#   �  �      �  �              �   �  �  �        �t�bhhK ��h��R�(KK��h�C,�     �     #      &   ~  �        �t�bhhK ��h��R�(KK��h�C@   #      &   �  �     �     �     �  .  K        �t�bhhK ��h��R�(KK��h�C #      -      �  �        �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C8  ?   �  �  .   �  	   �     �     #         �t�bhhK ��h��R�(KK��h�C,�  "   �     �  �     �          �t�bhhK ��h��R�(KK��h�CH&   "   �  �     �  �     �   e   �  �     �     �        �t�bhhK ��h��R�(KK��h�CT�  �  �     �  �  �     �  	   �  	   L     �  u   -   �  �        �t�bhhK ��h��R�(KK��h�CP�     �  	      �   [  K     �    	   �       �     Z        �t�bhhK ��h��R�(KK��h�Ch&   �  �  �  �  �  �  �  �  �     �     �  &   �  �     �     �  �              �t�bhhK ��h��R�(KK��h�C<�  �  u   �      �  �     �  a   �     �        �t�bhhK ��h��R�(KK��h�C8�  5  �  �   #      K        �     �        �t�bhhK ��h��R�(KK��h�C0�  �  �   e      �  	   �     �        �t�bhhK ��h��R�(KK��h�CP�  �  B   x           �  	     #      �     4   �            �t�bhhK ��h��R�(KK��h�C`I       �     	     �          	   �  M  N  &            	  �        �t�bhhK ��h��R�(KK��h�CX#   �   s     
        �          Z  M  N    �     �             �t�bhhK ��h��R�(KK��h�CPH       �            &   	   O                          �t�bhhK ��h��R�(KK	��h�C$#     u   ?     �   P        �t�bhhK ��h��R�(KK��h�Cd&     Q  �                 Z  	   5           �       M  N          �t�bhhK ��h��R�(KK��h�C4#   �      K    �  M  N               �t�bhhK ��h��R�(KK��h�C�                   �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C#   "   R          �t�bhhK ��h��R�(KK	��h�C$M   #      !  �     r        �t�bhhK ��h��R�(KK��h�C"        H   I        �t�bhhK ��h��R�(KK��h�C,#     �     9        �   �        �t�bhhK ��h��R�(KK��h�C8        �     x  �  $  %  U   #   I        �t�bhhK ��h��R�(KK��h�CH&    -   '   '  	   �  	   (     )  �     &   *  	        �t�bhhK ��h��R�(KK��h�C,#   "   +         �  ,     -        �t�bhhK ��h��R�(KK��h�C,.  /  :   >   0     �      \        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C1     
           �t�bhhK ��h��R�(KK��h�C2           �t�bhhK ��h��R�(KK��h�C3        �t�bhhK ��h��R�(KK��h�C 4                 E      �t�bhhK ��h��R�(KK��h�C5                 �t�bhhK ��h��R�(KK��h�C,�  U   #      �  6                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK	��h�C$   #      ^   >     S        �t�bhhK ��h��R�(KK��h�CH   q   �  �     7     1            
     S  6          �t�bhhK ��h��R�(KK��h�CD&   �      �   �  "   �   �  �        �  �     #         �t�bhhK ��h��R�(KK	��h�C$         #   �   �  2         �t�bhhK ��h��R�(KK��h�C    #         �  �        �t�bhhK ��h��R�(KK��h�CD      
   &   �   8  +     #         �  �   �  2         �t�bhhK ��h��R�(KK
��h�C(         T     �     1         �t�bhhK ��h��R�(KK��h�CU  �   �        �t�bhhK ��h��R�(KK��h�C #   �   �                 �t�bhhK ��h��R�(KK��h�C9  �   �        �t�bhhK ��h��R�(KK��h�C �  �   :           E      �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C0&   ;    <     #      =     �        �t�bhhK ��h��R�(KK��h�C0>     �  ?  �     �  �  �  I         �t�bhhK ��h��R�(KK��h�C0   H   2         
   �     �  �        �t�bhhK ��h��R�(KK��h�C,     �  H       �   �  @        �t�bhhK ��h��R�(KK��h�C8   
   >   �      �      �        H   2         �t�bhhK ��h��R�(KK��h�CPt  |   "   6  A  �       �   �   B     ]     �      V  �  +        �t�bhhK ��h��R�(KK��h�C@   #      C  	   D     E  \   '   f      F  G        �t�bhhK ��h��R�(KK��h�C0         �   H  	        I     1      �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C4�  �     4      .   k         "           �t�bhhK ��h��R�(KK��h�C  �   e   k         �t�bhhK ��h��R�(KK��h�C)      �t�bhhK ��h��R�(KK��h�C4�  �     4      .   k         "           �t�bhhK ��h��R�(KK��h�C  �   e   k         �t�bhhK ��h��R�(KK��h�C)      �t�bhhK ��h��R�(KK��h�C4�  �     4      .   k         "           �t�bhhK ��h��R�(KK��h�C  �   e   k         �t�bhhK ��h��R�(KK��h�C)      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C    �   a      �      �t�bhhK ��h��R�(KK��h�C�      7     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�     $      L      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C<#         �  J     T   �  �     K             �t�bhhK ��h��R�(KK��h�C\Y   L       �  �     
   �  ?   M  �    �   a      �   �     �          �t�bhhK ��h��R�(KK��h�C,^   �       �  �  �     �        �t�bhhK ��h��R�(KK��h�CT�      �  \   N     �  W  T   �      �     �  \   �  k      �        �t�bhhK ��h��R�(KK��h�C@   O     P        H     Q    �     �  �        �t�bhhK ��h��R�(KK#��h�C�R  �      #      �   e   S  T     �     �  	   �  U     V  	   W  #   X  	   �  Y  \   Z     #      [  #   \        �t�bhhK ��h��R�(KK��h�C4      
   ]     #         #   Q   2         �t�bhhK ��h��R�(KK��h�CL   H   2      -           ^     _     
   H   �     `        �t�bhhK ��h��R�(KK��h�C         X        �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C #   �        H   I        �t�bhhK ��h��R�(KK��h�C<a        b  	   8  	   �  \   Y  c     d        �t�bhhK ��h��R�(KK��h�C0   
     �     ;         �  2         �t�bhhK ��h��R�(KK��h�C     -              �t�bhhK ��h��R�(KK��h�Ctv      Q  e         	   f  Z  	   g  �  �  	   �  h     [       9  ?      \     �         �t�bhhK ��h��R�(KK��h�CPM  N  .   i  j     1      k     �  l         m     #         �t�bhhK ��h��R�(KK��h�C#   �  �  n     �t�bhhK ��h��R�(KK��h�Co  :  	   �   #      �t�bhhK ��h��R�(KK��h�C]      p  	   q     �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�Cr                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK	��h�C$   #      �    �  �         �t�bhhK ��h��R�(KK��h�C,�   �    �     s  t     u        �t�bhhK ��h��R�(KK
��h�C(�      .   �     ^   >   �        �t�bhhK ��h��R�(KK��h�C4�  v     �         w  x     y          �t�bhhK ��h��R�(KK��h�CT�   z  {  	     	   |  	     	     	   }     ~  \                �t�bhhK ��h��R�(KK��h�C0   �   �           
   ]  �  �        �t�bhhK ��h��R�(KK��h�CH   #      �     �  �     >   �  \   �      !  �  �         �t�bhhK ��h��R�(KK��h�C4      
        #         #   Q   2         �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�     "     �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�C    �   a      �      �t�bhhK ��h��R�(KK��h�CP    �   a      �         �     �  �     �     #  ?      �        �t�bhhK ��h��R�(KK��h�Cl   1      B      V      �  �  �     �     �     �   a      �  	      �     �  �        �t�bhhK ��h��R�(KK��h�C0.      4   �      �  �  �  �   �        �t�bhhK ��h��R�(KK��h�C4   L  �  �  	      $     �     �        �t�bhhK ��h��R�(KK��h�C-   �  �  �        �t�bhhK ��h��R�(KK"��h�C��  p   4   �       �  �     �   	   %  �     �  	   �     %  �     �  	   �  �  �   �  >     &  �  �  �        �t�bhhK ��h��R�(KK��h�C\      
   �  	   �  	   �     L     �  \   �  �     #         H   2         �t�bhhK ��h��R�(KK��h�CT�     �  	   �  	   �  	   �       '     #         (             �t�bhhK ��h��R�(KK��h�C0   (  �  -   u   P  )     �           �t�bhhK ��h��R�(KK��h�CD      �   �  ;  #   d   #   �     �  �  	   �   #         �t�bhhK ��h��R�(KK
��h�C(             �   a      �         �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C �                 E      �t�bhhK ��h��R�(KK��h�C�  ;  �           �t�bhhK ��h��R�(KK��h�C     �           �t�bhhK ��h��R�(KK��h�C�      7     �t�bhhK ��h��R�(KK��h�CX#         �     �  �  	      T   �     �  *  �     �  +     �        �t�bhhK ��h��R�(KK��h�C4#   �        .   �  �     ,  �           �t�bhhK ��h��R�(KK��h�C<      �     
   �  +     �  2         �        �t�bhhK ��h��R�(KK��h�CH   #      �  -  .  	   �  <  �  �  �     �     /        �t�bhhK ��h��R�(KK
��h�C(-  .  �     ?   0  �  �        �t�bhhK ��h��R�(KK��h�C          �      7        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C1     �t�bhhK ��h��R�(KK
��h�C(�      �     �                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C@   �     �   	      .   �  �  �  	      �  �        �t�bhhK ��h��R�(KK��h�CT#      �  �  �  2  U      �     �  �  �  �     �     �           �t�bhhK ��h��R�(KK��h�CL   �     3  �     4  ^  U   �     �  �        �  5        �t�bhhK ��h��R�(KK��h�CH-      �    �     �  
   H   �     �     �     ^        �t�bhhK ��h��R�(KK��h�CD   �  �  2            
   �  ;   	   �  \   6  +        �t�bhhK ��h��R�(KK$��h�C�7  �  �  8  .   a       �   .   �  �  �     �     �  z  ^     �     �     \   :   Z   �       :   �  �     9        �t�bhhK ��h��R�(KK��h�C8�     �     �     �  �  �  �  �  �        �t�bhhK ��h��R�(KK��h�CD   8  	   �  =  �  :  U   #   	      �  �     �        �t�bhhK ��h��R�(KK��h�C0      
   �  �      ?   ;  �  �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C �      �                 �t�bhhK ��h��R�(KK��h�C0�  3  �  �   t   3   �                 �t�bhhK ��h��R�(KK
��h�C(�  	   #   �  �                 �t�bhhK ��h��R�(KK��h�C�  �     �        �t�bhhK ��h��R�(KK
��h�C(�  �     �  )                  �t�bhhK ��h��R�(KK��h�C^  �     �t�bhhK ��h��R�(KK��h�C�     $      L      �t�bhhK ��h��R�(KK��h�C,^   �       �  �  �     �        �t�bhhK ��h��R�(KK��h�CT^   >   �   \   �  W  p   L   �      �   �     �  \   �  k      �        �t�bhhK ��h��R�(KK��h�CH$      L      �      [   s      �   	   �  	   �     �        �t�bhhK ��h��R�(KK��h�C �   T   H   <     �        �t�bhhK ��h��R�(KK��h�C,H   <  =  >  �  �   
      #         �t�bhhK ��h��R�(KK��h�Cx:   �     �  �  T   �  +     $      �  :     �     L      �  r     _  I      >   ?     #         �t�bhhK ��h��R�(KK��h�C4   
   �     $      L         H   2         �t�bhhK ��h��R�(KK��h�CXL     �  @  p   6     
   �  �  	   R  	    	  	   G   	   �     �         �t�bhhK ��h��R�(KK��h�CH�   W  T   $      L   >   �     �  	   �     �     �         �t�bhhK ��h��R�(KK��h�C,�  _  �         �     ]  	        �t�bhhK ��h��R�(KK��h�C\#   �      �   �  T   -   �     $      L   	   �  	  	   �  	   	     A        �t�bhhK ��h��R�(KK��h�C,      
   �        #   �  2         �t�bhhK ��h��R�(KK��h�C�  @     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK
��h�C(         �     $      L         �t�bhhK ��h��R�(KK��h�C�  s      �           �t�bhhK ��h��R�(KK��h�C	                 �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�CU  �   �        �t�bhhK ��h��R�(KK��h�C #   �   �                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8#   "   '   	     	  	     |         �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C    �   a      �      �t�bhhK ��h��R�(KK��h�C�      7     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�     $      L      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C<#         �  J     T   �  �     K             �t�bhhK ��h��R�(KK��h�C\Y   L       �  �     
   �  ?   M  �    �   a      �   �     �          �t�bhhK ��h��R�(KK��h�C,^   �       �  �  �     �        �t�bhhK ��h��R�(KK��h�CT�      �  \   N     �  W  T   �      �     �  \   �  k      �        �t�bhhK ��h��R�(KK��h�C@   O     P        H     Q    �     �  �        �t�bhhK ��h��R�(KK#��h�C�R  �      #      �   e   S  T     �     �  	   �  U     V  	   W  #   X  	   �  Y  \   Z     #      [  #   \        �t�bhhK ��h��R�(KK��h�C4      
   ]     #         #   Q   2         �t�bhhK ��h��R�(KK��h�CL   H   2      -           ^     _     
   H   �     `        �t�bhhK ��h��R�(KK��h�C         X        �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C #   �        H   I        �t�bhhK ��h��R�(KK��h�C<a        b  	   8  	   �  \   Y  c     d        �t�bhhK ��h��R�(KK��h�C0   
     �     ;         �  2         �t�bhhK ��h��R�(KK��h�C     -              �t�bhhK ��h��R�(KK��h�Ctv      Q  e         	   f  Z  	   g  �  �  	   �  h     [       9  ?      \     �         �t�bhhK ��h��R�(KK��h�CPM  N  .   i  j     1      k     �  l         m     #         �t�bhhK ��h��R�(KK��h�C#   �  �  n     �t�bhhK ��h��R�(KK��h�Co  :  	   �   #      �t�bhhK ��h��R�(KK��h�C]      p  	   q     �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�Cr                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK	��h�C$   #      �    �  �         �t�bhhK ��h��R�(KK��h�C,�   �    �     s  t     u        �t�bhhK ��h��R�(KK
��h�C(�      .   �     ^   >   �        �t�bhhK ��h��R�(KK��h�C4�  v     �         w  x     y          �t�bhhK ��h��R�(KK��h�CT�   z  {  	     	   |  	     	     	   }     ~  \                �t�bhhK ��h��R�(KK��h�C0   �   �           
   ]  �  �        �t�bhhK ��h��R�(KK��h�CH   #      �     �  �     >   �  \   �      !  �  �         �t�bhhK ��h��R�(KK��h�C4      
        #         #   Q   2         �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�     "     �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�C    �   a      �      �t�bhhK ��h��R�(KK��h�CP    �   a      �         �     �  �     �     #  ?      �        �t�bhhK ��h��R�(KK��h�Cl   1      B      V      �  �  �     �     �     �   a      �  	      �     �  �        �t�bhhK ��h��R�(KK��h�C0.      4   �      �  �  �  �   �        �t�bhhK ��h��R�(KK��h�C4   L  �  �  	      $     �     �        �t�bhhK ��h��R�(KK��h�C-   �  �  �        �t�bhhK ��h��R�(KK"��h�C��  p   4   �       �  �     �   	   %  �     �  	   �     %  �     �  	   �  �  �   �  >     &  �  �  �        �t�bhhK ��h��R�(KK��h�C\      
   �  	   �  	   �     L     �  \   �  �     #         H   2         �t�bhhK ��h��R�(KK��h�CT�     �  	   �  	   �  	   �       '     #         (             �t�bhhK ��h��R�(KK��h�C0   (  �  -   u   P  )     �           �t�bhhK ��h��R�(KK��h�CD      �   �  ;  #   d   #   �     �  �  	   �   #         �t�bhhK ��h��R�(KK
��h�C(             �   a      �         �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C �                 E      �t�bhhK ��h��R�(KK��h�C�  ;  �           �t�bhhK ��h��R�(KK��h�C     �           �t�bhhK ��h��R�(KK��h�C�      7     �t�bhhK ��h��R�(KK��h�CX#         �     �  �  	      T   �     �  *  �     �  +     �        �t�bhhK ��h��R�(KK��h�C4#   �        .   �  �     ,  �           �t�bhhK ��h��R�(KK��h�C<      �     
   �  +     �  2         �        �t�bhhK ��h��R�(KK��h�CH   #      �  -  .  	   �  <  �  �  �     �     /        �t�bhhK ��h��R�(KK
��h�C(-  .  �     ?   0  �  �        �t�bhhK ��h��R�(KK��h�C          �      7        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C1     �t�bhhK ��h��R�(KK
��h�C(�      �     �                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C@   �     �   	      .   �  �  �  	      �  �        �t�bhhK ��h��R�(KK��h�CT#      �  �  �  2  U      �     �  �  �  �     �     �           �t�bhhK ��h��R�(KK��h�CL   �     3  �     4  ^  U   �     �  �        �  5        �t�bhhK ��h��R�(KK��h�CH-      �    �     �  
   H   �     �     �     ^        �t�bhhK ��h��R�(KK��h�CD   �  �  2            
   �  ;   	   �  \   6  +        �t�bhhK ��h��R�(KK$��h�C�7  �  �  8  .   a       �   .   �  �  �     �     �  z  ^     �     �     \   :   Z   �       :   �  �     9        �t�bhhK ��h��R�(KK��h�C8�     �     �     �  �  �  �  �  �        �t�bhhK ��h��R�(KK��h�CD   8  	   �  =  �  :  U   #   	      �  �     �        �t�bhhK ��h��R�(KK��h�C0      
   �  �      ?   ;  �  �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C �      �                 �t�bhhK ��h��R�(KK��h�C0�  3  �  �   t   3   �                 �t�bhhK ��h��R�(KK
��h�C(�  	   #   �  �                 �t�bhhK ��h��R�(KK��h�C�  �     �        �t�bhhK ��h��R�(KK
��h�C(�  �     �  )                  �t�bhhK ��h��R�(KK��h�C^  �     �t�bhhK ��h��R�(KK��h�C�     $      L      �t�bhhK ��h��R�(KK��h�C,^   �       �  �  �     �        �t�bhhK ��h��R�(KK��h�CT^   >   �   \   �  W  p   L   �      �   �     �  \   �  k      �        �t�bhhK ��h��R�(KK��h�CH$      L      �      [   s      �   	   �  	   �     �        �t�bhhK ��h��R�(KK��h�C �   T   H   <     �        �t�bhhK ��h��R�(KK��h�C,H   <  =  >  �  �   
      #         �t�bhhK ��h��R�(KK��h�Cx:   �     �  �  T   �  +     $      �  :     �     L      �  r     _  I      >   ?     #         �t�bhhK ��h��R�(KK��h�C4   
   �     $      L         H   2         �t�bhhK ��h��R�(KK��h�CXL     �  @  p   6     
   �  �  	   R  	    	  	   G   	   �     �         �t�bhhK ��h��R�(KK��h�CH�   W  T   $      L   >   �     �  	   �     �     �         �t�bhhK ��h��R�(KK��h�C,�  _  �         �     ]  	        �t�bhhK ��h��R�(KK��h�C\#   �      �   �  T   -   �     $      L   	   �  	  	   �  	   	     A        �t�bhhK ��h��R�(KK��h�C,      
   �        #   �  2         �t�bhhK ��h��R�(KK��h�C�  @     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK
��h�C(         �     $      L         �t�bhhK ��h��R�(KK��h�C�  s      �           �t�bhhK ��h��R�(KK��h�C	                 �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�CU  �   �        �t�bhhK ��h��R�(KK��h�C #   �   �                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8#   "   '   	     	  	     |         �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C    �   a      �      �t�bhhK ��h��R�(KK��h�C�      7     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�     $      L      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C<#         �  J     T   �  �     K             �t�bhhK ��h��R�(KK��h�C\Y   L       �  �     
   �  ?   M  �    �   a      �   �     �          �t�bhhK ��h��R�(KK��h�C,^   �       �  �  �     �        �t�bhhK ��h��R�(KK��h�CT�      �  \   N     �  W  T   �      �     �  \   �  k      �        �t�bhhK ��h��R�(KK��h�C@   O     P        H     Q    �     �  �        �t�bhhK ��h��R�(KK#��h�C�R  �      #      �   e   S  T     �     �  	   �  U     V  	   W  #   X  	   �  Y  \   Z     #      [  #   \        �t�bhhK ��h��R�(KK��h�C4      
   ]     #         #   Q   2         �t�bhhK ��h��R�(KK��h�CL   H   2      -           ^     _     
   H   �     `        �t�bhhK ��h��R�(KK��h�C         X        �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C #   �        H   I        �t�bhhK ��h��R�(KK��h�C<a        b  	   8  	   �  \   Y  c     d        �t�bhhK ��h��R�(KK��h�C0   
     �     ;         �  2         �t�bhhK ��h��R�(KK��h�C     -              �t�bhhK ��h��R�(KK��h�Ctv      Q  e         	   f  Z  	   g  �  �  	   �  h     [       9  ?      \     �         �t�bhhK ��h��R�(KK��h�CPM  N  .   i  j     1      k     �  l         m     #         �t�bhhK ��h��R�(KK��h�C#   �  �  n     �t�bhhK ��h��R�(KK��h�Co  :  	   �   #      �t�bhhK ��h��R�(KK��h�C]      p  	   q     �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�Cr                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK	��h�C$   #      �    �  �         �t�bhhK ��h��R�(KK��h�C,�   �    �     s  t     u        �t�bhhK ��h��R�(KK
��h�C(�      .   �     ^   >   �        �t�bhhK ��h��R�(KK��h�C4�  v     �         w  x     y          �t�bhhK ��h��R�(KK��h�CT�   z  {  	     	   |  	     	     	   }     ~  \                �t�bhhK ��h��R�(KK��h�C0   �   �           
   ]  �  �        �t�bhhK ��h��R�(KK��h�CH   #      �     �  �     >   �  \   �      !  �  �         �t�bhhK ��h��R�(KK��h�C4      
        #         #   Q   2         �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�     "     �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�C    �   a      �      �t�bhhK ��h��R�(KK��h�CP    �   a      �         �     �  �     �     #  ?      �        �t�bhhK ��h��R�(KK��h�Cl   1      B      V      �  �  �     �     �     �   a      �  	      �     �  �        �t�bhhK ��h��R�(KK��h�C0.      4   �      �  �  �  �   �        �t�bhhK ��h��R�(KK��h�C4   L  �  �  	      $     �     �        �t�bhhK ��h��R�(KK��h�C-   �  �  �        �t�bhhK ��h��R�(KK"��h�C��  p   4   �       �  �     �   	   %  �     �  	   �     %  �     �  	   �  �  �   �  >     &  �  �  �        �t�bhhK ��h��R�(KK��h�C\      
   �  	   �  	   �     L     �  \   �  �     #         H   2         �t�bhhK ��h��R�(KK��h�CT�     �  	   �  	   �  	   �       '     #         (             �t�bhhK ��h��R�(KK��h�C0   (  �  -   u   P  )     �           �t�bhhK ��h��R�(KK��h�CD      �   �  ;  #   d   #   �     �  �  	   �   #         �t�bhhK ��h��R�(KK
��h�C(             �   a      �         �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C �                 E      �t�bhhK ��h��R�(KK��h�C�  ;  �           �t�bhhK ��h��R�(KK��h�C     �           �t�bhhK ��h��R�(KK��h�C�      7     �t�bhhK ��h��R�(KK��h�CX#         �     �  �  	      T   �     �  *  �     �  +     �        �t�bhhK ��h��R�(KK��h�C4#   �        .   �  �     ,  �           �t�bhhK ��h��R�(KK��h�C<      �     
   �  +     �  2         �        �t�bhhK ��h��R�(KK��h�CH   #      �  -  .  	   �  <  �  �  �     �     /        �t�bhhK ��h��R�(KK
��h�C(-  .  �     ?   0  �  �        �t�bhhK ��h��R�(KK��h�C          �      7        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C1     �t�bhhK ��h��R�(KK
��h�C(�      �     �                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C@   �     �   	      .   �  �  �  	      �  �        �t�bhhK ��h��R�(KK��h�CT#      �  �  �  2  U      �     �  �  �  �     �     �           �t�bhhK ��h��R�(KK��h�CL   �     3  �     4  ^  U   �     �  �        �  5        �t�bhhK ��h��R�(KK��h�CH-      �    �     �  
   H   �     �     �     ^        �t�bhhK ��h��R�(KK��h�CD   �  �  2            
   �  ;   	   �  \   6  +        �t�bhhK ��h��R�(KK$��h�C�7  �  �  8  .   a       �   .   �  �  �     �     �  z  ^     �     �     \   :   Z   �       :   �  �     9        �t�bhhK ��h��R�(KK��h�C8�     �     �     �  �  �  �  �  �        �t�bhhK ��h��R�(KK��h�CD   8  	   �  =  �  :  U   #   	      �  �     �        �t�bhhK ��h��R�(KK��h�C0      
   �  �      ?   ;  �  �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C �      �                 �t�bhhK ��h��R�(KK��h�C0�  3  �  �   t   3   �                 �t�bhhK ��h��R�(KK
��h�C(�  	   #   �  �                 �t�bhhK ��h��R�(KK��h�C�  �     �        �t�bhhK ��h��R�(KK
��h�C(�  �     �  )                  �t�bhhK ��h��R�(KK��h�C^  �     �t�bhhK ��h��R�(KK��h�C�     $      L      �t�bhhK ��h��R�(KK��h�C,^   �       �  �  �     �        �t�bhhK ��h��R�(KK��h�CT^   >   �   \   �  W  p   L   �      �   �     �  \   �  k      �        �t�bhhK ��h��R�(KK��h�CH$      L      �      [   s      �   	   �  	   �     �        �t�bhhK ��h��R�(KK��h�C �   T   H   <     �        �t�bhhK ��h��R�(KK��h�C,H   <  =  >  �  �   
      #         �t�bhhK ��h��R�(KK��h�Cx:   �     �  �  T   �  +     $      �  :     �     L      �  r     _  I      >   ?     #         �t�bhhK ��h��R�(KK��h�C4   
   �     $      L         H   2         �t�bhhK ��h��R�(KK��h�CXL     �  @  p   6     
   �  �  	   R  	    	  	   G   	   �     �         �t�bhhK ��h��R�(KK��h�CH�   W  T   $      L   >   �     �  	   �     �     �         �t�bhhK ��h��R�(KK��h�C,�  _  �         �     ]  	        �t�bhhK ��h��R�(KK��h�C\#   �      �   �  T   -   �     $      L   	   �  	  	   �  	   	     A        �t�bhhK ��h��R�(KK��h�C,      
   �        #   �  2         �t�bhhK ��h��R�(KK��h�C�  @     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK
��h�C(         �     $      L         �t�bhhK ��h��R�(KK��h�C�  s      �           �t�bhhK ��h��R�(KK��h�C	                 �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�CU  �   �        �t�bhhK ��h��R�(KK��h�C #   �   �                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8#   "   '   	     	  	     |         �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C,      {      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�C`     �     �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C,      &   `  a     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C0      �        �   B     �  �         �t�bhhK ��h��R�(KK
��h�C(:   	     �  /   ^     		        �t�bhhK ��h��R�(KK��h�CP   6   x  �   B     �   �  	   v   C  	   D     
	        E        �t�bhhK ��h��R�(KK��h�C,      {      �t�bhhK ��h��R�(KK��h�C<
      "   ,      �     r   {         =   �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CF  G     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C          ,      {         �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CD
      �   5   +      H        M  6      �   �   �         �t�bhhK ��h��R�(KK��h�C4�   4   �   
   .   4      �   
      M        �t�bhhK ��h��R�(KK	��h�C$      �      I             �t�bhhK ��h��R�(KK��h�C             	  2         �t�bhhK ��h��R�(KK��h�C@      -   �  �   	          �   �   &      �        �t�bhhK ��h��R�(KK��h�C#   	     �t�bhhK ��h��R�(KK��h�C�  	     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C	                 �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�CD
      �   5   +      H        M  6      �   �   �         �t�bhhK ��h��R�(KK��h�C         l         �t�bhhK ��h��R�(KK��h�C`     �     �t�bhhK ��h��R�(KK��h�Cl
      u         �  b     `  �      	  �         J  6      �  w   y  �     J   �        �t�bhhK ��h��R�(KK��h�CP
   	  4      	     J  6      =   	     �     �      �  1         �t�bhhK ��h��R�(KK��h�Cc        �t�bhhK ��h��R�(KK��h�C�     �      �  1      �t�bhhK ��h��R�(KK��h�C	  K     �t�bhhK ��h��R�(KK��h�C	  �     �t�bhhK ��h��R�(KK��h�C]      	     �t�bhhK ��h��R�(KK��h�C8
      	     `        >  
   +      	        �t�bhhK ��h��R�(KK��h�CP
      	  �     '   	  	  �         �      I          �        �t�bhhK ��h��R�(KK��h�C          `     �        �t�bhhK ��h��R�(KK��h�C 	     �      �  1         �t�bhhK ��h��R�(KK��h�C,�     �      �  �                 �t�bhhK ��h��R�(KK'��h�C�+            Y      	     	  	                 E      s     �      �      /     v     �     �      �     �     �     L     �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�ChM  ;      �  5  
      "   �      	  �  	         @   !	     N  �  �  U   �          �t�bhhK ��h��R�(KK��h�Ct   3      3        �t�bhhK ��h��R�(KK��h�C#   �     �t�bhhK ��h��R�(KK
��h�C(c     "	  	   ,  #	  	   �   #      �t�bhhK ��h��R�(KK��h�C]      O     �t�bhhK ��h��R�(KK��h�C4   
   P  Q     �   e      �   $	  2         �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�C�   %	        �t�bhhK ��h��R�(KK��h�C�   &	                 �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C4&   �      �   �  �  �  '	     �  �        �t�bhhK ��h��R�(KK��h�C4v      -   �     4      �     �  R        �t�bhhK ��h��R�(KK��h�C,:      �  N        |      �         �t�bhhK ��h��R�(KK
��h�C(            #   �   �  2         �t�bhhK ��h��R�(KK��h�Cd
      �  �  S        g   �     J   �   �   	      T  (	     U     t   3   V        �t�bhhK ��h��R�(KK��h�C0:   �      �   W     �  T   -   )	        �t�bhhK ��h��R�(KK	��h�C$-   *	  +	  T   X     ,	        �t�bhhK ��h��R�(KK��h�C         �        �t�bhhK ��h��R�(KK��h�CU  �   �        �t�bhhK ��h��R�(KK��h�C #   �   �                 �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Ct           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK��h�Ct   ,      m      �   O      +      t   3   Y     -	     #   �   �     t   3   0      K   �  �        �t�bhhK ��h��R�(KK��h�C.	     �t�bhhK ��h��R�(KK��h�C]      /	        �t�bhhK ��h��R�(KK��h�C#   �     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C�     Z     �t�bhhK ��h��R�(KK
��h�C(         ,      m      �         �t�bhhK ��h��R�(KK��h�CP   3   0	        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C<b      [     d  	      e        \  �  ?        �t�bhhK ��h��R�(KK��h�C B   �   
   b      ]        �t�bhhK ��h��R�(KK
��h�C(       f     �     ^  g        �t�bhhK ��h��R�(KK��h�C3   h  #   �     �t�bhhK ��h��R�(KK��h�C c     �  i  	   �   #      �t�bhhK ��h��R�(KK��h�C]      _     �t�bhhK ��h��R�(KK��h�C         b         �t�bhhK ��h��R�(KK��h�CH?     �  p   f      �      V  �  n   G   	   �     �        �t�bhhK ��h��R�(KK��h�C0�  p      
        T   +      �        �t�bhhK ��h��R�(KK��h�C8   ,   d   L      �   x   �  j  0     1	        �t�bhhK ��h��R�(KK	��h�C$         n      _   ,         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C`           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Ca           �t�bhhK ��h��R�(KK��h�CD      w   y  ,      ?     @     2	     �      �        �t�bhhK ��h��R�(KK��h�C4            t   3   0      K   �  2         �t�bhhK ��h��R�(KK	��h�C$�     L   �     =   �         �t�bhhK ��h��R�(KK��h�C4v      B   �  
   ,      @   +      V         �t�bhhK ��h��R�(KK��h�C4            t   3   0      K   �  2         �t�bhhK ��h��R�(KK��h�Cb  w     Z        �t�bhhK ��h��R�(KK	��h�C$         n      _   ,         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C3	           �t�bhhK ��h��R�(KK��h�C�     4	  )            �t�bhhK ��h��R�(KK��h�C,      &   `  a     �t�bhhK ��h��R�(KK��h�CL
      5   +      V      J   `  G         �      {     �         �t�bhhK ��h��R�(KK��h�Cc  |  d        �t�bhhK ��h��R�(KK��h�C,   �  e  c     5	     6	  7	        �t�bhhK ��h��R�(KK��h�C         �   G         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C8	           �t�bhhK ��h��R�(KK ��h�C�
      "   Q  ,         >  
   f   d   t   3   0      K   �  9	     :	     �  	   (   ;	     <	  	   (   f        �t�bhhK ��h��R�(KK��h�C,
      "   ,      �  	   =   =	        �t�bhhK ��h��R�(KK��h�C4      �  ,     a    >	     J   S        �t�bhhK ��h��R�(KK��h�Ct   3      3        �t�bhhK ��h��R�(KK��h�C#   �     �t�bhhK ��h��R�(KK��h�C]      O     �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C?	           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK ��h�C�
      "   ,      @	  	   A	  	   -     B	        @   o      g     C	  	   t   3   0      K   �  D	     �         �t�bhhK ��h��R�(KK��h�Cx      w   y  E	     +  �   �     F	  	         G	  /   ^     H	  	      .  =   �  I	  	   (   J	        �t�bhhK ��h��R�(KK��h�CH   K	     L	  M	     N	  O	  -      P	  	   x  g     �        �t�bhhK ��h��R�(KK��h�C4-   #   �      �   �  Q	  T   X     �         �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CR	  1     �t�bhhK ��h��R�(KK��h�C�  #      �t�bhhK ��h��R�(KK��h�C]      S	     �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�     h           �t�bhhK ��h��R�(KK��h�CU  �      �   i        �t�bhhK ��h��R�(KK��h�C,#   �      �   �  �   �   h           �t�bhhK ��h��R�(KK��h�C,      {      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�C`     �     �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C,      &   `  a     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C0      �        �   B     �  �         �t�bhhK ��h��R�(KK
��h�C(:   	     �  /   ^     		        �t�bhhK ��h��R�(KK��h�CP   6   x  �   B     �   �  	   v   C  	   D     
	        E        �t�bhhK ��h��R�(KK��h�C,      {      �t�bhhK ��h��R�(KK��h�C<
      "   ,      �     r   {         =   �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CF  G     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C          ,      {         �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CD
      �   5   +      H        M  6      �   �   �         �t�bhhK ��h��R�(KK��h�C4�   4   �   
   .   4      �   
      M        �t�bhhK ��h��R�(KK	��h�C$      �      I             �t�bhhK ��h��R�(KK��h�C             	  2         �t�bhhK ��h��R�(KK��h�C@      -   �  �   	          �   �   &      �        �t�bhhK ��h��R�(KK��h�C#   	     �t�bhhK ��h��R�(KK��h�C�  	     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C	                 �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�CD
      �   5   +      H        M  6      �   �   �         �t�bhhK ��h��R�(KK��h�C         l         �t�bhhK ��h��R�(KK��h�C`     �     �t�bhhK ��h��R�(KK��h�Cl
      u         �  b     `  �      	  �         J  6      �  w   y  �     J   �        �t�bhhK ��h��R�(KK��h�CP
   	  4      	     J  6      =   	     �     �      �  1         �t�bhhK ��h��R�(KK��h�Cc        �t�bhhK ��h��R�(KK��h�C�     �      �  1      �t�bhhK ��h��R�(KK��h�C	  K     �t�bhhK ��h��R�(KK��h�C	  �     �t�bhhK ��h��R�(KK��h�C]      	     �t�bhhK ��h��R�(KK��h�C8
      	     `        >  
   +      	        �t�bhhK ��h��R�(KK��h�CP
      	  �     '   	  	  �         �      I          �        �t�bhhK ��h��R�(KK��h�C          `     �        �t�bhhK ��h��R�(KK��h�C 	     �      �  1         �t�bhhK ��h��R�(KK��h�C,�     �      �  �                 �t�bhhK ��h��R�(KK'��h�C�+            Y      	     	  	                 E      s     �      �      /     v     �     �      �     �     �     L     �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�ChM  ;      �  5  
      "   �      	  �  	         @   !	     N  �  �  U   �          �t�bhhK ��h��R�(KK��h�Ct   3      3        �t�bhhK ��h��R�(KK��h�C#   �     �t�bhhK ��h��R�(KK
��h�C(c     "	  	   ,  #	  	   �   #      �t�bhhK ��h��R�(KK��h�C]      O     �t�bhhK ��h��R�(KK��h�C4   
   P  Q     �   e      �   $	  2         �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�C�   %	        �t�bhhK ��h��R�(KK��h�C�   &	                 �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C4&   �      �   �  �  �  '	     �  �        �t�bhhK ��h��R�(KK��h�C4v      -   �     4      �     �  R        �t�bhhK ��h��R�(KK��h�C,:      �  N        |      �         �t�bhhK ��h��R�(KK
��h�C(            #   �   �  2         �t�bhhK ��h��R�(KK��h�Cd
      �  �  S        g   �     J   �   �   	      T  (	     U     t   3   V        �t�bhhK ��h��R�(KK��h�C0:   �      �   W     �  T   -   )	        �t�bhhK ��h��R�(KK	��h�C$-   *	  +	  T   X     ,	        �t�bhhK ��h��R�(KK��h�C         �        �t�bhhK ��h��R�(KK��h�CU  �   �        �t�bhhK ��h��R�(KK��h�C #   �   �                 �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Ct           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK��h�Ct   ,      m      �   O      +      t   3   Y     -	     #   �   �     t   3   0      K   �  �        �t�bhhK ��h��R�(KK��h�C.	     �t�bhhK ��h��R�(KK��h�C]      /	        �t�bhhK ��h��R�(KK��h�C#   �     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C�     Z     �t�bhhK ��h��R�(KK
��h�C(         ,      m      �         �t�bhhK ��h��R�(KK��h�CP   3   0	        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C<b      [     d  	      e        \  �  ?        �t�bhhK ��h��R�(KK��h�C B   �   
   b      ]        �t�bhhK ��h��R�(KK
��h�C(       f     �     ^  g        �t�bhhK ��h��R�(KK��h�C3   h  #   �     �t�bhhK ��h��R�(KK��h�C c     �  i  	   �   #      �t�bhhK ��h��R�(KK��h�C]      _     �t�bhhK ��h��R�(KK��h�C         b         �t�bhhK ��h��R�(KK��h�CH?     �  p   f      �      V  �  n   G   	   �     �        �t�bhhK ��h��R�(KK��h�C0�  p      
        T   +      �        �t�bhhK ��h��R�(KK��h�C8   ,   d   L      �   x   �  j  0     1	        �t�bhhK ��h��R�(KK	��h�C$         n      _   ,         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C`           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Ca           �t�bhhK ��h��R�(KK��h�CD      w   y  ,      ?     @     2	     �      �        �t�bhhK ��h��R�(KK��h�C4            t   3   0      K   �  2         �t�bhhK ��h��R�(KK	��h�C$�     L   �     =   �         �t�bhhK ��h��R�(KK��h�C4v      B   �  
   ,      @   +      V         �t�bhhK ��h��R�(KK��h�C4            t   3   0      K   �  2         �t�bhhK ��h��R�(KK��h�Cb  w     Z        �t�bhhK ��h��R�(KK	��h�C$         n      _   ,         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C3	           �t�bhhK ��h��R�(KK��h�C�     4	  )            �t�bhhK ��h��R�(KK��h�C,      &   `  a     �t�bhhK ��h��R�(KK��h�CL
      5   +      V      J   `  G         �      {     �         �t�bhhK ��h��R�(KK��h�Cc  |  d        �t�bhhK ��h��R�(KK��h�C,   �  e  c     5	     6	  7	        �t�bhhK ��h��R�(KK��h�C         �   G         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C8	           �t�bhhK ��h��R�(KK ��h�C�
      "   Q  ,         >  
   f   d   t   3   0      K   �  9	     :	     �  	   (   ;	     <	  	   (   f        �t�bhhK ��h��R�(KK��h�C,
      "   ,      �  	   =   =	        �t�bhhK ��h��R�(KK��h�C4      �  ,     a    >	     J   S        �t�bhhK ��h��R�(KK��h�Ct   3      3        �t�bhhK ��h��R�(KK��h�C#   �     �t�bhhK ��h��R�(KK��h�C]      O     �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C?	           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK ��h�C�
      "   ,      @	  	   A	  	   -     B	        @   o      g     C	  	   t   3   0      K   �  D	     �         �t�bhhK ��h��R�(KK��h�Cx      w   y  E	     +  �   �     F	  	         G	  /   ^     H	  	      .  =   �  I	  	   (   J	        �t�bhhK ��h��R�(KK��h�CH   K	     L	  M	     N	  O	  -      P	  	   x  g     �        �t�bhhK ��h��R�(KK��h�C4-   #   �      �   �  Q	  T   X     �         �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CR	  1     �t�bhhK ��h��R�(KK��h�C�  #      �t�bhhK ��h��R�(KK��h�C]      S	     �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�     h           �t�bhhK ��h��R�(KK��h�CU  �      �   i        �t�bhhK ��h��R�(KK��h�C,#   �      �   �  �   �   h           �t�bhhK ��h��R�(KK��h�C,      {      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�C`     �     �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C,      &   `  a     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C0      �        �   B     �  �         �t�bhhK ��h��R�(KK
��h�C(:   	     �  /   ^     		        �t�bhhK ��h��R�(KK��h�CP   6   x  �   B     �   �  	   v   C  	   D     
	        E        �t�bhhK ��h��R�(KK��h�C,      {      �t�bhhK ��h��R�(KK��h�C<
      "   ,      �     r   {         =   �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CF  G     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C          ,      {         �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CD
      �   5   +      H        M  6      �   �   �         �t�bhhK ��h��R�(KK��h�C4�   4   �   
   .   4      �   
      M        �t�bhhK ��h��R�(KK	��h�C$      �      I             �t�bhhK ��h��R�(KK��h�C             	  2         �t�bhhK ��h��R�(KK��h�C@      -   �  �   	          �   �   &      �        �t�bhhK ��h��R�(KK��h�C#   	     �t�bhhK ��h��R�(KK��h�C�  	     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C	                 �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�CD
      �   5   +      H        M  6      �   �   �         �t�bhhK ��h��R�(KK��h�C         l         �t�bhhK ��h��R�(KK��h�C`     �     �t�bhhK ��h��R�(KK��h�Cl
      u         �  b     `  �      	  �         J  6      �  w   y  �     J   �        �t�bhhK ��h��R�(KK��h�CP
   	  4      	     J  6      =   	     �     �      �  1         �t�bhhK ��h��R�(KK��h�Cc        �t�bhhK ��h��R�(KK��h�C�     �      �  1      �t�bhhK ��h��R�(KK��h�C	  K     �t�bhhK ��h��R�(KK��h�C	  �     �t�bhhK ��h��R�(KK��h�C]      	     �t�bhhK ��h��R�(KK��h�C8
      	     `        >  
   +      	        �t�bhhK ��h��R�(KK��h�CP
      	  �     '   	  	  �         �      I          �        �t�bhhK ��h��R�(KK��h�C          `     �        �t�bhhK ��h��R�(KK��h�C 	     �      �  1         �t�bhhK ��h��R�(KK��h�C,�     �      �  �                 �t�bhhK ��h��R�(KK'��h�C�+            Y      	     	  	                 E      s     �      �      /     v     �     �      �     �     �     L     �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�ChM  ;      �  5  
      "   �      	  �  	         @   !	     N  �  �  U   �          �t�bhhK ��h��R�(KK��h�Ct   3      3        �t�bhhK ��h��R�(KK��h�C#   �     �t�bhhK ��h��R�(KK
��h�C(c     "	  	   ,  #	  	   �   #      �t�bhhK ��h��R�(KK��h�C]      O     �t�bhhK ��h��R�(KK��h�C4   
   P  Q     �   e      �   $	  2         �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�C�   %	        �t�bhhK ��h��R�(KK��h�C�   &	                 �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C4&   �      �   �  �  �  '	     �  �        �t�bhhK ��h��R�(KK��h�C4v      -   �     4      �     �  R        �t�bhhK ��h��R�(KK��h�C,:      �  N        |      �         �t�bhhK ��h��R�(KK
���7      h�C(            #   �   �  2         �t�bhhK ��h��R�(KK��h�Cd
      �  �  S        g   �     J   �   �   	      T  (	     U     t   3   V        �t�bhhK ��h��R�(KK��h�C0:   �      �   W     �  T   -   )	        �t�bhhK ��h��R�(KK	��h�C$-   *	  +	  T   X     ,	        �t�bhhK ��h��R�(KK��h�C         �        �t�bhhK ��h��R�(KK��h�CU  �   �        �t�bhhK ��h��R�(KK��h�C #   �   �                 �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Ct           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK��h�Ct   ,      m      �   O      +      t   3   Y     -	     #   �   �     t   3   0      K   �  �        �t�bhhK ��h��R�(KK��h�C.	     �t�bhhK ��h��R�(KK��h�C]      /	        �t�bhhK ��h��R�(KK��h�C#   �     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C�     Z     �t�bhhK ��h��R�(KK
��h�C(         ,      m      �         �t�bhhK ��h��R�(KK��h�CP   3   0	        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C<b      [     d  	      e        \  �  ?        �t�bhhK ��h��R�(KK��h�C B   �   
   b      ]        �t�bhhK ��h��R�(KK
��h�C(       f     �     ^  g        �t�bhhK ��h��R�(KK��h�C3   h  #   �     �t�bhhK ��h��R�(KK��h�C c     �  i  	   �   #      �t�bhhK ��h��R�(KK��h�C]      _     �t�bhhK ��h��R�(KK��h�C         b         �t�bhhK ��h��R�(KK��h�CH?     �  p   f      �      V  �  n   G   	   �     �        �t�bhhK ��h��R�(KK��h�C0�  p      
        T   +      �        �t�bhhK ��h��R�(KK��h�C8   ,   d   L      �   x   �  j  0     1	        �t�bhhK ��h��R�(KK	��h�C$         n      _   ,         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C`           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Ca           �t�bhhK ��h��R�(KK��h�CD      w   y  ,      ?     @     2	     �      �        �t�bhhK ��h��R�(KK��h�C4            t   3   0      K   �  2         �t�bhhK ��h��R�(KK	��h�C$�     L   �     =   �         �t�bhhK ��h��R�(KK��h�C4v      B   �  
   ,      @   +      V         �t�bhhK ��h��R�(KK��h�C4            t   3   0      K   �  2         �t�bhhK ��h��R�(KK��h�Cb  w     Z        �t�bhhK ��h��R�(KK	��h�C$         n      _   ,         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C3	           �t�bhhK ��h��R�(KK��h�C�     4	  )            �t�bhhK ��h��R�(KK��h�C,      &   `  a     �t�bhhK ��h��R�(KK��h�CL
      5   +      V      J   `  G         �      {     �         �t�bhhK ��h��R�(KK��h�Cc  |  d        �t�bhhK ��h��R�(KK��h�C,   �  e  c     5	     6	  7	        �t�bhhK ��h��R�(KK��h�C         �   G         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C8	           �t�bhhK ��h��R�(KK ��h�C�
      "   Q  ,         >  
   f   d   t   3   0      K   �  9	     :	     �  	   (   ;	     <	  	   (   f        �t�bhhK ��h��R�(KK��h�C,
      "   ,      �  	   =   =	        �t�bhhK ��h��R�(KK��h�C4      �  ,     a    >	     J   S        �t�bhhK ��h��R�(KK��h�Ct   3      3        �t�bhhK ��h��R�(KK��h�C#   �     �t�bhhK ��h��R�(KK��h�C]      O     �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C?	           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK ��h�C�
      "   ,      @	  	   A	  	   -     B	        @   o      g     C	  	   t   3   0      K   �  D	     �         �t�bhhK ��h��R�(KK��h�Cx      w   y  E	     +  �   �     F	  	         G	  /   ^     H	  	      .  =   �  I	  	   (   J	        �t�bhhK ��h��R�(KK��h�CH   K	     L	  M	     N	  O	  -      P	  	   x  g     �        �t�bhhK ��h��R�(KK��h�C4-   #   �      �   �  Q	  T   X     �         �t�bhhK ��h��R�(KK��h�C�      �t�be(hhK ��h��R�(KK��h�CR	  1     �t�bhhK ��h��R�(KK��h�C�  #      �t�bhhK ��h��R�(KK��h�C]      S	     �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�     h           �t�bhhK ��h��R�(KK��h�CU  �      �   i        �t�bhhK ��h��R�(KK��h�C,#   �      �   �  �   �   h           �t�bhhK ��h��R�(KK��h�Cm      �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C$      b      �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�Co      z      �t�bhhK ��h��R�(KK��h�Co      z      �      �t�bhhK ��h��R�(KK��h�Cm      �t�bhhK ��h��R�(KK��h�C4  �  T	  6      U	  >  
   �     V	        �t�bhhK ��h��R�(KK��h�CLW	  �     �            �   �   `   
   �     ,  �     a        �t�bhhK ��h��R�(KK��h�CX	  j  Y	     �         �t�bhhK ��h��R�(KK��h�C�      �   1      �t�bhhK ��h��R�(KK��h�C#   �     �t�bhhK ��h��R�(KK��h�C�  i  	   �  Z	     �t�bhhK ��h��R�(KK��h�Ck  #      �t�bhhK ��h��R�(KK��h�C]      l     �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�Cm         �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C<b      [     d  	      e        \  �  ?        �t�bhhK ��h��R�(KK��h�C B   �   
   b      ]        �t�bhhK ��h��R�(KK
��h�C(       f     �     ^  g        �t�bhhK ��h��R�(KK��h�C3   h  #   �     �t�bhhK ��h��R�(KK��h�C c     �  i  	   �   #      �t�bhhK ��h��R�(KK��h�C]      _     �t�bhhK ��h��R�(KK��h�C         b         �t�bhhK ��h��R�(KK��h�C$      b      �t�bhhK ��h��R�(KK��h�CD
      "   $      �  [	     b   6      w   �      �        �t�bhhK ��h��R�(KK��h�CH�  �  \	  
   u   k  6   �  	   �     k  	   �     �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C]	     b     �t�bhhK ��h��R�(KK��h�C�     ^	     �t�bhhK ��h��R�(KK��h�C          $      b         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C_	           �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�C4w   �      L  �      m            �        �t�bhhK ��h��R�(KK��h�C@   L  n  B      �  	   �      �  A  �  ?   �        �t�bhhK ��h��R�(KK��h�C4      >  
   f   �   ]      �      �        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�CN      u  $         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Co           �t�bhhK ��h��R�(KK��h�Co      z      �t�bhhK ��h��R�(KK��h�C4   #      H   �   	   �  	   l  \   �        �t�bhhK ��h��R�(KK��h�CP�      .   �      p     �     	   '   �   �      �   l     #         �t�bhhK ��h��R�(KK��h�Cp      i   
      �   �     r   $   m  M   q   `	           �     H   2      `   
   1           �t�bhhK ��h��R�(KK��h�C8`   6   �  �   �   n       5      �   �        �t�bhhK ��h��R�(KK��h�CT.      c      @         q  
   &   r            �  s  �      �         �t�bhhK ��h��R�(KK��h�C\`      �     t     1  	   �     1     �     u     &   v  w     �        �t�bhhK ��h��R�(KK��h�CH      i   
            H   �     �           H   2         �t�bhhK ��h��R�(KK��h�C,`      -   �  �        y  �         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C;      1     �t�bhhK ��h��R�(KK��h�Cx     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C�      W   y           �t�bhhK ��h��R�(KK��h�Cz           �t�bhhK ��h��R�(KK��h�C{           �t�bhhK ��h��R�(KK��h�C     i   
   |  �           �t�bhhK ��h��R�(KK��h�Co      z      �      �t�bhhK ��h��R�(KK��h�CT
   A  }  $      ~  B     I      a	  @   o     o      z      �         �t�bhhK ��h��R�(KK��h�C<
      "   �      �        i   
   �  d           �t�bhhK ��h��R�(KK��h�C@           `             &   �                �t�bhhK ��h��R�(KK��h�C       -   �   2          �t�bhhK ��h��R�(KK��h�CP#      �  �  b	     :        �   �   
   $   ?      I      �         �t�bhhK ��h��R�(KK��h�CT      i   
   �  
   &   �        �  3     A  $   ?   �      �         �t�bhhK ��h��R�(KK��h�C@
   J   �  �  c	  	   d	  �          e	     f	        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK	��h�C$V      o      $      �         �t�bhhK ��h��R�(KK��h�Cg	           �t�bhhK ��h��R�(KK	��h�C$   
   2  �                 �t�bhhK ��h��R�(KK��h�C  �                  �t�bhhK ��h��R�(KK��h�Cm      �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C$      b      �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�Co      z      �t�bhhK ��h��R�(KK��h�Co      z      �      �t�bhhK ��h��R�(KK��h�Cm      �t�bhhK ��h��R�(KK��h�C4  �  T	  6      U	  >  
   �     V	        �t�bhhK ��h��R�(KK��h�CLW	  �     �            �   �   `   
   �     ,  �     a        �t�bhhK ��h��R�(KK��h�CX	  j  Y	     �         �t�bhhK ��h��R�(KK��h�C�      �   1      �t�bhhK ��h��R�(KK��h�C#   �     �t�bhhK ��h��R�(KK��h�C�  i  	   �  Z	     �t�bhhK ��h��R�(KK��h�Ck  #      �t�bhhK ��h��R�(KK��h�C]      l     �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�Cm         �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C<b      [     d  	      e        \  �  ?        �t�bhhK ��h��R�(KK��h�C B   �   
   b      ]        �t�bhhK ��h��R�(KK
��h�C(       f     �     ^  g        �t�bhhK ��h��R�(KK��h�C3   h  #   �     �t�bhhK ��h��R�(KK��h�C c     �  i  	   �   #      �t�bhhK ��h��R�(KK��h�C]      _     �t�bhhK ��h��R�(KK��h�C         b         �t�bhhK ��h��R�(KK��h�C$      b      �t�bhhK ��h��R�(KK��h�CD
      "   $      �  [	     b   6      w   �      �        �t�bhhK ��h��R�(KK��h�CH�  �  \	  
   u   k  6   �  	   �     k  	   �     �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C]	     b     �t�bhhK ��h��R�(KK��h�C�     ^	     �t�bhhK ��h��R�(KK��h�C          $      b         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C_	           �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�C4w   �      L  �      m            �        �t�bhhK ��h��R�(KK��h�C@   L  n  B      �  	   �      �  A  �  ?   �        �t�bhhK ��h��R�(KK��h�C4      >  
   f   �   ]      �      �        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�CN      u  $         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Co           �t�bhhK ��h��R�(KK��h�Co      z      �t�bhhK ��h��R�(KK��h�C4   #      H   �   	   �  	   l  \   �        �t�bhhK ��h��R�(KK��h�CP�      .   �      p     �     	   '   �   �      �   l     #         �t�bhhK ��h��R�(KK��h�Cp      i   
      �   �     r   $   m  M   q   `	           �     H   2      `   
   1           �t�bhhK ��h��R�(KK��h�C8`   6   �  �   �   n       5      �   �        �t�bhhK ��h��R�(KK��h�CT.      c      @         q  
   &   r            �  s  �      �         �t�bhhK ��h��R�(KK��h�C\`      �     t     1  	   �     1     �     u     &   v  w     �        �t�bhhK ��h��R�(KK��h�CH      i   
            H   �     �           H   2         �t�bhhK ��h��R�(KK��h�C,`      -   �  �        y  �         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C;      1     �t�bhhK ��h��R�(KK��h�Cx     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C�      W   y           �t�bhhK ��h��R�(KK��h�Cz           �t�bhhK ��h��R�(KK��h�C{           �t�bhhK ��h��R�(KK��h�C     i   
   |  �           �t�bhhK ��h��R�(KK��h�Co      z      �      �t�bhhK ��h��R�(KK��h�CT
   A  }  $      ~  B     I      a	  @   o     o      z      �         �t�bhhK ��h��R�(KK��h�C<
      "   �      �        i   
   �  d           �t�bhhK ��h��R�(KK��h�C@           `             &   �                �t�bhhK ��h��R�(KK��h�C       -   �   2          �t�bhhK ��h��R�(KK��h�CP#      �  �  b	     :        �   �   
   $   ?      I      �         �t�bhhK ��h��R�(KK��h�CT      i   
   �  
   &   �        �  3     A  $   ?   �      �         �t�bhhK ��h��R�(KK��h�C@
   J   �  �  c	  	   d	  �          e	     f	        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK	��h�C$V      o      $      �         �t�bhhK ��h��R�(KK��h�Cg	           �t�bhhK ��h��R�(KK	��h�C$   
   2  �                 �t�bhhK ��h��R�(KK��h�C  �                  �t�bhhK ��h��R�(KK��h�Cm      �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C$      b      �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�Co      z      �t�bhhK ��h��R�(KK��h�Co      z      �      �t�bhhK ��h��R�(KK��h�Cm      �t�bhhK ��h��R�(KK��h�C4  �  T	  6      U	  >  
   �     V	        �t�bhhK ��h��R�(KK��h�CLW	  �     �            �   �   `   
   �     ,  �     a        �t�bhhK ��h��R�(KK��h�CX	  j  Y	     �         �t�bhhK ��h��R�(KK��h�C�      �   1      �t�bhhK ��h��R�(KK��h�C#   �     �t�bhhK ��h��R�(KK��h�C�  i  	   �  Z	     �t�bhhK ��h��R�(KK��h�Ck  #      �t�bhhK ��h��R�(KK��h�C]      l     �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�Cm         �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C<b      [     d  	      e        \  �  ?        �t�bhhK ��h��R�(KK��h�C B   �   
   b      ]        �t�bhhK ��h��R�(KK
��h�C(       f     �     ^  g        �t�bhhK ��h��R�(KK��h�C3   h  #   �     �t�bhhK ��h��R�(KK��h�C c     �  i  	   �   #      �t�bhhK ��h��R�(KK��h�C]      _     �t�bhhK ��h��R�(KK��h�C         b         �t�bhhK ��h��R�(KK��h�C$      b      �t�bhhK ��h��R�(KK��h�CD
      "   $      �  [	     b   6      w   �      �        �t�bhhK ��h��R�(KK��h�CH�  �  \	  
   u   k  6   �  	   �     k  	   �     �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C]	     b     �t�bhhK ��h��R�(KK��h�C�     ^	     �t�bhhK ��h��R�(KK��h�C          $      b         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C_	           �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�C4w   �      L  �      m            �        �t�bhhK ��h��R�(KK��h�C@   L  n  B      �  	   �      �  A  �  ?   �        �t�bhhK ��h��R�(KK��h�C4      >  
   f   �   ]      �      �        �t�bhhK ��h��R�(KK��h�C          �     T        �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Co           �t�bhhK ��h��R�(KK��h�Co      z      �t�bhhK ��h��R�(KK��h�C4   #      H   �   	   �  	   l  \   �        �t�bhhK ��h��R�(KK��h�CP�      .   �      p     �     	   '   �   �      �   l     #         �t�bhhK ��h��R�(KK��h�Cp      i   
      �   �     r   $   m  M   q   `	           �     H   2      `   
   1           �t�bhhK ��h��R�(KK��h�C8`   6   �  �   �   n       5      �   �        �t�bhhK ��h��R�(KK��h�CT.      c      @         q  
   &   r            �  s  �      �         �t�bhhK ��h��R�(KK��h�C\`      �     t     1  	   �     1     �     u     &   v  w     �        �t�bhhK ��h��R�(KK��h�CH      i   
            H   �     �           H   2         �t�bhhK ��h��R�(KK��h�C,`      -   �  �        y  �         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C;      1     �t�bhhK ��h��R�(KK��h�Cx     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�Co      z         �t�bhhK ��h��R�(KK��h�C�      W   y           �t�bhhK ��h��R�(KK��h�Cz           �t�bhhK ��h��R�(KK��h�C{           �t�bhhK ��h��R�(KK��h�C     i   
   |  �           �t�bhhK ��h��R�(KK��h�Co      z      �      �t�bhhK ��h��R�(KK��h�CT
   A  }  $      ~  B     I      a	  @   o     o      z      �         �t�bhhK ��h��R�(KK��h�C<
      "   �      �        i   
   �  d           �t�bhhK ��h��R�(KK��h�C@           `             &   �                �t�bhhK ��h��R�(KK��h�C       -   �   2          �t�bhhK ��h��R�(KK��h�CP#      �  �  b	     :        �   �   
   $   ?      I      �         �t�bhhK ��h��R�(KK��h�CT      i   
   �  
   &   �        �  3     A  $   ?   �      �         �t�bhhK ��h��R�(KK��h�C@
   J   �  �  c	  	   d	  �          e	     f	        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK	��h�C$V      o      $      �         �t�bhhK ��h��R�(KK��h�Cg	           �t�bhhK ��h��R�(KK	��h�C$   
   2  �                 �t�bhhK ��h��R�(KK��h�C  �                  �t�bhhK ��h��R�(KK��h�C�      #      �t�bhhK ��h��R�(KK��h�C�   �  G      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�   G      �t�bhhK ��h��R�(KK��h�C4  G      �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�CT     �t�bhhK ��h��R�(KK��h�C-     �t�bhhK ��h��R�(KK��h�C�   Y      �t�bhhK ��h��R�(KK��h�C'   �  $      �t�bhhK ��h��R�(KK��h�C�      #      �t�bhhK ��h��R�(KK��h�C,   #      5     >   ?     �         �t�bhhK ��h��R�(KK��h�C\d  �   "   '   �   w     b  	      B      �          �   }      �     @        �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C#   h	     �t�bhhK ��h��R�(KK��h�Cp  �     �t�bhhK ��h��R�(KK��h�C�  #      �t�bhhK ��h��R�(KK��h�C]         �      �     �t�bhhK ��h��R�(KK��h�CD   #   �  �  i	     �     j	     �  z  �  k	           �t�bhhK ��h��R�(KK��h�C<l	  O      }      m	  	   �     n	  R      �        �t�bhhK ��h��R�(KK��h�C@�     �  �     '        w  	      �      o	        �t�bhhK ��h��R�(KK��h�C�  #      �t�bhhK ��h��R�(KK��h�C]         �      �     �t�bhhK ��h��R�(KK��h�C  �  8     �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C�  8     �t�bhhK ��h��R�(KK��h�C]         �      p	     �t�bhhK ��h��R�(KK��h�C  �  �     �t�bhhK ��h��R�(KK��h�C]         �      q	     �t�bhhK ��h��R�(KK��h�C  �  Y     �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C�  Y     �t�bhhK ��h��R�(KK��h�C]         �      r	     �t�bhhK ��h��R�(KK��h�CH
      U          1   6      �  s	  
      t	     u	        �t�bhhK ��h��R�(KK��h�C         G         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Ct           �t�bhhK ��h��R�(KK	��h�C$?   �          �  �        �t�bhhK ��h��R�(KK
��h�C(�   �  v	  �     w	     e        �t�bhhK ��h��R�(KK��h�C8e     �     x	  �  {  y	  �   z	     o         �t�bhhK ��h��R�(KK
��h�C(   {	    6      �   �   �         �t�bhhK ��h��R�(KK��h�CP
      �  e  �     ?     6      �  �   �  |	     �      }	        �t�bhhK ��h��R�(KK��h�C~	  �         �t�bhhK ��h��R�(KK��h�Ct   3   V     �t�bhhK ��h��R�(KK��h�C4p  /     O     �     	  	   �	  �	        �t�bhhK ��h��R�(KK��h�C�  #      �t�bhhK ��h��R�(KK��h�C         �      1      �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Cn   G      �t�bhhK ��h��R�(KK��h�C0
   r   $   q  6      =   �      �        �t�bhhK ��h��R�(KK��h�C,�	  T   ;      �	     $   ?   �         �t�bhhK ��h��R�(KK
��h�C(   �  �  �	     $      �         �t�bhhK ��h��R�(KK��h�C8      =   L  M   &   r  s     �      �        �t�bhhK ��h��R�(KK��h�C<2  �	       �  6  �   G   	   �     �  y        �t�bhhK ��h��R�(KK��h�Cd   L    4   $      q  �  	   5        >  
   f   M   &   r  s     �      �        �t�bhhK ��h��R�(KK��h�C �  "   �   
   �	  G         �t�bhhK ��h��R�(KK��h�C4            t   3   0      K   �  2         �t�bhhK ��h��R�(KK��h�C         n   G         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Ca           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�	           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C`           �t�bhhK ��h��R�(KK��h�C�   �  G      �t�bhhK ��h��R�(KK��h�CP   �	  �	  V       c      Y   ;  A  I   
   �	  	   �      �	        �t�bhhK ��h��R�(KK��h�C,�	     Y   ;  A  I   �     �	        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C�   �  G         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�  �	           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C<
      5   �	     �   �   6      �   �	  r          �t�bhhK ��h��R�(KK
��h�C(�	  b  �   ]         �      �	     �t�bhhK ��h��R�(KK��h�C�	       �t�bhhK ��h��R�(KK��h�Cp  �  	   �  #      �t�bhhK ��h��R�(KK��h�C�	       �t�bhhK ��h��R�(KK��h�C�	       �t�bhhK ��h��R�(KK��h�C�	  �  	   �   #      �t�bhhK ��h��R�(KK��h�C8       �t�bhhK ��h��R�(KK��h�C�  �  	   �  	   8     �t�bhhK ��h��R�(KK��h�C�       �t�bhhK ��h��R�(KK��h�CY       �t�bhhK ��h��R�(KK��h�C�  �  	   �  Y     �t�bhhK ��h��R�(KK��h�C4\     \     �  �	  6  �	     3  �        �t�bhhK ��h��R�(KK��h�C@�   �   �  �  �     �  	   �  	   �	     �           �t�bhhK ��h��R�(KK��h�C4   �  O      �  �     �	  �	     �	        �t�bhhK ��h��R�(KK7��h�Cܝ	     �  	   �     �	     �      t     �	     �	     t   3   0      K   R   	   p  /     O  	   �  #      �  C  	     �	     	   �	  y      	     �  \   B     �  y      u     �        �t�bhhK ��h��R�(KK��h�C@         �	  �     �   2      �  =   e  M   ]         �t�bhhK ��h��R�(KK��h�C4   �   �  e  �   �        �      �	        �t�bhhK ��h��R�(KK��h�CPN      U     �   6      w      �	  	   �	     4   "      �	  }         �t�bhhK ��h��R�(KK
��h�C(�   �   �  �  �     �           �t�bhhK ��h��R�(KK��h�Cd�	  �     �	  �	  �	     �	  �	  �  �	     y      �  �	  u  	   �        �     �	     �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�	           �t�bhhK ��h��R�(KK��h�C�   G      �t�bhhK ��h��R�(KK��h�CP   ,      J   `  G   6         �  �   =   J   �   �      �	          �t�bhhK ��h��R�(KK	��h�C$   �   ,   	   =   �	  �	        �t�bhhK ��h��R�(KK��h�C         �   G         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Ct           �t�bhhK ��h��R�(KK��h�C4  G      �t�bhhK ��h��R�(KK��h�CL
      �	         5      
   �     �        =   J   �   �         �t�bhhK ��h��R�(KK��h�C`�   }      �   
      5   
  	   �      �      �     u         �	        �        �t�bhhK ��h��R�(KK��h�CD      -   �      }   d      �        �	     �	  �        �t�bhhK ��h��R�(KK��h�C8   �	        =   &   r  s     �      �        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Ct           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�	           �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�C4w   �      L  �      m            �        �t�bhhK ��h��R�(KK��h�C@   L  n  B      �  	   �      �  A  �  ?   �        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�CN      u  $         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Co           �t�bhhK ��h��R�(KK��h�CT     �t�bhhK ��h��R�(KK��h�C�     x  �   �         �t�bhhK ��h��R�(KK��h�CT
      �        �   �	  �   J   T  �	  �     
      �   �   
   f         �t�bhhK ��h��R�(KK��h�Ct�      U       6      �   �	  �	  y      �     O       \  �     �   &   �  �  �  �	  �	        �t�bhhK ��h��R�(KK��h�C�      �        �t�bhhK ��h��R�(KK��h�Cp  /     O  	      �t�bhhK ��h��R�(KK��h�C�  #      �t�bhhK ��h��R�(KK��h�C ]         �      �	        �t�bhhK ��h��R�(KK��h�C         T        �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�	           �t�bhhK ��h��R�(KK��h�C-     �t�bhhK ��h��R�(KK��h�C       �   -     �        �t�bhhK ��h��R�(KK	��h�C$      �     �     a        �t�bhhK ��h��R�(KK��h�C8      -   �   �     4         J   �   �        �t�bhhK ��h��R�(KK��h�C         -        �t�bhhK ��h��R�(KK��h�C�   Y      �t�bhhK ��h��R�(KK��h�Cl   �  �  �	     #   "   �       �	  :   ;          5        �	     :          ]        �t�bhhK ��h��R�(KK��h�C\�	     �     �     v  �     �  {  -   �	  �  ;      �          D  �        �t�bhhK ��h��R�(KK��h�C`   �      �      #     t   3   0      K   R   	   v   B      i   
   ;      �	        �t�bhhK ��h��R�(KK��h�C8;      ^   >   �    -      Y      �	  �        �t�bhhK ��h��R�(KK��h�C�  ;   �	  �   e         �t�bhhK ��h��R�(KK��h�C�	     �t�bhhK ��h��R�(KK��h�C�	     �	  �     �      �t�bhhK ��h��R�(KK��h�C�	     �     �t�bhhK ��h��R�(KK��h�C  +      �     �t�bhhK ��h��R�(KK��h�C�	     �t�bhhK ��h��R�(KK��h�C,V      |     Y   ?   A     �	        �t�bhhK ��h��R�(KK��h�CT�      .   c      i   
   �	  	   �	       o   \     d   &   �   �        �t�bhhK ��h��R�(KK��h�CX      
   ;      �   O      U   t   3   0      K   �  �	  �   ]      �	        �t�bhhK ��h��R�(KK��h�C         �   Y         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C;      �           �t�bhhK ��h��R�(KK��h�C�     �           �t�bhhK ��h��R�(KK��h�C�      &   [   �     �t�bhhK ��h��R�(KK��h�C'   �  $      �t�bhhK ��h��R�(KK��h�C0.  V     $      �  �   �     @        �t�bhhK ��h��R�(KK
��h�C(=   #   Q   �         
   �	        �t�bhhK ��h��R�(KK��h�C8      >  �	  
         
   ;      @  T         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK	��h�C$�  /     �  �     �        �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C]      �	     �t�bhhK ��h��R�(KK��h�C          '   �  $         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C;      �           �t�bhhK ��h��R�(KK��h�C�     �           �t�bhhK ��h��R�(KK��h�C�      &   [   �     �t�bhhK ��h��R�(KK��h�C�      #      �t�bhhK ��h��R�(KK��h�C�   �  G      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�   G      �t�bhhK ��h��R�(KK��h�C4  G      �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�CT     �t�bhhK ��h��R�(KK��h�C-     �t�bhhK ��h��R�(KK��h�C�   Y      �t�bhhK ��h��R�(KK��h�C'   �  $      �t�bhhK ��h��R�(KK��h�C�      #      �t�bhhK ��h��R�(KK��h�C,   #      5     >   ?     �         �t�bhhK ��h��R�(KK��h�C\d  �   "   '   �   w     b  	      B      �          �   }      �     @        �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C#   h	     �t�bhhK ��h��R�(KK��h�Cp  �     �t�bhhK ��h��R�(KK��h�C�  #      �t�bhhK ��h��R�(KK��h�C]         �      �     �t�bhhK ��h��R�(KK��h�CD   #   �  �  i	     �     j	     �  z  �  k	           �t�bhhK ��h��R�(KK��h�C<l	  O      }      m	  	   �     n	  R      �        �t�bhhK ��h��R�(KK��h�C@�     �  �     '        w  	      �      o	        �t�bhhK ��h��R�(KK��h�C�  #      �t�bhhK ��h��R�(KK��h�C]         �      �     �t�bhhK ��h��R�(KK��h�C  �  8     �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C�  8     �t�bhhK ��h��R�(KK��h�C]         �      p	     �t�bhhK ��h��R�(KK��h�C  �  �     �t�bhhK ��h��R�(KK��h�C]         �      q	     �t�bhhK ��h��R�(KK��h�C  �  Y     �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C�  Y     �t�bhhK ��h��R�(KK��h�C]         �      r	     �t�bhhK ��h��R�(KK��h�CH
      U          1   6      �  s	  
      t	     u	        �t�bhhK ��h��R�(KK��h�C         G         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Ct           �t�bhhK ��h��R�(KK	��h�C$?   �          �  �        �t�bhhK ��h��R�(KK
��h�C(�   �  v	  �     w	     e        �t�bhhK ��h��R�(KK��h�C8e     �     x	  �  {  y	  �   z	     o         �t�bhhK ��h��R�(KK
��h�C(   {	    6      �   �   �         �t�bhhK ��h��R�(KK��h�CP
      �  e  �     ?     6      �  �   �  |	     �      }	        �t�bhhK ��h��R�(KK��h�C~	  �         �t�bhhK ��h��R�(KK��h�Ct   3   V     �t�bhhK ��h��R�(KK��h�C4p  /     O     �     	  	   �	  �	        �t�bhhK ��h��R�(KK��h�C�  #      �t�bhhK ��h��R�(KK��h�C         �      1      �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Cn   G      �t�bhhK ��h��R�(KK��h�C0
   r   $   q  6      =   �      �        �t�bhhK ��h��R�(KK��h�C,�	  T   ;      �	     $   ?   �         �t�bhhK ��h��R�(KK
��h�C(   �  �  �	     $      �         �t�bhhK ��h��R�(KK��h�C8      =   L  M   &   r  s     �      �        �t�bhhK ��h��R�(KK��h�C<2  �	       �  6  �   G   	   �     �  y        �t�bhhK ��h��R�(KK��h�Cd   L    4   $      q  �  	   5        >  
   f   M   &   r  s     �      �        �t�bhhK ��h��R�(KK��h�C �  "   �   
   �	  G         �t�bhhK ��h��R�(KK��h�C4            t   3   0      K   �  2         �t�bhhK ��h��R�(KK��h�C         n   G         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Ca           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�	           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C`           �t�bhhK ��h��R�(KK��h�C�   �  G      �t�bhhK ��h��R�(KK��h�CP   �	  �	  V       c      Y   ;  A  I   
   �	  	   �      �	        �t�bhhK ��h��R�(KK��h�C,�	     Y   ;  A  I   �     �	        �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�  �	           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C<
      5   �	     �   �   6      �   �	  r          �t�bhhK ��h��R�(KK
��h�C(�	  b  �   ]         �      �	     �t�bhhK ��h��R�(KK��h�C�	       �t�bhhK ��h��R�(KK��h�Cp  �  	   �  #      �t�bhhK ��h��R�(KK��h�C�	       �t�bhhK ��h��R�(KK��h�C�	       �t�bhhK ��h��R�(KK��h�C�	  �  	   �   #      �t�bhhK ��h��R�(KK��h�C8       �t�bhhK ��h��R�(KK��h�C�  �  	   �  	   8     �t�bhhK ��h��R�(KK��h�C�       �t�bhhK ��h��R�(KK��h�CY       �t�bhhK ��h��R�(KK��h�C�  �  	   �  Y     �t�bhhK ��h��R�(KK��h�C4\     \     �  �	  6  �	     3  �        �t�bhhK ��h��R�(KK��h�C@�   �   �  �  �     �  	   �  	   �	     �           �t�bhhK ��h��R�(KK��h�C4   �  O      �  �     �	  �	     �	        �t�bhhK ��h��R�(KK7��h�Cܝ	     �  	   �     �	     �      t     �	     �	     t   3   0      K   R   	   p  /     O  	   �  #      �  C  	     �	     	   �	  y      	     �  \   B     �  y      u     �        �t�bhhK ��h��R�(KK��h�C@         �	  �     �   2      �  =   e  M   ]         �t�bhhK ��h��R�(KK��h�C4   �   �  e  �   �        �      �	        �t�bhhK ��h��R�(KK��h�CPN      U     �   6      w      �	  	   �	     4   "      �	  }         �t�bhhK ��h��R�(KK
��h�C(�   �   �  �  �     �           �t�bhhK ��h��R�(KK��h�Cd�	  �     �	  �	  �	     �	  �	  �  �	     y      �  �	  u  	   �        �     �	     �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�	           �t�bhhK ��h��R�(KK��h�C�   G      �t�bhhK ��h��R�(KK��h�CP   ,      J   `  G   6         �  �   =   J   �   �      �	          �t�bhhK ��h��R�(KK	��h�C$   �   ,   	   =   �	  �	        �t�bhhK ��h��R�(KK��h�C         �   G         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Ct           �t�bhhK ��h��R�(KK��h�C4  G      �t�bhhK ��h��R�(KK��h�CL
      �	         5      
   �     �        =   J   �   �         �t�bhhK ��h��R�(KK��h�C`�   }      �   
      5   
  	   �      �      �     u         �	        �        �t�bhhK ��h��R�(KK��h�CD      -   �      }   d      �        �	     �	  �        �t�bhhK ��h��R�(KK��h�C8   �	        =   &   r  s     �      �        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Ct           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�	           �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�C4w   �      L  �      m            �        �t�bhhK ��h��R�(KK��h�C@   L  n  B      �  	   �      �  A  �  ?   �        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�CN      u  $         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Co           �t�bhhK ��h��R�(KK��h�CT     �t�bhhK ��h��R�(KK��h�C�     x  �   �         �t�bhhK ��h��R�(KK��h�CT
      �        �   �	  �   J   T  �	  �     
      �   �   
   f         �t�bhhK ��h��R�(KK��h�Ct�      U       6      �   �	  �	  y      �     O       \  �     �   &   �  �  �  �	  �	        �t�bhhK ��h��R�(KK��h�C�      �        �t�bhhK ��h��R�(KK��h�Cp  /     O  	      �t�bhhK ��h��R�(KK��h�C�  #      �t�bhhK ��h��R�(KK��h�C ]         �      �	        �t�bhhK ��h��R�(KK��h�C         T        �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�	           �t�bhhK ��h��R�(KK��h�C-     �t�bhhK ��h��R�(KK��h�C       �   -     �        �t�bhhK ��h��R�(KK	��h�C$      �     �     a        �t�bhhK ��h��R�(KK��h�C8      -   �   �     4         J   �   �        �t�bhhK ��h��R�(KK��h�C         -        �t�bhhK ��h��R�(KK��h�C�   Y      �t�bhhK ��h��R�(KK��h�Cl   �  �  �	     #   "   �       �	  :   ;          5        �	     :          ]        �t�bhhK ��h��R�(KK��h�C\�	     �     �     v  �     �  {  -   �	  �  ;      �          D  �        �t�bhhK ��h��R�(KK��h�C`   �      �      #     t   3   0      K   R   	   v   B      i   
   ;      �	        �t�bhhK ��h��R�(KK��h�C8;      ^   >   �    -      Y      �	  �        �t�bhhK ��h��R�(KK��h�C�  ;   �	  �   e         �t�bhhK ��h��R�(KK��h�C�	     �t�bhhK ��h��R�(KK��h�C�	     �	  �     �      �t�bhhK ��h��R�(KK��h�C�	     �     �t�bhhK ��h��R�(KK��h�C  +      �     �t�bhhK ��h��R�(KK��h�C�	     �t�bhhK ��h��R�(KK��h�C,V      |     Y   ?   A     �	        �t�bhhK ��h��R�(KK��h�CT�      .   c      i   
   �	  	   �	       o   \     d   &   �   �        �t�bhhK ��h��R�(KK��h�CX      
   ;      �   O      U   t   3   0      K   �  �	  �   ]      �	        �t�bhhK ��h��R�(KK��h�C         �   Y         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C;      �           �t�bhhK ��h��R�(KK��h�C�     �           �t�bhhK ��h��R�(KK��h�C�      &   [   �     �t�bhhK ��h��R�(KK��h�C'   �  $      �t�bhhK ��h��R�(KK��h�C0.  V     $      �  �   �     @        �t�bhhK ��h��R�(KK
��h�C(=   #   Q   �         
   �	        �t�bhhK ��h��R�(KK��h�C8      >  �	  
         
   ;      @  T         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK	��h�C$�  /     �  �     �        �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C]      �	     �t�bhhK ��h��R�(KK��h�C          '   �  $         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C;      �           �t�bhhK ��h��R�(KK��h�C�     �           �t�bhhK ��h��R�(KK��h�C�      &   [   �     �t�bhhK ��h��R�(KK��h�C�      #      �t�bhhK ��h��R�(KK��h�C�   �  G      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�   G      �t�bhhK ��h��R�(KK��h�C4  G      �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�CT     �t�bhhK ��h��R�(KK��h�C-     �t�bhhK ��h��R�(KK��h�C�   Y      �t�bhhK ��h��R�(KK��h�C'   �  $      �t�bhhK ��h��R�(KK��h�C�      #      �t�bhhK ��h��R�(KK��h�C,   #      5     >   ?     �         �t�bhhK ��h��R�(KK��h�C\d  �   "   '   �   w     b  	      B      �          �   }      �     @        �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C#   h	     �t�bhhK ��h��R�(KK��h�Cp  �     �t�bhhK ��h��R�(KK��h�C�  #      �t�bhhK ��h��R�(KK��h�C]         �      �     �t�bhhK ��h��R�(KK��h�CD   #   �  �  i	     �     j	     �  z  �  k	           �t�bhhK ��h��R�(KK��h�C<l	  O      }      m	  	   �     n	  R      �        �t�bhhK ��h��R�(KK��h�C@�     �  �     '        w  	      �      o	        �t�bhhK ��h��R�(KK��h�C�  #      �t�bhhK ��h��R�(KK��h�C]         �      �     �t�bhhK ��h��R�(KK��h�C  �  8     �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C�  8     �t�bhhK ��h��R�(KK��h�C]         �      p	     �t�bhhK ��h��R�(KK��h�C  �  �     �t�bhhK ��h��R�(KK��h�C]         �      q	     �t�bhhK ��h��R�(KK��h�C  �  Y     �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C�  Y     �t�bhhK ��h��R�(KK��h�C]         �      r	     �t�bhhK ��h��R�(KK��h�CH
      U          1   6      �  s	  
      t	     u	        �t�bhhK ��h��R�(KK��h�C         G         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Ct           �t�bhhK ��h��R�(KK	��h�C$?   �          �  �        �t�bhhK ��h��R�(KK
��h�C(�   �  v	  �     w	     e        �t�bhhK ��h��R�(KK��h�C8e     �     x	  �  {  y	  �   z	     o         �t�bhhK ��h��R�(KK
��h�C(   {	    6      �   �   �         �t�bhhK ��h��R�(KK��h�CP
      �  e  �     ?     6      �  �   �  |	     �      }	        �t�bhhK ��h��R�(KK��h�C~	  �         �t�bhhK ��h��R�(KK��h�Ct   3   V     �t�bhhK ��h��R�(KK��h�C4p  /     O     �     	  	   �	  �	        �t�bhhK ��h��R�(KK��h�C�  #      �t�bhhK ��h��R�(KK��h�C         �      1      �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Cn   G      �t�bhhK ��h��R�(KK��h�C0
   r   $   q  6      =   �      �        �t�bhhK ��h��R�(KK��h�C,�	  T   ;      �	     $   ?   �         �t�bhhK ��h��R�(KK
��h�C(   �  �  �	     $      �         �t�bhhK ��h��R�(KK��h�C8      =   L  M   &   r  s     �      �        �t�bhhK ��h��R�(KK��h�C<2  �	       �  6  �   G   	   �     �  y        �t�bhhK ��h��R�(KK��h�Cd   L    4   $      q  �  	   5        >  
   f   M   &   r  s     �      �        �t�bhhK ��h��R�(KK��h�C �  "   �   
   �	  G         �t�bhhK ��h��R�(KK��h�C4            t   3   0      K   �  2         �t�bhhK ��h��R�(KK��h�C         n   G         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Ca           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�	           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C`           �t�bhhK ��h��R�(KK��h�C�   �  G      �t�bhhK ��h��R�(KK��h�CP   �	  �	  V       c      Y   ;  A  I   
   �	  	   �      �	        �t�bhhK ��h��R�(KK��h�C,�	     Y   ;  A  I   �     �	        �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�  �	           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C<
      5   �	     �   �   6      �   �	  r          �t�bhhK ��h��R�(KK
��h�C(�	  b  �   ]         �      �	     �t�bhhK ��h��R�(KK��h�C�	       �t�bhhK ��h��R�(KK��h�Cp  �  	   �  #      �t�bhhK ��h��R�(KK��h�C�	       �t�bhhK ��h��R�(KK��h�C�	       �t�bhhK ��h��R�(KK��h�C�	  �  	   �   #      �t�bhhK ��h��R�(KK��h�C8       �t�bhhK ��h��R�(KK��h�C�  �  	   �  	   8     �t�bhhK ��h��R�(KK��h�C�       �t�bhhK ��h��R�(KK��h�CY       �t�bhhK ��h��R�(KK��h�C�  �  	   �  Y     �t�bhhK ��h��R�(KK��h�C4\     \     �  �	  6  �	     3  �        �t�bhhK ��h��R�(KK��h�C@�   �   �  �  �     �  	   �  	   �	     �           �t�bhhK ��h��R�(KK��h�C4   �  O      �  �     �	  �	     �	        �t�bhhK ��h��R�(KK7��h�Cܝ	     �  	   �     �	     �      t     �	     �	     t   3   0      K   R   	   p  /     O  	   �  #      �  C  	     �	     	   �	  y      	     �  \   B     �  y      u     �        �t�bhhK ��h��R�(KK��h�C@         �	  �     �   2      �  =   e  M   ]         �t�bhhK ��h��R�(KK��h�C4   �   �  e  �   �        �      �	        �t�bhhK ��h��R�(KK��h�CPN      U     �   6      w      �	  	   �	     4   "      �	  }         �t�bhhK ��h��R�(KK
��h�C(�   �   �  �  �     �           �t�bhhK ��h��R�(KK��h�Cd�	  �     �	  �	  �	     �	  �	  �  �	     y      �  �	  u  	   �        �     �	     �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�	           �t�bhhK ��h��R�(KK��h�C�   G      �t�bhhK ��h��R�(KK��h�CP   ,      J   `  G   6         �  �   =   J   �   �      �	          �t�bhhK ��h��R�(KK	��h�C$   �   ,   	   =   �	  �	        �t�bhhK ��h��R�(KK��h�C         �   G         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Ct           �t�bhhK ��h��R�(KK��h�C4  G      �t�bhhK ��h��R�(KK��h�CL
      �	         5      
   �     �        =   J   �   �         �t�bhhK ��h��R�(KK��h�C`�   }      �   
      5   
  	   �      �      �     u         �	        �        �t�bhhK ��h��R�(KK��h�CD      -   �      }   d      �        �	     �	  �        �t�bhhK ��h��R�(KK��h�C8   �	        =   &   r  s     �      �        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C4  G      �        �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Ct           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�	           �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�C4w   �      L  �      m            �        �t�bhhK ��h��R�(KK��h�C@   L  n  B      �  	   �      �  A  �  ?   �        �t�bhhK ��h��R�(KK��h�C          �     T        �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Co           �t�bhhK ��h��R�(KK��h�CT     �t�bhhK ��h��R�(KK��h�C�     x  �   �         �t�bhhK ��h��R�(KK��h�CT
      �        �   �	  �   J   T  �	  �     
      �   �   
   f         �t�bhhK ��h��R�(KK��h�Ct�      U       6      �   �	  �	  y      �     O       \  �     �   &   �  �  �  �	  �	        �t�bhhK ��h��R�(KK��h�C�      �        �t�bhhK ��h��R�(KK��h�Cp  /     O  	      �t�bhhK ��h��R�(KK��h�C�  #      �t�bhhK ��h��R�(KK��h�C ]         �      �	        �t�bhhK ��h��R�(KK��h�C          �     T        �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�	           �t�bhhK ��h��R�(KK��h�C-     �t�bhhK ��h��R�(KK��h�C       �   -     �        �t�bhhK ��h��R�(KK	��h�C$      �     �     a        �t�bhhK ��h��R�(KK��h�C8      -   �   �     4         J   �   �        �t�bhhK ��h��R�(KK��h�C         -        �t�bhhK ��h��R�(KK��h�C�   Y      �t�bhhK ��h��R�(KK��h�Cl   �  �  �	     #   "   �       �	  :   ;          5        �	     :          ]        �t�bhhK ��h��R�(KK��h�C\�	     �     �     v  �     �  {  -   �	  �  ;      �          D  �        �t�bhhK ��h��R�(KK��h�C`   �      �      #     t   3   0      K   R   	   v   B      i   
   ;      �	        �t�bhhK ��h��R�(KK��h�C8;      ^   >   �    -      Y      �	  �        �t�bhhK ��h��R�(KK��h�C�  ;   �	  �   e         �t�bhhK ��h��R�(KK��h�C�	     �t�bhhK ��h��R�(KK��h�C�	     �	  �     �      �t�bhhK ��h��R�(KK��h�C�	     �     �t�bhhK ��h��R�(KK��h�C  +      �     �t�bhhK ��h��R�(KK��h�C�	     �t�bhhK ��h��R�(KK��h�C,V      |     Y   ?   A     �	        �t�bhhK ��h��R�(KK��h�CT�      .   c      i   
   �	  	   �	       o   \     d   &   �   �        �t�bhhK ��h��R�(KK��h�CX      
   ;      �   O      U   t   3   0      K   �  �	  �   ]      �	        �t�bhhK ��h��R�(KK��h�C         �   Y         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C;      �           �t�bhhK ��h��R�(KK��h�C�     �           �t�bhhK ��h��R�(KK��h�C�      &   [   �     �t�bhhK ��h��R�(KK��h�C'   �  $      �t�bhhK ��h��R�(KK��h�C0.  V     $      �  �   �     @        �t�bhhK ��h��R�(KK
��h�C(=   #   Q   �         
   �	        �t�bhhK ��h��R�(KK��h�C8      >  �	  
         
   ;      @  T         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK	��h�C$�  /     �  �     �        �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C]      �	     �t�bhhK ��h��R�(KK��h�C          '   �  $         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C;      �           �t�bhhK ��h��R�(KK��h�C�     �           �t�bhhK ��h��R�(KK��h�C�      &   [   �     �t�bhhK ��h��R�(KK��h�C1     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK��h�C s      .   �   �     C      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CL   �   �      �t�bhhK ��h��R�(KK��h�Cz     �t�bhhK ��h��R�(KK��h�CW   �     �t�bhhK ��h��R�(KK��h�C1     �t�bhhK ��h��R�(KK��h�C8   #      H   �   �   	   �  	   l  \   �        �t�bhhK ��h��R�(KK��h�CP�      .   �      p     �     	   '   �   �      �   l     #         �t�bhhK ��h��R�(KK��h�Cp      i   
      �   �     r   $   m  M   q   �	           �     H   2      `      �           �t�bhhK ��h��R�(KK��h�C8`   6   �  �   �   n       5      �   �        �t�bhhK ��h��R�(KK��h�CT.      c      @         q  
   &   r            �  s  �      �         �t�bhhK ��h��R�(KK��h�C\`      �     t     1  	   �     1     �     u     &   v  w     �        �t�bhhK ��h��R�(KK��h�CH      i   
            H   �     �           H   2         �t�bhhK ��h��R�(KK��h�C,`      -   �  �        y  �         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C;      1     �t�bhhK ��h��R�(KK��h�Cx     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C�      W   y           �t�bhhK ��h��R�(KK��h�Cz           �t�bhhK ��h��R�(KK��h�C{           �t�bhhK ��h��R�(KK��h�C     i   
   |  �           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C4#      T   �  �         �  I   �	  $         �t�bhhK ��h��R�(KK��h�Cl  V     �	     X      �	     w  �	  �  
   �  	       �   �  
   �	  	   6  j  �	        �t�bhhK ��h��R�(KK��h�C     �        �t�bhhK ��h��R�(KK��h�CX
   z   �   5     �	  +  �  �       x       	   �     $     �	        �t�bhhK ��h��R�(KK
��h�C(�	       y          �	        �t�bhhK ��h��R�(KK
��h�C(�  �	     �	        H   2         �t�bhhK ��h��R�(KK��h�C|
      4   �  '   �	  
   �     �   
   �  ?   z  }      �  	   w   �      �     1  �   ]      �  �	        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK��h�C\   1   "      $      �  �  I   �	  	     �      :   �   �      &   [            �t�bhhK ��h��R�(KK��h�C4�	  �	     �     .   �  �   z   �  _        �t�bhhK ��h��R�(KK��h�C8.            "   �	         z   �     @        �t�bhhK ��h��R�(KK
��h�C(�     �  y     �     �        �t�bhhK ��h��R�(KK��h�C4   H   2      �  �            
   �        �t�bhhK ��h��R�(KK��h�C@
      "   �   
   &   [            -   =   H   �        �t�bhhK ��h��R�(KK��h�C4d  $        �  "   �                    �t�bhhK ��h��R�(KK��h�CD
   z        #   ?   �            �	  f     @        �t�bhhK ��h��R�(KK%��h�C�
   z   �    �     )                �           �  �	         �     �   s         �            �  6  .   �   �	        �t�bhhK ��h��R�(KK��h�C`   #      {     &   �         �	     �	  �     �	  �        �	     �	          �t�bhhK ��h��R�(KK��h�C8�	     &   �    y  �     �  6    �	        �t�bhhK ��h��R�(KK��h�CLs           �	  )      W   k      �	       �	  �     �         �t�bhhK ��h��R�(KK��h�C@V      �	  �     C     �       �   f     @        �t�bhhK ��h��R�(KK��h�C<      
   &   �        C   O         H   �        �t�bhhK ��h��R�(KK��h�C         [   X         �t�bhhK ��h��R�(KK��h�C�      &   [   �     �t�bhhK ��h��R�(KK��h�C s      .   �   �     C      �t�bhhK ��h��R�(KK��h�Cps        �   f  �     #      ^   >   k   	      F   ?   �       �	  �	  s      �	  >   k         �t�bhhK ��h��R�(KK��h�C �	  6   �  w  �           �t�bhhK ��h��R�(KK��h�CH  y  �     :     v   .      �	         �      �         �t�bhhK ��h��R�(KK��h�CP     �   �   �	  �   e   �	  	    
     �  �   	   
     �          �t�bhhK ��h��R�(KK��h�CX   
   s        �   f     �   O         
          >   �     
        �t�bhhK ��h��R�(KK��h�C(   
     �t�bhhK ��h��R�(KK��h�CX      �      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CLt   3   
  T   �      #   	   8  	   
  	     	   
     �        �t�bhhK ��h��R�(KK��h�Cp�  �  -   
  X      [   �   	   	
     �     X   \   �   

     �   C      t   3   	     8        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�CP   3           �t�bhhK ��h��R�(KK��h�Ct   3   
           �t�bhhK ��h��R�(KK��h�CP   3           �t�bhhK ��h��R�(KK��h�CX      �            �t�bhhK ��h��R�(KK��h�CP   3   	        �t�bhhK ��h��R�(KK��h�C
  
     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C\   #   V  |     �      #   )   �      #      �   	   \      �      #   
        �t�bhhK ��h��R�(KK ��h�C�   |     �   �   B   ?   
  M   
  �          B      �  
  
   B      
  U   �  "   �  
  
     
        �t�bhhK ��h��R�(KK��h�C0      i      �  .  d   
  �  �         �t�bhhK ��h��R�(KK��h�C4#   )   �   T   �   s      �  -      C         �t�bhhK ��h��R�(KK��h�Cp&   �        �     '   �          &          �  
          '   e   f      D     �        �t�bhhK ��h��R�(KK��h�C,d  I   
  '   
  �  
   
  
        �t�bhhK ��h��R�(KK	��h�C$   d      '   �   
        �t�bhhK ��h��R�(KK��h�C8B   �      �   s      �  ?   �     
  
        �t�bhhK ��h��R�(KK��h�CL
        #   )   �      #   
     )            #      �         �t�bhhK ��h��R�(KK��h�C<   #   )   �   �  s      )      �     C   C         �t�bhhK ��h��R�(KK��h�CL         
  6   D     �     g  �  �  g   a      �  R        �t�bhhK ��h��R�(KK��h�C@      
    
     &   �        �  �     H   �        �t�bhhK ��h��R�(KK
��h�C(P             H   !
  2         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK	��h�C$�  /     �  �     �        �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C]      "
     �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C#
                �t�bhhK ��h��R�(KK��h�CL   �   �      �t�bhhK ��h��R�(KK��h�C<L      �  �      �      @   +      .     �        �t�bhhK ��h��R�(KK��h�C`.     �  x   L      �  h     �  I   E  �   ;      V      X   	   �      $
        �t�bhhK ��h��R�(KK"��h�C�:     �     %
  x          D  y  &   _   &
  	   '
  �  �   	   �    d   >   {  	      p       6  &   _   (
        �t�bhhK ��h��R�(KK��h�C  )
           �t�bhhK ��h��R�(KK��h�Cz     �t�bhhK ��h��R�(KK��h�CD   �  �     B   �   �     /  	   *
  	   0      �        �t�bhhK ��h��R�(KK��h�C0B      -   �      	  �   +
     ,
        �t�bhhK ��h��R�(KK��h�C0.      �   c      �      &   �   �        �t�bhhK ��h��R�(KK��h�C8   #   -
  �     B   �   
  .
  �     /
        �t�bhhK ��h��R�(KK��h�C,   �  �  -   0
     1
  2
  �        �t�bhhK ��h��R�(KK��h�C         z        �t�bhhK ��h��R�(KK��h�C3
     4
     �t�bhhK ��h��R�(KK��h�C5
  �        �t�bhhK ��h��R�(KK��h�C�                   �t�bhhK ��h��R�(KK��h�C6
  7
                 �t�bhhK ��h��R�(KK��h�CW   �     �t�bhhK ��h��R�(KK��h�CX�   W  	           8
     #      	      '   9
     )                    �t�bhhK ��h��R�(KK��h�CX  T   s      :
  	   �   	   �     �  	   �  	   �  	        �  �        �t�bhhK ��h��R�(KK��h�Cp  T   -   s      ^   >   k   	   �   e   )   	      	      	   }  	   �   	   E   	   /             �t�bhhK ��h��R�(KK��h�CP;
  <
  U   I      I   	   i  .   8  a       �  �  �      ]  2         �t�bhhK ��h��R�(KK��h�C C   V  �     �  �         �t�bhhK ��h��R�(KK��h�C8   =
  >
  
   .      c      @   �     ?
        �t�bhhK ��h��R�(KK��h�C,�     ]  2   _  �         �        �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C]      @
  	   A
     �t�bhhK ��h��R�(KK��h�Ch   t   3   �        �  �      B
     .   �   �  	   �      C
  �   \   �  �     D
        �t�bhhK ��h��R�(KK��h�C0?   �     .   c      E
  F
     G
        �t�bhhK ��h��R�(KK��h�C8�      .   -   c      �  H
  I
     J
  K
        �t�bhhK ��h��R�(KK��h�C L
  �      �     M
        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�CR     �  	   N
     �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK	��h�C$�   �                       �t�bhhK ��h��R�(KK��h�CP   3   �        �t�bhhK ��h��R�(KK��h�Ct   3   O
     �t�bhhK ��h��R�(KK��h�C�  s      �           �t�bhhK ��h��R�(KK��h�C1     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK��h�C s      .   �   �     C      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CL   �   �      �t�bhhK ��h��R�(KK��h�Cz     �t�bhhK ��h��R�(KK��h�CW   �     �t�bhhK ��h��R�(KK��h�C1     �t�bhhK ��h��R�(KK��h�C8   #      H   �   �   	   �  	   l  \   �        �t�bhhK ��h��R�(KK��h�CP�      .   �      p     �     	   '   �   �      �   l     #         �t�bhhK ��h��R�(KK��h�Cp      i   
      �   �     r   $   m  M   q   �	           �     H   2      `      �           �t�bhhK ��h��R�(KK��h�C8`   6   �  �   �   n       5      �   �        �t�bhhK ��h��R�(KK��h�CT.      c      @         q  
   &   r            �  s  �      �         �t�bhhK ��h��R�(KK��h�C\`      �     t     1  	   �     1     �     u     &   v  w     �        �t�bhhK ��h��R�(KK��h�CH      i   
            H   �     �           H   2         �t�bhhK ��h��R�(KK��h�C,`      -   �  �        y  �         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C;      1     �t�bhhK ��h��R�(KK��h�Cx     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C�      W   y           �t�bhhK ��h��R�(KK��h�Cz           �t�bhhK ��h��R�(KK��h�C{           �t�bhhK ��h��R�(KK��h�C     i   
   |  �           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C4#      T   �  �         �  I   �	  $         �t�bhhK ��h��R�(KK��h�Cl  V     �	     X      �	     w  �	  �  
   �  	       �   �  
   �	  	   6  j  �	        �t�bhhK ��h��R�(KK��h�C     �        �t�bhhK ��h��R�(KK��h�CX
   z   �   5     �	  +  �  �       x       	   �     $     �	        �t�bhhK ��h��R�(KK
��h�C(�	       y          �	        �t�bhhK ��h��R�(KK
��h�C(�  �	     �	        H   2         �t�bhhK ��h��R�(KK��h�C|
      4   �  '   �	  
   �     �   
   �  ?   z  }      �  	   w   �      �     1  �   ]      �  �	        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK��h�C\   1   "      $      �  �  I   �	  	     �      :   �   �      &   [            �t�bhhK ��h��R�(KK��h�C4�	  �	     �     .   �  �   z   �  _        �t�bhhK ��h��R�(KK��h�C8.            "   �	         z   �     @        �t�bhhK ��h��R�(KK
��h�C(�     �  y     �     �        �t�bhhK ��h��R�(KK��h�C4   H   2      �  �            
   �        �t�bhhK ��h��R�(KK��h�C@
      "   �   
   &   [            -   =   H   �        �t�bhhK ��h��R�(KK��h�C4d  $        �  "   �                    �t�bhhK ��h��R�(KK��h�CD
   z        #   ?   �            �	  f     @        �t�bhhK ��h��R�(KK%��h�C�
   z   �    �     )                �           �  �	         �     �   s         �            �  6  .   �   �	        �t�bhhK ��h��R�(KK��h�C`   #      {     &   �         �	     �	  �     �	  �        �	     �	          �t�b�      hhK ��h��R�(KK��h�C8�	     &   �    y  �     �  6    �	        �t�bhhK ��h��R�(KK��h�CLs           �	  )      W   k      �	       �	  �     �         �t�bhhK ��h��R�(KK��h�C@V      �	  �     C     �       �   f     @        �t�bhhK ��h��R�(KK��h�C<      
   &   �        C   O         H   �        �t�bhhK ��h��R�(KK��h�C         [   X         �t�bhhK ��h��R�(KK��h�C�      &   [   �     �t�bhhK ��h��R�(KK��h�C s      .   �   �     C      �t�bhhK ��h��R�(KK��h�Cps        �   f  �     #      ^   >   k   	      F   ?   �       �	  �	  s      �	  >   k         �t�bhhK ��h��R�(KK��h�C �	  6   �  w  �           �t�bhhK ��h��R�(KK��h�CH  y  �     :     v   .      �	         �      �         �t�bhhK ��h��R�(KK��h�CP     �   �   �	  �   e   �	  	    
     �  �   	   
     �          �t�bhhK ��h��R�(KK��h�CX   
   s        �   f     �   O         
          >   �     
        �t�bhhK ��h��R�(KK��h�C(   
     �t�bhhK ��h��R�(KK��h�CX      �      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CLt   3   
  T   �      #   	   8  	   
  	     	   
     �        �t�bhhK ��h��R�(KK��h�Cp�  �  -   
  X      [   �   	   	
     �     X   \   �   

     �   C      t   3   	     8        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�CP   3           �t�bhhK ��h��R�(KK��h�Ct   3   
           �t�bhhK ��h��R�(KK��h�CP   3           �t�bhhK ��h��R�(KK��h�CX      �            �t�bhhK ��h��R�(KK��h�CP   3   	        �t�bhhK ��h��R�(KK��h�C
  
     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C\   #   V  |     �      #   )   �      #      �   	   \      �      #   
        �t�bhhK ��h��R�(KK ��h�C�   |     �   �   B   ?   
  M   
  �          B      �  
  
   B      
  U   �  "   �  
  
     
        �t�bhhK ��h��R�(KK��h�C0      i      �  .  d   
  �  �         �t�bhhK ��h��R�(KK��h�C4#   )   �   T   �   s      �  -      C         �t�bhhK ��h��R�(KK��h�Cp&   �        �     '   �          &          �  
          '   e   f      D     �        �t�bhhK ��h��R�(KK��h�C,d  I   
  '   
  �  
   
  
        �t�bhhK ��h��R�(KK	��h�C$   d      '   �   
        �t�bhhK ��h��R�(KK��h�C8B   �      �   s      �  ?   �     
  
        �t�bhhK ��h��R�(KK��h�CL
        #   )   �      #   
     )            #      �         �t�bhhK ��h��R�(KK��h�C<   #   )   �   �  s      )      �     C   C         �t�bhhK ��h��R�(KK��h�CL         
  6   D     �     g  �  �  g   a      �  R        �t�bhhK ��h��R�(KK��h�C@      
    
     &   �        �  �     H   �        �t�bhhK ��h��R�(KK
��h�C(P             H   !
  2         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK	��h�C$�  /     �  �     �        �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C]      "
     �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C#
                �t�bhhK ��h��R�(KK��h�CL   �   �      �t�bhhK ��h��R�(KK��h�C<L      �  �      �      @   +      .     �        �t�bhhK ��h��R�(KK��h�C`.     �  x   L      �  h     �  I   E  �   ;      V      X   	   �      $
        �t�bhhK ��h��R�(KK"��h�C�:     �     %
  x          D  y  &   _   &
  	   '
  �  �   	   �    d   >   {  	      p       6  &   _   (
        �t�bhhK ��h��R�(KK��h�C  )
           �t�bhhK ��h��R�(KK��h�Cz     �t�bhhK ��h��R�(KK��h�CD   �  �     B   �   �     /  	   *
  	   0      �        �t�bhhK ��h��R�(KK��h�C0B      -   �      	  �   +
     ,
        �t�bhhK ��h��R�(KK��h�C0.      �   c      �      &   �   �        �t�bhhK ��h��R�(KK��h�C8   #   -
  �     B   �   
  .
  �     /
        �t�bhhK ��h��R�(KK��h�C,   �  �  -   0
     1
  2
  �        �t�bhhK ��h��R�(KK��h�C         z        �t�bhhK ��h��R�(KK��h�C3
     4
     �t�bhhK ��h��R�(KK��h�C5
  �        �t�bhhK ��h��R�(KK��h�C�                   �t�bhhK ��h��R�(KK��h�C6
  7
                 �t�bhhK ��h��R�(KK��h�CW   �     �t�bhhK ��h��R�(KK��h�CX�   W  	           8
     #      	      '   9
     )                    �t�bhhK ��h��R�(KK��h�CX  T   s      :
  	   �   	   �     �  	   �  	   �  	        �  �        �t�bhhK ��h��R�(KK��h�Cp  T   -   s      ^   >   k   	   �   e   )   	      	      	   }  	   �   	   E   	   /             �t�bhhK ��h��R�(KK��h�CP;
  <
  U   I      I   	   i  .   8  a       �  �  �      ]  2         �t�bhhK ��h��R�(KK��h�C C   V  �     �  �         �t�bhhK ��h��R�(KK��h�C8   =
  >
  
   .      c      @   �     ?
        �t�bhhK ��h��R�(KK��h�C,�     ]  2   _  �         �        �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C]      @
  	   A
     �t�bhhK ��h��R�(KK��h�Ch   t   3   �        �  �      B
     .   �   �  	   �      C
  �   \   �  �     D
        �t�bhhK ��h��R�(KK��h�C0?   �     .   c      E
  F
     G
        �t�bhhK ��h��R�(KK��h�C8�      .   -   c      �  H
  I
     J
  K
        �t�bhhK ��h��R�(KK��h�C L
  �      �     M
        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�CR     �  	   N
     �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK	��h�C$�   �                       �t�bhhK ��h��R�(KK��h�CP   3   �        �t�bhhK ��h��R�(KK��h�Ct   3   O
     �t�bhhK ��h��R�(KK��h�C�  s      �           �t�bhhK ��h��R�(KK��h�C1     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK��h�C s      .   �   �     C      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�be(hhK ��h��R�(KK��h�CL   �   �      �t�bhhK ��h��R�(KK��h�Cz     �t�bhhK ��h��R�(KK��h�CW   �     �t�bhhK ��h��R�(KK��h�C1     �t�bhhK ��h��R�(KK��h�C8   #      H   �   �   	   �  	   l  \   �        �t�bhhK ��h��R�(KK��h�CP�      .   �      p     �     	   '   �   �      �   l     #         �t�bhhK ��h��R�(KK��h�Cp      i   
      �   �     r   $   m  M   q   �	           �     H   2      `      �           �t�bhhK ��h��R�(KK��h�C8`   6   �  �   �   n       5      �   �        �t�bhhK ��h��R�(KK��h�CT.      c      @         q  
   &   r            �  s  �      �         �t�bhhK ��h��R�(KK��h�C\`      �     t     1  	   �     1     �     u     &   v  w     �        �t�bhhK ��h��R�(KK��h�CH      i   
            H   �     �           H   2         �t�bhhK ��h��R�(KK��h�C,`      -   �  �        y  �         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C;      1     �t�bhhK ��h��R�(KK��h�Cx     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C1        �t�bhhK ��h��R�(KK��h�C�      W   y           �t�bhhK ��h��R�(KK��h�Cz           �t�bhhK ��h��R�(KK��h�C{           �t�bhhK ��h��R�(KK��h�C     i   
   |  �           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C4#      T   �  �         �  I   �	  $         �t�bhhK ��h��R�(KK��h�Cl  V     �	     X      �	     w  �	  �  
   �  	       �   �  
   �	  	   6  j  �	        �t�bhhK ��h��R�(KK��h�C     �        �t�bhhK ��h��R�(KK��h�CX
   z   �   5     �	  +  �  �       x       	   �     $     �	        �t�bhhK ��h��R�(KK
��h�C(�	       y          �	        �t�bhhK ��h��R�(KK
��h�C(�  �	     �	        H   2         �t�bhhK ��h��R�(KK��h�C|
      4   �  '   �	  
   �     �   
   �  ?   z  }      �  	   w   �      �     1  �   ]      �  �	        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK��h�C\   1   "      $      �  �  I   �	  	     �      :   �   �      &   [            �t�bhhK ��h��R�(KK��h�C4�	  �	     �     .   �  �   z   �  _        �t�bhhK ��h��R�(KK��h�C8.            "   �	         z   �     @        �t�bhhK ��h��R�(KK
��h�C(�     �  y     �     �        �t�bhhK ��h��R�(KK��h�C4   H   2      �  �            
   �        �t�bhhK ��h��R�(KK��h�C@
      "   �   
   &   [            -   =   H   �        �t�bhhK ��h��R�(KK��h�C4d  $        �  "   �                    �t�bhhK ��h��R�(KK��h�CD
   z        #   ?   �            �	  f     @        �t�bhhK ��h��R�(KK%��h�C�
   z   �    �     )                �           �  �	         �     �   s         �            �  6  .   �   �	        �t�bhhK ��h��R�(KK��h�C`   #      {     &   �         �	     �	  �     �	  �        �	     �	          �t�bhhK ��h��R�(KK��h�C8�	     &   �    y  �     �  6    �	        �t�bhhK ��h��R�(KK��h�CLs           �	  )      W   k      �	       �	  �     �         �t�bhhK ��h��R�(KK��h�C@V      �	  �     C     �       �   f     @        �t�bhhK ��h��R�(KK��h�C<      
   &   �        C   O         H   �        �t�bhhK ��h��R�(KK��h�C         [   X         �t�bhhK ��h��R�(KK��h�C�      &   [   �     �t�bhhK ��h��R�(KK��h�C s      .   �   �     C      �t�bhhK ��h��R�(KK��h�Cps        �   f  �     #      ^   >   k   	      F   ?   �       �	  �	  s      �	  >   k         �t�bhhK ��h��R�(KK��h�C �	  6   �  w  �           �t�bhhK ��h��R�(KK��h�CH  y  �     :     v   .      �	         �      �         �t�bhhK ��h��R�(KK��h�CP     �   �   �	  �   e   �	  	    
     �  �   	   
     �          �t�bhhK ��h��R�(KK��h�CX   
   s        �   f     �   O         
          >   �     
        �t�bhhK ��h��R�(KK��h�C(   
     �t�bhhK ��h��R�(KK��h�CX      �      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CLt   3   
  T   �      #   	   8  	   
  	     	   
     �        �t�bhhK ��h��R�(KK��h�Cp�  �  -   
  X      [   �   	   	
     �     X   \   �   

     �   C      t   3   	     8        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�CP   3           �t�bhhK ��h��R�(KK��h�Ct   3   
           �t�bhhK ��h��R�(KK��h�CP   3           �t�bhhK ��h��R�(KK��h�CX      �            �t�bhhK ��h��R�(KK��h�CP   3   	        �t�bhhK ��h��R�(KK��h�C
  
     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C\   #   V  |     �      #   )   �      #      �   	   \      �      #   
        �t�bhhK ��h��R�(KK ��h�C�   |     �   �   B   ?   
  M   
  �          B      �  
  
   B      
  U   �  "   �  
  
     
        �t�bhhK ��h��R�(KK��h�C0      i      �  .  d   
  �  �         �t�bhhK ��h��R�(KK��h�C4#   )   �   T   �   s      �  -      C         �t�bhhK ��h��R�(KK��h�Cp&   �        �     '   �          &          �  
          '   e   f      D     �        �t�bhhK ��h��R�(KK��h�C,d  I   
  '   
  �  
   
  
        �t�bhhK ��h��R�(KK	��h�C$   d      '   �   
        �t�bhhK ��h��R�(KK��h�C8B   �      �   s      �  ?   �     
  
        �t�bhhK ��h��R�(KK��h�CL
        #   )   �      #   
     )            #      �         �t�bhhK ��h��R�(KK��h�C<   #   )   �   �  s      )      �     C   C         �t�bhhK ��h��R�(KK��h�CL         
  6   D     �     g  �  �  g   a      �  R        �t�bhhK ��h��R�(KK��h�C@      
    
     &   �        �  �     H   �        �t�bhhK ��h��R�(KK
��h�C(P             H   !
  2         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK	��h�C$�  /     �  �     �        �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C]      "
     �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C#
                �t�bhhK ��h��R�(KK��h�CL   �   �      �t�bhhK ��h��R�(KK��h�C<L      �  �      �      @   +      .     �        �t�bhhK ��h��R�(KK��h�C`.     �  x   L      �  h     �  I   E  �   ;      V      X   	   �      $
        �t�bhhK ��h��R�(KK"��h�C�:     �     %
  x          D  y  &   _   &
  	   '
  �  �   	   �    d   >   {  	      p       6  &   _   (
        �t�bhhK ��h��R�(KK��h�C  )
           �t�bhhK ��h��R�(KK��h�Cz     �t�bhhK ��h��R�(KK��h�CD   �  �     B   �   �     /  	   *
  	   0      �        �t�bhhK ��h��R�(KK��h�C0B      -   �      	  �   +
     ,
        �t�bhhK ��h��R�(KK��h�C0.      �   c      �      &   �   �        �t�bhhK ��h��R�(KK��h�C8   #   -
  �     B   �   
  .
  �     /
        �t�bhhK ��h��R�(KK��h�C,   �  �  -   0
     1
  2
  �        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C}  	            �t�bhhK ��h��R�(KK��h�C3
     4
     �t�bhhK ��h��R�(KK��h�C5
  �        �t�bhhK ��h��R�(KK��h�C�                   �t�bhhK ��h��R�(KK��h�C6
  7
                 �t�bhhK ��h��R�(KK��h�CW   �     �t�bhhK ��h��R�(KK��h�CX�   W  	           8
     #      	      '   9
     )                    �t�bhhK ��h��R�(KK��h�CX  T   s      :
  	   �   	   �     �  	   �  	   �  	        �  �        �t�bhhK ��h��R�(KK��h�Cp  T   -   s      ^   >   k   	   �   e   )   	      	      	   }  	   �   	   E   	   /             �t�bhhK ��h��R�(KK��h�CP;
  <
  U   I      I   	   i  .   8  a       �  �  �      ]  2         �t�bhhK ��h��R�(KK��h�C C   V  �     �  �         �t�bhhK ��h��R�(KK��h�C8   =
  >
  
   .      c      @   �     ?
        �t�bhhK ��h��R�(KK��h�C,�     ]  2   _  �         �        �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C]      @
  	   A
     �t�bhhK ��h��R�(KK��h�Ch   t   3   �        �  �      B
     .   �   �  	   �      C
  �   \   �  �     D
        �t�bhhK ��h��R�(KK��h�C0?   �     .   c      E
  F
     G
        �t�bhhK ��h��R�(KK��h�C8�      .   -   c      �  H
  I
     J
  K
        �t�bhhK ��h��R�(KK��h�C L
  �      �     M
        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�CR     �  	   N
     �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK	��h�C$�   �                       �t�bhhK ��h��R�(KK��h�CP   3   �        �t�bhhK ��h��R�(KK��h�Ct   3   O
     �t�bhhK ��h��R�(KK��h�C�  s      �           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C  �      �t�bhhK ��h��R�(KK��h�Cj          �t�bhhK ��h��R�(KK��h�C7     �t�bhhK ��h��R�(KK��h�Ck     ~     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CD#   Q   �     `   
   �      P
        �  �              �t�bhhK ��h��R�(KK��h�CDQ
     �  6   R
  �   �     	   5     -   �  �            �t�bhhK ��h��R�(KK
��h�C(B      -   �   �   �     �        �t�bhhK ��h��R�(KK��h�C<S
     �  U      �  �              !        �t�bhhK ��h��R�(KK��h�C�  #      �t�bhhK ��h��R�(KK��h�C]      T
     �t�bhhK ��h��R�(KK��h�CHU
    �      V
  W
  	      T   X
  Y
  \   Z
     >   [
        �t�bhhK ��h��R�(KK��h�CD   \
        ]
  ^
     x    �      Y        _
        �t�bhhK ��h��R�(KK��h�C8
  `
     a
  �  b
  �     i   
      c
        �t�bhhK ��h��R�(KK��h�Cd
       �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C]      e
     �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C!           �t�bhhK ��h��R�(KK
��h�C(`   
   #   Q   f
                 �t�bhhK ��h��R�(KK��h�C�   6  g
           �t�bhhK ��h��R�(KK��h�Ch
           �t�bhhK ��h��R�(KK��h�C�   !           �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�CH:   �  #  �        i
  	   �        �      :   �  j        �t�bhhK ��h��R�(KK��h�CD   �  j
     .   O  "      �   �  �   �   B      k
        �t�bhhK ��h��R�(KK��h�CT�   e   d   l
  	      "          �     �  
   �           �        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C        �t�bhhK ��h��R�(KK��h�C  �      �t�bhhK ��h��R�(KK��h�C   �    >   m
        �t�bhhK ��h��R�(KK��h�CP     ?   ;  n
        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C  �         �t�bhhK ��h��R�(KK��h�C o
     �                 �t�bhhK ��h��R�(KK��h�CT
      �  �      �     �     �  6      =         �     �        �t�bhhK ��h��R�(KK��h�Ch
   J   �   "   �  	      F      �     �     �  	      �     �  �  �  :   �  �        �t�bhhK ��h��R�(KK
��h�C(=   r     .  N   �  "   �        �t�bhhK ��h��R�(KK��h�CL
           p
     �     l   	   w   �      #   D     �         �t�bhhK ��h��R�(KK��h�C,      �   #  ?      \     �         �t�bhhK ��h��R�(KK��h�C,   5   4     r   �  �      �        �t�bhhK ��h��R�(KK��h�C#   D     �      �t�bhhK ��h��R�(KK��h�C]      q
     �t�bhhK ��h��R�(KK��h�C!           �t�bhhK ��h��R�(KK��h�C#   D     �     �t�bhhK ��h��R�(KK��h�Cj          �t�bhhK ��h��R�(KK��h�CD�       �  �     t   3   0      K   R   \   �   r
        �t�bhhK ��h��R�(KK��h�CL     �      �     Y   ;  A  I      5   o        �   �         �t�bhhK ��h��R�(KK��h�CT     s
     Y      4   t
  �  a      �   �      ;      8     �         �t�bhhK ��h��R�(KK��h�C`      
   �  �     t   3   0      K   R   O         �   e   u
  v
  	   (   f        �t�bhhK ��h��R�(KK��h�CL   �      Y      w
  a   U   `  ,     �     x
  �  �  �        �t�bhhK ��h��R�(KK��h�CT      Y      "   �         D  �  �   +   	   �  �      �   Y         �t�bhhK ��h��R�(KK��h�C0;      �  �     �   e   y
     z
        �t�bhhK ��h��R�(KK��h�CP     {
         �    o        \   |
  �  }
  	   ~
     
        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�Cj             �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�
           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�  ;   	   �
           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK	��h�C$�  ;   	   �
     �
           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C �     �
     �           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�
           �t�bhhK ��h��R�(KK��h�C7     �t�bhhK ��h��R�(KK��h�C<
          �     =         �     �        �t�bhhK ��h��R�(KK��h�C!           �t�bhhK ��h��R�(KK��h�Ck     ~     �t�bhhK ��h��R�(KK��h�C   �  �  �        �t�bhhK ��h��R�(KK��h�C�
     �t�bhhK ��h��R�(KK��h�C�
     �
  �
     �t�bhhK ��h��R�(KK��h�C�
  U   �
     �
     �t�bhhK ��h��R�(KK��h�Cp$  �  �  �        �
  	      �
  �
        �
        �     �       O   �    �
          �t�bhhK ��h��R�(KK��h�C    �
  �
  6   �
  �
        �t�bhhK ��h��R�(KK��h�C   �  �  �        �t�bhhK ��h��R�(KK��h�C�
  	   �
     �
     �t�bhhK ��h��R�(KK
��h�C(�
     4   �
  	   �
     �
        �t�bhhK ��h��R�(KK��h�C0�  �
     �
     �
  �  �
     �
        �t�bhhK ��h��R�(KK��h�C,$  �  �  6   �     �     �
        �t�bhhK ��h��R�(KK��h�C,�       O   �      �          �t�bhhK ��h��R�(KK��h�C  �
  �
        �t�bhhK ��h��R�(KK��h�C@�     4   O   �
     .   �   �
  �
     �
     �
        �t�bhhK ��h��R�(KK��h�C0�     %  ,  �
     �  �
  �   �
        �t�bhhK ��h��R�(KK��h�CX      
   �
     �        #   Q           �
       �  �
     2         �t�bhhK ��h��R�(KK��h�C          k     &        �t�bhhK ��h��R�(KK��h�Ck     ~  )            �t�bhhK ��h��R�(KK��h�Ch'   �  �
                 E      s     �      �      �     �      L     �     �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C  �      �t�bhhK ��h��R�(KK��h�Cj          �t�bhhK ��h��R�(KK��h�C7     �t�bhhK ��h��R�(KK��h�Ck     ~     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CD#   Q   �     `   
   �      P
        �  �              �t�bhhK ��h��R�(KK��h�CDQ
     �  6   R
  �   �     	   5     -   �  �            �t�bhhK ��h��R�(KK
��h�C(B      -   �   �   �     �        �t�bhhK ��h��R�(KK��h�C<S
     �  U      �  �              !        �t�bhhK ��h��R�(KK��h�C�  #      �t�bhhK ��h��R�(KK��h�C]      T
     �t�bhhK ��h��R�(KK��h�CHU
    �      V
  W
  	      T   X
  Y
  \   Z
     >   [
        �t�bhhK ��h��R�(KK��h�CD   \
        ]
  ^
     x    �      Y        _
        �t�bhhK ��h��R�(KK��h�C8
  `
     a
  �  b
  �     i   
      c
        �t�bhhK ��h��R�(KK��h�Cd
       �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C]      e
     �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C!           �t�bhhK ��h��R�(KK
��h�C(`   
   #   Q   f
                 �t�bhhK ��h��R�(KK��h�C�   6  g
           �t�bhhK ��h��R�(KK��h�Ch
           �t�bhhK ��h��R�(KK��h�C�   !           �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�CH:   �  #  �        i
  	   �        �      :   �  j        �t�bhhK ��h��R�(KK��h�CD   �  j
     .   O  "      �   �  �   �   B      k
        �t�bhhK ��h��R�(KK��h�CT�   e   d   l
  	      "          �     �  
   �           �        �t�bhhK ��h��R�(KK��h�C         �   �         �t�bhhK ��h��R�(KK��h�C  �      �t�bhhK ��h��R�(KK��h�C   �    >   m
        �t�bhhK ��h��R�(KK��h�CP     ?   ;  n
        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C  �         �t�bhhK ��h��R�(KK��h�C o
     �                 �t�bhhK ��h��R�(KK��h�CT
      �  �      �     �     �  6      =         �     �        �t�bhhK ��h��R�(KK��h�Ch
   J   �   "   �  	      F      �     �     �  	      �     �  �  �  :   �  �        �t�bhhK ��h��R�(KK
��h�C(=   r     .  N   �  "   �        �t�bhhK ��h��R�(KK��h�CL
           p
     �     l   	   w   �      #   D     �         �t�bhhK ��h��R�(KK��h�C,      �   #  ?      \     �         �t�bhhK ��h��R�(KK��h�C,   5   4     r   �  �      �        �t�bhhK ��h��R�(KK��h�C#   D     �      �t�bhhK ��h��R�(KK��h�C]      q
     �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C!           �t�bhhK ��h��R�(KK��h�C#   D     �     �t�bhhK ��h��R�(KK��h�Cj          �t�bhhK ��h��R�(KK��h�CD�       �  �     t   3   0      K   R   \   �   r
        �t�bhhK ��h��R�(KK��h�CL     �      �     Y   ;  A  I      5   o        �   �         �t�bhhK ��h��R�(KK��h�CT     s
     Y      4   t
  �  a      �   �      ;      8     �         �t�bhhK ��h��R�(KK��h�C`      
   �  �     t   3   0      K   R   O         �   e   u
  v
  	   (   f        �t�bhhK ��h��R�(KK��h�CL   �      Y      w
  a   U   `  ,     �     x
  �  �  �        �t�bhhK ��h��R�(KK��h�CT      Y      "   �         D  �  �   +   	   �  �      �   Y         �t�bhhK ��h��R�(KK��h�C0;      �  �     �   e   y
     z
        �t�bhhK ��h��R�(KK��h�CP     {
         �    o        \   |
  �  }
  	   ~
     
        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�Cj             �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�
           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�  ;   	   �
           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK	��h�C$�  ;   	   �
     �
           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C �     �
     �           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�
           �t�bhhK ��h��R�(KK��h�C7     �t�bhhK ��h��R�(KK��h�C<
          �     =         �     �        �t�bhhK ��h��R�(KK��h�C         7        �t�bhhK ��h��R�(KK��h�C!           �t�bhhK ��h��R�(KK��h�Ck     ~     �t�bhhK ��h��R�(KK��h�C   �  �  �        �t�bhhK ��h��R�(KK��h�C�
     �t�bhhK ��h��R�(KK��h�C�
     �
  �
     �t�bhhK ��h��R�(KK��h�C�
  U   �
     �
     �t�bhhK ��h��R�(KK��h�Cp$  �  �  �        �
  	      �
  �
        �
        �     �       O   �    �
          �t�bhhK ��h��R�(KK��h�C    �
  �
  6   �
  �
        �t�bhhK ��h��R�(KK��h�C   �  �  �        �t�bhhK ��h��R�(KK��h�C�
  	   �
     �
     �t�bhhK ��h��R�(KK
��h�C(�
     4   �
  	   �
     �
        �t�bhhK ��h��R�(KK��h�C0�  �
     �
     �
  �  �
     �
        �t�bhhK ��h��R�(KK��h�C,$  �  �  6   �     �     �
        �t�bhhK ��h��R�(KK��h�C,�       O   �      �          �t�bhhK ��h��R�(KK��h�C  �
  �
        �t�bhhK ��h��R�(KK��h�C@�     4   O   �
     .   �   �
  �
     �
     �
        �t�bhhK ��h��R�(KK��h�C0�     %  ,  �
     �  �
  �   �
        �t�bhhK ��h��R�(KK��h�CX      
   �
     �        #   Q           �
       �  �
     2         �t�bhhK ��h��R�(KK��h�C          k     &        �t�bhhK ��h��R�(KK��h�Ck     ~  )            �t�bhhK ��h��R�(KK��h�Ch'   �  �
                 E      s     �      �      �     �      L     �     �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C  �      �t�bhhK ��h��R�(KK��h�Cj          �t�bhhK ��h��R�(KK��h�C7     �t�bhhK ��h��R�(KK��h�Ck     ~     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CD#   Q   �     `   
   �      P
        �  �              �t�bhhK ��h��R�(KK��h�CDQ
     �  6   R
  �   �     	   5     -   �  �            �t�bhhK ��h��R�(KK
��h�C(B      -   �   �   �     �        �t�bhhK ��h��R�(KK��h�C<S
     �  U      �  �              !        �t�bhhK ��h��R�(KK��h�C�  #      �t�bhhK ��h��R�(KK��h�C]      T
     �t�bhhK ��h��R�(KK��h�CHU
    �      V
  W
  	      T   X
  Y
  \   Z
     >   [
        �t�bhhK ��h��R�(KK��h�CD   \
        ]
  ^
     x    �      Y        _
        �t�bhhK ��h��R�(KK��h�C8
  `
     a
  �  b
  �     i   
      c
        �t�bhhK ��h��R�(KK��h�Cd
       �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C]      e
     �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C!           �t�bhhK ��h��R�(KK
��h�C(`   
   #   Q   f
                 �t�bhhK ��h��R�(KK��h�C�   6  g
           �t�bhhK ��h��R�(KK��h�Ch
           �t�bhhK ��h��R�(KK��h�C�   !           �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�CH:   �  #  �        i
  	   �        �      :   �  j        �t�bhhK ��h��R�(KK��h�CD   �  j
     .   O  "      �   �  �   �   B      k
        �t�bhhK ��h��R�(KK��h�CT�   e   d   l
  	      "          �     �  
   �           �        �t�bhhK ��h��R�(KK��h�C         �   �         �t�bhhK ��h��R�(KK��h�C  �      �t�bhhK ��h��R�(KK��h�C   �    >   m
        �t�bhhK ��h��R�(KK��h�CP     ?   ;  n
        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C  �         �t�bhhK ��h��R�(KK��h�C o
     �                 �t�bhhK ��h��R�(KK��h�CT
      �  �      �     �     �  6      =         �     �        �t�bhhK ��h��R�(KK��h�Ch
   J   �   "   �  	      F      �     �     �  	      �     �  �  �  :   �  �        �t�bhhK ��h��R�(KK
��h�C(=   r     .  N   �  "   �        �t�bhhK ��h��R�(KK��h�CL
           p
     �     l   	   w   �      #   D     �         �t�bhhK ��h��R�(KK��h�C,      �   #  ?      \     �         �t�bhhK ��h��R�(KK��h�C,   5   4     r   �  �      �        �t�bhhK ��h��R�(KK��h�C#   D     �      �t�bhhK ��h��R�(KK��h�C]      q
     �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C!           �t�bhhK ��h��R�(KK��h�C#   D     �     �t�bhhK ��h��R�(KK��h�Cj          �t�bhhK ��h��R�(KK��h�CD�       �  �     t   3   0      K   R   \   �   r
        �t�bhhK ��h��R�(KK��h�CL     �      �     Y   ;  A  I      5   o        �   �         �t�bhhK ��h��R�(KK��h�CT     s
     Y      4   t
  �  a      �   �      ;      8     �         �t�bhhK ��h��R�(KK��h�C`      
   �  �     t   3   0      K   R   O         �   e   u
  v
  	   (   f        �t�bhhK ��h��R�(KK��h�CL   �      Y      w
  a   U   `  ,     �     x
  �  �  �        �t�bhhK ��h��R�(KK��h�CT      Y      "   �         D  �  �   +   	   �  �      �   Y         �t�bhhK ��h��R�(KK��h�C0;      �  �     �   e   y
     z
        �t�bhhK ��h��R�(KK��h�CP     {
         �    o        \   |
  �  }
  	   ~
     
        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�Cj             �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�
           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�  ;   	   �
           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK	��h�C$�  ;   	   �
     �
           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C �     �
     �           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�
           �t�bhhK ��h��R�(KK��h�C7     �t�bhhK ��h��R�(KK��h�C<
          �     =         �     �        �t�bhhK ��h��R�(KK��h�C         7        �t�bhhK ��h��R�(KK��h�C!           �t�bhhK ��h��R�(KK��h�Ck     ~     �t�bhhK ��h��R�(KK��h�C   �  �  �        �t�bhhK ��h��R�(KK��h�C�
     �t�bhhK ��h��R�(KK��h�C�
     �
  �
     �t�bhhK ��h��R�(KK��h�C�
  U   �
     �
     �t�bhhK ��h��R�(KK��h�Cp$  �  �  �        �
  	      �
  �
        �
        �     �       O   �    �
          �t�bhhK ��h��R�(KK��h�C    �
  �
  6   �
  �
        �t�bhhK ��h��R�(KK��h�C   �  �  �        �t�bhhK ��h��R�(KK��h�C�
  	   �
     �
     �t�bhhK ��h��R�(KK
��h�C(�
     4   �
  	   �
     �
        �t�bhhK ��h��R�(KK��h�C0�  �
     �
     �
  �  �
     �
        �t�bhhK ��h��R�(KK��h�C,$  �  �  6   �     �     �
        �t�bhhK ��h��R�(KK��h�C,�       O   �      �          �t�bhhK ��h��R�(KK��h�C  �
  �
        �t�bhhK ��h��R�(KK��h�C@�     4   O   �
     .   �   �
  �
     �
     �
        �t�bhhK ��h��R�(KK��h�C0�     %  ,  �
     �  �
  �   �
        �t�bhhK ��h��R�(KK��h�CX      
   �
     �        #   Q           �
       �  �
     2         �t�bhhK ��h��R�(KK��h�C          k     &        �t�bhhK ��h��R�(KK��h�Ck     ~  )            �t�bhhK ��h��R�(KK��h�Ch'   �  �
                 E      s     �      �      �     �      L     �     �     �t�bhhK ��h��R�(KK��h�C�      �   )            �t�bhhK ��h��R�(KK��h�C0�   W  T   s      )         U   �
        �t�bhhK ��h��R�(KK0��h�C�t   3     T   �      )      t   3   	     8  �         �
     �
     &   �         �   C      .   �  D       �   )   �         '     �      �        t   3   �
        �t�bhhK ��h��R�(KK��h�C@�  �  -   �   X      �   C      t   3   	     8        �t�bhhK ��h��R�(KK��h�C<   �  	        �   )            �
     �
        �t�bhhK ��h��R�(KK��h�CD
         �
     �
  6      =   S      �        �         �t�bhhK ��h��R�(KK��h�CD      >  
      
   s      )            C   d   (        �t�bhhK ��h��R�(KK��h�C          )         �      �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�CP   3           �t�bhhK ��h��R�(KK��h�CX      �            �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�
  	        �t�bhhK ��h��R�(KK��h�C�  �
                 �t�bhhK ��h��R�(KK��h�C�      �   )            �t�bhhK ��h��R�(KK��h�C0�   W  T   s      )         U   �
        �t�bhhK ��h��R�(KK0��h�C�t   3     T   �      )      t   3   	     8  �         �
     �
     &   �         �   C      .   �  D       �   )   �         '     �      �        t   3   �
        �t�bhhK ��h��R�(KK��h�C@�  �  -   �   X      �   C      t   3   	     8        �t�bhhK ��h��R�(KK��h�C<   �  	        �   )            �
     �
        �t�bhhK ��h��R�(KK��h�CD
         �
     �
  6      =   S      �        �         �t�bhhK ��h��R�(KK��h�CD      >  
      
   s      )            C   d   (        �t�bhhK ��h��R�(KK��h�C          )         �      �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�CP   3           �t�bhhK ��h��R�(KK��h�CX      �            �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�
  	        �t�bhhK ��h��R�(KK��h�C�  �
                 �t�bhhK ��h��R�(KK��h�C�      �   )            �t�bhhK ��h��R�(KK��h�C0�   W  T   s      )         U   �
        �t�bhhK ��h��R�(KK0��h�C�t   3     T   �      )      t   3   	     8  �         �
     �
     &   �         �   C      .   �  D       �   )   �         '     �      �        t   3   �
        �t�bhhK ��h��R�(KK��h�C@�  �  -   �   X      �   C      t   3   	     8        �t�bhhK ��h��R�(KK��h�C<   �  	        �   )            �
     �
        �t�bhhK ��h��R�(KK��h�CD
         �
     �
  6      =   S      �        �         �t�bhhK ��h��R�(KK��h�CD      >  
      
   s      )            C   d   (        �t�bhhK ��h��R�(KK��h�C          )         �      �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�CP   3           �t�bhhK ��h��R�(KK��h�CX      �            �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�
  	        �t�bhhK ��h��R�(KK��h�C�  �
                 �t�bhhK ��h��R�(KK��h�Cu   7   F  �   h      �t�bhhK ��h��R�(KK��h�C    �  '   �      �t�bhhK ��h��R�(KK��h�CG     �t�bhhK ��h��R�(KK��h�C
        �     �t�bhhK ��h��R�(KK��h�Cu   7   F  �   h      �t�bhhK ��h��R�(KK��h�C,      g   )     "        �        �t�bhhK ��h��R�(KK��h�CT   "  7      �  N      e  �  �
  �
  �     *  �         �
  �
        �t�bhhK ��h��R�(KK��h�CT   Z   �        �
  J   �     �
     �     i      �     �  #        �t�bhhK ��h��R�(KK��h�CP   3   S      �     �      +     O      +          E     �        �t�bhhK ��h��R�(KK��h�C8   5   4     �   }          �   S      �         �t�bhhK ��h��R�(KK��h�Ch   �       ;              �  �              �  �
     �     �
  
   �
        �t�bhhK ��h��R�(KK��h�Cl
      5   �      }      S      �   6      =   S      �   .  �   ]      �      }               �t�bhhK ��h��R�(KK��h�CDu   -   .     �      S      �   
      �  �     b        �t�bhhK ��h��R�(KK��h�C\      �   S      �  �      5      
   S      �  ;           �              �t�bhhK ��h��R�(KK��h�C\l     S      �           )   	   �        	   �           �     E         �t�bhhK ��h��R�(KK��h�CPS      �      �  �      #   	     	   �  	   �  	   �     �        �t�bhhK ��h��R�(KK��h�C0      ,  �  ,  S      �     �        �t�bhhK ��h��R�(KK	��h�C$�     S      �      #         �t�bhhK ��h��R�(KK��h�C�   #         �t�bhhK ��h��R�(KK��h�C8   S      �  �
     �
  )  �   
      1         �t�bhhK ��h��R�(KK��h�CL   7   *  )     J   �  2      �  t  �     �
  �  �
  �        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�Cu   7   F  �   h      �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK	��h�C$�   �                       �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK��h�C3   S      �           �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK
��h�C(S      �                 E      �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK��h�C�        �
           �t�bhhK ��h��R�(KK��h�C    �  '   �      �t�bhhK ��h��R�(KK��h�C`�
     �   -       T   ;      �
  �
  ?   �  �  �
  	   U             H  �
        �t�bhhK ��h��R�(KK��h�C@�  �  x   �   e          �
     �
         i   �        �t�bhhK ��h��R�(KK��h�C�      v        �t�bhhK ��h��R�(KK��h�C<�     t   3   �
  �
  �
             �  ;         �t�bhhK ��h��R�(KK��h�CD      �   �   -    
      5      
       �  '   �         �t�bhhK ��h��R�(KK��h�C�     �  �
     �t�bhhK ��h��R�(KK��h�C�
     �t�bhhK ��h��R�(KK��h�C�
          �t�bhhK ��h��R�(KK��h�C�
     �t�bhhK ��h��R�(KK��h�C�
     �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C    �  '   �         �t�bhhK ��h��R�(KK��h�C�
  �
        �t�bhhK ��h��R�(KK��h�C�
  �
     �t�bhhK ��h��R�(KK��h�C �   -  �                 �t�bhhK ��h��R�(KK��h�CG     �t�bhhK ��h��R�(KK��h�C<
      5   '   �     �        �   �   �   !        �t�bhhK ��h��R�(KK��h�C�
  �         �t�bhhK ��h��R�(KK��h�C�  �
  	   �
  #      �t�bhhK ��h��R�(KK��h�Cc     �  i  	   #      �t�bhhK ��h��R�(KK��h�C�    �     �
     �t�bhhK ��h��R�(KK��h�C         G        �t�bhhK ��h��R�(KK��h�C
        �     �t�bhhK ��h��R�(KK��h�Ch�     �
     �
     �     �   a      "          S      �  �  �       ;   �        �t�bhhK ��h��R�(KK��h�Cl      �   S      �   
      4      �   /                
         �     �   e   #        �t�bhhK ��h��R�(KK��h�Ch      �        �
  
      5   +          �        �            
   S      �  ;         �t�bhhK ��h��R�(KK��h�CT.     �
           )   	   �        	   �           �     E         �t�bhhK ��h��R�(KK��h�CPS      �      �  �      #   	     	   �  	   �  	   �     �        �t�bhhK ��h��R�(KK��h�C0      ,  �  ,  S      �     �        �t�bhhK ��h��R�(KK��h�CS      �  �      #      �t�bhhK ��h��R�(KK��h�C         �        �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK	��h�C$�   �                       �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK��h�C3   S      �           �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK
��h�C(S      �                 E      �t�bhhK ��h��R�(KK	��h�C$�  �
  �
  �  C     .        �t�bhhK ��h��R�(KK��h�CL/  �
     �
  �
  �  	   '   �
     $     &   E   �
     �
        �t�bhhK ��h��R�(KK��h�C46  &   �
  �
  U  /      �
  �
  I   �
        �t�bhhK ��h��R�(KK��h�CH�
     �
     /     '   �  %     �     =  I       �
        �t�bhhK ��h��R�(KK��h�CL?   �
  /  �
  U     �  y     �
     �
  Y       0     �        �t�bhhK ��h��R�(KK��h�CX�  !  �
     �
     �
  	      B   �
  g      �
  �
  i  �  �
     c        �t�bhhK ��h��R�(KK��h�C0   �
         '          Y         �t�bhhK ��h��R�(KK��h�CL   .     .     �  "   B     a      �       ^      }         �t�bhhK ��h��R�(KK��h�CX   
   �  "     �     �     �          )   	      	         E         �t�bhhK ��h��R�(KK
��h�C(&       �        	  2         �t�bhhK ��h��R�(KK��h�C0&   
  �                  �        �t�bhhK ��h��R�(KK��h�CX                �          
   �      �     �    �     '        �t�bhhK ��h��R�(KK	��h�C$      
          .        �t�bhhK ��h��R�(KK��h�C�             �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C@   
             9                     E      �t�bhhK ��h��R�(KK��h�C �   -  �                 �t�bhhK ��h��R�(KK��h�C  �        �t�bhhK ��h��R�(KK��h�C.                   �t�bhhK ��h��R�(KK��h�C0   
                         E      �t�bhhK ��h��R�(KK��h�Cu   7   F  �   h      �t�bhhK ��h��R�(KK��h�C    �  '   �      �t�bhhK ��h��R�(KK��h�CG     �t�bhhK ��h��R�(KK��h�C
        �     �t�bhhK ��h��R�(KK��h�Cu   7   F  �   h      �t�bhhK ��h��R�(KK��h�C,      g   )     "        �        �t�bhhK ��h��R�(KK��h�CT   "  7      �  N      e  �  �
  �
  �     *  �         �
  �
        �t�bhhK ��h��R�(KK��h�CT   Z   �        �
  J   �     �
     �     i      �     �  #        �t�bhhK ��h��R�(KK��h�CP   3   S      �     �      +     O      +          E     �        �t�bhhK ��h��R�(KK��h�C8   5   4     �   }          �   S      �         �t�bhhK ��h��R�(KK��h�Ch   �       ;              �  �              �  �
     �     �
  
   �
        �t�bhhK ��h��R�(KK��h�Cl
      5   �      }      S      �   6      =   S      �   .  �   ]      �      }               �t�bhhK ��h��R�(KK��h�CDu   -   .     �      S      �   
      �  �     b        �t�bhhK ��h��R�(KK��h�C\      �   S      �  �      5      
   S      �  ;           �              �t�bhhK ��h��R�(KK��h�C\l     S      �           )   	   �        	   �           �     E         �t�bhhK ��h��R�(KK��h�CPS      �      �  �      #   	     	   �  	   �  	   �     �        �t�bhhK ��h��R�(KK��h�C0      ,  �  ,  S      �     �        �t�bhhK ��h��R�(KK	��h�C$�     S      �      #         �t�bhhK ��h��R�(KK��h�C�   #         �t�bhhK ��h��R�(KK��h�C8   S      �  �
     �
  )  �   
      1         �t�bhhK ��h��R�(KK��h�CL   7   *  )     J   �  2      �  t  �     �
  �  �
  �        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�Cu   7   F  �   h      �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK	��h�C$�   �                       �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK��h�C3   S      �           �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK
��h�C(S      �                 E      �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK��h�C�        �
           �t�bhhK ��h��R�(KK��h�C    �  '   �      �t�bhhK ��h��R�(KK��h�C`�
     �   -       T   ;      �
  �
  ?   �  �  �
  	   U             H  �
        �t�bhhK ��h��R�(KK��h�C@�  �  x   �   e          �
     �
         i   �        �t�bhhK ��h��R�(KK��h�C�      v        �t�bhhK ��h��R�(KK��h�C<�     t   3   �
  �
  �
             �  ;         �t�bhhK ��h��R�(KK��h�CD      �   �   -    
      5      
       �  '   �         �t�bhhK ��h��R�(KK��h�C�     �  �
     �t�bhhK ��h��R�(KK��h�C�
     �t�bhhK ��h��R�(KK��h�C�
          �t�bhhK ��h��R�(KK��h�C�
     �t�bhhK ��h��R�(KK��h�C�
     �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C    �  '   �         �t�bhhK ��h��R�(KK��h�C�
  �
        �t�bhhK ��h��R�(KK��h�C�
  �
     �t�bhhK ��h��R�(KK��h�C �   -  �                 �t�bhhK ��h��R�(KK��h�CG     �t�bhhK ��h��R�(KK��h�C<
      5   '   �     �        �   �   �   !        �t�bhhK ��h��R�(KK��h�C�
  �         �t�bhhK ��h��R�(KK��h�C�  �
  	   �
  #      �t�bhhK ��h��R�(KK��h�Cc     �  i  	   #      �t�bhhK ��h��R�(KK��h�C�    �     �
     �t�bhhK ��h��R�(KK��h�C         G        �t�bhhK ��h��R�(KK��h�C
        �     �t�bhhK ��h��R�(KK��h�Ch�     �
     �
     �     �   a      "          S      �  �  �       ;   �        �t�bhhK ��h��R�(KK��h�Cl      �   S      �   
      4      �   /                
         �     �   e   #        �t�bhhK ��h��R�(KK��h�Ch      �        �
  
      5   +          �        �            
   S      �  ;         �t�bhhK ��h��R�(KK��h�CT.     �
           )   	   �        	   �           �     E         �t�bhhK ��h��R�(KK��h�CPS      �      �  �      #   	     	   �  	   �  	   �     �        �t�bhhK ��h��R�(KK��h�C0      ,  �  ,  S      �     �        �t�bhhK ��h��R�(KK��h�CS      �  �      #      �t�bhhK ��h��R�(KK��h�C         �        �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK	��h�C$�   �                       �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK��h�C3   S      �           �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK
��h�C(S      �                 E      �t�bhhK ��h��R�(KK	��h�C$�  �
  �
  �  C     .        �t�bhhK ��h��R�(KK��h�CL/  �
     �
  �
  �  	   '   �
     $     &   E   �
     �
        �t�bhhK ��h��R�(KK��h�C46  &   �
  �
  U  /      �
  �
  I   �
        �t�bhhK ��h��R�(KK��h�CH�
     �
     /     '   �  %     �     =  I       �
        �t�bhhK ��h��R�(KK��h�CL?   �
  /  �
  U     �  y     �
     �
  Y       0     �        �t�bhhK ��h��R�(KK��h�CX�  !  �
     �
     �
  	      B   �
  g      �
  �
  i  �  �
     c        �t�bhhK ��h��R�(KK��h�C0   �
         '          Y         �t�bhhK ��h��R�(KK��h�CL   .     .     �  "   B     a      �       ^      }         �t�bhhK ��h��R�(KK��h�CX   
   �  "     �     �     �          )   	      	         E         �t�bhhK ��h��R�(KK
��h�C(&       �        	  2         �t�bhhK ��h��R�(KK��h�C0&   
  �                  �        �t�bhhK ��h��R�(KK��h�CX                �          
   �      �     �    �     '        �t�bhhK ��h��R�(KK	��h�C$      
          .        �t�bhhK ��h��R�(KK��h�C�             �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C@   
             9                     E      �t�bhhK ��h��R�(KK��h�C �   -  �                 �t�bhhK ��h��R�(KK��h�C  �        �t�bhhK ��h��R�(KK��h�C.                   �t�bhhK ��h��R�(KK��h�C0   
                         E      �t�bhhK ��h��R�(KK��h�Cu   7   F  �   h      �t�bhhK ��h��R�(KK��h�C    �  '   �      �t�bhhK ��h��R�(KK��h�CG     �t�bhhK ��h��R�(KK��h�C
        �     �t�bhhK ��h��R�(KK��h�Cu   7   F  �   h      �t�bhhK ��h��R�(KK��h�C,      g   )     "        �        �t�bhhK ��h��R�(KK��h�CT   "  7      �  N      e  �  �
  �
  �     *  �         �
  �
        �t�bhhK ��h��R�(KK��h�CT   Z   �        �
  J   �     �
     �     i      �     �  #        �t�bhhK ��h��R�(KK��h�CP   3   S      �     �      +     O      +          E     �        �t�bhhK ��h��R�(KK��h�C8   5   4     �   }          �   S      �         �t�bhhK ��h��R�(KK��h�Ch   �       ;              �  �              �  �
     �     �
  
   �
        �t�bhhK ��h��R�(KK��h�Cl
      5   �      }      S      �   6      =   S      �   .  �   ]      �      }               �t�bhhK ��h��R�(KK��h�CDu   -   .     �      S      �   
      �  �     b        �t�bhhK ��h��R�(KK��h�C\      �   S      �  �      5      
   S      �  ;           �              �t�bhhK ��h��R�(KK��h�C\l     S      �           )   	   �        	   �           �     E         �t�bhhK ��h��R�(KK��h�CPS      �      �  �      #   	     	   �  	   �  	   �     �        �t�bhhK ��h��R�(KK��h�C0      ,  �  ,  S      �     �        �t�bhhK ��h��R�(KK	��h�C$�     S      �      #         �t�bhhK ��h��R�(KK��h�C�   #         �t�bhhK ��h��R�(KK��h�C8   S      �  �
     �
  )  �   
      1         �t�bhhK ��h��R�(KK��h�CL   7   *  )     J   �  2      �  t  �     �
  �  �
  �        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�Cu   7   F  �   h      �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK	��h�C$�   �                       �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK��h�C3   S      �           �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK
��h�C(S      �                 E      �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK��h�C�        �
           �t�bhhK ��h��R�(KK��h�C    �  '   �      �t�bhhK ��h��R�(KK��h�C`�
     �   -       T   ;      �
  �
  ?   �  �  �
  	   U             H  �
        �t�bhhK ��h��R�(KK��h�C@�  �  x   �   e          �
     �
         i   �        �t�bhhK ��h��R�(KK��h�C�      v        �t�bhhK ��h��R�(KK��h�C<�     t   3   �
  �
  �
             �  ;         �t�bhhK ��h��R�(KK��h�CD      �   �   -    
      5      
       �  '   �         �t�bhhK ��h��R�(KK��h�C�     �  �
     �t�bhhK ��h��R�(KK��h�C�
     �t�bhhK ��h��R�(KK��h�C�
          �t�bhhK ��h��R�(KK��h�C�
     �t�bhhK ��h��R�(KK��h�C�
     �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C    �  '   �         �t�bhhK ��h��R�(KK��h�C�
  �
        �t�bhhK ��h��R�(KK��h�C�
  �
     �t�bhhK ��h��R�(KK��h�C �   -  �                 �t�bhhK ��h��R�(KK��h�CG     �t�bhhK ��h��R�(KK��h�C<
      5   '   �     �        �   �   �   !        �t�bhhK ��h��R�(KK��h�C�
  �         �t�bhhK ��h��R�(KK��h�C�  �
  	   �
  #      �t�bhhK ��h��R�(KK��h�Cc     �  i  	   #      �t�bhhK ��h��R�(KK��h�C�    �     �
     �t�bhhK ��h��R�(KK��h�C         G        �t�bhhK ��h��R�(KK��h�C
        �     �t�bhhK ��h��R�(KK��h�Ch�     �
     �
     �     �   a      "          S      �  �  �       ;   �        �t�bhhK ��h��R�(KK��h�Cl      �   S      �   
      4      �   /                
         �     �   e   #        �t�bhhK ��h��R�(KK��h�Ch      �        �
  
      5   +          �        �            
   S      �  ;         �t�bhhK ��h��R�(KK��h�CT.     �
           )   	   �        	   �           �     E         �t�bhhK ��h��R�(KK��h�CPS      �      �  �      #   	     	   �  	   �  	   �     �        �t�bhhK ��h��R�(KK��h�C0      ,  �  ,  S      �     �        �t�bhhK ��h��R�(KK��h�CS      �  �      #      �t�bhhK ��h��R�(KK��h�C         �        �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK	��h�C$�   �                       �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK��h�C3   S      �           �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK
��h�C(S      �                 E      �t�bhhK ��h��R�(KK	��h�C$�  �
  �
  �  C     .        �t�bhhK ��h��R�(KK��h�CL/  �
     �
  �
  �  	   '   �
     $     &   E   �
     �
        �t�bhhK ��h��R�(KK��h�C46  &   �
  �
  U  /      �
  �
  I   �
        �t�bhhK ��h��R�(KK��h�CH�
     �
     /     '   �  %     �     =  I       �
        �t�bhhK ��h��R�(KK��h�CL?   �
  /  �
  U     �  y     �
     �
  Y       0     �        �t�bhhK ��h��R�(KK��h�CX�  !  �
     �
     �
  	      B   �
  g      �
  �
  i  �  �
     c        �t�bhhK ��h��R�(KK��h�C0   �
         '          Y         �t�bhhK ��h��R�(KK��h�CL   .     .     �  "   B     a      �       ^      }         �t�bhhK ��h��R�(KK��h�CX   
   �  "     �     �     �          )   	      	         E         �t�bhhK ��h��R�(KK
��h�C(&       �        	  2         �t�bhhK ��h��R�(KK��h�C0&   
  �                  �        �t�bhhK ��h��R�(KK��h�CX                �          
   �      �     �    �     '        �t�bhhK ��h��R�(KK	��h�C$      
          .        �t�bhhK ��h��R�(KK��h�C�             �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C@   
             9                     E      �t�bhhK ��h��R�(KK��h�C �   -  �                 �t�bhhK ��h��R�(KK��h�C  �        �t�bhhK ��h��R�(KK��h�C.                   �t�bhhK ��h��R�(KK��h�C0   
                         E      �t�bhhK ��h��R�(KK��h�Cc      $     C      �t�bhhK ��h��R�(KK��h�C�   �      �     �t�bhhK ��h��R�(KK��h�C5         �   h      �t�bhhK ��h��R�(KK��h�Cc      $     C      �t�bhhK ��h��R�(KK"��h�C��           1         �   /      S      �     �           ;      x   /       �   /        1      E     �        �t�bhhK ��h��R�(KK��h�C ;   .  N     C            �t�bhhK ��h��R�(KK��h�C     c      C      �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C3   S      �     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C<#   �      �   �    (         .   �          �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK��h�C�   �                 �t�bhhK ��h��R�(KK��h�C�      w        �t�bhhK ��h��R�(KK��h�Cl�  ~     �                 E      s     �      �      /     v     �     �     �      �t�bhhK ��h��R�(KK��h�CU  �      �   i        �t�bhhK ��h��R�(KK��h�C4#   �      �   �                    E      �t�bhhK ��h��R�(KK��h�C�   �      �     �t�bhhK ��h��R�(KK��h�CH   �   �      �       /      �           
      !        �t�bhhK ��h��R�(KK��h�C<1             �   �      �     /      (        �t�bhhK ��h��R�(KK��h�C@      �      
   �     )     (     S      �         �t�bhhK ��h��R�(KK��h�C(     �t�bhhK ��h��R�(KK��h�C�  �       �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C5         �   h      �t�bhhK ��h��R�(KK)��h�C�
      �   9  �      �  {  	   5  4      )            .   4        �   e   k      �            	            �  �  �  �      "        �t�bhhK ��h��R�(KK��h�C<      
         %  #         5      �         �t�bhhK ��h��R�(KK��h�C<   �  �     .   �     /       �   /      �         �t�bhhK ��h��R�(KK��h�CH      �     N      %  �  
      �  �         %        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C5         �   h      �t�bhhK ��h��R�(KK��h�Cc      $     C      �t�bhhK ��h��R�(KK��h�C�   �      �     �t�bhhK ��h��R�(KK��h�C5         �   h      �t�bhhK ��h��R�(KK��h�Cc      $     C      �t�bhhK ��h��R�(KK"��h�C��           1         �   /      S      �     �           ;      x   /       �   /        1      E     �        �t�bhhK ��h��R�(KK��h�C ;   .  N     C            �t�bhhK ��h��R�(KK��h�C     c      C      �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C3   S      �     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C<#   �      �   �    (         .   �          �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK��h�C�   �                 �t�bhhK ��h��R�(KK��h�C�      w        �t�bhhK ��h��R�(KK��h�Cl�  ~     �                 E      s     �      �      /     v     �     �     �      �t�bhhK ��h��R�(KK��h�CU  �      �   i        �t�bhhK ��h��R�(KK��h�C4#   �      �   �                    E      �t�bhhK ��h��R�(KK��h�C�   �      �     �t�bhhK ��h��R�(KK��h�CH   �   �      �       /      �           
      !        �t�bhhK ��h��R�(KK��h�C<1             �   �      �     /      (        �t�bhhK ��h��R�(KK��h�C@      �      
   �     )     (     S      �         �t�bhhK ��h��R�(KK��h�C(     �t�bhhK ��h��R�(KK��h�C�  �       �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C5         �   h      �t�bhhK ��h��R�(KK)��h�C�
      �   9  �      �  {  	   5  4      )            .   4        �   e   k      �            	            �  �  �  �      "        �t�bhhK ��h��R�(KK��h�C<      
         %  #         5      �         �t�bhhK ��h��R�(KK��h�C<   �  �     .   �     /       �   /      �         �t�bhhK ��h��R�(KK��h�CH      �     N      %  �  
      �  �         %        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C5         �   h      �t�bhhK ��h��R�(KK��h�Cc      $     C      �t�bhhK ��h��R�(KK��h�C�   �      �     �t�bhhK ��h��R�(KK��h�C5         �   h      �t�bhhK ��h��R�(KK��h�Cc      $     C      �t�bhhK ��h��R�(KK"��h�C��           1         �   /      S      �     �           ;      x   /       �   /        1      E     �        �t�bhhK ��h��R�(KK��h�C ;   .  N     C            �t�bhhK ��h��R�(KK��h�C     c      C      �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C3   S      �     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C<#   �      �   �    (         .   �          �t�bhhK ��h��R�(KK��h�C�        ;         �t�bhhK ��h��R�(KK��h�C�   �                 �t�bhhK ��h��R�(KK��h�C�      w        �t�bhhK ��h��R�(KK��h�Cl�  ~     �                 E      s     �      �      /     v     �     �     �      �t�bhhK ��h��R�(KK��h�CU  �      �   i        �t�bhhK ��h��R�(KK��h�C4#   �      �   �                    E      �t�bhhK ��h��R�(KK��h�C�   �      �     �t�bhhK ��h��R�(KK��h�CH   �   �      �       /      �           
      !        �t�bhhK ��h��R�(KK��h�C<1             �   �      �     /      (        �t�bhhK ��h��R�(KK��h�C@      �      
   �     )     (     S      �         �t�bhhK ��h��R�(KK��h�C(     �t�bhhK ��h��R�(KK��h�C�  �       �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C5         �   h      �t�bhhK ��h��R�(KK)��h�C�
      �   9  �      �  {  	   5  4      )            .   4        �   e   k      �            	            �  �  �  �      "        �t�bhhK ��h��R�(KK��h�C<      
         %  #         5      �         �t�b�      hhK ��h��R�(KK��h�C<   �  �     .   �     /       �   /      �         �t�bhhK ��h��R�(KK��h�CH      �     N      %  �  
      �  �         %        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C5         �   h      �t�bhhK ��h��R�(KK��h�C     |      �t�bhhK ��h��R�(KK��h�C4
      �   �     1   5      �  '   {         �t�bhhK ��h��R�(KK��h�C,$  �     �   %          �        �t�bhhK ��h��R�(KK��h�C          �     1         �t�bhhK ��h��R�(KK��h�CH�           #      �     6      I  /      |      ]        �t�bhhK ��h��R�(KK��h�C<      1  I  /      #   2     &     �   1         �t�bhhK ��h��R�(KK��h�C�      �   1      �t�bhhK ��h��R�(KK��h�C#   �     �t�bhhK ��h��R�(KK��h�C�  i     �t�bhhK ��h��R�(KK��h�Ck  #      �t�bhhK ��h��R�(KK��h�C]      l     �t�bhhK ��h��R�(KK��h�C,N      �     �   6      w      /      �t�bhhK ��h��R�(KK��h�C4{      *     
      5   '   {      1         �t�bhhK ��h��R�(KK��h�C@+  ;  ,     m     �     
         m     �        �t�bhhK ��h��R�(KK��h�C'     �t�bhhK ��h��R�(KK��h�C-       $      �t�bhhK ��h��R�(KK��h�Cd3        �     (     U     6   �  .        )  \        )   	                  �t�bhhK ��h��R�(KK��h�CL      
   *     �  O      d   �      d   r   +  ,     1         �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C     |         �t�bhhK ��h��R�(KK��h�C	  �                  �t�bhhK ��h��R�(KK��h�C4  {      �t�bhhK ��h��R�(KK��h�C8   6   i   
   4  {     r      {   �  �         �t�bhhK ��h��R�(KK	��h�C$   �   
   -     �  .        �t�bhhK ��h��R�(KK��h�C,      x  i   
   4  {      1         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CF  G     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C         4  {         �t�bhhK ��h��R�(KK��h�C     |      �t�bhhK ��h��R�(KK��h�C4
      �   �     1   5      �  '   {         �t�bhhK ��h��R�(KK��h�C,$  �     �   %          �        �t�bhhK ��h��R�(KK��h�C          �     1         �t�bhhK ��h��R�(KK��h�CH�           #      �     6      I  /      |      ]        �t�bhhK ��h��R�(KK��h�C<      1  I  /      #   2     &     �   1         �t�bhhK ��h��R�(KK��h�C�      �   1      �t�bhhK ��h��R�(KK��h�C#   �     �t�bhhK ��h��R�(KK��h�C�  i     �t�bhhK ��h��R�(KK��h�Ck  #      �t�bhhK ��h��R�(KK��h�C]      l     �t�bhhK ��h��R�(KK��h�C,N      �     �   6      w      /      �t�bhhK ��h��R�(KK��h�C4{      *     
      5   '   {      1         �t�bhhK ��h��R�(KK��h�C@+  ;  ,     m     �     
         m     �        �t�bhhK ��h��R�(KK��h�C'     �t�bhhK ��h��R�(KK��h�C-       $      �t�bhhK ��h��R�(KK��h�Cd3        �     (     U     6   �  .        )  \        )   	                  �t�bhhK ��h��R�(KK��h�CL      
   *     �  O      d   �      d   r   +  ,     1         �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C     |         �t�bhhK ��h��R�(KK��h�C	  �                  �t�bhhK ��h��R�(KK��h�C4  {      �t�bhhK ��h��R�(KK��h�C8   6   i   
   4  {     r      {   �  �         �t�bhhK ��h��R�(KK	��h�C$   �   
   -     �  .        �t�bhhK ��h��R�(KK��h�C,      x  i   
   4  {      1         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CF  G     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C         4  {         �t�bhhK ��h��R�(KK��h�C     |      �t�bhhK ��h��R�(KK��h�C4
      �   �     1   5      �  '   {         �t�bhhK ��h��R�(KK��h�C,$  �     �   %          �        �t�bhhK ��h��R�(KK��h�C          �     1         �t�bhhK ��h��R�(KK��h�CH�           #      �     6      I  /      |      ]        �t�bhhK ��h��R�(KK��h�C<      1  I  /      #   2     &     �   1         �t�bhhK ��h��R�(KK��h�C�      �   1      �t�bhhK ��h��R�(KK��h�C#   �     �t�bhhK ��h��R�(KK��h�C�  i     �t�bhhK ��h��R�(KK��h�Ck  #      �t�bhhK ��h��R�(KK��h�C]      l     �t�bhhK ��h��R�(KK��h�C,N      �     �   6      w      /      �t�bhhK ��h��R�(KK��h�C4{      *     
      5   '   {      1         �t�bhhK ��h��R�(KK��h�C@+  ;  ,     m     �     
         m     �        �t�bhhK ��h��R�(KK��h�C'     �t�bhhK ��h��R�(KK��h�C-       $      �t�bhhK ��h��R�(KK��h�Cd3        �     (     U     6   �  .        )  \        )   	                  �t�bhhK ��h��R�(KK��h�CL      
   *     �  O      d   �      d   r   +  ,     1         �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C     |         �t�bhhK ��h��R�(KK��h�C	  �                  �t�bhhK ��h��R�(KK��h�C4  {      �t�bhhK ��h��R�(KK��h�C8   6   i   
   4  {     r      {   �  �         �t�bhhK ��h��R�(KK	��h�C$   �   
   -     �  .        �t�bhhK ��h��R�(KK��h�C,      x  i   
   4  {      1         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CF  G     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C         4  {         �t�bhhK ��h��R�(KK��h�C �  /     0     
        �t�bhhK ��h��R�(KK��h�CX         u   �    �      w  	   /     5  	     	        0        �t�bhhK ��h��R�(KK��h�C �  1     2     3        �t�bhhK ��h��R�(KK��h�C|&      1      �     1      +        7        
       4  	   �  	   0     �      1      Z   >   k         �t�bhhK ��h��R�(KK��h�C
     �t�bhhK ��h��R�(KK��h�C�      w     �t�bhhK ��h��R�(KK��h�CH�      w       5     �      �          C      1         �t�bhhK ��h��R�(KK��h�CL6     $     C   (  �      7       C   8  	   9             �t�bhhK ��h��R�(KK��h�C�      w        �t�bhhK ��h��R�(KK��h�C $     �                  �t�bhhK ��h��R�(KK��h�C/     5     �t�bhhK ��h��R�(KK��h�C\/     5       �        .   ~    �   :  	   ;  	   �  	   <     =        �t�bhhK ��h��R�(KK��h�C>     5        �t�bhhK ��h��R�(KK��h�C6                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C?        �t�bhhK ��h��R�(KK��h�C6                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C@  2  @     >   A     3     #     �     1         �t�bhhK ��h��R�(KK��h�CP2  B        Y      �     1      C        D     E     1         �t�bhhK ��h��R�(KK��h�CD     0  T         4         �  �  1      9         �t�bhhK ��h��R�(KK
��h�C(F        U   �                 �t�bhhK ��h��R�(KK��h�C0     �t�bhhK ��h��R�(KK��h�C5        �t�bhhK ��h��R�(KK��h�C6                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C9         �t�bhhK ��h��R�(KK��h�CG     H  �        �t�bhhK ��h��R�(KK��h�C6              I     �t�bhhK ��h��R�(KK��h�Cj   7     �t�bhhK ��h��R�(KK��h�Cxj     "   J  '   7       B   K  
   L          M       �                               �t�bhhK ��h��R�(KK ��h�C�  �    N     C      Y      1      �     1         {  �   O     '   �     D   (  �                   �t�bhhK ��h��R�(KK��h�Cp.               '   P  �  E  Q     
   $     C      
       �     1      '   x  	   R        �t�bhhK ��h��R�(KK��h�C S  =       q   ?        �t�bhhK ��h��R�(KK��h�Ct:   �   �   T  j     U  	   i      .      c       6     W   �        a      q   D      V        �t�bhhK ��h��R�(KK	��h�C$W  X  Y  2  U   �  |         �t�bhhK ��h��R�(KK
��h�C(     8  6  y        Z        �t�bhhK ��h��R�(KK��h�CL  [           \  &   ]  9     C        a      j   7        �t�bhhK ��h��R�(KK��h�C|�     
   �  B   ^  a      8  p   j   _  `  a     b  	   c     d     e     f     g  	   (   h        �t�bhhK ��h��R�(KK��h�C �  /     0     
        �t�bhhK ��h��R�(KK��h�CX         u   �    �      w  	   /     5  	     	        0        �t�bhhK ��h��R�(KK��h�C �  1     2     3        �t�bhhK ��h��R�(KK��h�C|&      1      �     1      +        7        
       4  	   �  	   0     �      1      Z   >   k         �t�bhhK ��h��R�(KK��h�C
     �t�bhhK ��h��R�(KK��h�C�      w     �t�bhhK ��h��R�(KK��h�CH�      w       5     �      �          C      1         �t�bhhK ��h��R�(KK��h�CL6     $     C   (  �      7       C   8  	   9             �t�bhhK ��h��R�(KK��h�C�      w        �t�bhhK ��h��R�(KK��h�C $     �                  �t�bhhK ��h��R�(KK��h�C/     5     �t�bhhK ��h��R�(KK��h�C\/     5       �        .   ~    �   :  	   ;  	   �  	   <     =        �t�bhhK ��h��R�(KK��h�C>     5        �t�bhhK ��h��R�(KK��h�C6                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C?        �t�bhhK ��h��R�(KK��h�C6                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C@  2  @     >   A     3     #     �     1         �t�bhhK ��h��R�(KK��h�CP2  B        Y      �     1      C        D     E     1         �t�bhhK ��h��R�(KK��h�CD     0  T         4         �  �  1      9         �t�bhhK ��h��R�(KK
��h�C(F        U   �                 �t�bhhK ��h��R�(KK��h�C0     �t�bhhK ��h��R�(KK��h�C5        �t�bhhK ��h��R�(KK��h�C6                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C9         �t�bhhK ��h��R�(KK��h�CG     H  �        �t�bhhK ��h��R�(KK��h�C6              I     �t�bhhK ��h��R�(KK��h�Cj   7     �t�bhhK ��h��R�(KK��h�Cxj     "   J  '   7       B   K  
   L          M       �                               �t�bhhK ��h��R�(KK ��h�C�  �    N     C      Y      1      �     1         {  �   O     '   �     D   (  �                   �t�bhhK ��h��R�(KK��h�Cp.               '   P  �  E  Q     
   $     C      
       �     1      '   x  	   R        �t�bhhK ��h��R�(KK��h�C S  =       q   ?        �t�bhhK ��h��R�(KK��h�Ct:   �   �   T  j     U  	   i      .      c       6     W   �        a      q   D      V        �t�bhhK ��h��R�(KK	��h�C$W  X  Y  2  U   �  |         �t�bhhK ��h��R�(KK
��h�C(     8  6  y        Z        �t�bhhK ��h��R�(KK��h�CL  [           \  &   ]  9     C        a      j   7        �t�bhhK ��h��R�(KK��h�C|�     
   �  B   ^  a      8  p   j   _  `  a     b  	   c     d     e     f     g  	   (   h        �t�bhhK ��h��R�(KK��h�C �  /     0     
        �t�bhhK ��h��R�(KK��h�CX         u   �    �      w  	   /     5  	     	        0        �t�bhhK ��h��R�(KK��h�C �  1     2     3        �t�bhhK ��h��R�(KK��h�C|&      1      �     1      +        7        
       4  	   �  	   0     �      1      Z   >   k         �t�bhhK ��h��R�(KK��h�C
     �t�bhhK ��h��R�(KK��h�C�      w     �t�bhhK ��h��R�(KK��h�CH�      w       5     �      �          C      1         �t�bhhK ��h��R�(KK��h�CL6     $     C   (  �      7       C   8  	   9             �t�bhhK ��h��R�(KK��h�C�      w        �t�bhhK ��h��R�(KK��h�C $     �                  �t�bhhK ��h��R�(KK��h�C/     5     �t�bhhK ��h��R�(KK��h�C\/     5       �        .   ~    �   :  	   ;  	   �  	   <     =        �t�bhhK ��h��R�(KK��h�C>     5        �t�bhhK ��h��R�(KK��h�C6                 �t�be(hhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C?        �t�bhhK ��h��R�(KK��h�C6                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C@  2  @     >   A     3     #     �     1         �t�bhhK ��h��R�(KK��h�CP2  B        Y      �     1      C        D     E     1         �t�bhhK ��h��R�(KK��h�CD     0  T         4         �  �  1      9         �t�bhhK ��h��R�(KK
��h�C(F        U   �                 �t�bhhK ��h��R�(KK��h�C0     �t�bhhK ��h��R�(KK��h�C5        �t�bhhK ��h��R�(KK��h�C6                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C9         �t�bhhK ��h��R�(KK��h�CG     H  �        �t�bhhK ��h��R�(KK��h�C6              I     �t�bhhK ��h��R�(KK��h�Cj   7     �t�bhhK ��h��R�(KK��h�Cxj     "   J  '   7       B   K  
   L          M       �                               �t�bhhK ��h��R�(KK ��h�C�  �    N     C      Y      1      �     1         {  �   O     '   �     D   (  �                   �t�bhhK ��h��R�(KK��h�Cp.               '   P  �  E  Q     
   $     C      
       �     1      '   x  	   R        �t�bhhK ��h��R�(KK��h�C S  =       q   ?        �t�bhhK ��h��R�(KK��h�Ct:   �   �   T  j     U  	   i      .      c       6     W   �        a      q   D      V        �t�bhhK ��h��R�(KK	��h�C$W  X  Y  2  U   �  |         �t�bhhK ��h��R�(KK
��h�C(     8  6  y        Z        �t�bhhK ��h��R�(KK��h�CL  [           \  &   ]  9     C        a      j   7        �t�bhhK ��h��R�(KK��h�C|�     
   �  B   ^  a      8  p   j   _  `  a     b  	   c     d     e     f     g  	   (   h        �t�bhhK ��h��R�(KK��h�C\   i          j   2         k      ,            :  j  k  ;  <        �t�bhhK ��h��R�(KK��h�C   "   >            �t�bhhK ��h��R�(KK��h�C,l  �   m     n    o  p     �     �t�bhhK ��h��R�(KK��h�CLq  �   r  	   s  	      &  ^             t  	   -   u        �t�bhhK ��h��R�(KK��h�C   y  v        �t�bhhK ��h��R�(KK��h�C0;          �     �   w  x  �        �t�bhhK ��h��R�(KK��h�C8          =  �     y  :  z    <        �t�bhhK ��h��R�(KK��h�C  
   {     |        �t�bhhK ��h��R�(KK��h�Ct   5   �   i          }  ~  	      4      '   �     p               �    /      r   �        �t�bhhK ��h��R�(KK��h�Ch�      �     O   4   �  �       �  �     �  �  W   U       �  �      :  �        �t�bhhK ��h��R�(KK��h�Cx;  <  �                 E      �      /     v     �     �     �      }     �     �     �     �t�bhhK ��h��R�(KK��h�C4   �     �     �     �     �          �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C<7  T   �  �     �  M   '   �                    �t�bhhK ��h��R�(KK��h�CH   +      �        �  j   �     W   �     8  >   �        �t�bhhK ��h��R�(KK��h�C   
   �           �t�bhhK ��h��R�(KK��h�C�   �     �t�bhhK ��h��R�(KK��h�C\   i          j   2         k      ,            :  j  k  ;  <        �t�bhhK ��h��R�(KK��h�C   "   >            �t�bhhK ��h��R�(KK��h�C,l  �   m     n    o  p     �     �t�bhhK ��h��R�(KK��h�CLq  �   r  	   s  	      &  ^             t  	   -   u        �t�bhhK ��h��R�(KK��h�C   y  v        �t�bhhK ��h��R�(KK��h�C0;          �     �   w  x  �        �t�bhhK ��h��R�(KK��h�C8          =  �     y  :  z    <        �t�bhhK ��h��R�(KK��h�C  
   {     |        �t�bhhK ��h��R�(KK��h�Ct   5   �   i          }  ~  	      4      '   �     p               �    /      r   �        �t�bhhK ��h��R�(KK��h�Ch�      �     O   4   �  �       �  �     �  �  W   U       �  �      :  �        �t�bhhK ��h��R�(KK��h�Cx;  <  �                 E      �      /     v     �     �     �      }     �     �     �     �t�bhhK ��h��R�(KK��h�C4   �     �     �     �     �          �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C<7  T   �  �     �  M   '   �                    �t�bhhK ��h��R�(KK��h�CH   +      �        �  j   �     W   �     8  >   �        �t�bhhK ��h��R�(KK��h�C   
   �           �t�bhhK ��h��R�(KK��h�C�   �     �t�bhhK ��h��R�(KK	��h�C$      �     �     W        �t�bhhK ��h��R�(KK
��h�C(�        �        y  ;         �t�bhhK ��h��R�(KK��h�C�      w        �t�bhhK ��h��R�(KK"��h�C��  ~     1      �  	      �     )                  E      s     �      �      /     v     �     �     �      �t�bhhK ��h��R�(KK��h�C\   i          j   2         k      ,            :  j  k  ;  <        �t�bhhK ��h��R�(KK��h�C   "   >            �t�bhhK ��h��R�(KK��h�C,l  �   m     n    o  p     �     �t�bhhK ��h��R�(KK��h�CLq  �   r  	   s  	      &  ^             t  	   -   u        �t�bhhK ��h��R�(KK��h�C   y  v        �t�bhhK ��h��R�(KK��h�C0;          �     �   w  x  �        �t�bhhK ��h��R�(KK��h�C8          =  �     y  :  z    <        �t�bhhK ��h��R�(KK��h�C  
   {     |        �t�bhhK ��h��R�(KK��h�Ct   5   �   i          }  ~  	      4      '   �     p               �    /      r   �        �t�bhhK ��h��R�(KK��h�Ch�      �     O   4   �  �       �  �     �  �  W   U       �  �      :  �        �t�bhhK ��h��R�(KK��h�Cx;  <  �                 E      �      /     v     �     �     �      }     �     �     �     �t�bhhK ��h��R�(KK��h�C4   �     �     �     �     �          �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C<7  T   �  �     �  M   '   �                    �t�bhhK ��h��R�(KK��h�CH   +      �        �  j   �     W   �     8  >   �        �t�bhhK ��h��R�(KK��h�C   
   �           �t�bhhK ��h��R�(KK��h�C�   �     �t�bhhK ��h��R�(KK	��h�C$      �     �     W        �t�bhhK ��h��R�(KK
��h�C(�        �        y  ;         �t�bhhK ��h��R�(KK��h�C�      w        �t�bhhK ��h��R�(KK"��h�C��  ~     1      �  	      �     )                  E      s     �      �      /     v     �     �     �      �t�bhhK ��h��R�(KK��h�C0   "   %  �   
         :              �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C�        )         �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C�        )         �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C�        )         �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�   "   R          �t�bhhK ��h��R�(KK��h�C4   8         �        �      Z   >        �t�bhhK ��h��R�(KK��h�C,      g      
   �     q   !        �t�bhhK ��h��R�(KK��h�C<q   p   /   "     >     U   '   x     '   e         �t�bhhK ��h��R�(KK��h�C ?                 E      �t�bhhK ��h��R�(KK��h�C,�   J        �     9     &        �t�bhhK ��h��R�(KK
��h�C(   :  �      �   @     �        �t�bhhK ��h��R�(KK	��h�C$      �   ;     8   A        �t�bhhK ��h��R�(KK��h�C@      -   �      B     <        C        �        �t�bhhK ��h��R�(KK��h�CD     �t�bhhK ��h��R�(KK��h�C=  =     �t�bhhK ��h��R�(KK��h�CTC       y      u     �  �  �  	   �  	   #  -   y      �     �     �t�bhhK ��h��R�(KK
��h�C(&   |  �     9      !   >        �t�bhhK ��h��R�(KK
��h�C($                 E      �     �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C	     1         �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C    8   E  �      �        �t�bhhK ��h��R�(KK��h�C0   �  F  K  G     H  >   �  {        �t�bhhK ��h��R�(KK	��h�C$I  �  u   �  I   2  �        �t�bhhK ��h��R�(KK��h�C0   8   Q   2           %     �        �t�bhhK ��h��R�(KK��h�CH      D   �   �     &  �   \   �  �      )                  �t�bhhK ��h��R�(KK��h�C-   �  �   �        �t�bhhK ��h��R�(KK��h�C�      J           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C,Z     S     ?     *      9         �t�bhhK ��h��R�(KK��h�C@   q   �  �        g      6  .     K     L        �t�bhhK ��h��R�(KK��h�C  M           �t�bhhK ��h��R�(KK��h�C�   �   �        �t�bhhK ��h��R�(KK��h�C�   N     E      �t�bhhK ��h��R�(KK��h�CL   8         �      �  �     <  �  	      �        �        �t�bhhK ��h��R�(KK��h�CO           �t�bhhK ��h��R�(KK
��h�C(         T     �     1         �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK��h�C,8            :   �        �         �t�bhhK ��h��R�(KK��h�C4&   �   '     *   	   h  �  �  U   9         �t�bhhK ��h��R�(KK��h�Cd8   "     �  |   	   @  (  �  "   )   	   �  �        1  �  '   e   k      f        �t�bhhK ��h��R�(KK��h�C)  *     �  �        �t�bhhK ��h��R�(KK��h�C    
   +                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C@I   �  �  '   �     8      �  �          �         �t�bhhK ��h��R�(KK	��h�C$�  A     .  �     9         �t�bhhK ��h��R�(KK��h�C I   �  �   �     ,        �t�bhhK ��h��R�(KK��h�C,      �  u   P  )       �        �t�bhhK ��h��R�(KK��h�CI   P  �  �  �        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�   "   R          �t�bhhK ��h��R�(KK��h�C4   8         �        �      Z   >        �t�bhhK ��h��R�(KK��h�C,      g      
   �     q   !        �t�bhhK ��h��R�(KK��h�C<q   p   /   "     >     U   '   x     '   e         �t�bhhK ��h��R�(KK��h�C ?                 E      �t�bhhK ��h��R�(KK��h�C,�   J        �     9     &        �t�bhhK ��h��R�(KK
��h�C(   :  �      �   @     �        �t�bhhK ��h��R�(KK	��h�C$      �   ;     8   A        �t�bhhK ��h��R�(KK��h�C@      -   �      B     <        C        �        �t�bhhK ��h��R�(KK��h�CD     �t�bhhK ��h��R�(KK��h�C=  =     �t�bhhK ��h��R�(KK��h�CTC       y      u     �  �  �  	   �  	   #  -   y      �     �     �t�bhhK ��h��R�(KK
��h�C(&   |  �     9      !   >        �t�bhhK ��h��R�(KK
��h�C($                 E      �     �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C	     1         �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C    8   E  �      �        �t�bhhK ��h��R�(KK��h�C0   �  F  K  G     H  >   �  {        �t�bhhK ��h��R�(KK	��h�C$I  �  u   �  I   2  �        �t�bhhK ��h��R�(KK��h�C0   8   Q   2           %     �        �t�bhhK ��h��R�(KK��h�CH      D   �   �     &  �   \   �  �      )                  �t�bhhK ��h��R�(KK��h�C-   �  �   �        �t�bhhK ��h��R�(KK��h�C�      J           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C,Z     S     ?     *      9         �t�bhhK ��h��R�(KK��h�C@   q   �  �        g      6  .     K     L        �t�bhhK ��h��R�(KK��h�C  M           �t�bhhK ��h��R�(KK��h�C�   �   �        �t�bhhK ��h��R�(KK��h�C�   N     E      �t�bhhK ��h��R�(KK��h�CL   8         �      �  �     <  �  	      �        �        �t�bhhK ��h��R�(KK��h�CO           �t�bhhK ��h��R�(KK
��h�C(         T     �     1         �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK��h�C,8            :   �        �         �t�bhhK ��h��R�(KK��h�C4&   �   '     *   	   h  �  �  U   9         �t�bhhK ��h��R�(KK��h�Cd8   "     �  |   	   @  (  �  "   )   	   �  �        1  �  '   e   k      f        �t�bhhK ��h��R�(KK��h�C)  *     �  �        �t�bhhK ��h��R�(KK��h�C    
   +                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C@I   �  �  '   �     8      �  �          �         �t�bhhK ��h��R�(KK	��h�C$�  A     .  �     9         �t�bhhK ��h��R�(KK��h�C I   �  �   �     ,        �t�bhhK ��h��R�(KK��h�C,      �  u   P  )       �        �t�bhhK ��h��R�(KK��h�CI   P  �  �  �        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�   "   R          �t�bhhK ��h��R�(KK��h�C4   8         �        �      Z   >        �t�bhhK ��h��R�(KK��h�C,      g      
   �     q   !        �t�bhhK ��h��R�(KK��h�C<q   p   /   "     >     U   '   x     '   e         �t�bhhK ��h��R�(KK��h�C?                 �t�bhhK ��h��R�(KK��h�C,�   J        �     9     &        �t�bhhK ��h��R�(KK
��h�C(   :  �      �   @     �        �t�bhhK ��h��R�(KK	��h�C$      �   ;     8   A        �t�bhhK ��h��R�(KK��h�C@      -   �      B     <        C        �        �t�bhhK ��h��R�(KK��h�CD     �t�bhhK ��h��R�(KK��h�C=  =     �t�bhhK ��h��R�(KK��h�CTC       y      u     �  �  �  	   �  	   #  -   y      �     �     �t�bhhK ��h��R�(KK
��h�C(&   |  �     9      !   >        �t�bhhK ��h��R�(KK
��h�C($                 E      �     �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C	     1         �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C    8   E  �      �        �t�bhhK ��h��R�(KK��h�C0   �  F  K  G     H  >   �  {        �t�bhhK ��h��R�(KK	��h�C$I  �  u   �  I   2  �        �t�bhhK ��h��R�(KK��h�C0   8   Q   2           %     �        �t�bhhK ��h��R�(KK��h�CH      D   �   �     &  �   \   �  �      )                  �t�bhhK ��h��R�(KK��h�C-   �  �   �        �t�bhhK ��h��R�(KK��h�C�      J           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C,Z     S     ?     *      9         �t�bhhK ��h��R�(KK��h�C@   q   �  �        g      6  .     K     L        �t�bhhK ��h��R�(KK��h�C  M           �t�bhhK ��h��R�(KK��h�C�   �   �        �t�bhhK ��h��R�(KK��h�C�   N     E      �t�bhhK ��h��R�(KK��h�CL   8         �      �  �     <  �  	      �        �        �t�bhhK ��h��R�(KK��h�CO           �t�bhhK ��h��R�(KK
��h�C(         T     �     1         �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK��h�C,8            :   �        �         �t�bhhK ��h��R�(KK��h�C4&   �   '     *   	   h  �  �  U   9         �t�bhhK ��h��R�(KK��h�Cd8   "     �  |   	   @  (  �  "   )   	   �  �        1  �  '   e   k      f        �t�bhhK ��h��R�(KK��h�C)  *     �  �        �t�bhhK ��h��R�(KK��h�C    
   +                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C@I   �  �  '   �     8      �  �          �         �t�bhhK ��h��R�(KK	��h�C$�  A     .  �     9         �t�bhhK ��h��R�(KK��h�C I   �  �   �     ,        �t�bhhK ��h��R�(KK��h�C,      �  u   P  )       �        �t�bhhK ��h��R�(KK��h�CI   P  �  �  �        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cn     $      L      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C �      �                 �t�bhhK ��h��R�(KK��h�CP   �     B      F   8  ^  	   �   Q  	   R  S  	   T     -        �t�bhhK ��h��R�(KK��h�CB      -   �   k         �t�bhhK ��h��R�(KK��h�CU                 �t�bhhK ��h��R�(KK��h�C   �     B   �        �t�bhhK ��h��R�(KK��h�C   
   .           �t�bhhK ��h��R�(KK��h�C8      �   �  �        �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK��h�C    �      D   Z   �        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C .         �     8         �t�bhhK ��h��R�(KK��h�C�  V        �t�bhhK ��h��R�(KK��h�C1     �t�bhhK ��h��R�(KK��h�C         X        �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CP   8   �        [  9  	   �  	   �   	   W  	   X     [  e         �t�bhhK ��h��R�(KK	��h�C$           D   �   B        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C8�  �  /                 �      �     �      �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C�       �t�bhhK ��h��R�(KK��h�C �    �           9      �t�bhhK ��h��R�(KK��h�CD�     9  	   �   	   �     0  \   1     ^   >   k         �t�bhhK ��h��R�(KK��h�C8                �  Z     r   �   2        �t�bhhK ��h��R�(KK��h�C�   �        �t�bhhK ��h��R�(KK��h�C�  Y                 �t�bhhK ��h��R�(KK��h�C�     $      L      �t�bhhK ��h��R�(KK��h�C@$      �      �   �      8   3     �     8   4        �t�bhhK ��h��R�(KK��h�C0   8      B   D   -     Z   >   �        �t�bhhK ��h��R�(KK
��h�C(   8   �  �   Z   >   �  �        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK	��h�C$         �     $      L      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8   8      Z   >   �   	      F   Z             �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C         X     *      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cn     $      L      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C �      �                 �t�bhhK ��h��R�(KK��h�CP   �     B      F   8  ^  	   �   Q  	   R  S  	   T     -        �t�bhhK ��h��R�(KK��h�CB      -   �   k         �t�bhhK ��h��R�(KK��h�CU                 �t�bhhK ��h��R�(KK��h�C   �     B   �        �t�bhhK ��h��R�(KK��h�C   
   .           �t�bhhK ��h��R�(KK��h�C8      �   �  �        �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK��h�C    �      D   Z   �        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C .         �     8         �t�bhhK ��h��R�(KK��h�C�  V        �t�bhhK ��h��R�(KK��h�C1     �t�bhhK ��h��R�(KK��h�C         X        �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CP   8   �        [  9  	   �  	   �   	   W  	   X     [  e         �t�bhhK ��h��R�(KK	��h�C$           D   �   B        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C8�  �  /                 �      �     �      �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C�       �t�bhhK ��h��R�(KK��h�C �    �           9      �t�bhhK ��h��R�(KK��h�CD�     9  	   �   	   �     0  \   1     ^   >   k         �t�bhhK ��h��R�(KK��h�C8                �  Z     r   �   2        �t�bhhK ��h��R�(KK��h�C�   �        �t�bhhK ��h��R�(KK��h�C�  Y                 �t�bhhK ��h��R�(KK��h�C�     $      L      �t�bhhK ��h��R�(KK��h�C@$      �      �   �      8   3     �     8   4        �t�bhhK ��h��R�(KK��h�C0   8      B   D   -     Z   >   �        �t�bhhK ��h��R�(KK
��h�C(   8   �  �   Z   >   �  �        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK	��h�C$         �     $      L      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8   8      Z   >   �   	      F   Z             �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C         X     *      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cn     $      L      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C �      �                 �t�bhhK ��h��R�(KK��h�CP   �     B      F   8  ^  	   �   Q  	   R  S  	   T     -        �t�bhhK ��h��R�(KK��h�CB      -   �   k         �t�bhhK ��h��R�(KK��h�CU                 �t�bhhK ��h��R�(KK��h�C   �     B   �        �t�bhhK ��h��R�(KK��h�C   
   .           �t�bhhK ��h��R�(KK��h�C8      �   �  �        �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK��h�C    �      D   Z   �        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C .         �     8         �t�bhhK ��h��R�(KK��h�C�  V        �t�bhhK ��h��R�(KK��h�C1     �t�bhhK ��h��R�(KK��h�C         X        �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CP   8   �        [  9  	   �  	   �   	   W  	   X     [  e         �t�bhhK ��h��R�(KK	��h�C$           D   �   B        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C8�  �  /                 �      �     �      �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C�       �t�bhhK ��h��R�(KK��h�C �    �           9      �t�bhhK ��h��R�(KK��h�CD�     9  	   �   	   �     0  \   1     ^   >   k         �t�bhhK ��h��R�(KK��h�C8                �  Z     r   �   2        �t�bhhK ��h��R�(KK��h�C�   �        �t�bhhK ��h��R�(KK��h�C�  Y                 �t�bhhK ��h��R�(KK��h�C�     $      L      �t�bhhK ��h��R�(KK��h�C@$      �      �   �      8   3     �     8   4        �t�bhhK ��h��R�(KK��h�C0   8      B   D   -     Z   >   �        �t�bhhK ��h��R�(KK
��h�C(   8   �  �   Z   >   �  �        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK	��h�C$         �     $      L      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8   8      Z   >   �   	      F   Z             �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C         X     *      �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C,      {      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK	��h�C$5      �  h   n      _   ,      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C0�   �   �   
   .      �   
      M        �t�bhhK ��h��R�(KK��h�C0M   �         5  6  	   7     8        �t�bhhK ��h��R�(KK��h�C,�   4   �   
   .   4         M        �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK$��h�C�0      �      W  �      *   x   �   �   
         J   �  5   +           �  	      F      l   	   ,      k     C  ,         �t�bhhK ��h��R�(KK��h�C,   o        �           e        �t�bhhK ��h��R�(KK��h�C*   0           �t�bhhK ��h��R�(KK��h�C W  �   	   �  �  	   *      �t�bhhK ��h��R�(KK��h�C(      <      D     �t�bhhK ��h��R�(KK��h�C<\  y      h     �  	        [     �  �   �      �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C 0                       �t�bhhK ��h��R�(KK��h�C 9     �   G      1         �t�bhhK ��h��R�(KK��h�C@�     �                  E      �      �      �     �t�bhhK ��h��R�(KK��h�C,      {      �t�bhhK ��h��R�(KK��h�Cl
      "   ,         .   �  �  :  �        w   �      �  	   :     9   Q   0     ;        �t�bhhK ��h��R�(KK��h�C         ,      {      �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C<  =        �t�bhhK ��h��R�(KK��h�C �     >                 �t�bhhK ��h��R�(KK��h�C 9      ?                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C<
        b     '   �   	   �        d   �        �t�bhhK ��h��R�(KK��h�C       �         "        �t�bhhK ��h��R�(KK��h�C<      -           �     �   &      *   E        �t�bhhK ��h��R�(KK��h�C*   E     �t�bhhK ��h��R�(KK��h�C�  1     �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C�                  �t�bhhK ��h��R�(KK��h�C'  \                 �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK	��h�C$�   ~     �        8         �t�bhhK ��h��R�(KK��h�C�   ~        �t�bhhK ��h��R�(KK��h�C�  C  �     �t�bhhK ��h��R�(KK��h�C(   @        �t�bhhK ��h��R�(KK��h�CF  ~           �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�C<
      5   �   +      �     �  	   �   �   �         �t�bhhK ��h��R�(KK��h�CP
        J   �  G  l   p  /      �  /      l   	   =   '   �         �t�bhhK ��h��R�(KK	��h�C$(      <      ]     �        �t�bhhK ��h��R�(KK��h�C+      �     �     �t�bhhK ��h��R�(KK��h�CD�  H     ^  A  "      �     �     �  �     l         �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�CP+      V      I           E      �      �      �      �     �     �t�bhhK ��h��R�(KK��h�C<_     "   ,      l      @   +   M   q   �  `        �t�bhhK ��h��R�(KK��h�C(      <      a     �t�bhhK ��h��R�(KK��h�C+      B           �t�bhhK ��h��R�(KK��h�C         l      �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK��h�C8   ,      m      �         @   +      �         �t�bhhK ��h��R�(KK��h�C�   �        8         �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK��h�Cn      _   ,      �t�bhhK ��h��R�(KK��h�C0   ,      V  $   ?   �   	   =   J        �t�bhhK ��h��R�(KK��h�CJ     �t�bhhK ��h��R�(KK��h�C,(      <      �        <      �     �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C8   ,      V  $      �   x      F   j  0        �t�bhhK ��h��R�(KK��h�CK           �t�bhhK ��h��R�(KK��h�CX
      5   f      �   :  n   C  �     �  	         �      }   d   �         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�CH      L  
     ,      j     �  0     :   �      �        �t�bhhK ��h��R�(KK��h�C,&   L   %           D   =   �         �t�bhhK ��h��R�(KK��h�CP        4           v  �   M     =   �   	  
  !  _   (        �t�bhhK ��h��R�(KK��h�C"        �        �t�bhhK ��h��R�(KK��h�C:   _   (     �t�bhhK ��h��R�(KK��h�C(      <      C     �t�bhhK ��h��R�(KK��h�C�   	  
        �t�bhhK ��h��R�(KK��h�C:   _   #     �t�bhhK ��h��R�(KK��h�C          n      _   ,      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C\
      �  N     /   b  D  	         @   V      )        �  	   (   �        �t�bhhK ��h��R�(KK
��h�C(8      "      �   c     �        �t�bhhK ��h��R�(KK��h�C &      �     H   |         �t�bhhK ��h��R�(KK��h�C         �     �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C,      {      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK	��h�C$5      �  h   n      _   ,      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C0�   �   �   
   .      �   
      M        �t�bhhK ��h��R�(KK��h�C0M   �         5  6  	   7     8        �t�bhhK ��h��R�(KK��h�C,�   4   �   
   .   4         M        �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK$��h�C�0      �      W  �      *   x   �   �   
         J   �  5   +           �  	      F      l   	   ,      k     C  ,         �t�bhhK ��h��R�(KK��h�C,   o        �           e        �t�bhhK ��h��R�(KK��h�C*   0           �t�bhhK ��h��R�(KK��h�C W  �   	   �  �  	   *      �t�bhhK ��h��R�(KK��h�C(      <      D     �t�bhhK ��h��R�(KK��h�C<\  y      h     �  	        [     �  �   �      �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C 0                       �t�bhhK ��h��R�(KK��h�C 9     �   G      1         �t�bhhK ��h��R�(KK��h�C@�     �                  E      �      �      �     �t�bhhK ��h��R�(KK��h�C,      {      �t�bhhK ��h��R�(KK��h�Cl
      "   ,         .   �  �  :  �        w   �      �  	   :     9   Q   0     ;        �t�bhhK ��h��R�(KK��h�C         ,      {      �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C<  =        �t�bhhK ��h��R�(KK��h�C �     >                 �t�bhhK ��h��R�(KK��h�C 9      ?                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C<
        b     '   �   	   �        d   �        �t�bhhK ��h��R�(KK��h�C       �         "        �t�bhhK ��h��R�(KK��h�C<      -           �     �   &      *   E        �t�bhhK ��h��R�(KK��h�C*   E     �t�bhhK ��h��R�(KK��h�C�  1     �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C�                  �t�bhhK ��h��R�(KK��h�C'  \                 �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK	��h�C$�   ~     �        8         �t�bhhK ��h��R�(KK��h�C�   ~        �t�bhhK ��h��R�(KK��h�C�  C  �     �t�bhhK ��h��R�(KK��h�C(   @        �t�bhhK ��h��R�(KK��h�CF  ~           �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�C<
      5   �   +      �     �  	   �   �   �         �t�bhhK ��h��R�(KK��h�CP
        J   �  G  l   p  /      �  /      l   	   =   '   �         �t�bhhK ��h��R�(KK	��h�C$(      <      ]     �        �t�bhhK ��h��R�(KK��h�C+      �     �     �t�bhhK ��h��R�(KK��h�CD�  H     ^  A  "      �     �     �  �     l         �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�CP+      V      I           E      �      �      �      �     �     �t�bhhK ��h��R�(KK��h�C<_     "   ,      l      @   +   M   q   �  `        �t�bhhK ��h��R�(KK��h�C(      <      a     �t�bhhK ��h��R�(KK��h�C+      B           �t�bhhK ��h��R�(KK��h�C         l      �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK��h�C8   ,      m      �         @   +      �         �t�bhhK ��h��R�(KK��h�C�   �        8         �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK��h�Cn      _   ,      �t�bhhK ��h��R�(KK��h�C0   ,      V  $   ?   �   	   =   J        �t�bhhK ��h��R�(KK��h�CJ     �t�bhhK ��h��R�(KK��h�C,(      <      �        <      �     �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C8   ,      V  $      �   x      F   j  0        �t�bhhK ��h��R�(KK��h�CK           �t�bhhK ��h��R�(KK��h�CX
      5   f      �   :  n   C  �     �  	         �      }   d   �         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�CH      L  
     ,      j     �  0     :   �      �        �t�bhhK ��h��R�(KK��h�C,&   L   %           D   =   �         �t�bhhK ��h��R�(KK��h�CP        4           v  �   M     =   �   	  
  !  _   (        �t�bhhK ��h��R�(KK��h�C"        �        �t�bhhK ��h��R�(KK��h�C:   _   (     �t�bhhK ��h��R�(KK��h�C(      <      C     �t�bhhK ��h��R�(KK��h�C�   	  
        �t�bhhK ��h��R�(KK��h�C:   _   #     �t�bhhK ��h��R�(KK��h�C          n      _   ,      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C\
      �  N     /   b  D  	         @   V      )        �  	   (   �        �t�bhhK ��h��R�(KK
��h�C(8      "      �   c     �        �t�bhhK ��h��R�(KK��h�C &      �     H   |         �t�bhhK ��h��R�(KK��h�C         �     �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C,      {      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK	��h�C$5      �  h   n      _   ,      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C0�   �   �   
   .      �   
      M        �t�bhhK ��h��R�(KK��h�C0M   �         5  6  	   7     8        �t�bhhK ��h��R�(KK��h�C,�   4   �   
   .   4         M        �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK$��h�C�0      �      W  �      *   x   �   �   
         J   �  5   +           �  	      F      l   	   ,      k     C  ,         �t�bhhK ��h��R�(KK��h�C,   o        �           e        �t�bhhK ��h��R�(KK��h�C*   0           �t�bhhK ��h��R�(KK��h�C W  �   	   �  �  	   *      �t�bhhK ��h��R�(KK��h�C(      <      D     �t�bhhK ��h��R�(KK��h�C<\  y      h     �  	        [     �  �   �      �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C 0                       �t�bhhK ��h��R�(KK��h�C 9     �   G      1         �t�bhhK ��h��R�(KK��h�C@�     �                  E      �      �      �     �t�bhhK ��h��R�(KK��h�C,      {      �t�bhhK ��h��R�(KK��h�Cl
      "   ,         .   �  �  :  �        w   �      �  	   :     9   Q   0     ;        �t�bhhK ��h��R�(KK��h�C         ,      {      �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C<  =        �t�bhhK ��h��R�(KK��h�C �     >                 �t�bhhK ��h��R�(KK��h�C 9      ?                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C<
        b     '   �   	   �        d   �        �t�bhhK ��h��R�(KK��h�C       �         "        �t�bhhK ��h��R�(KK��h�C<      -           �     �   &      *   E        �t�bhhK ��h��R�(KK��h�C*   E     �t�bhhK ��h��R�(KK��h�C�  1     �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C�                  �t�bhhK ��h��R�(KK��h�C'  \                 �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK	��h�C$�   ~     �        8         �t�bhhK ��h��R�(KK��h�C�   ~        �t�bhhK ��h��R�(KK��h�C�  C  �     �t�bhhK ��h��R�(KK��h�C(   @        �t�bhhK ��h��R�(KK��h�CF  ~           �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�C<
      5   �   +      �     �  	   �   �   �         �t�bhhK ��h��R�(KK��h�CP
        J   �  G  l   p  /      �  /      l   	   =   '   �         �t�bhhK ��h��R�(KK	��h�C$(      <      ]     �        �t�bhhK ��h��R�(KK��h�C+      �     �     �t�bhhK ��h��R�(KK��h�CD�  H     ^  A  "      �     �     �  �     l         �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�CP+      V      I           E      �      �      �      �     �     �t�bhhK ��h��R�(KK��h�C<_     "   ,      l      @   +   M   q   �  `        �t�bhhK ��h��R�(KK��h�C(      <      a     �t�bhhK ��h��R�(KK��h�C+      B           �t�bhhK ��h��R�(KK��h�C         l      �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK��h�C8   ,      m      �         @   +      �         �t�bhhK ��h��R�(KK��h�C�   �        8         �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK��h�Cn      _   ,      �t�bhhK ��h��R�(KK��h�C0   ,      V  $   ?   �   	   =   J        �t�bhhK ��h��R�(KK��h�CJ     �t�bhhK ��h��R�(KK��h�C,(      <      �        <      �     �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C8   ,      V  $      �   x      F   j  0        �t�bhhK ��h��R�(KK��h�CK           �t�bhhK ��h��R�(KK��h�CX
      5   f      �   :  n   C  �     �  	         �      }   d   �         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�CH      L  
     ,      j     �  0     :   �      �        �t�bhhK ��h��R�(KK��h�C,&   L   %           D   =   �         �t�bhhK ��h��R�(KK��h�CP        4           v  �   M     =   �   	  
  !  _   (        �t�bhhK ��h��R�(KK��h�C"        �        �t�bhhK ��h��R�(KK��h�C:   _   (     �t�bhhK ��h��R�(KK��h�C(      <      C     �t�bhhK ��h��R�(KK��h�C�   	  
        �t�bhhK ��h��R�(KK��h�C:   _   #     �t�bhhK ��h��R�(KK��h�C          n      _   ,      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C\
      �  N     /   b  D  	         @   V      )        �  	   (   �        �t�bhhK ��h��R�(KK
��h�C(8      "      �   c     �        �t�bhhK ��h��R�(KK��h�C &      �     H   |         �t�bhhK ��h��R�(KK��h�C         �     �t�bhhK ��h��R�(KK��h�Cm      �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C$      b      �t�bhhK ��h��R�(KK��h�Co      z      �t�bhhK ��h��R�(KK��h�Cm      �t�bhhK ��h��R�(KK��h�C4�  �  6      d  $  �     O  p  m         �t�bhhK ��h��R�(KK��h�Ce  �     �         �t�bhhK ��h��R�(KK��h�C,         �     O  p  m   	   �     �t�bhhK ��h��R�(KK��h�C �      �                 �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C8d     e     �   �   g     �   ~   f  �        �t�bhhK ��h��R�(KK��h�C<      D   g   b   g  	   �   J   E     F  G        �t�bhhK ��h��R�(KK��h�CL        �   `      h  �  �     	   i     M                �t�bhhK ��h��R�(KK��h�C�   ~   h     �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�C         b      �t�bhhK ��h��R�(KK��h�CF  ~   h        �t�bhhK ��h��R�(KK��h�C�            �t�bhhK ��h��R�(KK��h�C$      b      �t�bhhK ��h��R�(KK��h�C<
      "   $      6   j  /   	   w   �      �        �t�bhhK ��h��R�(KK��h�C<H  �  '   k  
   �  �   	   l  	   �     �        �t�bhhK ��h��R�(KK��h�C         $      b      �t�bhhK ��h��R�(KK��h�C l  
   $      �           �t�bhhK ��h��R�(KK��h�Co      z      �t�bhhK ��h��R�(KK��h�C8   j   �   P     8         
   �      $         �t�bhhK ��h��R�(KK��h�Co      z      �      �t�bhhK ��h��R�(KK��h�C\
      2  r   $   �        �      8   Q   �   �     v         I  W   J        �t�bhhK ��h��R�(KK��h�C,         V      o      $      �      �t�bhhK ��h��R�(KK��h�Cx  �           �t�bhhK ��h��R�(KK��h�C V      �     �           �t�bhhK ��h��R�(KK��h�Cm      �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C$      b      �t�bhhK ��h��R�(KK��h�Co      z      �t�bhhK ��h��R�(KK��h�Cm      �t�bhhK ��h��R�(KK��h�C4�  �  6      d  $  �     O  p  m         �t�bhhK ��h��R�(KK��h�Ce  �     �         �t�bhhK ��h��R�(KK��h�C,         �     O  p  m   	   �     �t�bhhK ��h��R�(KK��h�C �      �                 �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C8d     e     �   �   g     �   ~   f  �        �t�bhhK ��h��R�(KK��h�C<      D   g   b   g  	   �   J   E     F  G        �t�bhhK ��h��R�(KK��h�CL        �   `      h  �  �     	   i     M                �t�bhhK ��h��R�(KK��h�C�   ~   h     �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�C         b      �t�bhhK ��h��R�(KK��h�CF  ~   h        �t�bhhK ��h��R�(KK��h�C�            �t�bhhK ��h��R�(KK��h�C$      b      �t�bhhK ��h��R�(KK��h�C<
      "   $      6   j  /   	   w   �      �        �t�bhhK ��h��R�(KK��h�C<H  �  '   k  
   �  �   	   l  	   �     �        �t�bhhK ��h��R�(KK��h�C         $      b      �t�bhhK ��h��R�(KK��h�C l  
   $      �           �t�bhhK ��h��R�(KK��h�Co      z      �t�bhhK ��h��R�(KK��h�C8   j   �   P     8         
   �      $         �t�bhhK ��h��R�(KK��h�Co      z      �      �t�bhhK ��h��R�(KK��h�C\
      2  r   $   �        �      8   Q   �   �     v         I  W   J        �t�bhhK ��h��R�(KK��h�C,         V      o      $      �      �t�bhhK ��h��R�(KK��h�Cx  �           �t�bhhK ��h��R�(KK��h�C V      �     �           �t�bhhK ��h��R�(KK��h�Cm      �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C$      b      �t�bhhK ��h��R�(KK��h�Co      z      �t�bhhK ��h��R�(KK��h�Cm      �t�bhhK ��h��R�(KK��h�C4�  �  6      d  $  �     O  p  m         �t�bhhK ��h��R�(KK��h�Ce  �     �         �t�bhhK ��h��R�(KK��h�C,         �     O  p  m   	   �     �t�bhhK ��h��R�(KK��h�C �      �                 �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C8d     e     �   �   g     �   ~   f  �        �t�bhhK ��h��R�(KK��h�C<      D   g   b   g  	   �   J   E     F  G        �t�bhhK ��h��R�(KK��h�CL        �   `      h  �  �     	   i     M                �t�bhhK ��h��R�(KK��h�C�   ~   h     �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�C         b      �t�bhhK ��h��R�(KK��h�CF  ~   h        �t�bhhK ��h��R�(KK��h�C�            �t�bhhK ��h��R�(KK��h�C$      b      �t�bhhK ��h��R�(KK��h�C<
      "   $      6   j  /   	   w   �      �        �t�bhhK ��h��R�(KK��h�C<H  �  '   k  
   �  �   	   l  	   �     �        �t�bhhK ��h��R�(KK��h�C         $      b      �t�bhhK ��h��R�(KK��h�C l  
   $      �           �t�bhhK ��h��R�(KK��h�Co      z      �t�bhhK ��h��R�(KK��h�C8   j   �   P     8         
   �      $         �t�bhhK ��h��R�(KK��h�Co      z      �      �t�bhhK ��h��R�(KK��h�C\
      2  r   $   �        �      8   Q   �   �     v         I  W   J        �t�bhhK ��h��R�(KK��h�C,         V      o      $      �      �t�bhhK ��h��R�(KK��h�Cx  �           �t�bhhK ��h��R�(KK��h�C V      �     �           �t�bhhK ��h��R�(KK��h�C�     8      �t�bhhK ��h��R�(KK��h�Cn   G      �t�bhhK ��h��R�(KK��h�C�   �  G      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�   G      �t�bhhK ��h��R�(KK��h�CK     �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�C�   Y      �t�bhhK ��h��R�(KK��h�C4�   �   �   
   .      �   
      �   M        �t�bhhK ��h��R�(KK��h�CD�   �      F         �  �     N     �        L        �t�bhhK ��h��R�(KK��h�C,�   4   �   
   .   4         M        �t�bhhK ��h��R�(KK��h�CH
      "   J   S     8   	         �  :   �   �     }        �t�bhhK ��h��R�(KK��h�CD�   �     M  8     F      5  	   �  	   Q     �         �t�bhhK ��h��R�(KK��h�C\
      4   "   �       �   :   �   �     }  	         g   /         �   �        �t�bhhK ��h��R�(KK��h�C0      �   �  �      �  3  ~  %        �t�bhhK ��h��R�(KK��h�C         G      �t�bhhK ��h��R�(KK��h�C�     8      �t�bhhK ��h��R�(KK��h�C,   8   8  �   �     M     �         �t�bhhK ��h��R�(KK��h�C,   �      N  	   O     P  Q        �t�bhhK ��h��R�(KK��h�C,�   "   �   \  y      u     	        �t�bhhK ��h��R�(KK��h�CL
      5   o   ?     E  6      =   �   .     �  N   �   m        �t�bhhK ��h��R�(KK��h�C8   �      �t�bhhK ��h��R�(KK��h�Cn  %     �t�bhhK ��h��R�(KK��h�C�  8      �t�bhhK ��h��R�(KK��h�C(      <      R     �t�bhhK ��h��R�(KK��h�Co                 �t�bhhK ��h��R�(KK��h�C�   �     �t�bhhK ��h��R�(KK��h�CD   
   �   �  7         S  T     *      T     9         �t�bhhK ��h��R�(KK��h�C-     �t�bhhK ��h��R�(KK��h�C       �   -     �        �t�bhhK ��h��R�(KK��h�C0�     �     8      �  h  	   8         �t�bhhK ��h��R�(KK��h�C         -        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�CU        �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�CL   9      3  X  	   v   Y      �     1   �   >     @   �        �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�C8�            E      �      �      �     �     �t�bhhK ��h��R�(KK��h�C         �      1      �t�bhhK ��h��R�(KK	��h�C$�     ?   B  "   �   �        �t�bhhK ��h��R�(KK
��h�C(�     z  �     �     �         �t�bhhK ��h��R�(KK��h�C,&   |  �         W  �      *         �t�bhhK ��h��R�(KK��h�C8�   &   R  �     (          U     �         �t�bhhK ��h��R�(KK��h�Ce     W  �      �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C�      ~   q  �        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C         �      1      �t�bhhK ��h��R�(KK��h�Cn   G      �t�bhhK ��h��R�(KK��h�CH   �     �     $   ?   �   O   B   +      �  0     @        �t�bhhK ��h��R�(KK��h�CD#        �   
   f      @   V      �     �     $         �t�bhhK ��h��R�(KK	��h�C$   �  6  �   G      �        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C4N   z     �  6         �  =   8   �         �t�bhhK ��h��R�(KK��h�C8   �      �t�bhhK ��h��R�(KK��h�Cn  %     �t�bhhK ��h��R�(KK��h�C�  8      �t�bhhK ��h��R�(KK��h�C(      <      R     �t�bhhK ��h��R�(KK��h�Co                 �t�bhhK ��h��R�(KK��h�C �  �   �   
   �  G         �t�bhhK ��h��R�(KK��h�CK           �t�bhhK ��h��R�(KK��h�C\?   �     B     �      $   ?   /  I      W  �      *         �     9         �t�bhhK ��h��R�(KK��h�C�      ~   q  �        �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK��h�C         n   G      �t�bhhK ��h��R�(KK��h�C�   �  G      �t�bhhK ��h��R�(KK��h�C<
         ;  A  I         =   ;     8   �         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C4�     S     �  	      �     )            �t�bhhK ��h��R�(KK��h�C�      �t�b�       hhK ��h��R�(KK��h�C,�     V     8   �   C             �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C\�      W    "   �   \  y      p     F     �     [  y      �     F        �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C�     �           �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C    8      D   �   �        �t�bhhK ��h��R�(KK��h�C\
   
      4   "   �       �   :   �   �     }  	                 �   �        �t�bhhK ��h��R�(KK	��h�C$�   �      �  B  X  �         �t�bhhK ��h��R�(KK��h�C�   Y           �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C�   G      �t�bhhK ��h��R�(KK��h�C8
      5   q  +      �  V         =   �         �t�bhhK ��h��R�(KK��h�C8   �      �t�bhhK ��h��R�(KK��h�Cn  %     �t�bhhK ��h��R�(KK��h�C�  8      �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�C<*   0           W  �   �   Y      �     8         �t�bhhK ��h��R�(KK��h�C,   o        �           e        �t�bhhK ��h��R�(KK��h�C*   0           �t�bhhK ��h��R�(KK��h�C W  �   	   �  �  	   *      �t�bhhK ��h��R�(KK��h�C(      <      D     �t�bhhK ��h��R�(KK��h�C<\  y      h     �  	        [     �  �   �      �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C         �   G      �t�bhhK ��h��R�(KK��h�CK     �t�bhhK ��h��R�(KK��h�C4   D     �  O      +      �     �        �t�bhhK ��h��R�(KK��h�C8�  Z     �         t     �     9            �t�bhhK ��h��R�(KK��h�Co                 �t�bhhK ��h��R�(KK��h�C�      ~   q  �        �t�bhhK ��h��R�(KK��h�C t     [                 �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�C8   \  6  �  	   ]     �  A  ^  ?   �        �t�bhhK ��h��R�(KK��h�C,=   �  N      _            �        �t�bhhK ��h��R�(KK��h�C b  \  y      J     r     �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK
��h�C(.   |  �     W  �      *         �t�bhhK ��h��R�(KK��h�CX
      �         -   �  z      �   e   �   �   9      ~   q     �           �t�bhhK ��h��R�(KK��h�C�      ~   q  �        �t�bhhK ��h��R�(KK��h�C      �                 �t�bhhK ��h��R�(KK��h�C�      ~   q        �t�bhhK ��h��R�(KK��h�C`  a                 �t�bhhK ��h��R�(KK��h�C         T     �t�bhhK ��h��R�(KK��h�C�   Y      �t�bhhK ��h��R�(KK��h�C<8      T   >   ;      �   	      F   �     �        �t�bhhK ��h��R�(KK��h�C8      �   
   �      �   d   �     r   �        �t�bhhK ��h��R�(KK��h�C;   �   �           �t�bhhK ��h��R�(KK��h�C         �   Y      �t�bhhK ��h��R�(KK��h�C�     8      �t�bhhK ��h��R�(KK��h�Cn   G      �t�bhhK ��h��R�(KK��h�C�   �  G      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�   G      �t�bhhK ��h��R�(KK��h�CK     �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�C�   Y      �t�bhhK ��h��R�(KK��h�C4�   �   �   
   .      �   
      �   M        �t�bhhK ��h��R�(KK��h�CD�   �      F         �  �     N     �        L        �t�bhhK ��h��R�(KK��h�C,�   4   �   
   .   4         M        �t�bhhK ��h��R�(KK��h�CH
      "   J   S     8   	         �  :   �   �     }        �t�bhhK ��h��R�(KK��h�CD�   �     M  8     F      5  	   �  	   Q     �         �t�bhhK ��h��R�(KK��h�C\
      4   "   �       �   :   �   �     }  	         g   /         �   �        �t�bhhK ��h��R�(KK��h�C0      �   �  �      �  3  ~  %        �t�bhhK ��h��R�(KK��h�C         G      �t�bhhK ��h��R�(KK��h�C�     8      �t�bhhK ��h��R�(KK��h�C,   8   8  �   �     M     �         �t�bhhK ��h��R�(KK��h�C,   �      N  	   O     P  Q        �t�bhhK ��h��R�(KK��h�C,�   "   �   \  y      u     	        �t�bhhK ��h��R�(KK��h�CL
      5   o   ?     E  6      =   �   .     �  N   �   m        �t�bhhK ��h��R�(KK��h�C8   �      �t�bhhK ��h��R�(KK��h�Cn  %     �t�bhhK ��h��R�(KK��h�C�  8      �t�bhhK ��h��R�(KK��h�C(      <      R     �t�bhhK ��h��R�(KK��h�Co                 �t�bhhK ��h��R�(KK��h�C�   �     �t�bhhK ��h��R�(KK��h�CD   
   �   �  7         S  T     *      T     9         �t�bhhK ��h��R�(KK��h�C-     �t�bhhK ��h��R�(KK��h�C       �   -     �        �t�bhhK ��h��R�(KK��h�C0�     �     8      �  h  	   8         �t�bhhK ��h��R�(KK��h�C         -        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�CU        �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�CL   9      3  X  	   v   Y      �     1   �   >     @   �        �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�C8�            E      �      �      �     �     �t�bhhK ��h��R�(KK��h�C         �      1      �t�bhhK ��h��R�(KK	��h�C$�     ?   B  "   �   �        �t�bhhK ��h��R�(KK
��h�C(�     z  �     �     �         �t�bhhK ��h��R�(KK��h�C,&   |  �         W  �      *         �t�bhhK ��h��R�(KK��h�C8�   &   R  �     (          U     �         �t�bhhK ��h��R�(KK��h�Ce     W  �      �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C�      ~   q  �        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C         �      1      �t�bhhK ��h��R�(KK��h�Cn   G      �t�bhhK ��h��R�(KK��h�CH   �     �     $   ?   �   O   B   +      �  0     @        �t�bhhK ��h��R�(KK��h�CD#        �   
   f      @   V      �     �     $         �t�bhhK ��h��R�(KK	��h�C$   �  6  �   G      �        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C4N   z     �  6         �  =   8   �         �t�bhhK ��h��R�(KK��h�C8   �      �t�bhhK ��h��R�(KK��h�Cn  %     �t�bhhK ��h��R�(KK��h�C�  8      �t�bhhK ��h��R�(KK��h�C(      <      R     �t�bhhK ��h��R�(KK��h�Co                 �t�bhhK ��h��R�(KK��h�C �  �   �   
   �  G         �t�bhhK ��h��R�(KK��h�CK           �t�bhhK ��h��R�(KK��h�C\?   �     B     �      $   ?   /  I      W  �      *         �     9         �t�bhhK ��h��R�(KK��h�C�      ~   q  �        �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK��h�C         n   G      �t�bhhK ��h��R�(KK��h�C�   �  G      �t�bhhK ��h��R�(KK��h�C<
         ;  A  I         =   ;     8   �         �t�bhhK ��h��R�(KK��h�C    
   ;      "           �t�bhhK ��h��R�(KK��h�C4�     S     �  	      �     )            �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C,�     V     8   �   C             �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C\�      W    "   �   \  y      p     F     �     [  y      �     F        �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C�     �           �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C    8      D   �   �        �t�bhhK ��h��R�(KK��h�C\
   
      4   "   �       �   :   �   �     }  	                 �   �        �t�bhhK ��h��R�(KK	��h�C$�   �      �  B  X  �         �t�bhhK ��h��R�(KK��h�C�   Y           �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C�   G      �t�bhhK ��h��R�(KK��h�C8
      5   q  +      �  V         =   �         �t�bhhK ��h��R�(KK��h�C8   �      �t�bhhK ��h��R�(KK��h�Cn  %     �t�bhhK ��h��R�(KK��h�C�  8      �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�C<*   0           W  �   �   Y      �     8         �t�bhhK ��h��R�(KK��h�C,   o        �           e        �t�bhhK ��h��R�(KK��h�C*   0           �t�bhhK ��h��R�(KK��h�C W  �   	   �  �  	   *      �t�bhhK ��h��R�(KK��h�C(      <      D     �t�bhhK ��h��R�(KK��h�C<\  y      h     �  	        [     �  �   �      �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C         �   G      �t�bhhK ��h��R�(KK��h�CK     �t�bhhK ��h��R�(KK��h�C4   D     �  O      +      �     �        �t�bhhK ��h��R�(KK��h�C8�  Z     �         t     �     9            �t�bhhK ��h��R�(KK��h�Co                 �t�bhhK ��h��R�(KK��h�C�      ~   q  �        �t�bhhK ��h��R�(KK��h�C t     [                 �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�C8   \  6  �  	   ]     �  A  ^  ?   �        �t�bhhK ��h��R�(KK��h�C,=   �  N      _            �        �t�bhhK ��h��R�(KK��h�C b  \  y      J     r     �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK
��h�C(.   |  �     W  �      *         �t�bhhK ��h��R�(KK��h�CX
      �         -   �  z      �   e   �   �   9      ~   q     �           �t�bhhK ��h��R�(KK��h�C�      ~   q  �        �t�bhhK ��h��R�(KK��h�C      �                 �t�bhhK ��h��R�(KK��h�C�      ~   q        �t�bhhK ��h��R�(KK��h�C`  a                 �t�bhhK ��h��R�(KK��h�C         T     �t�bhhK ��h��R�(KK��h�C�   Y      �t�bhhK ��h��R�(KK��h�C<8      T   >   ;      �   	      F   �     �        �t�bhhK ��h��R�(KK��h�C8      �   
   �      �   d   �     r   �        �t�bhhK ��h��R�(KK��h�C;   �   �           �t�bhhK ��h��R�(KK��h�C         �   Y      �t�bhhK ��h��R�(KK��h�C�     8      �t�bhhK ��h��R�(KK��h�Cn   G      �t�bhhK ��h��R�(KK��h�C�   �  G      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�   G      �t�bhhK ��h��R�(KK��h�CK     �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�C�   Y      �t�bhhK ��h��R�(KK��h�C4�   �   �   
   .      �   
      �   M        �t�bhhK ��h��R�(KK��h�CD�   �      F         �  �     N     �        L        �t�bhhK ��h��R�(KK��h�C,�   4   �   
   .   4         M        �t�bhhK ��h��R�(KK��h�CH
      "   J   S     8   	         �  :   �   �     }        �t�bhhK ��h��R�(KK��h�CD�   �     M  8     F      5  	   �  	   Q     �         �t�bhhK ��h��R�(KK��h�C\
      4   "   �       �   :   �   �     }  	         g   /         �   �        �t�bhhK ��h��R�(KK��h�C0      �   �  �      �  3  ~  %        �t�be(hhK ��h��R�(KK��h�C         G      �t�bhhK ��h��R�(KK��h�C�     8      �t�bhhK ��h��R�(KK��h�C,   8   8  �   �     M     �         �t�bhhK ��h��R�(KK��h�C,   �      N  	   O     P  Q        �t�bhhK ��h��R�(KK��h�C,�   "   �   \  y      u     	        �t�bhhK ��h��R�(KK��h�CL
      5   o   ?     E  6      =   �   .     �  N   �   m        �t�bhhK ��h��R�(KK��h�C8   �      �t�bhhK ��h��R�(KK��h�Cn  %     �t�bhhK ��h��R�(KK��h�C�  8      �t�bhhK ��h��R�(KK��h�C(      <      R     �t�bhhK ��h��R�(KK��h�Co           �t�bhhK ��h��R�(KK��h�C�   �     �t�bhhK ��h��R�(KK��h�CD   
   �   �  7         S  T     *      T     9         �t�bhhK ��h��R�(KK��h�C-     �t�bhhK ��h��R�(KK��h�C       �   -     �        �t�bhhK ��h��R�(KK��h�C0�     �     8      �  h  	   8         �t�bhhK ��h��R�(KK��h�C         -        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�CU        �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�CL   9      3  X  	   v   Y      �     1   �   >     @   �        �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�C8�            E      �      �      �     �     �t�bhhK ��h��R�(KK��h�C         �      1      �t�bhhK ��h��R�(KK	��h�C$�     ?   B  "   �   �        �t�bhhK ��h��R�(KK
��h�C(�     z  �     �     �         �t�bhhK ��h��R�(KK��h�C,&   |  �         W  �      *         �t�bhhK ��h��R�(KK��h�C8�   &   R  �     (          U     �         �t�bhhK ��h��R�(KK��h�Ce     W  �      �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C�      ~   q  �        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C         �      1      �t�bhhK ��h��R�(KK��h�Cn   G      �t�bhhK ��h��R�(KK��h�CH   �     �     $   ?   �   O   B   +      �  0     @        �t�bhhK ��h��R�(KK��h�CD#        �   
   f      @   V      �     �     $         �t�bhhK ��h��R�(KK	��h�C$   �  6  �   G      �        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C4N   z     �  6         �  =   8   �         �t�bhhK ��h��R�(KK��h�C8   �      �t�bhhK ��h��R�(KK��h�Cn  %     �t�bhhK ��h��R�(KK��h�C�  8      �t�bhhK ��h��R�(KK��h�C(      <      R     �t�bhhK ��h��R�(KK��h�Co           �t�bhhK ��h��R�(KK��h�C �  �   �   
   �  G         �t�bhhK ��h��R�(KK��h�CK           �t�bhhK ��h��R�(KK��h�C\?   �     B     �      $   ?   /  I      W  �      *         �     9         �t�bhhK ��h��R�(KK��h�C�      ~   q  �        �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK��h�C         n   G      �t�bhhK ��h��R�(KK��h�C�   �  G      �t�bhhK ��h��R�(KK��h�C<
         ;  A  I         =   ;     8   �         �t�bhhK ��h��R�(KK��h�C    
   ;      "           �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C,�     V     8   �   C             �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C\�      W    "   �   \  y      p     F     �     [  y      �     F        �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C�     �           �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C    8      D   �   �        �t�bhhK ��h��R�(KK��h�C\
   
      4   "   �       �   :   �   �     }  	                 �   �        �t�bhhK ��h��R�(KK	��h�C$�   �      �  B  X  �         �t�bhhK ��h��R�(KK��h�C�   Y           �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C�   G      �t�bhhK ��h��R�(KK��h�C8
      5   q  +      �  V         =   �         �t�bhhK ��h��R�(KK��h�C8   �      �t�bhhK ��h��R�(KK��h�Cn  %     �t�bhhK ��h��R�(KK��h�C�  8      �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�C<*   0           W  �   �   Y      �     8         �t�bhhK ��h��R�(KK��h�C,   o        �           e        �t�bhhK ��h��R�(KK��h�C*   0           �t�bhhK ��h��R�(KK��h�C W  �   	   �  �  	   *      �t�bhhK ��h��R�(KK��h�C(      <      D     �t�bhhK ��h��R�(KK��h�C<\  y      h     �  	        [     �  �   �      �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C         �   G      �t�bhhK ��h��R�(KK��h�CK     �t�bhhK ��h��R�(KK��h�C4   D     �  O      +      �     �        �t�bhhK ��h��R�(KK��h�C8�  Z     �         t     �     9            �t�bhhK ��h��R�(KK��h�Co           �t�bhhK ��h��R�(KK��h�C�      ~   q  �        �t�bhhK ��h��R�(KK��h�C t     [                 �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�C8   \  6  �  	   ]     �  A  ^  ?   �        �t�bhhK ��h��R�(KK��h�C,=   �  N      _            �        �t�bhhK ��h��R�(KK��h�C b  \  y      J     r     �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK
��h�C(.   |  �     W  �      *         �t�bhhK ��h��R�(KK��h�CX
      �         -   �  z      �   e   �   �   9      ~   q     �           �t�bhhK ��h��R�(KK��h�C�      ~   q  �        �t�bhhK ��h��R�(KK��h�C      �                 �t�bhhK ��h��R�(KK��h�C�      ~   q        �t�bhhK ��h��R�(KK��h�C`  a                 �t�bhhK ��h��R�(KK��h�C         T     �t�bhhK ��h��R�(KK��h�C�   Y      �t�bhhK ��h��R�(KK��h�C<8      T   >   ;      �   	      F   �     �        �t�bhhK ��h��R�(KK��h�C8      �   
   �      �   d   �     r   �        �t�bhhK ��h��R�(KK��h�C;   �   �           �t�bhhK ��h��R�(KK��h�C         �   Y      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cz     �t�bhhK ��h��R�(KK��h�CW   �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8   8      H   �   �   	   �   �      �   l        �t�bhhK ��h��R�(KK	��h�C$�   �     )                  �t�bhhK ��h��R�(KK	��h�C$   8      D   '   �  �         �t�bhhK ��h��R�(KK��h�CD�  
   �     r   $   w  �   n    z   6   f     &        �t�bhhK ��h��R�(KK��h�C@
      �   
   �     �  �  6      �   &   &  `         �t�bhhK ��h��R�(KK��h�C8      D   b  �     T        9     D        �t�bhhK ��h��R�(KK	��h�C$�   �   `      T     D        �t�bhhK ��h��R�(KK��h�CP     �     8      D   g   �     v  $      *   	   9      !         �t�bhhK ��h��R�(KK��h�C,   6   c  �   �   J   `      8         �t�bhhK ��h��R�(KK��h�C             q            �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C �                       �t�bhhK ��h��R�(KK��h�C`   
   d           �t�bhhK ��h��R�(KK��h�C     e  r           �t�bhhK ��h��R�(KK��h�C                   �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C    8   �       U        �t�bhhK ��h��R�(KK��h�C,            f                �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C    
   g                 �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK��h�CX   8      �             �  h     �     �  6        �     �        �t�bhhK ��h��R�(KK��h�C8
      "   �   
   &   [            =   i        �t�bhhK ��h��R�(KK��h�Ci     �t�bhhK ��h��R�(KK��h�C8   A     �t�bhhK ��h��R�(KK��h�C=  =     �t�bhhK ��h��R�(KK��h�C�  8      �t�bhhK ��h��R�(KK	��h�C$(      <      j     k        �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK	��h�C$[   X      l                 �t�bhhK ��h��R�(KK��h�C~            �t�bhhK ��h��R�(KK��h�C	        �t�bhhK ��h��R�(KK��h�C~       
     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK
��h�C(:   |          *      9         �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C       �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C4   8      <    	   '   e     '           �t�bhhK ��h��R�(KK��h�C8   *      '   
  v   �      �   �             �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK	��h�C$[   X      l                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�Cz     �t�bhhK ��h��R�(KK��h�C`   �     m  s  n     8         �     o    	   v         �                �t�bhhK ��h��R�(KK��h�C@             *      9         �   �   Z   p        �t�bhhK ��h��R�(KK��h�C<      
        *      9   7           �        �t�bhhK ��h��R�(KK��h�C         z     �t�bhhK ��h��R�(KK��h�C  �        �t�bhhK ��h��R�(KK��h�C   
   o             �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cq           �t�bhhK ��h��R�(KK��h�Cq     �t�bhhK ��h��R�(KK��h�CW   �     �t�bhhK ��h��R�(KK��h�CP   8           �      F   k   	   t          �      r  �         �t�bhhK ��h��R�(KK��h�CU                 �t�bhhK ��h��R�(KK��h�CT   8   4     $      L   �   �        8   3     $      �   �   �         �t�bhhK ��h��R�(KK��h�C   
              �t�bhhK ��h��R�(KK��h�C   
   .           �t�bhhK ��h��R�(KK��h�C   8   �   V          �t�bhhK ��h��R�(KK��h�C@           �   P  �      �           ]          �t�bhhK ��h��R�(KK��h�C,�       s     C       I         �t�bhhK ��h��R�(KK��h�C8        -               .  �     C         �t�bhhK ��h��R�(KK��h�C!  "           �t�bhhK ��h��R�(KK��h�CPm  s  n  u  s   �   Z   #  $  \   %     #     �   �     t        �t�bhhK ��h��R�(KK��h�C   
   s  &           �t�bhhK ��h��R�(KK��h�C         W   �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cz     �t�bhhK ��h��R�(KK��h�CW   �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8   8      H   �   �   	   �   �      �   l        �t�bhhK ��h��R�(KK	��h�C$�   �     )                  �t�bhhK ��h��R�(KK	��h�C$   8      D   '   �  �         �t�bhhK ��h��R�(KK��h�CD�  
   �     r   $   w  �   n    z   6   f     &        �t�bhhK ��h��R�(KK��h�C@
      �   
   �     �  �  6      �   &   &  `         �t�bhhK ��h��R�(KK��h�C8      D   b  �     T        9     D        �t�bhhK ��h��R�(KK	��h�C$�   �   `      T     D        �t�bhhK ��h��R�(KK��h�CP     �     8      D   g   �     v  $      *   	   9      !         �t�bhhK ��h��R�(KK��h�C,   6   c  �   �   J   `      8         �t�bhhK ��h��R�(KK��h�C             q            �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C �                       �t�bhhK ��h��R�(KK��h�C`   
   d           �t�bhhK ��h��R�(KK��h�C     e  r           �t�bhhK ��h��R�(KK��h�C                   �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C    8   �       U        �t�bhhK ��h��R�(KK��h�C,            f                �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C    
   g                 �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK��h�CX   8      �             �  h     �     �  6        �     �        �t�bhhK ��h��R�(KK��h�C8
      "   �   
   &   [            =   i        �t�bhhK ��h��R�(KK��h�Ci     �t�bhhK ��h��R�(KK��h�C8   A     �t�bhhK ��h��R�(KK��h�C=  =     �t�bhhK ��h��R�(KK��h�C�  8      �t�bhhK ��h��R�(KK	��h�C$(      <      j     k        �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK	��h�C$[   X      l                 �t�bhhK ��h��R�(KK��h�C~            �t�bhhK ��h��R�(KK��h�C	        �t�bhhK ��h��R�(KK��h�C~       
     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK
��h�C(:   |          *      9         �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C       �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C4   8      <    	   '   e     '           �t�bhhK ��h��R�(KK��h�C8   *      '   
  v   �      �   �             �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK	��h�C$[   X      l                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�Cz     �t�bhhK ��h��R�(KK��h�C`   �     m  s  n     8         �     o    	   v         �                �t�bhhK ��h��R�(KK��h�C@             *      9         �   �   Z   p        �t�bhhK ��h��R�(KK��h�C<      
        *      9   7           �        �t�bhhK ��h��R�(KK��h�C         z     �t�bhhK ��h��R�(KK��h�C  �        �t�bhhK ��h��R�(KK��h�C   
   o             �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cq           �t�bhhK ��h��R�(KK��h�Cq     �t�bhhK ��h��R�(KK��h�CW   �     �t�bhhK ��h��R�(KK��h�CP   8           �      F   k   	   t          �      r  �         �t�bhhK ��h��R�(KK��h�CU                 �t�bhhK ��h��R�(KK��h�CT   8   4     $      L   �   �        8   3     $      �   �   �         �t�bhhK ��h��R�(KK��h�C   
              �t�bhhK ��h��R�(KK��h�C   
   .           �t�bhhK ��h��R�(KK��h�C   8   �   V          �t�bhhK ��h��R�(KK��h�C@           �   P  �      �           ]          �t�bhhK ��h��R�(KK��h�C,�       s     C       I         �t�bhhK ��h��R�(KK��h�C8        -               .  �     C         �t�bhhK ��h��R�(KK��h�C!  "           �t�bhhK ��h��R�(KK��h�CPm  s  n  u  s   �   Z   #  $  \   %     #     �   �     t        �t�bhhK ��h��R�(KK��h�C   
   s  &           �t�bhhK ��h��R�(KK��h�C         W   �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cz     �t�bhhK ��h��R�(KK��h�CW   �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8   8      H   �   �   	   �   �      �   l        �t�bhhK ��h��R�(KK	��h�C$�   �     )                  �t�bhhK ��h��R�(KK	��h�C$   8      D   '   �  �         �t�bhhK ��h��R�(KK��h�CD�  
   �     r   $   w  �   n    z   6   f     &        �t�bhhK ��h��R�(KK��h�C@
      �   
   �     �  �  6      �   &   &  `         �t�bhhK ��h��R�(KK��h�C8      D   b  �     T        9     D        �t�bhhK ��h��R�(KK	��h�C$�   �   `      T     D        �t�bhhK ��h��R�(KK��h�CP     �     8      D   g   �     v  $      *   	   9      !         �t�bhhK ��h��R�(KK��h�C,   6   c  �   �   J   `      8         �t�bhhK ��h��R�(KK��h�C             q            �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C �                       �t�bhhK ��h��R�(KK��h�C`   
   d           �t�bhhK ��h��R�(KK��h�C     e  r           �t�bhhK ��h��R�(KK��h�C                   �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C    8   �       U        �t�bhhK ��h��R�(KK��h�C,            f                �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C    
   g                 �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK��h�CX   8      �             �  h     �     �  6        �     �        �t�bhhK ��h��R�(KK��h�C8
      "   �   
   &   [            =   i        �t�bhhK ��h��R�(KK��h�Ci     �t�bhhK ��h��R�(KK��h�C8   A     �t�bhhK ��h��R�(KK��h�C=  =     �t�bhhK ��h��R�(KK��h�C�  8      �t�bhhK ��h��R�(KK	��h�C$(      <      j     k        �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK	��h�C$[   X      l                 �t�bhhK ��h��R�(KK��h�C~            �t�bhhK ��h��R�(KK��h�C	        �t�bhhK ��h��R�(KK��h�C~       
     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK
��h�C(:   |          *      9         �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C       �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C4   8      <    	   '   e     '           �t�bhhK ��h��R�(KK��h�C8   *      '   
  v   �      �   �             �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK	��h�C$[   X      l                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�Cz     �t�bhhK ��h��R�(KK��h�C`   �     m  s  n     8         �     o    	   v         �                �t�bhhK ��h��R�(KK��h�C@             *      9         �   �   Z   p        �t�bhhK ��h��R�(KK��h�C<      
        *      9   7           �        �t�bhhK ��h��R�(KK��h�C         z     �t�bhhK ��h��R�(KK��h�C  �        �t�bhhK ��h��R�(KK��h�C   
   o             �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cq           �t�bhhK ��h��R�(KK��h�Cq     �t�bhhK ��h��R�(KK��h�CW   �     �t�bhhK ��h��R�(KK��h�CP   8           �      F   k   	   t          �      r  �         �t�bhhK ��h��R�(KK��h�CU                 �t�bhhK ��h��R�(KK��h�CT   8   4     $      L   �   �        8   3     $      �   �   �         �t�bhhK ��h��R�(KK��h�C   
              �t�bhhK ��h��R�(KK��h�C   
   .           �t�bhhK ��h��R�(KK��h�C   8   �   V          �t�bhhK ��h��R�(KK��h�C@           �   P  �      �           ]          �t�bhhK ��h��R�(KK��h�C,�       s     C       I         �t�bhhK ��h��R�(KK��h�C8        -               .  �     C         �t�bhhK ��h��R�(KK��h�C!  "           �t�bhhK ��h��R�(KK��h�CPm  s  n  u  s   �   Z   #  $  \   %     #     �   �     t        �t�bhhK ��h��R�(KK��h�C   
   s  &           �t�bhhK ��h��R�(KK��h�C         W   �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�Cj          �t�bhhK ��h��R�(KK��h�Ck     ~     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cu     v     �         �t�bhhK ��h��R�(KK��h�C<H   �      "  B  �       �      �      w        �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C@   7   �       �      �      w  M   '     "        �t�bhhK ��h��R�(KK��h�Cv     !     �t�bhhK ��h��R�(KK��h�Cv     !           �t�bhhK ��h��R�(KK��h�CH   �      �t�bhhK ��h��R�(KK��h�CH
      �   g         H   �   6              x     �         �t�bhhK ��h��R�(KK��h�CL�  O      w     9     8   A  	      W        8   Q   2         �t�bhhK ��h��R�(KK��h�C8   H   2   7      D   �  
   �     �  �         �t�bhhK ��h��R�(KK��h�C  J   `      �        �t�bhhK ��h��R�(KK��h�C�  (     �t�bhhK ��h��R�(KK��h�C)  8      �t�bhhK ��h��R�(KK��h�CH   !                 �t�bhhK ��h��R�(KK��h�C<
                 @      �   M   X  x  y        �t�bhhK ��h��R�(KK��h�Cy        �t�bhhK ��h��R�(KK��h�C �      z                 �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C4   "     Z   �  
   �           �        �t�bhhK ��h��R�(KK��h�C {     8      *  v        �t�bhhK ��h��R�(KK��h�C4   
   �     �   7         j   �           �t�bhhK ��h��R�(KK��h�CL
             �        �        �  	   6      =   W        �t�bhhK ��h��R�(KK��h�CX
        J   �  G  l   p  /      �  /      l   	         =   '   �         �t�bhhK ��h��R�(KK��h�Cz  O     �t�bhhK ��h��R�(KK��h�C0      �   #  �   �   	   l     +        �t�bhhK ��h��R�(KK��h�C,   5   4     r   �  N      �        �t�bhhK ��h��R�(KK��h�CP
              "   ,   �  	         =   �   	  
  !  _   (        �t�bhhK ��h��R�(KK��h�C .   |  "        *         �t�bhhK ��h��R�(KK��h�C:   _   (     �t�bhhK ��h��R�(KK��h�C(   ,     �t�bhhK ��h��R�(KK��h�C+      �     �     �t�bhhK ��h��R�(KK��h�C|     D     �         �t�bhhK ��h��R�(KK��h�C   
   �      -     �t�bhhK ��h��R�(KK��h�C�   	  
        �t�bhhK ��h��R�(KK��h�C :   _   #                 �t�bhhK ��h��R�(KK��h�Cj          �t�bhhK ��h��R�(KK��h�CxY      "   {      D     :   |  }  �   +   	      F   �      Y      .  	      @   w                  �t�bhhK ��h��R�(KK��h�C@   �     4      �     �   �      �        ~        �t�bhhK ��h��R�(KK��h�C@   8           �      
          �      ~        �t�bhhK ��h��R�(KK��h�C8        �t�bhhK ��h��R�(KK��h�C}  V     �t�bhhK ��h��R�(KK��h�C=  /  8      �t�bhhK ��h��R�(KK��h�C(   0     �t�bhhK ��h��R�(KK��h�C         j          �t�bhhK ��h��R�(KK��h�C   
     �           �t�bhhK ��h��R�(KK��h�C    
   �      1           �t�bhhK ��h��R�(KK��h�Ck     &     �t�bhhK ��h��R�(KK��h�C4   j   �   2     &  7         
   3        �t�bhhK ��h��R�(KK��h�C4  5        �t�bhhK ��h��R�(KK��h�C6                 �t�bhhK ��h��R�(KK��h�C7     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�Cj          �t�bhhK ��h��R�(KK��h�Ck     ~     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cu     v     �         �t�bhhK ��h��R�(KK��h�C<H   �      "  B  �       �      �      w        �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C@   7   �       �      �      w  M   '     "        �t�bhhK ��h��R�(KK��h�Cv     !     �t�bhhK ��h��R�(KK��h�Cv     !           �t�bhhK ��h��R�(KK��h�CH   �      �t�bhhK ��h��R�(KK��h�CH
      �   g         H   �   6              x     �         �t�bhhK ��h��R�(KK��h�CL�  O      w     9     8   A  	      W        8   Q   2         �t�bhhK ��h��R�(KK��h�C8   H   2   7      D   �  
   �     �  �         �t�bhhK ��h��R�(KK��h�C  J   `      �        �t�bhhK ��h��R�(KK��h�C�  (     �t�bhhK ��h��R�(KK��h�C)  8      �t�bhhK ��h��R�(KK��h�CH   !                 �t�bhhK ��h��R�(KK��h�C<
                 @      �   M   X  x  y        �t�bhhK ��h��R�(KK��h�Cy        �t�bhhK ��h��R�(KK��h�C �      z                 �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C4   "     Z   �  
   �           �        �t�bhhK ��h��R�(KK��h�C {     8      *  v        �t�bhhK ��h��R�(KK��h�C4   
   �     �   7         j   �           �t�bhhK ��h��R�(KK��h�CL
             �        �        �  	   6      =   W        �t�bhhK ��h��R�(KK��h�CX
        J   �  G  l   p  /      �  /      l   	         =   '   �         �t�bhhK ��h��R�(KK��h�Cz  O     �t�bhhK ��h��R�(KK��h�C0      �   #  �   �   	   l     +        �t�bhhK ��h��R�(KK��h�C,   5   4     r   �  N      �        �t�bhhK ��h��R�(KK��h�CP
              "   ,   �  	         =   �   	  
  !  _   (        �t�bhhK ��h��R�(KK��h�C .   |  "        *         �t�bhhK ��h��R�(KK��h�C:   _   (     �t�bhhK ��h��R�(KK��h�C(   ,     �t�bhhK ��h��R�(KK��h�C+      �     �     �t�bhhK ��h��R�(KK��h�C|     D     �         �t�bhhK ��h��R�(KK��h�C   
   �      -     �t�bhhK ��h��R�(KK��h�C�   	  
        �t�bhhK ��h��R�(KK��h�C :   _   #                 �t�bhhK ��h��R�(KK��h�Cj          �t�bhhK ��h��R�(KK��h�CxY      "   {      D     :   |  }  �   +   	      F   �      Y      .  	      @   w                  �t�bhhK ��h��R�(KK��h�C@   �     4      �     �   �      �        ~        �t�bhhK ��h��R�(KK��h�C@   8           �      
          �      ~        �t�bhhK ��h��R�(KK��h�C8        �t�bhhK ��h��R�(KK��h�C}  V     �t�bhhK ��h��R�(KK��h�C=  /  8      �t�bhhK ��h��R�(KK��h�C(   0     �t�bhhK ��h��R�(KK��h�C         j          �t�bhhK ��h��R�(KK��h�C   
     �           �t�bhhK ��h��R�(KK��h�C    
   �      1           �t�bhhK ��h��R�(KK��h�Ck     &     �t�bhhK ��h��R�(KK��h�C4   j   �   2     &  7         
   3        �t�bhhK ��h��R�(KK��h�C4  5        �t�bhhK ��h��R�(KK��h�C6                 �t�bhhK ��h��R�(KK��h�C7     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�Cj          �t�bhhK ��h��R�(KK��h�Ck     ~     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cu     v     �         �t�bhhK ��h��R�(KK��h�C<H   �      "  B  �       �      �      w        �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C@   7   �       �      �      w  M   '     "        �t�bhhK ��h��R�(KK��h�Cv     !     �t�bhhK ��h��R�(KK��h�Cv     !           �t�bhhK ��h��R�(KK��h�CH   �      �t�bhhK ��h��R�(KK��h�CH
      �   g         H   �   6              x     �         �t�bhhK ��h��R�(KK��h�CL�  O      w     9     8   A  	      W        8   Q   2         �t�bhhK ��h��R�(KK��h�C8   H   2   7      D   �  
   �     �  �         �t�bhhK ��h��R�(KK��h�C  J   `      �        �t�bhhK ��h��R�(KK��h�C�  (     �t�bhhK ��h��R�(KK��h�C)  8      �t�bhhK ��h��R�(KK��h�CH   !                 �t�bhhK ��h��R�(KK��h�C<
                 @      �   M   X  x  y        �t�bhhK ��h��R�(KK��h�Cy        �t�bhhK ��h��R�(KK��h�C �      z                 �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C4   "     Z   �  
   �           �        �t�bhhK ��h��R�(KK��h�C {     8      *  v        �t�bhhK ��h��R�(KK��h�C4   
   �     �   7         j   �           �t�bhhK ��h��R�(KK��h�CL
             �        �        �  	   6      =   W        �t�bhhK ��h��R�(KK��h�CX
        J   �  G  l   p  /      �  /      l   	         =   '   �         �t�bhhK ��h��R�(KK��h�Cz  O     �t�bhhK ��h��R�(KK��h�C0      �   #  �   �   	   l     +        �t�bhhK ��h��R�(KK��h�C,   5   4     r   �  N      �        �t�bhhK ��h��R�(KK��h�CP
              "   ,   �  	         =   �   	  
  !  _   (        �t�bhhK ��h��R�(KK��h�C .   |  "        *         �t�bhhK ��h��R�(KK��h�C:   _   (     �t�bhhK ��h��R�(KK��h�C(   ,     �t�bhhK ��h��R�(KK��h�C+      �     �     �t�bhhK ��h��R�(KK��h�C|     D     �         �t�bhhK ��h��R�(KK��h�C   
   �      -     �t�bhhK ��h��R�(KK��h�C�   	  
        �t�bhhK ��h��R�(KK��h�C :   _   #                 �t�bhhK ��h��R�(KK��h�Cj          �t�bhhK ��h��R�(KK��h�CxY      "   {      D     :   |  }  �   +   	      F   �      Y      .  	      @   w                  �t�bhhK ��h��R�(KK��h�C@   �     4      �     �   �      �        ~        �t�bhhK ��h��R�(KK��h�C@   8           �      
          �      ~        �t�bhhK ��h��R�(KK��h�C8        �t�bhhK ��h��R�(KK��h�C}  V     �t�bhhK ��h��R�(KK��h�C=  /  8      �t�bhhK ��h��R�(KK��h�C(   0     �t�bhhK ��h��R�(KK��h�C         j          �t�bhhK ��h��R�(KK��h�C   
     �           �t�bhhK ��h��R�(KK��h�C    
   �      1           �t�bhhK ��h��R�(KK��h�Ck     &     �t�bhhK ��h��R�(KK��h�C4   j   �   2     &  7         
   3        �t�bhhK ��h��R�(KK��h�C4  5        �t�bhhK ��h��R�(KK��h�C6                 �t�bhhK ��h��R�(KK��h�C7     �t�bhhK ��h��R�(KK��h�C~     �t�bhhK ��h��R�(KK��h�C\   +      q           g      Y  �     )      9   	   !   	   *      8         �t�bhhK ��h��R�(KK��h�C,   q      D      
   �               �t�bhhK ��h��R�(KK��h�C,�      )         �           E      �t�bhhK ��h��R�(KK��h�C4   8   �   �      )            8           �t�bhhK ��h��R�(KK��h�C8      �   /      8  �   �   ]      M   "        �t�bhhK ��h��R�(KK��h�CU                 �t�bhhK ��h��R�(KK	��h�C$         R     )            �t�bhhK ��h��R�(KK��h�C   �      1         �t�bhhK ��h��R�(KK��h�C�     )      �t�bhhK ��h��R�(KK��h�Cp   
   9  :     W   )   ;  7         j   '  V        �      *      V        �      9         �t�bhhK ��h��R�(KK��h�C'  �     �t�bhhK ��h��R�(KK��h�CD      �   '  �     )            F      *      9         �t�bhhK ��h��R�(KK��h�CP   <  2         �     ,        �  u      N         �   	        �t�bhhK ��h��R�(KK	��h�C$         �  �     �        �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C�  =                 �t�bhhK ��h��R�(KK��h�C~     �t�bhhK ��h��R�(KK��h�C\   +      q           g      Y  �     )      9   	   !   	   *      8         �t�bhhK ��h��R�(KK��h�C,   q      D      
   �               �t�bhhK ��h��R�(KK��h�C,�      )         �           E      �t�bhhK ��h��R�(KK��h�C4   8   �   �      )            8           �t�bhhK ��h��R�(KK��h�C8      �   /      8  �   �   ]      M   "        �t�bhhK ��h��R�(KK��h�CU                 �t�bhhK ��h��R�(KK	��h�C$         R     )            �t�bhhK ��h��R�(KK��h�C   �      1         �t�bhhK ��h��R�(KK��h�C�     )      �t�bhhK ��h��R�(KK��h�Cp   
   9  :     W   )   ;  7         j   '  V        �      *      V        �      9         �t�bhhK ��h��R�(KK��h�C'  �     �t�bhhK ��h��R�(KK��h�CD      �   '  �     )            F      *      9         �t�bhhK ��h��R�(KK��h�CP   <  2         �     ,        �  u      N         �   	        �t�bhhK ��h��R�(KK	��h�C$         �  �     �        �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C�  =                 �t�bhhK ��h��R�(KK��h�C~     �t�bhhK ��h��R�(KK��h�C\   +      q           g      Y  �     )      9   	   !   	   *      8         �t�bhhK ��h��R�(KK��h�C,   q      D      
   �               �t�bhhK ��h��R�(KK��h�C,�      )         �           E      �t�bhhK ��h��R�(KK��h�C4   8   �   �      )            8           �t�bhhK ��h��R�(KK��h�C8      �   /      8  �   �   ]      M   "        �t�bhhK ��h��R�(KK��h�CU                 �t�bhhK ��h��R�(KK	��h�C$         R     )            �t�bhhK ��h��R�(KK��h�C   �      1         �t�bhhK ��h��R�(KK��h�C�     )      �t�bhhK ��h��R�(KK��h�Cp   
   9  :     W   )   ;  7         j   '  V        �      *      V        �      9         �t�bhhK ��h��R�(KK��h�C'  �     �t�bhhK ��h��R�(KK��h�CD      �   '  �     )            F      *      9         �t�bhhK ��h��R�(KK��h�CP   <  2         �     ,        �  u      N         �   	        �t�bhhK ��h��R�(KK	��h�C$         �  �     �        �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C�  =                 �t�bhhK ��h��R�(KK��h�Cu   7   F  �   h      �t�bhhK ��h��R�(KK��h�C    �  '   �      �t�bhhK ��h��R�(KK��h�CG     �t�bhhK ��h��R�(KK��h�Cu   7   F  �   h      �t�bhhK ��h��R�(KK��h�C4~   �      +  x   |      8       g   �         �t�bhhK ��h��R�(KK��h�C &   |  �         *         �t�bhhK ��h��R�(KK��h�C~   �      +  	   *      �t�bhhK ��h��R�(KK	��h�C$         �      �     *      �t�bhhK ��h��R�(KK��h�CD   
   �        ;   7         j   �   �       �        �t�bhhK ��h��R�(KK��h�C@   
   �     1   7         j   �   �  7   F  �   h      �t�bhhK ��h��R�(KK��h�C<>  T   ?  �      9   	   !   	   *      8   @        �t�bhhK ��h��R�(KK��h�C0A        F        	   �      �         �t�bhhK ��h��R�(KK��h�C)     B           �t�bhhK ��h��R�(KK��h�C*  �                 �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C8   
       i   
   �  7         j   �   �        �t�bhhK ��h��R�(KK��h�C    �  '   �      �t�bhhK ��h��R�(KK��h�CP   j   �     �  '   �   7         
   �  B   C  '   �      1         �t�bhhK ��h��R�(KK��h�CTD  /      :     �      S  �     �     *      �     �     9         �t�bhhK ��h��R�(KK��h�Cd
         �        �  �     �  �  8   �  �     T   �  �  X   	   �     c         �t�bhhK ��h��R�(KK��h�C      E     �t�bhhK ��h��R�(KK��h�CG     �t�bhhK ��h��R�(KK��h�C0�  !  �      �  �     �     9         �t�bhhK ��h��R�(KK��h�C5        �t�bhhK ��h��R�(KK��h�C �      F                 �t�bhhK ��h��R�(KK��h�CL      -   �     �  �  1            9          �   
   �        �t�bhhK ��h��R�(KK��h�CP  �   C      U     1          0     �      �  G     (  Z        �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C�     G     �t�bhhK ��h��R�(KK��h�Cu   7   F  �   h      �t�bhhK ��h��R�(KK��h�C    �  '   �      �t�bhhK ��h��R�(KK��h�CG     �t�bhhK ��h��R�(KK��h�Cu   7   F  �   h      �t�bhhK ��h��R�(KK��h�C4~   �      +  x   |      8       g   �         �t�bhhK ��h��R�(KK��h�C &   |  �         *         �t�bhhK ��h��R�(KK��h�C~   �      +  	   *      �t�bhhK ��h��R�(KK	��h�C$         �      �     *      �t�bhhK ��h��R�(KK��h�CD   
   �        ;   7         j   �   �       �        �t�bhhK ��h��R�(KK��h�C@   
   �     1   7         j   �   �  7   F  �   h      �t�bhhK ��h��R�(KK��h�C<>  T   ?  �      9   	   !   	   *      8   @        �t�bhhK ��h��R�(KK��h�C0A        F        	   �      �         �t�bhhK ��h��R�(KK��h�C)     B           �t�bhhK ��h��R�(KK��h�C*  �                 �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C8   
       i   
   �  7         j   �   �        �t�bhhK ��h��R�(KK��h�C    �  '   �      �t�bhhK ��h��R�(KK��h�CP   j   �     �  '   �   7         
   �  B   C  '   �      1         �t�bhhK ��h��R�(KK��h�CTD  /      :     �      S  �     �     *      �     �     9         �t�bhhK ��h��R�(KK��h�Cd
         �        �  �     �  �  8   �  �     T   �  �  X   	   �     c         �t�bhhK ��h��R�(KK��h�C      E     �t�bhhK ��h��R�(KK��h�CG     �t�bhhK ��h��R�(KK��h�C0�  !  �      �  �     �     9         �t�bhhK ��h��R�(KK��h�C5        �t�bhhK ��h��R�(KK��h�C �      F                 �t�bhhK ��h��R�(KK��h�C0C      -   9  �        <  =  0        �t�bhhK ��h��R�(KK��h�Cd     x   2     �  �  C      U     1          0     �      �  G     (  Z        �t�bhhK ��h��R�(KK��h�C�     G     �t�bhhK ��h��R�(KK��h�Cu   7   F  �   h      �t�bhhK ��h��R�(KK��h�C    �  '   �      �t�bhhK ��h��R�(KK��h�CG     �t�bhhK ��h��R�(KK��h�Cu   7   F  �   h      �t�bhhK ��h��R�(KK��h�C4~   �      +  x   |      8       g   �         �t�bhhK ��h��R�(KK��h�C &   |  �         *         �t�bhhK ��h��R�(KK��h�C~   �      +  	   *      �t�bhhK ��h��R�(KK	��h�C$         �      �     *      �t�bhhK ��h��R�(KK��h�CD   
   �        ;   7         j   �   �       �        �t�bhhK ��h��R�(KK��h�C@   
   �     1   7         j   �   �  7   F  �   h      �t�bhhK ��h��R�(KK��h�C<>  T   ?  �      9   	   !   	   *      8   @        �t�bhhK ��h��R�(KK��h�C0A        F        	   �      �         �t�bhhK ��h��R�(KK��h�C )     B                 �t�bhhK ��h��R�(KK��h�C*  �                 �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C8   
       i   
   �  7         j   �   �        �t�bhhK ��h��R�(KK��h�C    �  '   �      �t�bhhK ��h��R�(KK��h�CP   j   �     �  '   �   7         
   �  B   C  '   �      1         �t�bhhK ��h��R�(KK��h�CTD  /      :     �      S  �     �     *      �     �     9         �t�bhhK ��h��R�(KK��h�Cd
         �        �  �     �  �  8   �  �     T   �  �  X   	   �     c         �t�bhhK ��h��R�(KK��h�C      E     �t�bhhK ��h��R�(KK��h�CG     �t�bhhK ��h��R�(KK��h�C0�  !  �      �  �     �     9         �t�bhhK ��h��R�(KK��h�C5        �t�bhhK ��h��R�(KK��h�C �      F                 �t�bhhK ��h��R�(KK��h�C0C      -   9  �        <  =  0        �t�bhhK ��h��R�(KK��h�Cd     x   2     �  �  C      U     1          0     �      �  G     (  Z        �t�bhhK ��h��R�(KK��h�C,4  �   �     /           1         �t�bhhK ��h��R�(KK��h�C�     G     �t�bhhK ��h��R�(KK��h�Cc         $     C      �t�bhhK ��h��R�(KK��h�C�   �      �     �t�bhhK ��h��R�(KK��h�C5         �   h      �t�bhhK ��h��R�(KK��h�Cc         $     C      �t�bhhK ��h��R�(KK��h�Cl
      "   �   
   �      8            =   H   �  M             �  H     �     I        �t�bhhK ��h��R�(KK��h�C,      �     )   	                  �t�bhhK ��h��R�(KK��h�CD9   Q   c      C   	   9      ;  	   �      C      �         �t�bhhK ��h��R�(KK��h�C 9      ?                 �t�bhhK ��h��R�(KK��h�Cp
      "   �     �   �  	            <  =  0     4     @   c      �     '                �t�bhhK ��h��R�(KK��h�C,4  �   �     /           1         �t�bhhK ��h��R�(KK��h�C�   �      �     �t�bhhK ��h��R�(KK ��h�C�?        J     �           S      �      �        �   �         �                 K  /              �t�bhhK ��h��R�(KK��h�C�      w        �t�bhhK ��h��R�(KK��h�C �      L     M           �t�bhhK ��h��R�(KK��h�CL
      4      N  d   �        �  &   �   �     )     W        �t�bhhK ��h��R�(KK��h�C�      W        �t�bhhK ��h��R�(KK��h�C}  V     �t�bhhK ��h��R�(KK��h�C=  �     �t�bhhK ��h��R�(KK��h�C�  8      �t�bhhK ��h��R�(KK��h�C(      <      j     �t�bhhK ��h��R�(KK��h�CO           �t�bhhK ��h��R�(KK��h�C5         �   h      �t�bhhK ��h��R�(KK��h�CP
      4      )               �     �   N      2  �      {        �t�bhhK ��h��R�(KK��h�CH      �     �   N      a  
      �       �  �  %        �t�bhhK ��h��R�(KK��h�C,   �  �  O         �   M           �t�bhhK ��h��R�(KK��h�C �      P  �     /         �t�bhhK ��h��R�(KK	��h�C$         5         �   h      �t�bhhK ��h��R�(KK��h�C�   �     �        �t�bhhK ��h��R�(KK	��h�C$�  �      �                 �t�bhhK ��h��R�(KK��h�Cc         $     C      �t�bhhK ��h��R�(KK��h�C�   �      �     �t�bhhK ��h��R�(KK��h�C5         �   h      �t�bhhK ��h��R�(KK��h�Cc         $     C      �t�bhhK ��h��R�(KK��h�Cl
      "   �   
   �      8            =   H   �  M             �  H     �     I        �t�bhhK ��h��R�(KK��h�C,      �     )   	                  �t�bhhK ��h��R�(KK��h�CD9   Q   c      C   	   9      ;  	   �      C      �         �t�bhhK ��h��R�(KK��h�C 9      ?                 �t�bhhK ��h��R�(KK��h�Cp
      "   �     �   �  	            <  =  0     4     @   c      �     '                �t�bhhK ��h��R�(KK��h�C,4  �   �     /           1         �t�bhhK ��h��R�(KK��h�C�   �      �     �t�bhhK ��h��R�(KK ��h�C�?        J     �           S      �      �        �   �         �                 K  /              �t�bhhK ��h��R�(KK��h�C�      w        �t�bhhK ��h��R�(KK��h�C �      L     M           �t�bhhK ��h��R�(KK��h�CL
      4      N  d   �        �  &   �   �     )     W        �t�bhhK ��h��R�(KK��h�C�      W        �t�bhhK ��h��R�(KK��h�C}  V     �t�bhhK ��h��R�(KK��h�C=  �     �t�bhhK ��h��R�(KK��h�C�  8      �t�bhhK ��h��R�(KK��h�C(      <      j     �t�bhhK ��h��R�(KK��h�CO           �t�bhhK ��h��R�(KK��h�C5         �   h      �t�bhhK ��h��R�(KK��h�CP
      4      )               �     �   N      2  �      {        �t�bhhK ��h��R�(KK��h�CH      �     �   N      a  
      �       �  �  %        �t�bhhK ��h��R�(KK��h�C,   �  �  O         �   M           �t�bhhK ��h��R�(KK��h�C �      P  �     /         �t�bhhK ��h��R�(KK	��h�C$         5         �   h      �t�bhhK ��h��R�(KK��h�C�   �     �        �t�bhhK ��h��R�(KK	��h�C$�  �      �                 �t�bhhK ��h��R�(KK��h�Cc         $     C      �t�bhhK ��h��R�(KK��h�C�   �      �     �t�bhhK ��h��R�(KK��h�C5         �   h      �t�bhhK ��h��R�(KK��h�Cc         $     C      �t�bhhK ��h��R�(KK��h�Cl
      "   �   
   �      8            =   H   �  M             �  H     �     I        �t�bhhK ��h��R�(KK��h�C,      �     )   	                  �t�bhhK ��h��R�(KK��h�CD9   Q   c      C   	   9      ;  	   �      C      �         �t�bhhK ��h��R�(KK��h�C 9      ?                 �t�bhhK ��h��R�(KK��h�Cp
      "   �     �   �  	            <  =  0     4     @   c      �     '                �t�bhhK ��h��R�(KK��h�C,4  �   �     /           1         �t�bhhK ��h��R�(KK��h�C�   �      �     �t�bhhK ��h��R�(KK ��h�C�?        J     �           S      �      �        �   �         �                 K  /              �t�bhhK ��h��R�(KK��h�C�      w        �t�bhhK ��h��R�(KK��h�C �      L     M           �t�bhhK ��h��R�(KK��h�CL
      4      N  d   �        �  &   �   �     )     W        �t�bhhK ��h��R�(KK��h�C�      W        �t�bhhK ��h��R�(KK��h�C}  V     �t�bhhK ��h��R�(KK��h�C=  �     �t�bhhK ��h��R�(KK��h�C�  8      �t�bhhK ��h��R�(KK��h�C(      <      j     �t�bhhK ��h��R�(KK��h�CO           �t�bhhK ��h��R�(KK��h�C5         �   h      �t�bhhK ��h��R�(KK��h�CP
      4      )               �     �   N      2  �      {        �t�bhhK ��h��R�(KK��h�CH      �     �   N      a  
      �       �  �  %        �t�bhhK ��h��R�(KK��h�C,   �  �  O         �   M           �t�bhhK ��h��R�(KK��h�C �      P  �     /         �t�bhhK ��h��R�(KK	��h�C$         5         �   h      �t�bhhK ��h��R�(KK��h�C�   �     �        �t�bhhK ��h��R�(KK	��h�C$�  �      �                 �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CH   �  �     9         i   
   {      I  m     �  ,        �t�bhhK ��h��R�(KK��h�C�      }      �        �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C'  �                 �t�bhhK ��h��R�(KK��h�CP      D   i   
   Z   �  {      m          "     q   �  1         �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C'  �                 �t�bhhK ��h��R�(KK��h�C          �     1         �t�bhhK ��h��R�(KK��h�C     |      �t�bhhK ��h��R�(KK��h�CL
        r   �  �      8   	   6      I  /      |      ]        �t�bhhK ��h��R�(KK��h�C4      I  /      9   �     �      �        �t�bhhK ��h��R�(KK��h�C9   �     �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�C,N      �     �   6      w      /      �t�bhhK ��h��R�(KK��h�C[        F   �        �t�bhhK ��h��R�(KK��h�C0{      *     
      5   {      1         �t�bhhK ��h��R�(KK��h�C0+  ;  �     
         m     �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C  n   -        �t�bhhK ��h��R�(KK��h�C<3      4  �  6   �  .  \        )               �t�bhhK ��h��R�(KK��h�C              |      �t�bhhK ��h��R�(KK��h�CS     1      �t�bhhK ��h��R�(KK��h�C      �                 �t�bhhK ��h��R�(KK��h�C,4  �   �     /           1         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CH   �  �     9         i   
   {      I  m     �  ,        �t�bhhK ��h��R�(KK��h�C�      }      �        �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C'  �                 �t�bhhK ��h��R�(KK��h�CP      D   i   
   Z   �  {      m          "     q   �  1         �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C'  �                 �t�bhhK ��h��R�(KK��h�C          �     1         �t�bhhK ��h��R�(KK��h�C     |      �t�bhhK ��h��R�(KK��h�CL
        r   �  �      8   	   6      I  /      |      ]        �t�bhhK ��h��R�(KK��h�C4      I  /      9   �     �      �        �t�bhhK ��h��R�(KK��h�C9   �     �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�C,N      �     �   6      w      /      �t�bhhK ��h��R�(KK��h�C[        F   �        �t�bhhK ��h��R�(KK��h�C0{      *     
      5   {      1         �t�bhhK ��h��R�(KK��h�C0+  ;  �     
         m     �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C  n   -        �t�bhhK ��h��R�(KK��h�C<3      4  �  6   �  .  \        )               �t�bhhK ��h��R�(KK��h�C              |      �t�bhhK ��h��R�(KK��h�CS     1      �t�bhhK ��h��R�(KK��h�C      �                 �t�bhhK ��h��R�(KK��h�C,4  �   �     /           1         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CH   �  �     9         i   
   {      I  m     �  ,        �t�bhhK ��h��R�(KK��h�C�      }      �        �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C'  �                 �t�bhhK ��h��R�(KK��h�CP      D   i   
   Z   �  {      m          "     q   �  1         �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C'  �                 �t�bhhK ��h��R�(KK��h�C          �     1         �t�bhhK ��h��R�(KK��h�C     |      �t�bhhK ��h��R�(KK��h�CL
        r   �  �      8   	   6      I  /      |      ]        �t�bhhK ��h��R�(KK��h�C4      I  /      9   �     �      �        �t�bhhK ��h��R�(KK��h�C9   �     �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�C,N      �     �   6      w      /      �t�bhhK ��h��R�(KK��h�C[        F   �        �t�bhhK ��h��R�(KK��h�C0{      *     
      5   {      1         �t�bhhK ��h��R�(KK��h�C0+  ;  �     
         m     �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C  n   -        �t�bhhK ��h��R�(KK��h�C<3      4  �  6   �  .  \        )               �t�bhhK ��h��R�(KK��h�C              |      �t�bhhK ��h��R�(KK��h�CS     1      �t�bhhK ��h��R�(KK��h�C      �                 �t�bhhK ��h��R�(KK��h�C,4  �   �     /           1         �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CJ     �t�bhhK ��h��R�(KK	��h�C$!      �  �   "   R          �t�bhhK ��h��R�(KK
��h�C(�  Q     R  S     ^   T        �t�bhhK ��h��R�(KK��h�C   �      ^   >        �t�bhhK ��h��R�(KK��h�Cd!   �  �  X  �      �        �  �  U  V     �        	      �   J     �         �t�bhhK ��h��R�(KK	��h�C$      7         �  2         �t�bhhK ��h��R�(KK��h�C4      g      
   �     !     �           �t�bhhK ��h��R�(KK��h�C<q   p   /   "     >     U   '   x     '   e         �t�bhhK ��h��R�(KK��h�C,   J        �     9     &        �t�bhhK ��h��R�(KK
��h�C(   :  �      �   @     �        �t�bhhK ��h��R�(KK��h�C@      -   �      B     <        C        �        �t�bhh�       K ��h��R�(KK��h�C ?                 E      �t�bhhK ��h��R�(KK��h�C&     �t�bhhK ��h��R�(KK��h�C8   '   &     W     X     "  B     9        �t�bhhK ��h��R�(KK��h�C<;  V     Y  �  	   :  	   Z  	   [     \        �t�bhhK ��h��R�(KK��h�C.      <  �  &        �t�bhhK ��h��R�(KK	��h�C$.      .   ]  ^      �        �t�bhhK ��h��R�(KK��h�C4'   _     `  a        b     ^   Y         �t�bhhK ��h��R�(KK��h�C\     c  /   '   \  �  6      I  /      |             �   �     �        �t�bhhK ��h��R�(KK��h�CD      �   &     �  �     d        �     e           �t�bhhK ��h��R�(KK��h�C:      �     �         �t�bhhK ��h��R�(KK	��h�C$\  &        �      f        �t�bhhK ��h��R�(KK��h�C0w      /   �  
      6   �   \  &        �t�bhhK ��h��R�(KK��h�C@
      "   )   �        -   �   \  &     �  2         �t�bhhK ��h��R�(KK��h�CT      �     ;  N      g  �     �     h        �     i           �t�bhhK ��h��R�(KK��h�C,   �  �  }         F      j        �t�bhhK ��h��R�(KK��h�C�  �  k        �t�bhhK ��h��R�(KK��h�C<
      �  J  O  l            �  �     �        �t�bhhK ��h��R�(KK��h�CD      �  ;       �     &     m  n        a        �t�bhhK ��h��R�(KK	��h�C$   7            �  2         �t�bhhK ��h��R�(KK��h�C `   
   o                 �t�bhhK ��h��R�(KK
��h�C(      f      �                 �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK��h�C         ]     �t�bhhK ��h��R�(KK��h�CX
      �        ]     !         g      Y  �     �     �     �        �t�bhhK ��h��R�(KK��h�C4   p     q     !         b     ^        �t�bhhK ��h��R�(KK��h�C�     R        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK
��h�C(9      !   ~  >  �      !         �t�bhhK ��h��R�(KK��h�C8  "   R       F      �  	   r     �        �t�bhhK ��h��R�(KK��h�C8      �  �     Z   �     �  �     J        �t�bhhK ��h��R�(KK��h�C0s     �     �  7      t     �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK
��h�C($                 E      �     �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C,   !   E  �      �     u           �t�bhhK ��h��R�(KK��h�C0   �  F  v  G     H  >   �  {        �t�bhhK ��h��R�(KK��h�C0I  �  u   �  I   2  �     w           �t�bhhK ��h��R�(KK��h�C@     !      �  �     �     �      Z   >   �        �t�bhhK ��h��R�(KK��h�C<   x        y  z  �     @         
   �        �t�bhhK ��h��R�(KK��h�C\   !         �     �  �      {  |        }  ~       �      �  C         �t�bhhK ��h��R�(KK��h�C          !   Q   2         �t�bhhK ��h��R�(KK��h�CP   !      Z   �  �   	   �     W   �   M   _     D      �  �        �t�bhhK ��h��R�(KK��h�C,      
   �  7         �  �        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�      J     �t�bhhK ��h��R�(KK��h�C�  �     �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     �  �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C,Z     S     ?     !      9         �t�bhhK ��h��R�(KK��h�C@M   q   �  �        g      g  .     K     L        �t�bhhK ��h��R�(KK��h�CD&   �      �   �  "   �  �  �        �  �     !         �t�bhhK ��h��R�(KK	��h�C$         !   �   �  2         �t�bhhK ��h��R�(KK��h�C    �        �  �        �t�bhhK ��h��R�(KK��h�CL      
   �     &   �   �     !   7         9   �   �  2         �t�bhhK ��h��R�(KK
��h�C(         T     �     1         �t�bhhK ��h��R�(KK��h�C%   �   �        �t�bhhK ��h��R�(KK��h�C�      �   O     �t�bhhK ��h��R�(KK��h�C�   �   �        �t�bhhK ��h��R�(KK��h�C�   N     E      �t�bhhK ��h��R�(KK��h�C  M           �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK��h�C,!            :   �        �         �t�bhhK ��h��R�(KK��h�C &   �   �  *      9         �t�bhhK ��h��R�(KK��h�C!   I  �      �        �t�bhhK ��h��R�(KK��h�Cp_     .   W   �  �     !   	      F   �  	   �     �  	   �  	   �  	   �  	   �     �        �t�bhhK ��h��R�(KK��h�C!   "   �  �  |         �t�bhhK ��h��R�(KK��h�CP   #       �  �  �     �  �  "   �   e   f  B  )               �t�bhhK ��h��R�(KK��h�C<�       �  �  	   @      �  �     �        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C[   �                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C !   �  "   �  �  �        �t�bhhK ��h��R�(KK��h�C4B   "   �  y     �  I   �  �  g  �        �t�bhhK ��h��R�(KK��h�C8�  !   "   �     '   �     �  u   9   �        �t�bhhK ��h��R�(KK��h�C09   �    �  a   �     �     Z        �t�bhhK ��h��R�(KK��h�CT9   �  �   �  9   �  	   `  !   ,  I   P        �  !      I   �        �t�bhhK ��h��R�(KK��h�C4�     �     �  9   "   �  �     !         �t�bhhK ��h��R�(KK��h�C`�  �  	   �  �  U      M   9      �     �  �  :  U   9   	   "   �  2  !         �t�bhhK ��h��R�(KK��h�C4�     �     �  "   .   �  �     �        �t�bhhK ��h��R�(KK	��h�C$!      B  �     K  �        �t�bhhK ��h��R�(KK��h�C,   F   �   9      !   >     !         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CJ     �t�bhhK ��h��R�(KK	��h�C$!      �  �   "   R          �t�bhhK ��h��R�(KK
��h�C(�  Q     R  S     ^   T        �t�bhhK ��h��R�(KK��h�C   �      ^   >        �t�bhhK ��h��R�(KK��h�Cd!   �  �  X  �      �        �  �  U  V     �        	      �   J     �         �t�bhhK ��h��R�(KK	��h�C$      7         �  2         �t�bhhK ��h��R�(KK��h�C4      g      
   �     !     �           �t�bhhK ��h��R�(KK��h�C<q   p   /   "     >     U   '   x     '   e         �t�bhhK ��h��R�(KK��h�C,   J        �     9     &        �t�bhhK ��h��R�(KK
��h�C(   :  �      �   @     �        �t�bhhK ��h��R�(KK��h�C@      -   �      B     <        C        �        �t�bhhK ��h��R�(KK��h�C ?                 E      �t�bhhK ��h��R�(KK��h�C&     �t�bhhK ��h��R�(KK��h�C8   '   &     W     X     "  B     9        �t�bhhK ��h��R�(KK��h�C<;  V     Y  �  	   :  	   Z  	   [     \        �t�bhhK ��h��R�(KK��h�C.      <  �  &        �t�bhhK ��h��R�(KK	��h�C$.      .   ]  ^      �        �t�bhhK ��h��R�(KK��h�C4'   _     `  a        b     ^   Y         �t�bhhK ��h��R�(KK��h�C\     c  /   '   \  �  6      I  /      |             �   �     �        �t�bhhK ��h��R�(KK��h�CD      �   &     �  �     d        �     e           �t�bhhK ��h��R�(KK��h�C:      �     �         �t�bhhK ��h��R�(KK	��h�C$\  &        �      f        �t�bhhK ��h��R�(KK��h�C0w      /   �  
      6   �   \  &        �t�bhhK ��h��R�(KK��h�C@
      "   )   �        -   �   \  &     �  2         �t�bhhK ��h��R�(KK��h�CT      �     ;  N      g  �     �     h        �     i           �t�bhhK ��h��R�(KK��h�C,   �  �  }         F      j        �t�bhhK ��h��R�(KK��h�C�  �  k        �t�bhhK ��h��R�(KK��h�C<
      �  J  O  l            �  �     �        �t�bhhK ��h��R�(KK��h�CD      �  ;       �     &     m  n        a        �t�bhhK ��h��R�(KK	��h�C$   7            �  2         �t�bhhK ��h��R�(KK��h�C `   
   o                 �t�bhhK ��h��R�(KK
��h�C(      f      �                 �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK��h�C         ]     �t�bhhK ��h��R�(KK��h�CX
      �        ]     !         g      Y  �     �     �     �        �t�bhhK ��h��R�(KK��h�C4   p     q     !         b     ^        �t�bhhK ��h��R�(KK��h�C�     R        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK
��h�C(9      !   ~  >  �      !         �t�bhhK ��h��R�(KK��h�C8  "   R       F      �  	   r     �        �t�bhhK ��h��R�(KK��h�C8      �  �     Z   �     �  �     J        �t�bhhK ��h��R�(KK��h�C0s     �     �  7      t     �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK
��h�C($                 E      �     �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C,   !   E  �      �     u           �t�bhhK ��h��R�(KK��h�C0   �  F  v  G     H  >   �  {        �t�bhhK ��h��R�(KK��h�C0I  �  u   �  I   2  �     w           �t�bhhK ��h��R�(KK��h�C@     !      �  �     �     �      Z   >   �        �t�bhhK ��h��R�(KK��h�C<   x        y  z  �     @         
   �        �t�bhhK ��h��R�(KK��h�C\   !         �     �  �      {  |        }  ~       �      �  C         �t�bhhK ��h��R�(KK��h�C          !   Q   2         �t�bhhK ��h��R�(KK��h�CP   !      Z   �  �   	   �     W   �   M   _     D      �  �        �t�bhhK ��h��R�(KK��h�C,      
   �  7         �  �        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�      J     �t�bhhK ��h��R�(KK��h�C�  �     �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     �  �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C,Z     S     ?     !      9         �t�bhhK ��h��R�(KK��h�C@M   q   �  �        g      g  .     K     L        �t�bhhK ��h��R�(KK��h�CD&   �      �   �  "   �  �  �        �  �     !         �t�bhhK ��h��R�(KK	��h�C$         !   �   �  2         �t�bhhK ��h��R�(KK��h�C    �        �  �        �t�bhhK ��h��R�(KK��h�CL      
   �     &   �   �     !   7         9   �   �  2         �t�bhhK ��h��R�(KK
��h�C(         T     �     1         �t�bhhK ��h��R�(KK��h�C%   �   �        �t�bhhK ��h��R�(KK��h�C�      �   O     �t�bhhK ��h��R�(KK��h�C�   �   �        �t�bhhK ��h��R�(KK��h�C�   N     E      �t�bhhK ��h��R�(KK��h�C  M           �t�be(hhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK��h�C,!            :   �        �         �t�bhhK ��h��R�(KK��h�C &   �   �  *      9         �t�bhhK ��h��R�(KK��h�C!   I  �      �        �t�bhhK ��h��R�(KK��h�Cp_     .   W   �  �     !   	      F   �  	   �     �  	   �  	   �  	   �  	   �     �        �t�bhhK ��h��R�(KK��h�C!   "   �  �  |         �t�bhhK ��h��R�(KK��h�CP   #       �  �  �     �  �  "   �   e   f  B  )               �t�bhhK ��h��R�(KK��h�C<�       �  �  	   @      �  �     �        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C[   �                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C !   �  "   �  �  �        �t�bhhK ��h��R�(KK��h�C4B   "   �  y     �  I   �  �  g  �        �t�bhhK ��h��R�(KK��h�C8�  !   "   �     '   �     �  u   9   �        �t�bhhK ��h��R�(KK��h�C09   �    �  a   �     �     Z        �t�bhhK ��h��R�(KK��h�CT9   �  �   �  9   �  	   `  !   ,  I   P        �  !      I   �        �t�bhhK ��h��R�(KK��h�C4�     �     �  9   "   �  �     !         �t�bhhK ��h��R�(KK��h�C`�  �  	   �  �  U      M   9      �     �  �  :  U   9   	   "   �  2  !         �t�bhhK ��h��R�(KK��h�C4�     �     �  "   .   �  �     �        �t�bhhK ��h��R�(KK	��h�C$!      B  �     K  �        �t�bhhK ��h��R�(KK��h�C,   F   �   9      !   >     !         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CJ     �t�bhhK ��h��R�(KK	��h�C$!      �  �   "   R          �t�bhhK ��h��R�(KK
��h�C(�  Q     R  S     ^   T        �t�bhhK ��h��R�(KK��h�C   �      ^   >        �t�bhhK ��h��R�(KK��h�Cd!   �  �  X  �      �        �  �  U  V     �        	      �   J     �         �t�bhhK ��h��R�(KK	��h�C$      7         �  2         �t�bhhK ��h��R�(KK��h�C4      g      
   �     !     �           �t�bhhK ��h��R�(KK��h�C<q   p   /   "     >     U   '   x     '   e         �t�bhhK ��h��R�(KK��h�C,   J        �     9     &        �t�bhhK ��h��R�(KK
��h�C(   :  �      �   @     �        �t�bhhK ��h��R�(KK��h�C@      -   �      B     <        C        �        �t�bhhK ��h��R�(KK��h�C?                 �t�bhhK ��h��R�(KK��h�C&     �t�bhhK ��h��R�(KK��h�C8   '   &     W     X     "  B     9        �t�bhhK ��h��R�(KK��h�C<;  V     Y  �  	   :  	   Z  	   [     \        �t�bhhK ��h��R�(KK��h�C.      <  �  &        �t�bhhK ��h��R�(KK	��h�C$.      .   ]  ^      �        �t�bhhK ��h��R�(KK��h�C4'   _     `  a        b     ^   Y         �t�bhhK ��h��R�(KK��h�C\     c  /   '   \  �  6      I  /      |             �   �     �        �t�bhhK ��h��R�(KK��h�CD      �   &     �  �     d        �     e           �t�bhhK ��h��R�(KK��h�C:      �     �         �t�bhhK ��h��R�(KK	��h�C$\  &        �      f        �t�bhhK ��h��R�(KK��h�C0w      /   �  
      6   �   \  &        �t�bhhK ��h��R�(KK��h�C@
      "   )   �        -   �   \  &     �  2         �t�bhhK ��h��R�(KK��h�CT      �     ;  N      g  �     �     h        �     i           �t�bhhK ��h��R�(KK��h�C,   �  �  }         F      j        �t�bhhK ��h��R�(KK��h�C�  �  k        �t�bhhK ��h��R�(KK��h�C<
      �  J  O  l            �  �     �        �t�bhhK ��h��R�(KK��h�CD      �  ;       �     &     m  n        a        �t�bhhK ��h��R�(KK	��h�C$   7            �  2         �t�bhhK ��h��R�(KK��h�C `   
   o                 �t�bhhK ��h��R�(KK
��h�C(      f      �                 �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK��h�C         ]     �t�bhhK ��h��R�(KK��h�CX
      �        ]     !         g      Y  �     �     �     �        �t�bhhK ��h��R�(KK��h�C4   p     q     !         b     ^        �t�bhhK ��h��R�(KK��h�C�     R        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK
��h�C(9      !   ~  >  �      !         �t�bhhK ��h��R�(KK��h�C8  "   R       F      �  	   r     �        �t�bhhK ��h��R�(KK��h�C8      �  �     Z   �     �  �     J        �t�bhhK ��h��R�(KK��h�C0s     �     �  7      t     �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK
��h�C($                 E      �     �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C,   !   E  �      �     u           �t�bhhK ��h��R�(KK��h�C0   �  F  v  G     H  >   �  {        �t�bhhK ��h��R�(KK��h�C0I  �  u   �  I   2  �     w           �t�bhhK ��h��R�(KK��h�C@     !      �  �     �     �      Z   >   �        �t�bhhK ��h��R�(KK��h�C<   x        y  z  �     @         
   �        �t�bhhK ��h��R�(KK��h�C\   !         �     �  �      {  |        }  ~       �      �  C         �t�bhhK ��h��R�(KK��h�C          !   Q   2         �t�bhhK ��h��R�(KK��h�CP   !      Z   �  �   	   �     W   �   M   _     D      �  �        �t�bhhK ��h��R�(KK��h�C,      
   �  7         �  �        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�      J     �t�bhhK ��h��R�(KK��h�C�  �     �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     �  �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C,Z     S     ?     !      9         �t�bhhK ��h��R�(KK��h�C@M   q   �  �        g      g  .     K     L        �t�bhhK ��h��R�(KK��h�CD&   �      �   �  "   �  �  �        �  �     !         �t�bhhK ��h��R�(KK	��h�C$         !   �   �  2         �t�bhhK ��h��R�(KK��h�C    �        �  �        �t�bhhK ��h��R�(KK��h�CL      
   �     &   �   �     !   7         9   �   �  2         �t�bhhK ��h��R�(KK
��h�C(         T     �     1         �t�bhhK ��h��R�(KK��h�C%   �   �        �t�bhhK ��h��R�(KK��h�C�      �   O     �t�bhhK ��h��R�(KK��h�C�   �   �        �t�bhhK ��h��R�(KK��h�C�   N     E      �t�bhhK ��h��R�(KK��h�C  M           �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK��h�C,!            :   �        �         �t�bhhK ��h��R�(KK��h�C &   �   �  *      9         �t�bhhK ��h��R�(KK��h�C!   I  �      �        �t�bhhK ��h��R�(KK��h�Cp_     .   W   �  �     !   	      F   �  	   �     �  	   �  	   �  	   �  	   �     �        �t�bhhK ��h��R�(KK��h�C!   "   �  �  |         �t�bhhK ��h��R�(KK��h�CP   #       �  �  �     �  �  "   �   e   f  B  )               �t�bhhK ��h��R�(KK��h�C<�       �  �  	   @      �  �     �        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C[   �                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C !   �  "   �  �  �        �t�bhhK ��h��R�(KK��h�C4B   "   �  y     �  I   �  �  g  �        �t�bhhK ��h��R�(KK��h�C8�  !   "   �     '   �     �  u   9   �        �t�bhhK ��h��R�(KK��h�C09   �    �  a   �     �     Z        �t�bhhK ��h��R�(KK��h�CT9   �  �   �  9   �  	   `  !   ,  I   P        �  !      I   �        �t�bhhK ��h��R�(KK��h�C4�     �     �  9   "   �  �     !         �t�bhhK ��h��R�(KK��h�C`�  �  	   �  �  U      M   9      �     �  �  :  U   9   	   "   �  2  !         �t�bhhK ��h��R�(KK��h�C4�     �     �  "   .   �  �     �        �t�bhhK ��h��R�(KK	��h�C$!      B  �     K  �        �t�bhhK ��h��R�(KK��h�C,   F   �   9      !   >     !         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C    �   a      �      �t�bhhK ��h��R�(KK��h�C�      7     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cn     $      L      �t�bhhK ��h��R�(KK��h�Cn     S     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CX   !   )     �   �        B      F   8  ^  	   Q  	   R  S     T        �t�bhhK ��h��R�(KK��h�CB      -   �   k         �t�bhhK ��h��R�(KK��h�C4   !      <  �     �  �     �  �        �t�bhhK ��h��R�(KK��h�C �   �   �  �  Z   �         �t�bhhK ��h��R�(KK��h�CH�     $      L   �  	   �  �     �  �  �   �     $         �t�bhhK ��h��R�(KK��h�C         X        �t�bhhK ��h��R�(KK��h�C%   )        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C �     $      L   �        �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�C�     �           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�      �           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C@   !      =  �      �        <  �     �           �t�bhhK ��h��R�(KK��h�CL           [  9  	   �  	   �   	   W  	   X     [  e         �t�bhhK ��h��R�(KK��h�C,9     e   Z        ^   >   k         �t�bhhK ��h��R�(KK	��h�C$           D   �   B        �t�bhhK ��h��R�(KK��h�C8   �  �   �   -   �     .   )   �      C         �t�bhhK ��h��R�(KK��h�C,a     !            �  �  �        �t�bhhK ��h��R�(KK��h�CH      �  �     �     �     !   	   *   	   8      9         �t�bhhK ��h��R�(KK
��h�C(   9   �          �  �         �t�bhhK ��h��R�(KK��h�C,v   7   B   9     ;  (  >   k         �t�bhhK ��h��R�(KK��h�CH
      "   '   �     �  	         D   [  9     �          �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C�   �        �t�bhhK ��h��R�(KK��h�C�  Y                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C    !      �  �  �        �t�bhhK ��h��R�(KK��h�C4�     �  "   '   �   �     �     �        �t�bhhK ��h��R�(KK��h�C<   !      ^   �  	   �     W   �     >   �        �t�bhhK ��h��R�(KK��h�C8   �     B   �     �       �     �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�  �                  �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     I           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C    �   a      �      �t�bhhK ��h��R�(KK	��h�C$   !      Z   �     �        �t�bhhK ��h��R�(KK��h�C0      -   �   /      �      �  �        �t�bhhK ��h��R�(KK��h�CL      �     !   Q   �     !   �  	   �  �        V  �        �t�bhhK ��h��R�(KK
��h�C(             �   a      �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     �           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     �           �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�CL     �     �t�bhhK ��h��R�(KK��h�C�      7     �t�bhhK ��h��R�(KK	��h�C$   !      ^   �     �        �t�bhhK ��h��R�(KK��h�C   !      �   �        �t�bhhK ��h��R�(KK��h�C,      
   �  7         �  �        �t�bhhK ��h��R�(KK��h�C_  �   !      �        �t�bhhK ��h��R�(KK��h�C          �      7        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C 7  	   �     �           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C   !      ^   �         �t�bhhK ��h��R�(KK��h�C8   !   �  �   �  �     �     �  �  ^        �t�bhhK ��h��R�(KK��h�C4
   :     �  7            !   Q   2         �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�Cn     $      L      �t�bhhK ��h��R�(KK��h�CD   !      ^   �     p   �     ^  �     $      L         �t�bhhK ��h��R�(KK��h�CP>   �     �   	   �  	   �  	   �   	   �  	   �  	   t     �        �t�bhhK ��h��R�(KK��h�C<H   �     �         �      �  =     _  I         �t�bhhK ��h��R�(KK��h�C`�  �           �  �     �     �     	   �     A     $      �      �        �t�bhhK ��h��R�(KK��h�C,D   �        �   [  +     �         �t�bhhK ��h��R�(KK
��h�C(      7         !   Q   2         �t�bhhK ��h��R�(KK
��h�C(         n     $      L         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   �     �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK
��h�C(�     $      *                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   �           �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�      J           �t�bhhK ��h��R�(KK��h�Cn     S     �t�bhhK ��h��R�(KK%��h�C�
      "   �  �  I      !      J   S        �  �   !   Q   �     �        U  �  �      �  
      "   '   �     �           �t�bhhK ��h��R�(KK��h�C,      �  �  �     !      �        �t�bhhK ��h��R�(KK��h�C8w      /   �     '   �  N      �   
   �        �t�bhhK ��h��R�(KK��h�C`   �     �     O         
   �     ;      S     >   �  	   �      �   T         �t�bhhK ��h��R�(KK��h�C;     �t�bhhK ��h��R�(KK��h�C(         <      �     �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8   !      Z   >   �   	      F   Z             �t�bhhK ��h��R�(KK
��h�C(      7         !   Q   2         �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C    �   a      �      �t�bhhK ��h��R�(KK��h�C�      7     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cn     $      L      �t�bhhK ��h��R�(KK��h�Cn     S     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CX   !   )     �   �        B      F   8  ^  	   Q  	   R  S     T        �t�bhhK ��h��R�(KK��h�CB      -   �   k         �t�bhhK ��h��R�(KK��h�C4   !      <  �     �  �     �  �        �t�bhhK ��h��R�(KK��h�C �   �   �  �  Z   �         �t�bhhK ��h��R�(KK��h�CH�     $      L   �  	   �  �     �  �  �   �     $         �t�bhhK ��h��R�(KK��h�C         X        �t�bhhK ��h��R�(KK��h�C%   )        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C �     $      L   �        �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�C�     �           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�      �           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C@   !      =  �      �        <  �     �           �t�bhhK ��h��R�(KK��h�CL           [  9  	   �  	   �   	   W  	   X     [  e         �t�bhhK ��h��R�(KK��h�C,9     e   Z        ^   >   k         �t�bhhK ��h��R�(KK	��h�C$           D   �   B        �t�bhhK ��h��R�(KK��h�C8   �  �   �   -   �     .   )   �      C         �t�bhhK ��h��R�(KK��h�C,a     !            �  �  �        �t�bhhK ��h��R�(KK��h�CH      �  �     �     �     !   	   *   	   8      9         �t�bhhK ��h��R�(KK
��h�C(   9   �          �  �         �t�bhhK ��h��R�(KK��h�C,v   7   B   9     ;  (  >   k         �t�bhhK ��h��R�(KK��h�CH
      "   '   �     �  	         D   [  9     �          �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C�   �        �t�bhhK ��h��R�(KK��h�C�  Y                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C    !      �  �  �        �t�bhhK ��h��R�(KK��h�C4�     �  "   '   �   �     �     �        �t�bhhK ��h��R�(KK��h�C<   !      ^   �  	   �     W   �     >   �        �t�bhhK ��h��R�(KK��h�C8   �     B   �     �       �     �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�  �                  �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     I           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C    �   a      �      �t�bhhK ��h��R�(KK	��h�C$   !      Z   �     �        �t�bhhK ��h��R�(KK��h�C0      -   �   /      �      �  �        �t�bhhK ��h��R�(KK��h�CL      �     !   Q   �     !   �  	   �  �        V  �        �t�bhhK ��h��R�(KK
��h�C(             �   a      �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     �           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     �           �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�CL     �     �t�bhhK ��h��R�(KK��h�C�      7     �t�bhhK ��h��R�(KK	��h�C$   !      ^   �     �        �t�bhhK ��h��R�(KK��h�C   !      �   �        �t�bhhK ��h��R�(KK��h�C,      
   �  7         �  �        �t�bhhK ��h��R�(KK��h�C_  �   !      �        �t�bhhK ��h��R�(KK��h�C          �      7        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C 7  	   �     �           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C   !      ^   �         �t�bhhK ��h��R�(KK��h�C8   !   �  �   �  �     �     �  �  ^        �t�bhhK ��h��R�(KK��h�C4
   :     �  7            !   Q   2         �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�Cn     $      L      �t�bhhK ��h��R�(KK��h�CD   !      ^   �     p   �     ^  �     $      L         �t�bhhK ��h��R�(KK��h�CP>   �     �   	   �  	   �  	   �   	   �  	   �  	   t     �        �t�bhhK ��h��R�(KK��h�C<H   �     �         �      �  =     _  I         �t�bhhK ��h��R�(KK��h�C`�  �           �  �     �     �     	   �     A     $      �      �        �t�bhhK ��h��R�(KK��h�C,D   �        �   [  +     �         �t�bhhK ��h��R�(KK
��h�C(      7         !   Q   2         �t�bhhK ��h��R�(KK
��h�C(         n     $      L         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   �     �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK
��h�C(�     $      *                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   �           �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�      J           �t�bhhK ��h��R�(KK��h�Cn     S     �t�bhhK ��h��R�(KK%��h�C�
      "   �  �  I      !      J   S        �  �   !   Q   �     �        U  �  �      �  
      "   '   �     �           �t�bhhK ��h��R�(KK��h�C,      �  �  �     !      �        �t�bhhK ��h��R�(KK��h�C8w      /   �     '   �  N      �   
   �        �t�bhhK ��h��R�(KK��h�C`   �     �     O         
   �     ;      S     >   �  	   �      �   T         �t�bhhK ��h��R�(KK��h�C;     �t�bhhK ��h��R�(KK��h�C(         <      �     �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8   !      Z   >   �   	      F   Z             �t�bhhK ��h��R�(KK
��h�C(      7         !   Q   2         �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C    �   a      �      �t�bhhK ��h��R�(KK��h�C�      7     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cn     $      L      �t�bhhK ��h��R�(KK��h�Cn     S     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CX   !   )     �   �        B      F   8  ^  	   Q  	   R  S     T        �t�bhhK ��h��R�(KK��h�CB      -   �   k         �t�bhhK ��h��R�(KK��h�C4   !      <  �     �  �     �  �        �t�bhhK ��h��R�(KK��h�C �   �   �  �  Z   �         �t�bhhK ��h��R�(KK��h�CH�     $      L   �  	   �  �     �  �  �   �     $         �t�bhhK ��h��R�(KK��h�C         X        �t�bhhK ��h��R�(KK��h�C%   )        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C �     $      L   �        �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�C�     �           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�      �           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C@   !      =  �      �        <  �     �           �t�bhhK ��h��R�(KK��h�CL           [  9  	   �  	   �   	   W  	   X     [  e         �t�bhhK ��h��R�(KK��h�C,9     e   Z        ^   >   k         �t�bhhK ��h��R�(KK	��h�C$           D   �   B        �t�bhhK ��h��R�(KK��h�C8   �  �   �   -   �     .   )   �      C         �t�bhhK ��h��R�(KK��h�C,a     !            �  �  �        �t�bhhK ��h��R�(KK��h�CH      �  �     �     �     !   	   *   	   8      9         �t�bhhK ��h��R�(KK
��h�C(   9   �          �  �         �t�bhhK ��h��R�(KK��h�C,v   7   B   9     ;  (  >   k         �t�bhhK ��h��R�(KK��h�CH
      "   '   �     �  	         D   [  9     �          �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C�   �        �t�bhhK ��h��R�(KK��h�C�  Y                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C    !      �  �  �        �t�bhhK ��h��R�(KK��h�C4�     �  "   '   �   �     �     �        �t�bhhK ��h��R�(KK��h�C<   !      ^   �  	   �     W   �     >   �        �t�bhhK ��h��R�(KK��h�C8   �     B   �     �       �     �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�  �                  �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     I           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C    �   a      �      �t�bhhK ��h��R�(KK	��h�C$   !      Z   �     �        �t�bhhK ��h��R�(KK��h�C0      -   �   /      �      �  �        �t�bhhK ��h��R�(KK��h�CL      �     !   Q   �     !   �  	   �  �        V  �        �t�bhhK ��h��R�(KK
��h�C(             �   a      �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     �           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     �           �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�CL     �     �t�bhhK ��h��R�(KK��h�C�      7     �t�bhhK ��h��R�(KK	��h�C$   !      ^   �     �        �t�bhhK ��h��R�(KK��h�C   !      �   �        �t�bhhK ��h��R�(KK��h�C,      
   �  7         �  �        �t�bhhK ��h��R�(KK��h�C_  �   !      �        �t�bhhK ��h��R�(KK��h�C          �      7        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C 7  	   �     �           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C   !      ^   �         �t�bhhK ��h��R�(KK��h�C8   !   �  �   �  �     �     �  �  ^        �t�bhhK ��h��R�(KK��h�C4
   :     �  7            !   Q   2         �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�Cn     $      L      �t�bhhK ��h��R�(KK��h�CD   !      ^   �     p   �     ^  �     $      L         �t�bhhK ��h��R�(KK��h�CP>   �     �   	   �  	   �  	   �   	   �  	   �  	   t     �        �t�bhhK ��h��R�(KK��h�C<H   �     �         �      �  =     _  I         �t�bhhK ��h��R�(KK��h�C`�  �           �  �     �     �     	   �     A     $      �      �        �t�bhhK ��h��R�(KK��h�C,D   �        �   [  +     �         �t�bhhK ��h��R�(KK
��h�C(      7         !   Q   2         �t�bhhK ��h��R�(KK
��h�C(         n     $      L         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   �     �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK
��h�C(�     $      *                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   �           �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�      J           �t�bhhK ��h��R�(KK��h�Cn     S     �t�bhhK ��h��R�(KK%��h�C�
      "   �  �  I      !      J   S        �  �   !   Q   �     �        U  �  �      �  
      "   '   �     �           �t�bhhK ��h��R�(KK��h�C,      �  �  �     !      �        �t�bhhK ��h��R�(KK��h�C8w      /   �     '   �  N      �   
   �        �t�bhhK ��h��R�(KK��h�C`   �     �     O         
   �     ;      S     >   �  	   �      �   T         �t�bhhK ��h��R�(KK��h�C;     �t�bhhK ��h��R�(KK��h�C(         <      �     �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8   !      Z   >   �   	      F   Z             �t�bhhK ��h��R�(KK
��h�C(      7         !   Q   2         �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C,      �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�C�      �     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CD
      5   �   +      �  	   �     �  	   �   �   �         �t�bhhK ��h��R�(KK��h�CT   O   �   �   x     �   �  v   C  	   G   	   D     5        E        �t�bhhK ��h��R�(KK ��h�C�
      �          �  	   �         �  b        �     �  	         =   0      �      )  }  *           �t�bhhK ��h��R�(KK��h�C4      D   g   +                 �        �t�bhhK ��h��R�(KK��h�C,0      �   "   �   �   �   d  E        �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C(      <      +     �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�Cd�     �  �                 E      s     �      �      �      �     �     }     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C 0                       �t�bhhK ��h��R�(KK��h�C,      �     �t�bhhK ��h��R�(KK��h�C4
      "   ,      �     �  	   =   �        �t�bhhK ��h��R�(KK��h�C0      -   �   
   f      �     C         �t�bhhK ��h��R�(KK��h�C0   
   �         �  �  C      !         �t�bhhK ��h��R�(KK��h�C �  |  �        9         �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C         ,      �     �t�bhhK ��h��R�(KK��h�C>   �                 �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�CL   9      3  X  	   v   Y      �     1   �   >     @   �        �t�bhhK ��h��R�(KK
��h�C(�      3  X     v     Q        �t�bhhK ��h��R�(KK��h�C03  X  �  4   Q     �     W   {        �t�bhhK ��h��R�(KK��h�C4       �  Q  �  4   �  �      �  �        �t�bhhK ��h��R�(KK
��h�C(l     3  X     9      �        �t�bhhK ��h��R�(KK
��h�C(�  �        �        @        �t�bhhK ��h��R�(KK��h�C,     �     �     �     �        �t�bhhK ��h��R�(KK��h�C         ,      {      �t�bhhK ��h��R�(KK��h�C@�     �           E      �      �      �     �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8      �        �  �   ]      1     �        �t�bhhK ��h��R�(KK��h�C\      D   �         "  
   �     �      �         4   5   �  +      �        �t�bhhK ��h��R�(KK��h�C�  F     �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�            �t�bhhK ��h��R�(KK��h�C'  \                 �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�C<�  ~        �     �  �     �        !         �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�CP      D   g      
   �   Q        F   �   �     �  �     2         �t�bhhK ��h��R�(KK	��h�C$         5           h      �t�bhhK ��h��R�(KK��h�C�  ~           �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C�   �        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�C    �  �     �   �         �t�bhhK ��h��R�(KK��h�Cd   o  O   B   -   +      !   Q   0           )  }  *     	      "   �   �   �         �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C(      <      +     �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�Cd�     �  �                 E      s     �      �      �      �     �     }     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cd
        J   �  G  l   p  /      �  /      l   	         =   '   �      �           �t�bhhK ��h��R�(KK��h�C�  "   �  �   �         �t�bhhK ��h��R�(KK��h�CD#  �     �  �        '   �   �     �     �  $         �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�C�  �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CP      -        !   �      �   �        �  �      �  �           �t�bhhK ��h��R�(KK��h�C         <      �     �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�Cz  O     �t�bhhK ��h��R�(KK��h�C(      <      ]     �t�bhhK ��h��R�(KK��h�C+      �     �     �t�bhhK ��h��R�(KK��h�C+      �     �t�bhhK ��h��R�(KK��h�CL�  H     ^       H     ^  A     p   f      V      �        �t�bhhK ��h��R�(KK��h�CD�  "   '                !   v   B   O   V      f         �t�bhhK ��h��R�(KK��h�C(      <           �t�bhhK ��h��R�(KK��h�CP+      V      I           E      �      �      �      �     �     �t�bhhK ��h��R�(KK��h�C+      G     �t�bhhK ��h��R�(KK#��h�C�G     "     l   p  �  �     "   �  �  �     l      �   	      @   +   U   �          !      �   �                �t�bhhK ��h��R�(KK	��h�C$+      G      �     �  �     �t�bhhK ��h��R�(KK��h�C<�  `     �  `     x   _     "   ,      l         �t�bhhK ��h��R�(KK��h�C(      <      a     �t�bhhK ��h��R�(KK��h�C0+      G         �     �  �           �t�bhhK ��h��R�(KK��h�C+      L      �t�bhhK ��h��R�(KK��h�Cl�   	  
  !  _   (     �  �  �  �  �     p   V      +      o     J     %     �        �t�bhhK ��h��R�(KK��h�C<"  "   �   y      _     =  	   �  �   �   �         �t�bhhK ��h��R�(KK��h�C�  :     �  �        �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C�   	  
        �t�bhhK ��h��R�(KK��h�C :   _   #                 �t�bhhK ��h��R�(KK��h�C         l      �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK��h�CX�     $   ?   r  I         ,      m      �   @   +      �      �           �t�bhhK ��h��R�(KK	��h�C$P  7         !   Q   2         �t�bhhK ��h��R�(KK��h�C b  ;      �     v        �t�bhhK ��h��R�(KK��h�Ch   z  o  �   K        =   0      �      )  }  *     	      "   �   �   �   d  E        �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C(      <      +     �t�bhhK ��h��R�(KK��h�CX   ,      b     K  O   B   -   +      �      !   �     �     	           �t�bhhK ��h��R�(KK	��h�C$         ,      m      �      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�Cc           �t�bhhK ��h��R�(KK��h�C%   �   �        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C\
     �        �     �     p   f      �      �  n   G   	        �        �t�bhhK ��h��R�(KK��h�Ch   ,   d   $      �   O   B   +   d             	   �                             �t�bhhK ��h��R�(KK
��h�C(      7         !   Q   2         �t�bhhK ��h��R�(KK��h�C          n      _   ,      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�Cc           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C8   
   ;      $   	   �                       �t�bhhK ��h��R�(KK��h�Cl   @  O   :   L   +                  }       	   �                             �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
   K                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CTr     F     H  $      �   \   �       @   +   d   �     �           �t�bhhK ��h��R�(KK��h�C<   �           F   @   +      `  ,      �         �t�bhhK ��h��R�(KK��h�C +      *                 �t�bhhK ��h��R�(KK��h�CH
         ?     I   	         @   f        M   q   d        �t�bhhK ��h��R�(KK��h�C@�     d  x   /   
      4   "   �   �         �         �t�bhhK ��h��R�(KK��h�CD      -   >  
   f   �  W   �  	      F   �              �t�bhhK ��h��R�(KK��h�C:   _   (     �t�bhhK ��h��R�(KK��h�Cl�   	  
  !  _   (     �  �  �  �  �     p   V      +      o     J     %     �        �t�bhhK ��h��R�(KK��h�C<"  "   �   y      _     =  	   �  �   �   �         �t�bhhK ��h��R�(KK��h�C�  :     �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C          n      _   ,      �t�bhhK ��h��R�(KK��h�C�   	  
        �t�bhhK ��h��R�(KK��h�C :   _   #                 �t�bhhK ��h��R�(KK��h�C      V      *           �t�bhhK ��h��R�(KK��h�CT          p      
   �              W     
      "   Q  ,         �t�bhhK ��h��R�(KK��h�C(      <              �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�Ct!              �        "  #  �      4   "   $  W   �     %  	      
     �     [  �        �t�bhhK ��h��R�(KK��h�C`�        @   
      4   &  @     �  2  �   �   	   '          �   e   �        �t�bhhK ��h��R�(KK��h�CP      >  
   f   �  `   
   �  M   &   r  s  (      <      (        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
                    �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�CX
      4      �    )     �  �   :   *  	   6      =   +     ,           �t�bhhK ��h��R�(KK��h�C(      <               �t�bhhK ��h��R�(KK��h�C%   �     �        �t�bhhK ��h��R�(KK��h�C �                      �t�bhhK ��h��R�(KK��h�C(  -     �t�bhhK ��h��R�(KK��h�Cx
      "   �  �        .  \   "   {      @   �  	         i   
   �  M   &   �  /     0  1           �t�bhhK ��h��R�(KK��h�C0l     2             <      3        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK	��h�C$   
   (  4                 �t�bhhK ��h��R�(KK��h�C�      �     �t�bhhK ��h��R�(KK��h�C�     �   �     �     �t�bhhK ��h��R�(KK��h�C�  O    �        �t�bhhK ��h��R�(KK��h�C(      <      5     �t�bhhK ��h��R�(KK��h�C6     �   �     �     �t�bhhK ��h��R�(KK��h�C(      <      7     �t�bhhK ��h��R�(KK��h�C     �     �t�bhhK ��h��R�(KK��h�C8  �  e  	   �        �t�bhhK ��h��R�(KK��h�C(      <      9     �t�bhhK ��h��R�(KK��h�C4       "   D   !     �     �  5        �t�bhhK ��h��R�(KK��h�CT
      "   :        g   +      ;          	              9         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C(   <        �t�bhhK ��h��R�(KK��h�C@�  �     �  �     x   �      �   	   =     �        �t�bhhK ��h��R�(KK��h�CD�  p   D   V      �      >  a      ?  d     �  �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C +                       �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK
��h�C(   
   o      @                 �t�bhhK ��h��R�(KK��h�C+      A     �t�bhhK ��h��R�(KK��h�C +      *                 �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C8   !      �   �     �  :   �      �   W        �t�bhhK ��h��R�(KK��h�C`   B     !      �   �     9   �  c     �  Y      4   "   �  �     �           �t�bhhK ��h��R�(KK��h�C\   
   	  O         !   �  
     �   C             �   �                �t�bhhK ��h��R�(KK��h�C!   �  
     �t�bhhK ��h��R�(KK��h�CD  �     �t�bhhK ��h��R�(KK��h�C(      <      E     �t�bhhK ��h��R�(KK&��h�C�
   J   �  b  �  	         @   +          F  /   U   &   G  H     V          D  /   g  I     �  0           )  }  *           �t�bhhK ��h��R�(KK	��h�C$e  "   �   d  E  �   �         �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C(      <      +     �t�bhhK ��h��R�(KK��h�C         �     �t�bhhK ��h��R�(KK��h�C%   �   �        �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�   �   �        �t�bhhK ��h��R�(KK��h�CJ  K     �t�bhhK ��h��R�(KK��h�C�             �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK
��h�C(N      �  "   L                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C 0                       �t�bhhK ��h��R�(KK��h�C,      �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�C�      �     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CD
      5   �   +      �  	   �     �  	   �   �   �         �t�bhhK ��h��R�(KK��h�CT   O   �   �   x     �   �  v   C  	   G   	   D     5        E        �t�bhhK ��h��R�(KK ��h�C�
      �          �  	   �         �  b        �     �  	         =   0      �      )  }  *           �t�bhhK ��h��R�(KK��h�C4      D   g   +                 �        �t�bhhK ��h��R�(KK��h�C,0      �   "   �   �   �   d  E        �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C(      <      +     �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�Cd�     �  �                 E      s     �      �      �      �     �     }     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C 0                       �t�bhhK ��h��R�(KK��h�C,      �     �t�bhhK ��h��R�(KK��h�C4
      "   ,      �     �  	   =   �        �t�bhhK ��h��R�(KK��h�C0      -   �   
   f      �     C         �t�bhhK ��h��R�(KK��h�C0   
   �         �  �  C      !         �t�bhhK ��h��R�(KK��h�C �  |  �        9         �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C         ,      �     �t�bhhK ��h��R�(KK��h�C>   �                 �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�CL   9      3  X  	   v   Y      �     1   �   >     @   �        �t�bhhK ��h��R�(KK
��h�C(�      3  X     v     Q        �t�bhhK ��h��R�(KK��h�C03  X  �  4   Q     �     W   {        �t�bhhK ��h��R�(KK��h�C4       �  Q  �  4   �  �      �  �        �t�bhhK ��h��R�(KK
��h�C(l     3  X     9      �        �t�bhhK ��h��R�(KK
��h�C(�  �        �        @        �t�bhhK ��h��R�(KK��h�C,     �     �     �     �        �t�bhhK ��h��R�(KK��h�C         ,      {      �t�bhhK ��h��R�(KK��h�C@�     �           E      �      �      �     �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8      �        �  �   ]      1     �        �t�bhhK ��h��R�(KK��h�C\      D   �         "  
   �     �      �         4   5   �  +      �        �t�bhhK ��h��R�(KK��h�C�  F     �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�            �t�bhhK ��h��R�(KK��h�C'  \                 �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�C<�  ~        �     �  �     �        !         �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�CP      D   g      
   �   Q        F   �   �     �  �     2         �t�bhhK ��h��R�(KK	��h�C$         5           h      �t�bhhK ��h��R�(KK��h�C�  ~           �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C�   �        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�C    �  �     �   �         �t�bhhK ��h��R�(KK��h�Cd   o  O   B   -   +      !   Q   0           )  }  *     	      "   �   �   �         �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C(      <      +     �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�Cd�     �  �                 E      s     �      �      �      �     �     }     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cd
        J   �  G  l   p  /      �  /      l   	         =   '   �      �           �t�bhhK ��h��R�(KK��h�C�  "   �  �   �         �t�bhhK ��h��R�(KK��h�CD#  �     �  �        '   �   �     �     �  $         �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�C�  �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CP      -        !   �      �   �        �  �      �  �           �t�bhhK ��h��R�(KK��h�C         <      �     �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�Cz  O     �t�bhhK ��h��R�(KK��h�C(      <      ]     �t�bhhK ��h��R�(KK��h�C+      �     �     �t�bhhK ��h��R�(KK��h�C+      �     �t�bhhK ��h��R�(KK��h�CL�  H     ^       H     ^  A     p   f      V      �        �t�bhhK ��h��R�(KK��h�CD�  "   '                !   v   B   O   V      f         �t�bhhK ��h��R�(KK��h�C(      <           �t�bhhK ��h��R�(KK��h�CP+      V      I           E      �      �      �      �     �     �t�bhhK ��h��R�(KK��h�C+      G     �t�bhhK ��h��R�(KK#��h�C�G     "     l   p  �  �     "   �  �  �     l      �   	      @   +   U   �          !      �   �                �t�bhhK ��h��R�(KK	��h�C$+      G      �     �  �     �t�bhhK ��h��R�(KK��h�C<�  `     �  `     x   _     "   ,      l         �t�bhhK ��h��R�(KK��h�C(      <      a     �t�bhhK ��h��R�(KK��h�C0+      G         �     �  �           �t�bhhK ��h��R�(KK��h�C+      L      �t�bhhK ��h��R�(KK��h�Cl�   	  
  !  _   (     �  �  �  �  �     p   V      +      o     J     %     �        �t�bhhK ��h��R�(KK��h�C<"  "   �   y      _     =  	   �  �   �   �         �t�bhhK ��h��R�(KK��h�C�  :     �  �        �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C�   	  
        �t�bhhK ��h��R�(KK��h�C :   _   #                 �t�bhhK ��h��R�(KK��h�C         l      �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK��h�CX�     $   ?   r  I         ,      m      �   @   +      �      �           �t�bhhK ��h��R�(KK	��h�C$P  7         !   Q   2         �t�bhhK ��h��R�(KK��h�C b  ;      �     v        �t�bhhK ��h��R�(KK��h�Ch   z  o  �   K        =   0      �      )  }  *     	      "   �   �   �   d  E        �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C(      <      +     �t�bhhK ��h��R�(KK��h�CX   ,      b     K  O   B   -   +      �      !   �     �     	           �t�bhhK ��h��R�(KK	��h�C$         ,      m      �      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�Cc           �t�bhhK ��h��R�(KK��h�C%   �   �        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C\
     �        �     �     p   f      �      �  n   G   	        �        �t�bhhK ��h��R�(KK��h�Ch   ,   d   $      �   O   B   +   d             	   �                             �t�bhhK ��h��R�(KK
��h�C(      7         !   Q   2         �t�bhhK ��h��R�(KK��h�C          n      _   ,      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�Cc           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C8   
   ;      $   	   �                       �t�bhhK ��h��R�(KK��h�Cl   @  O   :   L   +                  }       	   �                             �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
   K                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C%            �t�bh�      hK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CTr     F     H  $      �   \   �       @   +   d   �     �           �t�bhhK ��h��R�(KK��h�C<   �           F   @   +      `  ,      �         �t�bhhK ��h��R�(KK��h�C +      *                 �t�bhhK ��h��R�(KK��h�CH
         ?     I   	         @   f        M   q   d        �t�bhhK ��h��R�(KK��h�C@�     d  x   /   
      4   "   �   �         �         �t�bhhK ��h��R�(KK��h�CD      -   >  
   f   �  W   �  	      F   �              �t�bhhK ��h��R�(KK��h�C:   _   (     �t�bhhK ��h��R�(KK��h�Cl�   	  
  !  _   (     �  �  �  �  �     p   V      +      o     J     %     �        �t�bhhK ��h��R�(KK��h�C<"  "   �   y      _     =  	   �  �   �   �         �t�bhhK ��h��R�(KK��h�C�  :     �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C          n      _   ,      �t�bhhK ��h��R�(KK��h�C�   	  
        �t�bhhK ��h��R�(KK��h�C :   _   #                 �t�bhhK ��h��R�(KK��h�C      V      *           �t�bhhK ��h��R�(KK��h�CT          p      
   �              W     
      "   Q  ,         �t�bhhK ��h��R�(KK��h�C(      <              �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�Ct!              �        "  #  �      4   "   $  W   �     %  	      
     �     [  �        �t�bhhK ��h��R�(KK��h�C`�        @   
      4   &  @     �  2  �   �   	   '          �   e   �        �t�bhhK ��h��R�(KK��h�CP      >  
   f   �  `   
   �  M   &   r  s  (      <      (        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
                    �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�CX
      4      �    )     �  �   :   *  	   6      =   +     ,           �t�bhhK ��h��R�(KK��h�C(      <               �t�bhhK ��h��R�(KK��h�C%   �     �        �t�bhhK ��h��R�(KK��h�C �                      �t�bhhK ��h��R�(KK��h�C(  -     �t�bhhK ��h��R�(KK��h�Cx
      "   �  �        .  \   "   {      @   �  	         i   
   �  M   &   �  /     0  1           �t�bhhK ��h��R�(KK��h�C0l     2             <      3        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK	��h�C$   
   (  4                 �t�bhhK ��h��R�(KK��h�C�      �     �t�bhhK ��h��R�(KK��h�C�     �   �     �     �t�bhhK ��h��R�(KK��h�C�  O    �        �t�bhhK ��h��R�(KK��h�C(      <      5     �t�bhhK ��h��R�(KK��h�C6     �   �     �     �t�bhhK ��h��R�(KK��h�C(      <      7     �t�bhhK ��h��R�(KK��h�C     �     �t�bhhK ��h��R�(KK��h�C8  �  e  	   �        �t�bhhK ��h��R�(KK��h�C(      <      9     �t�bhhK ��h��R�(KK��h�C4       "   D   !     �     �  5        �t�bhhK ��h��R�(KK��h�CT
      "   :        g   +      ;          	              9         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C(   <        �t�bhhK ��h��R�(KK��h�C@�  �     �  �     x   �      �   	   =     �        �t�bhhK ��h��R�(KK��h�CD�  p   D   V      �      >  a      ?  d     �  �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C +                       �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK
��h�C(   
   o      @                 �t�bhhK ��h��R�(KK��h�C+      A     �t�bhhK ��h��R�(KK��h�C +      *                 �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C8   !      �   �     �  :   �      �   W        �t�bhhK ��h��R�(KK��h�C`   B     !      �   �     9   �  c     �  Y      4   "   �  �     �           �t�bhhK ��h��R�(KK��h�C\   
   	  O         !   �  
     �   C             �   �                �t�bhhK ��h��R�(KK��h�C!   �  
     �t�bhhK ��h��R�(KK��h�CD  �     �t�bhhK ��h��R�(KK��h�C(      <      E     �t�bhhK ��h��R�(KK&��h�C�
   J   �  b  �  	         @   +          F  /   U   &   G  H     V          D  /   g  I     �  0           )  }  *           �t�bhhK ��h��R�(KK	��h�C$e  "   �   d  E  �   �         �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C(      <      +     �t�bhhK ��h��R�(KK��h�C         �     �t�bhhK ��h��R�(KK��h�C%   �   �        �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�   �   �        �t�bhhK ��h��R�(KK��h�CJ  K     �t�bhhK ��h��R�(KK��h�C�             �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK
��h�C(N      �  "   L                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C 0                       �t�bhhK ��h��R�(KK��h�C,      �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�C�      �     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CD
      5   �   +      �  	   �     �  	   �   �   �         �t�bhhK ��h��R�(KK��h�CT   O   �   �   x     �   �  v   C  	   G   	   D     5        E        �t�bhhK ��h��R�(KK ��h�C�
      �          �  	   �         �  b        �     �  	         =   0      �      )  }  *           �t�bhhK ��h��R�(KK��h�C4      D   g   +                 �        �t�bhhK ��h��R�(KK��h�C,0      �   "   �   �   �   d  E        �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C(      <      +     �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�Cd�     �  �                 E      s     �      �      �      �     �     }     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C 0                       �t�bhhK ��h��R�(KK��h�C,      �     �t�bhhK ��h��R�(KK��h�C4
      "   ,      �     �  	   =   �        �t�bhhK ��h��R�(KK��h�C0      -   �   
   f      �     C         �t�bhhK ��h��R�(KK��h�C0   
   �         �  �  C      !         �t�bhhK ��h��R�(KK��h�C �  |  �        9         �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C         ,      �     �t�bhhK ��h��R�(KK��h�C>   �                 �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�CL   9      3  X  	   v   Y      �     1   �   >     @   �        �t�bhhK ��h��R�(KK
��h�C(�      3  X     v     Q        �t�bhhK ��h��R�(KK��h�C03  X  �  4   Q     �     W   {        �t�bhhK ��h��R�(KK��h�C4       �  Q  �  4   �  �      �  �        �t�bhhK ��h��R�(KK
��h�C(l     3  X     9      �        �t�bhhK ��h��R�(KK
��h�C(�  �        �        @        �t�bhhK ��h��R�(KK��h�C,     �     �     �     �        �t�bhhK ��h��R�(KK��h�C         ,      {      �t�bhhK ��h��R�(KK��h�C@�     �           E      �      �      �     �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8      �        �  �   ]      1     �        �t�bhhK ��h��R�(KK��h�C\      D   �         "  
   �     �      �         4   5   �  +      �        �t�bhhK ��h��R�(KK��h�C�  F     �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�            �t�bhhK ��h��R�(KK��h�C'  \                 �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�C<�  ~        �     �  �     �        !         �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�CP      D   g      
   �   Q        F   �   �     �  �     2         �t�bhhK ��h��R�(KK	��h�C$         5           h      �t�bhhK ��h��R�(KK��h�C�  ~           �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C�   �        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�C    �  �     �   �         �t�bhhK ��h��R�(KK��h�Cd   o  O   B   -   +      !   Q   0           )  }  *     	      "   �   �   �         �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C(      <      +     �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�Cd�     �  �                 E      s     �      �      �      �     �     }     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cd
        J   �  G  l   p  /      �  /      l   	         =   '   �      �           �t�bhhK ��h��R�(KK��h�C�  "   �  �   �         �t�bhhK ��h��R�(KK��h�CD#  �     �  �        '   �   �     �     �  $         �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�C�  �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CP      -        !   �      �   �        �  �      �  �           �t�bhhK ��h��R�(KK��h�C         <      �     �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�Cz  O     �t�bhhK ��h��R�(KK��h�C(      <      ]     �t�bhhK ��h��R�(KK��h�C+      �     �     �t�bhhK ��h��R�(KK��h�C+      �     �t�bhhK ��h��R�(KK��h�CL�  H     ^       H     ^  A     p   f      V      �        �t�bhhK ��h��R�(KK��h�CD�  "   '                !   v   B   O   V      f         �t�bhhK ��h��R�(KK��h�C(      <           �t�bhhK ��h��R�(KK��h�CP+      V      I           E      �      �      �      �     �     �t�bhhK ��h��R�(KK��h�C+      G     �t�bhhK ��h��R�(KK#��h�C�G     "     l   p  �  �     "   �  �  �     l      �   	      @   +   U   �          !      �   �                �t�bhhK ��h��R�(KK	��h�C$+      G      �     �  �     �t�bhhK ��h��R�(KK��h�C<�  `     �  `     x   _     "   ,      l         �t�bhhK ��h��R�(KK��h�C(      <      a     �t�bhhK ��h��R�(KK��h�C0+      G         �     �  �           �t�bhhK ��h��R�(KK��h�C+      L      �t�bhhK ��h��R�(KK��h�Cl�   	  
  !  _   (     �  �  �  �  �     p   V      +      o     J     %     �        �t�bhhK ��h��R�(KK��h�C<"  "   �   y      _     =  	   �  �   �   �         �t�bhhK ��h��R�(KK��h�C�  :     �  �        �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C�   	  
        �t�bhhK ��h��R�(KK��h�C :   _   #                 �t�bhhK ��h��R�(KK��h�C         l      �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK��h�CX�     $   ?   r  I         ,      m      �   @   +      �      �           �t�bhhK ��h��R�(KK	��h�C$P  7         !   Q   2         �t�bhhK ��h��R�(KK��h�C b  ;      �     v        �t�bhhK ��h��R�(KK��h�Ch   z  o  �   K        =   0      �      )  }  *     	      "   �   �   �   d  E        �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C(      <      +     �t�bhhK ��h��R�(KK��h�CX   ,      b     K  O   B   -   +      �      !   �     �     	           �t�bhhK ��h��R�(KK	��h�C$         ,      m      �      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�Cc           �t�bhhK ��h��R�(KK��h�C%   �   �        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C\
     �        �     �     p   f      �      �  n   G   	        �        �t�be(hhK ��h��R�(KK��h�Ch   ,   d   $      �   O   B   +   d             	   �                             �t�bhhK ��h��R�(KK
��h�C(      7         !   Q   2         �t�bhhK ��h��R�(KK��h�C          n      _   ,      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�Cc           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C8   
   ;      $   	   �                       �t�bhhK ��h��R�(KK��h�Cl   @  O   :   L   +                  }       	   �                             �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
   K                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CTr     F     H  $      �   \   �       @   +   d   �     �           �t�bhhK ��h��R�(KK��h�C<   �           F   @   +      `  ,      �         �t�bhhK ��h��R�(KK��h�C +      *                 �t�bhhK ��h��R�(KK��h�CH
         ?     I   	         @   f        M   q   d        �t�bhhK ��h��R�(KK��h�C@�     d  x   /   
      4   "   �   �         �         �t�bhhK ��h��R�(KK��h�CD      -   >  
   f   �  W   �  	      F   �              �t�bhhK ��h��R�(KK��h�C:   _   (     �t�bhhK ��h��R�(KK��h�Cl�   	  
  !  _   (     �  �  �  �  �     p   V      +      o     J     %     �        �t�bhhK ��h��R�(KK��h�C<"  "   �   y      _     =  	   �  �   �   �         �t�bhhK ��h��R�(KK��h�C�  :     �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C          n      _   ,      �t�bhhK ��h��R�(KK��h�C�   	  
        �t�bhhK ��h��R�(KK��h�C :   _   #                 �t�bhhK ��h��R�(KK��h�C      V      *           �t�bhhK ��h��R�(KK��h�CT          p      
   �              W     
      "   Q  ,         �t�bhhK ��h��R�(KK��h�C(      <              �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�Ct!              �        "  #  �      4   "   $  W   �     %  	      
     �     [  �        �t�bhhK ��h��R�(KK��h�C`�        @   
      4   &  @     �  2  �   �   	   '          �   e   �        �t�bhhK ��h��R�(KK��h�CP      >  
   f   �  `   
   �  M   &   r  s  (      <      (        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
                    �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�CX
      4      �    )     �  �   :   *  	   6      =   +     ,           �t�bhhK ��h��R�(KK��h�C(            �t�bhhK ��h��R�(KK��h�C%   �     �        �t�bhhK ��h��R�(KK��h�C �                      �t�bhhK ��h��R�(KK��h�C(  -     �t�bhhK ��h��R�(KK��h�Cx
      "   �  �        .  \   "   {      @   �  	         i   
   �  M   &   �  /     0  1           �t�bhhK ��h��R�(KK��h�C0l     2             <      3        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK	��h�C$   
   (  4                 �t�bhhK ��h��R�(KK��h�C�      �     �t�bhhK ��h��R�(KK��h�C�     �   �     �     �t�bhhK ��h��R�(KK��h�C�  O    �        �t�bhhK ��h��R�(KK��h�C(      <      5     �t�bhhK ��h��R�(KK��h�C6     �   �     �     �t�bhhK ��h��R�(KK��h�C(      <      7     �t�bhhK ��h��R�(KK��h�C     �     �t�bhhK ��h��R�(KK��h�C8  �  e  	   �        �t�bhhK ��h��R�(KK��h�C(      <      9     �t�bhhK ��h��R�(KK��h�C4       "   D   !     �     �  5        �t�bhhK ��h��R�(KK��h�CT
      "   :        g   +      ;          	              9         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C(   <        �t�bhhK ��h��R�(KK��h�C@�  �     �  �     x   �      �   	   =     �        �t�bhhK ��h��R�(KK��h�CD�  p   D   V      �      >  a      ?  d     �  �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C +                       �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK
��h�C(   
   o      @                 �t�bhhK ��h��R�(KK��h�C+      A     �t�bhhK ��h��R�(KK��h�C +      *                 �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C8   !      �   �     �  :   �      �   W        �t�bhhK ��h��R�(KK��h�C`   B     !      �   �     9   �  c     �  Y      4   "   �  �     �           �t�bhhK ��h��R�(KK��h�C\   
   	  O         !   �  
     �   C             �   �                �t�bhhK ��h��R�(KK��h�C!   �  
     �t�bhhK ��h��R�(KK��h�CD  �     �t�bhhK ��h��R�(KK��h�C(      <      E     �t�bhhK ��h��R�(KK&��h�C�
   J   �  b  �  	         @   +          F  /   U   &   G  H     V          D  /   g  I     �  0           )  }  *           �t�bhhK ��h��R�(KK	��h�C$e  "   �   d  E  �   �         �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C(      <      +     �t�bhhK ��h��R�(KK��h�C         �     �t�bhhK ��h��R�(KK��h�C%   �   �        �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�   �   �        �t�bhhK ��h��R�(KK��h�CJ  K     �t�bhhK ��h��R�(KK��h�C�             �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK
��h�C(N      �  "   L                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C 0                       �t�bhhK ��h��R�(KK��h�Cm      �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C�   f     �t�bhhK ��h��R�(KK��h�Co      $      �t�bhhK ��h��R�(KK��h�C,      K     �t�bhhK ��h��R�(KK��h�Cm      �t�bhhK ��h��R�(KK��h�C8�  �  6      d  $  g                    �t�bhhK ��h��R�(KK	��h�C$e  �     �                 �t�bhhK ��h��R�(KK��h�C,      $  g     ,  �     a        �t�bhhK ��h��R�(KK	��h�C$      7         	  2         �t�bhhK ��h��R�(KK��h�C D   M  N  O     �         �t�bhhK ��h��R�(KK��h�C�  h  	   �  �      �t�bhhK ��h��R�(KK��h�CP  !      �t�bhhK ��h��R�(KK��h�C         m         �t�bhhK ��h��R�(KK
��h�C(  
   �     O  p  �           �t�bhhK ��h��R�(KK��h�C Q     �                 �t�bhhK ��h��R�(KK��h�C%   �        �t�bhhK ��h��R�(KK	��h�C$   
   R  �                 �t�bhhK ��h��R�(KK��h�C�   �   �        �t�bhhK ��h��R�(KK��h�C   
   �  �     E      �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C4d     e     �   �   g     !   f  �        �t�bhhK ��h��R�(KK��h�CD�     i   
   b   ?     D      &   �  S  �   .   g        �t�bhhK ��h��R�(KK��h�CP`      �     h  �     �  T  �     	   i     M                �t�bhhK ��h��R�(KK��h�C(   U     �t�bhhK ��h��R�(KK��h�C         b         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
              �t�bhhK ��h��R�(KK	��h�C$    i   
                    �t�bhhK ��h��R�(KK��h�CT
      "   $      6   j  /   �      �      �             !            �t�bhhK ��h��R�(KK��h�C<H  �  '   k  
   �  �   	   l  	   �     �        �t�bhhK ��h��R�(KK��h�C,�  p   -   f      �     6   V        �t�bhhK ��h��R�(KK��h�C,P     �  7         !   Q   2         �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C$      b         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C �                       �t�bhhK ��h��R�(KK��h�C�   f     �t�bhhK ��h��R�(KK��h�C4W  
   �   f  �  U        X     1         �t�bhhK ��h��R�(KK��h�Cl   6     �   �  	   f     W   Y       �      Z           $  �     �  M     /         �t�bhhK ��h��R�(KK��h�Cl      �     
        �   f  	   [     \  
   z      j   �      N   '   $   �     1         �t�bhhK ��h��R�(KK��h�Co      $      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CD   j   �   P     !   7         
   �      $      !         �t�bhhK ��h��R�(KK��h�Co     �t�bhhK ��h��R�(KK��h�CP
      �   �   
   '   ?     $   	         @   o       �           �t�bhhK ��h��R�(KK��h�C    �   
   h  d           �t�bhhK ��h��R�(KK��h�Cd!      �  �   '        h     $      :        �  '   ?   C  ]  ^  $      �         �t�bhhK ��h��R�(KK��h�CX   5   4   i   $  
   �  	   �     �  �   _     `     a        h        �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK	��h�C$   
   b  c                 �t�bhhK ��h��R�(KK��h�C�   �      ,     �t�bhhK ��h��R�(KK��h�C`�   �      �          N     $   ?   �      :   �     �     �   �   
   #        �t�bhhK ��h��R�(KK��h�CH,     d        N     $         �     �  �     �        �t�bhhK ��h��R�(KK��h�C8�  $      �      �  ?     �  �     �        �t�bhhK ��h��R�(KK��h�CH�     �   �      ,     �        5   4   �   /      %        �t�bhhK ��h��R�(KK��h�CD   �  $  e       �  	      F   �   	   �              �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C,     |      �   r                 �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CT!      �   -   �     f        g     �     H  $           �         �t�bhhK ��h��R�(KK��h�C     v        �t�bhhK ��h��R�(KK��h�CT      �  a   z   �  )   	   h              v      z   I  W   $         �t�bhhK ��h��R�(KK��h�C`      �      
           `   
   i     j     	      ,     -   �   
   �        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�Ck                 �t�bhhK ��h��R�(KK��h�C!     $      �t�bhhK ��h��R�(KK ��h�C�
      �  r   $      �      5        l     z   	      F   N      6   9  �   	         =   m     n           �t�bhhK ��h��R�(KK��h�Co             �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C!     �           �t�bhhK ��h��R�(KK��h�C  "     �t�bhhK ��h��R�(KK��h�CD
      5     "     �   	         =   #  �     i        �t�bhhK ��h��R�(KK��h�C&   �  p             �t�bhhK ��h��R�(KK��h�C         o      z      �t�bhhK ��h��R�(KK��h�C$  q        �t�bhhK ��h��R�(KK��h�Cr           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C<+      �      J     �  	   s  t     )            �t�bhhK ��h��R�(KK��h�C,      K     �t�bhhK ��h��R�(KK��h�C\
      u      r   $      J   u  5   v     w     +   	   6      =      %        �t�bhhK ��h��R�(KK��h�C(   x  y     �t�bhhK ��h��R�(KK	��h�C$C       y      z     	     �t�bhhK ��h��R�(KK��h�C�          �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C(   {     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C|           �t�bhhK ��h��R�(KK��h�Cl   j   �   &       !   7         
   u   }     !   .      +       @      n      _   ,         �t�bhhK ��h��R�(KK��h�CL   
   n      _   ,      -      j   '  '     _   ,      ~        �t�bhhK ��h��R�(KK��h�CX   j   �   �     m      �         
   u   B      @   +      ,              �t�bhhK ��h��R�(KK��h�Cm      �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C�   f     �t�bhhK ��h��R�(KK��h�Co      $      �t�bhhK ��h��R�(KK��h�C,      K     �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�Cm      �t�bhhK ��h��R�(KK��h�C8�  �  6      d  $  g                    �t�bhhK ��h��R�(KK	��h�C$e  �     �                 �t�bhhK ��h��R�(KK��h�C,      $  g     ,  �     a        �t�bhhK ��h��R�(KK	��h�C$      7         	  2         �t�bhhK ��h��R�(KK��h�C D   M  N  O     �         �t�bhhK ��h��R�(KK��h�C�  h  	   �  �      �t�bhhK ��h��R�(KK��h�CP  !      �t�bhhK ��h��R�(KK��h�C         m         �t�bhhK ��h��R�(KK
��h�C(  
   �     O  p  �           �t�bhhK ��h��R�(KK��h�C Q     �                 �t�bhhK ��h��R�(KK��h�C%   �        �t�bhhK ��h��R�(KK	��h�C$   
   R  �                 �t�bhhK ��h��R�(KK��h�C�   �   �        �t�bhhK ��h��R�(KK��h�C   
   �  �     E      �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C4d     e     �   �   g     !   f  �        �t�bhhK ��h��R�(KK��h�CD�     i   
   b   ?     D      &   �  S  �   .   g        �t�bhhK ��h��R�(KK��h�CP`      �     h  �     �  T  �     	   i     M                �t�bhhK ��h��R�(KK��h�C(   U     �t�bhhK ��h��R�(KK��h�C         b         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
              �t�bhhK ��h��R�(KK	��h�C$    i   
                    �t�bhhK ��h��R�(KK��h�CT
      "   $      6   j  /   �      �      �             !            �t�bhhK ��h��R�(KK��h�C<H  �  '   k  
   �  �   	   l  	   �     �        �t�bhhK ��h��R�(KK��h�C,�  p   -   f      �     6   V        �t�bhhK ��h��R�(KK��h�C,P     �  7         !   Q   2         �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C$      b         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C �                       �t�bhhK ��h��R�(KK��h�C�   f     �t�bhhK ��h��R�(KK��h�C4W  
   �   f  �  U        X     1         �t�bhhK ��h��R�(KK��h�Cl   6     �   �  	   f     W   Y       �      Z           $  �     �  M     /         �t�bhhK ��h��R�(KK��h�Cl      �     
        �   f  	   [     \  
   z      j   �      N   '   $   �     1         �t�bhhK ��h��R�(KK��h�Co      $      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CD   j   �   P     !   7         
   �      $      !         �t�bhhK ��h��R�(KK��h�Co     �t�bhhK ��h��R�(KK��h�CP
      �   �   
   '   ?     $   	         @   o       �           �t�bhhK ��h��R�(KK��h�C    �   
   h  d           �t�bhhK ��h��R�(KK��h�Cd!      �  �   '        h     $      :        �  '   ?   C  ]  ^  $      �         �t�bhhK ��h��R�(KK��h�CX   5   4   i   $  
   �  	   �     �  �   _     `     a        h        �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK	��h�C$   
   b  c                 �t�bhhK ��h��R�(KK��h�C�   �      ,     �t�bhhK ��h��R�(KK��h�C`�   �      �          N     $   ?   �      :   �     �     �   �   
   #        �t�bhhK ��h��R�(KK��h�CH,     d        N     $         �     �  �     �        �t�bhhK ��h��R�(KK��h�C8�  $      �      �  ?     �  �     �        �t�bhhK ��h��R�(KK��h�CH�     �   �      ,     �        5   4   �   /      %        �t�bhhK ��h��R�(KK��h�CD   �  $  e       �  	      F   �   	   �              �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C,     |      �   r                 �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CT!      �   -   �     f        g     �     H  $           �         �t�bhhK ��h��R�(KK��h�C     v        �t�bhhK ��h��R�(KK��h�CT      �  a   z   �  )   	   h              v      z   I  W   $         �t�bhhK ��h��R�(KK��h�C`      �      
           `   
   i     j     	      ,     -   �   
   �        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�Ck                 �t�bhhK ��h��R�(KK��h�C!     $      �t�bhhK ��h��R�(KK ��h�C�
      �  r   $      �      5        l     z   	      F   N      6   9  �   	         =   m     n           �t�bhhK ��h��R�(KK��h�Co             �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C!     �           �t�bhhK ��h��R�(KK��h�C  "     �t�bhhK ��h��R�(KK��h�CD
      5     "     �   	         =   #  �     i        �t�bhhK ��h��R�(KK��h�C&   �  p             �t�bhhK ��h��R�(KK��h�C         o      z      �t�bhhK ��h��R�(KK��h�C$  q        �t�bhhK ��h��R�(KK��h�Cr           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C<+      �      J     �  	   s  t     )            �t�bhhK ��h��R�(KK��h�C,      K     �t�bhhK ��h��R�(KK��h�C\
      u      r   $      J   u  5   v     w     +   	   6      =      %        �t�bhhK ��h��R�(KK��h�C(   x  y     �t�bhhK ��h��R�(KK	��h�C$C       y      z     	     �t�bhhK ��h��R�(KK��h�C�          �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C(   {     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C|           �t�bhhK ��h��R�(KK��h�Cl   j   �   &       !   7         
   u   }     !   .      +       @      n      _   ,         �t�bhhK ��h��R�(KK��h�CL   
   n      _   ,      -      j   '  '     _   ,      ~        �t�bhhK ��h��R�(KK��h�CX   j   �   �     m      �         
   u   B      @   +      ,              �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C0   !      ;         .  N     �         �t�bhhK ��h��R�(KK	��h�C$   O      
   #     ;        �t�bhhK ��h��R�(KK��h�C;  �           �t�bhhK ��h��R�(KK
��h�C(N      �   �   
      N     �      �t�bhhK ��h��R�(KK��h�ChN        5   �  +      �     �  �     �  	      .   �      @   V      |     ]        �t�bhhK ��h��R�(KK��h�C,;  |  �              �   �        �t�bhhK ��h��R�(KK��h�C         �           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�Cm      �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C�   f     �t�bhhK ��h��R�(KK��h�Co      $      �t�bhhK ��h��R�(KK��h�C,      K     �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�Cm      �t�bhhK ��h��R�(KK��h�C8�  �  6      d  $  g                    �t�bhhK ��h��R�(KK	��h�C$e  �     �                 �t�bhhK ��h��R�(KK��h�C,      $  g     ,  �     a        �t�bhhK ��h��R�(KK	��h�C$      7         	  2         �t�bhhK ��h��R�(KK��h�C D   M  N  O     �         �t�bhhK ��h��R�(KK��h�C�  h  	   �  �      �t�bhhK ��h��R�(KK��h�CP  !      �t�bhhK ��h��R�(KK��h�C         m         �t�bhhK ��h��R�(KK��h�C0  
   �     O  p  �                 �t�bhhK ��h��R�(KK��h�C Q     �                 �t�bhhK ��h��R�(KK��h�C%   �        �t�bhhK ��h��R�(KK	��h�C$   
   R  �                 �t�bhhK ��h��R�(KK��h�C�   �   �        �t�bhhK ��h��R�(KK��h�C   
   �  �     E      �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C4d     e     �   �   g     !   f  �        �t�bhhK ��h��R�(KK��h�CD�     i   
   b   ?     D      &   �  S  �   .   g        �t�bhhK ��h��R�(KK��h�CP`      �     h  �     �  T  �     	   i     M                �t�bhhK ��h��R�(KK��h�C(   U     �t�bhhK ��h��R�(KK��h�C         b         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
              �t�bhhK ��h��R�(KK	��h�C$    i   
                    �t�bhhK ��h��R�(KK��h�CT
      "   $      6   j  /   �      �      �             !            �t�bhhK ��h��R�(KK��h�C<H  �  '   k  
   �  �   	   l  	   �     �        �t�bhhK ��h��R�(KK��h�C,�  p   -   f      �     6   V        �t�bhhK ��h��R�(KK��h�C,P     �  7         !   Q   2         �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C$      b         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C �                       �t�bhhK ��h��R�(KK��h�C�   f     �t�bhhK ��h��R�(KK��h�C4W  
   �   f  �  U        X     1         �t�bhhK ��h��R�(KK��h�Cl   6     �   �  	   f     W   Y       �      Z           $  �     �  M     /         �t�bhhK ��h��R�(KK��h�Cl      �     
        �   f  	   [     \  
   z      j   �      N   '   $   �     1         �t�bhhK ��h��R�(KK��h�Co      $      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CD   j   �   P     !   7         
   �      $      !         �t�bhhK ��h��R�(KK��h�Co     �t�bhhK ��h��R�(KK��h�CP
      �   �   
   '   ?     $   	         @   o       �           �t�bhhK ��h��R�(KK��h�C    �   
   h  d           �t�bhhK ��h��R�(KK��h�Cd!      �  �   '        h     $      :        �  '   ?   C  ]  ^  $      �         �t�bhhK ��h��R�(KK��h�CX   5   4   i   $  
   �  	   �     �  �   _     `     a        h        �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK	��h�C$   
   b  c                 �t�bhhK ��h��R�(KK��h�C�   �      ,     �t�bhhK ��h��R�(KK��h�C`�   �      �          N     $   ?   �      :   �     �     �   �   
   #        �t�bhhK ��h��R�(KK��h�CH,     d        N     $         �     �  �     �        �t�bhhK ��h��R�(KK��h�C8�  $      �      �  ?     �  �     �        �t�bhhK ��h��R�(KK��h�CH�     �   �      ,     �        5   4   �   /      %        �t�bhhK ��h��R�(KK��h�CD   �  $  e       �  	      F   �   	   �              �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C,     |      �   r                 �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CT!      �   -   �     f        g     �     H  $           �         �t�bhhK ��h��R�(KK��h�C     v        �t�bhhK ��h��R�(KK��h�CT      �  a   z   �  )   	   h              v      z   I  W   $         �t�bhhK ��h��R�(KK��h�C`      �      
           `   
   i     j     	      ,     -   �   
   �        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�Ck                 �t�bhhK ��h��R�(KK��h�C!     $      �t�bhhK ��h��R�(KK ��h�C�
      �  r   $      �      5        l     z   	      F   N      6   9  �   	         =   m     n           �t�bhhK ��h��R�(KK��h�Co             �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C!     �           �t�bhhK ��h��R�(KK��h�C  "     �t�bhhK ��h��R�(KK��h�CD
      5     "     �   	         =   #  �     i        �t�bhhK ��h��R�(KK��h�C&   �  p             �t�bhhK ��h��R�(KK��h�C         o      z      �t�bhhK ��h��R�(KK��h�C$  q        �t�bhhK ��h��R�(KK��h�Cr           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C<+      �      J     �  	   s  t     )            �t�bhhK ��h��R�(KK��h�C,      K     �t�bhhK ��h��R�(KK��h�C\
      u      r   $      J   u  5   v     w     +   	   6      =      %        �t�bhhK ��h��R�(KK��h�C(   x  y     �t�bhhK ��h��R�(KK	��h�C$C       y      z     	     �t�bhhK ��h��R�(KK��h�C�          �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C(   {     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C|           �t�bhhK ��h��R�(KK��h�Cl   j   �   &       !   7         
   u   }     !   .      +       @      n      _   ,         �t�bhhK ��h��R�(KK��h�CL   
   n      _   ,      -      j   '  '     _   ,      ~        �t�bhhK ��h��R�(KK��h�CX   j   �   �     m      �         
   u   B      @   +      ,              �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C0   !      ;         .  N     �         �t�bhhK ��h��R�(KK	��h�C$   O      
   #     ;        �t�bhhK ��h��R�(KK��h�C;  �           �t�bhhK ��h��R�(KK
��h�C(N      �   �   
      N     �      �t�bhhK ��h��R�(KK��h�ChN        5   �  +      �     �  �     �  	      .   �      @   V      |     ]        �t�bhhK ��h��R�(KK��h�C,;  |  �              �   �        �t�bhhK ��h��R�(KK��h�C         �           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�     !      �t�bhhK ��h��R�(KK��h�C�   �     �t�bhhK ��h��R�(KK��h�Cn   G      �t�bhhK ��h��R�(KK��h�C�   �  G      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�   G      �t�bhhK ��h��R�(KK��h�C4  G      �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�     !      �t�bhhK ��h��R�(KK��h�Cp
      5      
   �  	         �         (      <         	   C       y      �     /        �t�bhhK ��h��R�(KK��h�C8M   q         D   �   
   �     o      �        �t�bhhK ��h��R�(KK
��h�C(      �  )   	                  �t�bhhK ��h��R�(KK��h�C         G         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C@
      "   J   S     !   	         �  :   �   �        �t�bhhK ��h��R�(KK��h�C<�   �   8     F      5  	   �  	   Q     �         �t�bhhK ��h��R�(KK��h�Ch
      q  �     
      �  �         �  	   O        (  -   
   J   S  4      !         �t�bhhK ��h��R�(KK��h�C8   !      >  5     )        u  �   �         �t�bhhK ��h��R�(KK��h�C,�  "   �   \  y      u     	        �t�bhhK ��h��R�(KK��h�Cp�        2      �            �   w        w     <               J   �                     �t�bhhK ��h��R�(KK��h�CH
      5     o     E  	   6      �   �   .  �   &   m        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C�  �   	      1     �t�bhhK ��h��R�(KK��h�C�  �   	      �     �t�bhhK ��h��R�(KK��h�C�  �   	      C     �t�bhhK ��h��R�(KK��h�C�  �   	      1     �t�bhhK ��h��R�(KK��h�C�  �   	   �  �     �t�bhhK ��h��R�(KK
��h�C(�     7            �   �        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�Ct                 �t�bhhK ��h��R�(KK��h�C�   �     �t�bhhK ��h��R�(KK��h�C,   !      ^   *     T   �   �         �t�bhhK ��h��R�(KK��h�C\              �   �  -   
      4   "   �       �   &   �   �  ;      1         �t�bhhK ��h��R�(KK��h�C0      �   �  �      �  3  ~  %        �t�bhhK ��h��R�(KK��h�C<   �  �  +  ,     �       �     �   (        �t�bhhK ��h��R�(KK��h�C�   �                 �t�bhhK ��h��R�(KK	��h�C$�   �                 E      �t�bhhK ��h��R�(KK��h�C�   �                 �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C�   �                 �t�bhhK ��h��R�(KK��h�C-     �t�bhhK ��h��R�(KK��h�C4   
   �     -  7         j   �   �        �t�bhhK ��h��R�(KK��h�CU        �t�bhhK ��h��R�(KK��h�C�  �      �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�CL   9      3  X  	   v   Y      �     1   �   >     @   �        �t�bhhK ��h��R�(KK
��h�C(�      3  X     v     Q        �t�bhhK ��h��R�(KK��h�C03  X  �  4   Q     �     W   {        �t�bhhK ��h��R�(KK��h�C4       �  Q  �  4   �  �      �  �        �t�bhhK ��h��R�(KK	��h�C$l     9   3  �     �        �t�bhhK ��h��R�(KK	��h�C$   �     @       <        �t�bhhK ��h��R�(KK��h�C          �      1         �t�bhhK ��h��R�(KK��h�C@�     �           E      �      �      �     �     �t�bhhK ��h��R�(KK��h�C,   �  	        �     �  �        �t�bhhK ��h��R�(KK��h�C4�     z        �     �      �           �t�bhhK ��h��R�(KK��h�C �      x        �   �      �t�bhhK ��h��R�(KK��h�C4   !      �      -  �      .  �           �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C�  C     �t�bhhK ��h��R�(KK��h�C(        �t�bhhK ��h��R�(KK��h�CD
          /  	         -   �     z  �     �         �t�bhhK ��h��R�(KK��h�C8      
   �  7         !   Q   2   
   �         �t�bhhK ��h��R�(KK
��h�C(   �  �     .   �  �   �         �t�bhhK ��h��R�(KK��h�C          �      1         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�Cn   G      �t�bhhK ��h��R�(KK��h�C@   �     $   ?   �   O   B   +      0     �           �t�bhhK ��h��R�(KK��h�CDv         �   
   f      @   V      �     �     $         �t�bhhK ��h��R�(KK��h�CD   �  6  �   G   	   �     �  y     v   V  -            �t�bhhK ��h��R�(KK
��h�C(P     0  7         !   2         �t�bhhK ��h��R�(KK��h�CTM   j  �        �   }      �     �   ?  
   f   �  �     n   G         �t�bhhK ��h��R�(KK
��h�C(�     s        <               �t�bhhK ��h��R�(KK��h�CP&      x  C     #  y      �     h       y      �     r        �t�bhhK ��h��R�(KK��h�C �  "   �   
   �  G         �t�bhhK ��h��R�(KK
��h�C(      7         !   Q   2         �t�bhhK ��h��R�(KK��h�CD
   '   $       �  	   6      w   �      �      �         �t�bhhK ��h��R�(KK
��h�C(   �  �     .   �  �   �         �t�bhhK ��h��R�(KK��h�C         n   G         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C b     �                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
   K                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�Ct                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�   �  G      �t�bhhK ��h��R�(KK
��h�C(�     �    �         W         �t�bhhK ��h��R�(KK��h�CT�      .      !   �  ;      �         O      
   M   ;     �           �t�bhhK ��h��R�(KK��h�C(         <      �     �t�bhhK ��h��R�(KK��h�C8      
   �      �   7         !   Q   2         �t�bhhK ��h��R�(KK��h�C,         �   �  G                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK
��h�C(   
   ;      "                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C,�     S     �  	   C  �     )      �t�bhhK ��h��R�(KK
��h�C(N      �   �   
      N     �      �t�bhhK ��h��R�(KK��h�ChN        5   �  +      �     �  �     �  	      .   �      @   V      |     ]        �t�bhhK ��h��R�(KK��h�C �     |     �   ;        �t�bhhK ��h��R�(KK��h�C(         <      �     �t�bhhK ��h��R�(KK��h�C4�     |     Y   ?   A  I      �   �        �t�bhhK ��h��R�(KK��h�C(         <      �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�CV      �           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CX  �      �t�bhhK ��h��R�(KK��h�C8�     !   �      �           <      �        �t�bhhK ��h��R�(KK��h�C        �         �t�bhhK ��h��R�(KK��h�CC     #  �     h     �t�bhhK ��h��R�(KK��h�C          �     p        �t�bhhK ��h��R�(KK��h�C8
   r      4      �   	   �   g  y      �        �t�bhhK ��h��R�(KK��h�CT
   q            	         �   '      
       �        '   �           �t�bhhK ��h��R�(KK��h�CL
      5     �            	   6      �     i  �  &   m        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�CD?   �     B     �     1  �        W       9         �t�bhhK ��h��R�(KK��h�C(      <      �        �t�bhhK ��h��R�(KK��h�C4�  �     1  �           2  �   3        �t�bhhK ��h��R�(KK	��h�C$2  �   3  	   �     �  �     �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK
��h�C(�  �  �     �                 �t�bhhK ��h��R�(KK��h�Cn   �      �t�bhhK ��h��R�(KK��h�CX
   �     $   ?   �   O            J     �           �     �           �t�bhhK ��h��R�(KK��h�C@$   ?   _  I   �     V     �       <     �        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   �     �     �t�bhhK ��h��R�(KK��h�C�   �     �t�bhhK ��h��R�(KK��h�C    !      D   �   �        �t�bhhK ��h��R�(KK��h�CT
      4   "   �       �   :   �   �  	         g   /         �   �        �t�bhhK ��h��R�(KK��h�C0d      �   �  �      �  3  ~  %        �t�bhhK ��h��R�(KK��h�C<   �  �  +  ,     �       �     �   �         �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�  Y     �t�bhhK ��h��R�(KK��h�C�   G      �t�bhhK ��h��R�(KK��h�CH
      5   q  +      V   	   6      =   J   �      )           �t�bhhK ��h��R�(KK	��h�C$   �   Z  :   �  C  �        �t�bhhK ��h��R�(KK��h�C,U   �         �  ^  �     �        �t�bhhK ��h��R�(KK��h�C`
   �   4   "   �      d       	   6      =   U     -  �      .  �  �           �t�bhhK ��h��R�(KK��h�C�  C     �t�bhhK ��h��R�(KK��h�C(      <            �t�bhhK ��h��R�(KK��h�CD
      5   �  �  	         D   w   �      0      �         �t�bhhK ��h��R�(KK��h�C&   "   �   �   �         �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C(      <      +     �t�bhhK ��h��R�(KK��h�C         �   G         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
   4                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�Ct                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C 0                       �t�bhhK ��h��R�(KK��h�C4  G      �t�bhhK ��h��R�(KK��h�Cp
      �   "      
   �  	   �  	   4  G      �  	         =   �     �        }              �t�bhhK ��h��R�(KK��h�C0�        �         G        �        �t�bhhK ��h��R�(KK��h�C    �   �  }      �        �t�bhhK ��h��R�(KK��h�C      v     Q        �t�bhhK ��h��R�(KK
��h�C(   
   �         !   Q   2         �t�bhhK ��h��R�(KK��h�Ch�      }   d      @     0  
      5   
                 
      �  �                 �t�bhhK ��h��R�(KK��h�CP�      }   d      �  
         F   "   ,                           �t�bhhK ��h��R�(KK
��h�C(   �    -   �                 �t�bhhK ��h��R�(KK��h�C,      -   �   t     �     9         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     5              �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�Ct                 �t�bhhK ��h��R�(KK��h�C�      ~   q  �        �t�bhhK ��h��R�(KK��h�C t     [                 �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�CD   \     �     6  �  	   ]     �  A  ^  ?   �        �t�bhhK ��h��R�(KK��h�C8=   �     �     N      _            �        �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C@C     #  y      �     h       y      �     r     �t�bhhK ��h��R�(KK��h�CPM   j  �        �   }      �     �   ?  
   f   �  �     T        �t�bhhK ��h��R�(KK��h�CT      
   �     T  7         !   Q   D           �                 �t�bhhK ��h��R�(KK	��h�C$         N      u  $         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     5           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C         T        �t�bhhK ��h��R�(KK��h�C�      ~   q  �        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�      ~   q        �t�bhhK ��h��R�(KK��h�C`  a                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK'��h�C�      @   ;      �      �     
            �     /   "      �        {     �  �  	   �  �      D  a   �        3  T  �         �t�bhhK ��h��R�(KK��h�CH;      �         F     �  	     	   �     �     ~        �t�bhhK ��h��R�(KK��h�CLw   �      �     �  r   �     V   	        ;   �  J   �        �t�bhhK ��h��R�(KK��h�C�  y      �     h     �t�bhhK ��h��R�(KK��h�C(         <      �     �t�bhhK ��h��R�(KK��h�C         �   Y         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C�     !      �t�bhhK ��h��R�(KK��h�Cn   G      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�   G      �t�bhhK ��h��R�(KK��h�C4  G      �     �t�bhhK ��h��R�(KK��h�C�     T     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�     !      �t�bhhK ��h��R�(KK��h�C.   �  �      �         �t�bhhK ��h��R�(KK��h�CD�   �   x  
   .      
   '   �  	      F        L        �t�bhhK ��h��R�(KK��h�C4
   J   S     !         �   t  �   �         �t�bhhK ��h��R�(KK��h�C<�   �   8     F      5  	   �  	   Q     �         �t�bhhK ��h��R�(KK��h�C\
      q       �  �         �  O        (  -   
   J   S  4      !         �t�bhhK ��h��R�(KK��h�C\
      4   "   �       �   :   �   �     }  	         �   }         �   �        �t�bhhK ��h��R�(KK��h�C          �      1         �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C4l     &   �  s     �     !               �t�bhhK ��h��R�(KK��h�C\      �   �  �  
      5   c               {     �   �      �     {        �t�bhhK ��h��R�(KK��h�C4q   "   �   �     �  y      �     /        �t�bhhK ��h��R�(KK��h�C,   !      >  5     u  �   �         �t�bhhK ��h��R�(KK��h�C,   �     N  	   O     P  Q        �t�bhhK ��h��R�(KK��h�C<
      q            .     ,     a  �         �t�bhhK ��h��R�(KK��h�C0.                  �   .     �        �t�bhhK ��h��R�(KK��h�C,�  "   �   \  y      u     	        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�Ct                 �t�bhhK ��h��R�(KK��h�C�   �     �t�bhhK ��h��R�(KK��h�C,   !      ^   *     T   �   �         �t�bhhK ��h��R�(KK��h�C\              �   �  -   
      4   "   �       �   &   �   �  ;      1         �t�bhhK ��h��R�(KK��h�C0      �   �  �      �  3  ~  %        �t�bhhK ��h��R�(KK��h�C<   �  �  +  ,     �       �     �   (        �t�bhhK ��h��R�(KK��h�C          �      1         �t�bhhK ��h��R�(KK��h�C�   �                 �t�bhhK ��h��R�(KK	��h�C$�   �                 E      �t�bhhK ��h��R�(KK��h�C�   �                 �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C�   �                 �t�bhhK ��h��R�(KK��h�C-     �t�bhhK ��h��R�(KK��h�C4   
   �     -  7         j   �   �        �t�bhhK ��h��R�(KK��h�CU        �t�bhhK ��h��R�(KK��h�C�  �      �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�CL   9      3  X  	   v   Y      �     1   �   >     @   �        �t�bhhK ��h��R�(KK
��h�C(�      3  X     v     Q        �t�bhhK ��h��R�(KK��h�C03  X  �  4   Q     �     W   {        �t�bhhK ��h��R�(KK��h�C4       �  Q  �  4   �  �      �  �        �t�bhhK ��h��R�(KK	��h�C$l     9   3  �     �        �t�bhhK ��h��R�(KK	��h�C$   �     @       <        �t�bhhK ��h��R�(KK��h�C@�     �           E      �      �      �     �     �t�bhhK ��h��R�(KK��h�C,   �  	        �     �  �        �t�bhhK ��h��R�(KK��h�CX
      q       �  �         �     4         z  �   m  	   =   �         �t�bhhK ��h��R�(KK��h�C4   !      �      -  �      .  �           �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C�  C     �t�bhhK ��h��R�(KK��h�C(        �t�bhhK ��h��R�(KK��h�CD
          /  	         -   �     z  �     �         �t�bhhK ��h��R�(KK��h�C8      
   �  7         !   Q   2   
   �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�Cn   G      �t�bhhK ��h��R�(KK��h�C@   �     $   ?   �   O   B   +      0     �           �t�bhhK ��h��R�(KK	��h�C$l     0     !               �t�bhhK ��h��R�(KK��h�CP      �      }      L     �   
   f   
      "   �   :  �   G         �t�bhhK ��h��R�(KK��h�C �  "   �   
   �  G         �t�bhhK ��h��R�(KK
��h�C(      7         !   Q   2         �t�bhhK ��h��R�(KK��h�C0
   '   $   q    	   6      =   �         �t�bhhK ��h��R�(KK��h�C4�  "   �   �     �  y      �     /        �t�bhhK ��h��R�(KK��h�C0N   �   "   �  6      =   �      �        �t�bhhK ��h��R�(KK��h�C,�   �   x  �   
   $      �            �t�bhhK ��h��R�(KK��h�Cl     �              �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C,      -   w   z         �   �        �t�bhhK ��h��R�(KK��h�C8   !      Z   �   *     -   �   �   
   $         �t�bhhK ��h��R�(KK��h�C         n   G         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C b     �                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
   K                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�Ct                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CX  �      �t�bhhK ��h��R�(KK��h�C8�     !   �      �           <      �        �t�bhhK ��h��R�(KK��h�C8
      4   5   �   �   	   �   g  y      �        �t�bhhK ��h��R�(KK��h�CL
      5   �   �   	   6      �     i  �  &   m  y      �        �t�bhhK ��h��R�(KK��h�CH�     �   o         �  �   �     �  y      �     p        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�CD?   �     B     �     1  �        W       9         �t�bhhK ��h��R�(KK��h�Cl              �t�bhhK ��h��R�(KK��h�CL  "   �   \  y      p     F        B  y      �     F        �t�bhhK ��h��R�(KK��h�C4�  �     1  �           2  �   3        �t�bhhK ��h��R�(KK	��h�C$2  �   3  	   �     �  �     �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK
��h�C(�  �  �     �                 �t�bhhK ��h��R�(KK��h�Cn   �      �t�bhhK ��h��R�(KK��h�CX
   �     $   ?   �   O            J     �           �     �           �t�bhhK ��h��R�(KK��h�C@$   ?   _  I   �     V     �       <     �        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   �     �     �t�bhhK ��h��R�(KK��h�C�   �     �t�bhhK ��h��R�(KK��h�C    !      D   �   �        �t�bhhK ��h��R�(KK��h�CT
      4   "   �       �   :   �   �  	         g   /         �   �        �t�bhhK ��h��R�(KK��h�C0d      �   �  �      �  3  ~  %        �t�bhhK ��h��R�(KK��h�C<   �  �  +  ,     �       �     �   �         �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�  Y     �t�bhhK ��h��R�(KK��h�C�   G      �t�bhhK ��h��R�(KK��h�CH
      5   q  +      V   	   6      =   J   �      )           �t�bhhK ��h��R�(KK	��h�C$   �   Z  :   �  C  �        �t�bhhK ��h��R�(KK��h�C,U   �         �  ^  �     �        �t�bhhK ��h��R�(KK��h�C`
   �   4   "   �      d       	   6      =   U     -  �      .  �  �           �t�bhhK ��h��R�(KK��h�C�  C     �t�bhhK ��h��R�(KK��h�C(        �t�bhhK ��h��R�(KK��h�CD
      5   �  �  	         D   w   �      0      �         �t�bhhK ��h��R�(KK��h�C&   "   �   �   �         �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C(      <      +     �t�bhhK ��h��R�(KK��h�C         �   G         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
   4                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�Ct                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C 0                       �t�bhhK ��h��R�(KK��h�C4  G      �     �t�bhhK ��h��R�(KK��h�CX
      5   
     �     u         "      �  	         =   �     �        �t�bhhK ��h��R�(KK��h�C       �   }   �   ]         �t�bhhK ��h��R�(KK��h�C�              �t�bhhK ��h��R�(KK��h�CL
      "      �        -   �   t     �     9         �         �t�bhhK ��h��R�(KK
��h�C(!   T   �   ?   O  I   �  
        �t�bhhK ��h��R�(KK��h�C\-   L   �   ?   �  I      @   �  
  
   :   �  �  
  �                       �t�bhhK ��h��R�(KK	��h�C$         4  G      �        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     5              �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�Ct                 �t�bhhK ��h��R�(KK��h�C�      ~   q  �        �t�bhhK ��h��R�(KK��h�C t     [                 �t�bhhK ��h��R�(KK��h�C�     T     �t�bhhK ��h��R�(KK��h�CD   \     �     6  �  	   ]     �  A  ^  ?   �        �t�bhhK ��h��R�(KK��h�C8=   �     �     N      _            �        �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�CPM   j  �        �   }      �     �   ?  
   f   �  �     T        �t�bhhK ��h��R�(KK��h�C<         �     T        '   $   �     1         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     5           �t�bhhK ��h��R�(KK��h�C�      ~   q  �        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�      ~   q        �t�bhhK ��h��R�(KK��h�C`  a                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK'��h�C�      @   ;      �      �     
            �     /   "      �        {     �  �  	   �  �      D  a   �        3  T  �         �t�bhhK ��h��R�(KK��h�CH;      �         F     �  	     	   �     �     ~        �t�bhhK ��h��R�(KK��h�CLw   �      �     �  r   �     V   	        ;   �  J   �        �t�bhhK ��h��R�(KK��h�C�  y      �     h     �t�bhhK ��h��R�(KK��h�C(         <      �     �t�bhhK ��h��R�(KK��h�C         �   Y         �t�b�       hhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C�     !      �t�bhhK ��h��R�(KK��h�Cn   G      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�   G      �t�bhhK ��h��R�(KK��h�C4  G      �     �t�bhhK ��h��R�(KK��h�C�     T     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�     !      �t�bhhK ��h��R�(KK��h�C.   �  �      �         �t�bhhK ��h��R�(KK��h�CD�   �   x  
   .      
   '   �  	      F        L        �t�bhhK ��h��R�(KK��h�C4
   J   S     !         �   t  �   �         �t�bhhK ��h��R�(KK��h�C<�   �   8     F      5  	   �  	   Q     �         �t�bhhK ��h��R�(KK��h�C\
      q       �  �         �  O        (  -   
   J   S  4      !         �t�bhhK ��h��R�(KK��h�C\
      4   "   �       �   :   �   �     }  	         �   }         �   �        �t�bhhK ��h��R�(KK��h�C          �      1         �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C4l     &   �  s     �     !               �t�bhhK ��h��R�(KK��h�C\      �   �  �  
      5   c               {     �   �      �     {        �t�bhhK ��h��R�(KK��h�C4q   "   �   �     �  y      �     /        �t�bhhK ��h��R�(KK��h�C,   !      >  5     u  �   �         �t�bhhK ��h��R�(KK��h�C,   �     N  	   O     P  Q        �t�bhhK ��h��R�(KK��h�C<
      q            .     ,     a  �         �t�bhhK ��h��R�(KK��h�C0.                  �   .     �        �t�bhhK ��h��R�(KK��h�C,�  "   �   \  y      u     	        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�Ct                 �t�bhhK ��h��R�(KK��h�C�   �     �t�bhhK ��h��R�(KK��h�C,   !      ^   *     T   �   �         �t�bhhK ��h��R�(KK��h�C\              �   �  -   
      4   "   �       �   &   �   �  ;      1         �t�bhhK ��h��R�(KK��h�C0      �   �  �      �  3  ~  %        �t�bhhK ��h��R�(KK��h�C<   �  �  +  ,     �       �     �   (        �t�bhhK ��h��R�(KK��h�C          �      1         �t�bhhK ��h��R�(KK��h�C�   �                 �t�bhhK ��h��R�(KK	��h�C$�   �                 E      �t�bhhK ��h��R�(KK��h�C�   �                 �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C�   �                 �t�bhhK ��h��R�(KK��h�C-     �t�bhhK ��h��R�(KK��h�C4   
   �     -  7         j   �   �        �t�bhhK ��h��R�(KK��h�CU        �t�bhhK ��h��R�(KK��h�C�  �      �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�CL   9      3  X  	   v   Y      �     1   �   >     @   �        �t�bhhK ��h��R�(KK
��h�C(�      3  X     v     Q        �t�bhhK ��h��R�(KK��h�C03  X  �  4   Q     �     W   {        �t�bhhK ��h��R�(KK��h�C4       �  Q  �  4   �  �      �  �        �t�bhhK ��h��R�(KK	��h�C$l     9   3  �     �        �t�bhhK ��h��R�(KK	��h�C$   �     @       <        �t�bhhK ��h��R�(KK��h�C@�     �           E      �      �      �     �     �t�bhhK ��h��R�(KK��h�C,   �  	        �     �  �        �t�bhhK ��h��R�(KK��h�CX
      q       �  �         �     4         z  �   m  	   =   �         �t�bhhK ��h��R�(KK��h�C4   !      �      -  �      .  �           �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C�  C     �t�bhhK ��h��R�(KK��h�C(        �t�bhhK ��h��R�(KK��h�CD
          /  	         -   �     z  �     �         �t�bhhK ��h��R�(KK��h�C8      
   �  7         !   Q   2   
   �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�Cn   G      �t�bhhK ��h��R�(KK��h�C@   �     $   ?   �   O   B   +      0     �           �t�bhhK ��h��R�(KK	��h�C$l     0     !               �t�bhhK ��h��R�(KK��h�CP      �      }      L     �   
   f   
      "   �   :  �   G         �t�bhhK ��h��R�(KK��h�C �  "   �   
   �  G         �t�bhhK ��h��R�(KK
��h�C(      7         !   Q   2         �t�bhhK ��h��R�(KK��h�C0
   '   $   q    	   6      =   �         �t�bhhK ��h��R�(KK��h�C4�  "   �   �     �  y      �     /        �t�bhhK ��h��R�(KK��h�C0N   �   "   �  6      =   �      �        �t�bhhK ��h��R�(KK��h�C,�   �   x  �   
   $      �            �t�bhhK ��h��R�(KK��h�Cl     �              �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C,      -   w   z         �   �        �t�bhhK ��h��R�(KK��h�C8   !      Z   �   *     -   �   �   
   $         �t�bhhK ��h��R�(KK��h�C         n   G         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C b     �                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
   K                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�Ct                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CX  �      �t�bhhK ��h��R�(KK��h�C8�     !   �      �           <      �        �t�bhhK ��h��R�(KK��h�C8
      4   5   �   �   	   �   g  y      �        �t�bhhK ��h��R�(KK��h�CL
      5   �   �   	   6      �     i  �  &   m  y      �        �t�bhhK ��h��R�(KK��h�CH�     �   o         �  �   �     �  y      �     p        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�CD?   �     B     �     1  �        W       9         �t�bhhK ��h��R�(KK��h�Cl              �t�bhhK ��h��R�(KK��h�CL  "   �   \  y      p     F        B  y      �     F        �t�bhhK ��h��R�(KK��h�C4�  �     1  �           2  �   3        �t�bhhK ��h��R�(KK	��h�C$2  �   3  	   �     �  �     �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK
��h�C(�  �  �     �                 �t�bhhK ��h��R�(KK��h�Cn   �      �t�bhhK ��h��R�(KK��h�CX
   �     $   ?   �   O            J     �           �     �           �t�bhhK ��h��R�(KK��h�C@$   ?   _  I   �     V     �       <     �        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   �     �     �t�bhhK ��h��R�(KK��h�C�   �     �t�bhhK ��h��R�(KK��h�C    !      D   �   �        �t�bhhK ��h��R�(KK��h�CT
      4   "   �       �   :   �   �  	         g   /         �   �        �t�bhhK ��h��R�(KK��h�C0d      �   �  �      �  3  ~  %        �t�bhhK ��h��R�(KK��h�C<   �  �  +  ,     �       �     �   �         �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�  Y     �t�bhhK ��h��R�(KK��h�C�   G      �t�bhhK ��h��R�(KK��h�CH
      5   q  +      V   	   6      =   J   �      )           �t�bhhK ��h��R�(KK	��h�C$   �   Z  :   �  C  �        �t�bhhK ��h��R�(KK��h�C,U   �         �  ^  �     �        �t�bhhK ��h��R�(KK��h�C`
   �   4   "   �      d       	   6      =   U     -  �      .  �  �           �t�bhhK ��h��R�(KK��h�C�  C     �t�bhhK ��h��R�(KK��h�C(        �t�bhhK ��h��R�(KK��h�CD
      5   �  �  	         D   w   �      0      �         �t�bhhK ��h��R�(KK��h�C&   "   �   �   �         �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C(      <      +     �t�bhhK ��h��R�(KK��h�C         �   G         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
   4                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�Ct                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C 0                       �t�bhhK ��h��R�(KK��h�C4  G      �     �t�bhhK ��h��R�(KK��h�CX
      5   
     �     u         "      �  	         =   �     �        �t�bhhK ��h��R�(KK��h�C       �   }   �   ]         �t�bhhK ��h��R�(KK��h�C�              �t�bhhK ��h��R�(KK��h�CL
      "      �        -   �   t     �     9         �         �t�bhhK ��h��R�(KK
��h�C(!   T   �   ?   O  I   �  
        �t�bhhK ��h��R�(KK��h�C\-   L   �   ?   �  I      @   �  
  
   :   �  �  
  �                       �t�bhhK ��h��R�(KK	��h�C$         4  G      �        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     5              �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�Ct                 �t�bhhK ��h��R�(KK��h�C�      ~   q  �        �t�bhhK ��h��R�(KK��h�C t     [                 �t�bhhK ��h��R�(KK��h�C�     T     �t�bhhK ��h��R�(KK��h�CD   \     �     6  �  	   ]     �  A  ^  ?   �        �t�bhhK ��h��R�(KK��h�C8=   �     �     N      _            �        �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�CPM   j  �        �   }      �     �   ?  
   f   �  �     T        �t�bhhK ��h��R�(KK��h�C<         �     T        '   $   �     1         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�     5           �t�bhhK ��h��R�(KK��h�C�      ~   q  �        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�      ~   q        �t�bhhK ��h��R�(KK��h�C`  a                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK'��h�C�      @   ;      �      �     
            �     /   "      �        {     �  �  	   �  �      D  a   �        3  T  �         �t�bhhK ��h��R�(KK��h�CH;      �         F     �  	     	   �     �     ~        �t�bhhK ��h��R�(KK��h�CLw   �      �     �  r   �     V   	        ;   �  J   �        �t�bhhK ��h��R�(KK��h�C�  y      �     h     �t�bhhK ��h��R�(KK��h�C(         <      �     �t�bhhK ��h��R�(KK��h�C         �   Y         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CV           L      �t�bhhK ��h��R�(KK��h�Cz     �t�bhhK ��h��R�(KK��h�C  �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK
��h�C(   !      �  �     �   �         �t�bhhK ��h��R�(KK��h�C ]  6  D   &   �   &        �t�bhhK ��h��R�(KK��h�C8   !   V  �      )   	      	   E               �t�bhhK ��h��R�(KK��h�C0�   &  V  -   s      )      W   k         �t�bhhK ��h��R�(KK
��h�C(�   �   D   �   �        �        �t�bhhK ��h��R�(KK��h�CLB   6   i   
   �     v  $   w  �   n    z   6   f     &        �t�bhhK ��h��R�(KK��h�CD      i   
         &   �  &  M   �           7        �t�bhhK ��h��R�(KK��h�C8      '  `   5      �   �        '  [        �t�bhhK ��h��R�(KK��h�C,�     �     F      ^     U        �t�bhhK ��h��R�(KK��h�C �   �  �  .     T        �t�bhhK ��h��R�(KK��h�C\�   :  �      `   
   �        &     �          �  �     �     �        �t�bhhK ��h��R�(KK��h�C,�  �   B   
   �     &   �   ]        �t�bhhK ��h��R�(KK��h�CL
   K  �  �  �     9      *   	         D   g   �     �        �t�bhhK ��h��R�(KK��h�C4   6   c  �   �   J   `      &   �   ]        �t�bhhK ��h��R�(KK	��h�C$      7      M   q   �        �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�   �                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�   �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C `   
   d                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK	��h�C$'  x     �                 �t�bhhK ��h��R�(KK	��h�C$   
   &  )                  �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CL�      �     �      �  �     �   �   \      �     �  �        �t�bhhK ��h��R�(KK��h�C8   !      B   @   �      )   	                  �t�bhhK ��h��R�(KK	��h�C$   �   i   
                 �t�bhhK ��h��R�(KK��h�C4`      �  m  M   H   2            7        �t�bhhK ��h��R�(KK��h�Chf          	   5  `      -   �  �     \  	   
   K     F        !   '  ?   �        �t�bhhK ��h��R�(KK��h�CP�   s   8     �     4   "     k     )          D  a              �t�bhhK ��h��R�(KK��h�C8&   �        �     �     H  $      �        �t�bhhK ��h��R�(KK��h�C&   �      �  �        �t�be(hhK ��h��R�(KK��h�C<T  8  z      &   �             �             �t�bhhK ��h��R�(KK��h�Cl   7         
     	   �          
   s      �     �      !   Q      �   9     2         �t�bhhK ��h��R�(KK��h�C,      -   �   
            U        �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C `                       �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
   &   �   �           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK	��h�C$'  x     g                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�      p              �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK��h�C0   !      �     �  �     �           �t�bhhK ��h��R�(KK��h�CD   !      -      �    	   v   B      �   �              �t�bhhK ��h��R�(KK��h�CH      
   �     !   7         !   Q      �   9     2         �t�bhhK ��h��R�(KK	��h�C$�     �  6   �     %        �t�bhhK ��h��R�(KK��h�C�     �             �t�bhhK ��h��R�(KK��h�C<   H   2   7      P     �           
   �        �t�bhhK ��h��R�(KK��h�C         [   X      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�  �      �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�   X   �  h     �t�bhhK ��h��R�(KK��h�Ct
   �   k     .   )   �   4      �  �     R     &   �  �  	      z   @   �   X      �  �           �t�bhhK ��h��R�(KK��h�C8   &   �      �  k  .   )   �      l  �        �t�bhhK ��h��R�(KK��h�C   s  �     '   I         �t�bhhK ��h��R�(KK��h�Cx
      "   �     1         �  }   `     "   $   ?   �   6      w   �      :     r   ;     <           �t�bhhK ��h��R�(KK��h�CD:  �  
   �    �      x   /      �      �  �   �        �t�bhhK ��h��R�(KK��h�C   
   &   �   �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C=     �t�bhhK ��h��R�(KK��h�C[   X      L   C      �t�bhhK ��h��R�(KK��h�CL   !   )     �   m        _     �     H  �  �   l  >        �t�bhhK ��h��R�(KK��h�CX
   B   "   �     �  	      B   �   l  �  D      �  
     �  �           �t�bhhK ��h��R�(KK��h�C[   X      �      �t�bhhK ��h��R�(KK��h�C�  
        �t�bhhK ��h��R�(KK��h�C�     ?     �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK*��h�C�      i      &   [   �  �  	   .   �   �        �  �     �     	   
      �  l  >    I      �    	   5  4   "   �     �      W   �        �t�bhhK ��h��R�(KK��h�CP   �  �        @    �  U   �        O      �     �  R        �t�bhhK ��h��R�(KK��h�CX�     !         �     �  !      �  !        �  �      A  n           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�CC      [   X      �t�bhhK ��h��R�(KK��h�C0   �     !   V  �     ^   >   k         �t�bhhK ��h��R�(KK+��h�C�   �  V  -   X      )      �     �  �  �             "   '   e   f  B  )   	         �  	      �  k     .   )   �   4         *     �        �t�bhhK ��h��R�(KK��h�CXN      �  /      @  	         �  �   /      �     s      J   �   �         �t�bhhK ��h��R�(KK��h�C\      -   �   /        2              �  	         O   U   J   �           �t�bhhK ��h��R�(KK
��h�C(&   �  �  �     &   �   @        �t�bhhK ��h��R�(KK��h�C@s      &   �   �     �   
   �  �     w             �t�bhhK ��h��R�(KK��h�C`      
   �     
   s        �   �   7         H   2      d   �     <           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�Cs      &   �   �     �t�bhhK ��h��R�(KK	��h�C$)      W   k      &   [   �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C=     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CT   !   �   �      �  �   �  �  	   �  �  \   �  B  C  �     !         �t�bhhK ��h��R�(KK��h�C<   �  �   -   �  s   \   �  �  .  N     C         �t�bhhK ��h��R�(KK��h�C�  �   �      �         �t�bhhK ��h��R�(KK��h�C<   !      -   �  �  �     p   X      >   �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�CD  �     !         �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C    B  C  �     !         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK	��h�C$X      '     �      �        �t�bhhK ��h��R�(KK��h�ChX      '     [   �                   �     �     #     �   �      [   �         �t�bhhK ��h��R�(KK��h�CL?   �        O           �     x   /        �    R        �t�bhhK ��h��R�(KK��h�C<      -   �  J              D   @    	        �t�bhhK ��h��R�(KK
��h�C(   !   �   �     X      �        �t�bhhK ��h��R�(KK��h�C@      
   �           j   �   P     '     �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   �     
     �t�bhhK ��h��R�(KK��h�CD  �     !         �t�bhhK ��h��R�(KK��h�CH   !         �      �     n        )   	                  �t�bhhK ��h��R�(KK��h�C8s                            n        �t�bhhK ��h��R�(KK��h�C    !      -   '   
        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   E           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�   |     �        �t�bhhK ��h��R�(KK��h�Ch
      �   �    k     )              �     '   �   	         g         �   |        �t�bhhK ��h��R�(KK��h�C&      �     C         �t�bhhK ��h��R�(KK��h�C,   !   �   �     X      A  n        �t�bhhK ��h��R�(KK��h�C4      
   �           j   �     |        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�   E     �t�bhhK ��h��R�(KK��h�CV           L      �t�bhhK ��h��R�(KK��h�CL
         ?     I   �        @   f        M        q         �t�bhhK ��h��R�(KK��h�C<    x   /   
      4   "   '   �         �         �t�bhhK ��h��R�(KK��h�CD      -   �   
   W   �  	         F   �      Q  �         �t�bhhK ��h��R�(KK��h�C        �t�bhhK ��h��R�(KK��h�C V           *           �t�bhhK ��h��R�(KK��h�C  o     �t�bhhK ��h��R�(KK��h�Cx
         ?     I   �  	   �     !      4   "   '   �         �   	         @   f           o        �t�bhhK ��h��R�(KK	��h�C$�      �      }      �        �t�bhhK ��h��R�(KK��h�CD�   b        �   o          F  y                   �t�bhhK ��h��R�(KK��h�C       7         =        �t�bhhK ��h��R�(KK��h�Co     �t�bhhK ��h��R�(KK��h�CG    	   �     �t�bhhK ��h��R�(KK��h�C(        �t�bhhK ��h��R�(KK��h�C      V      *           �t�bhhK ��h��R�(KK��h�Cz     �t�bhhK ��h��R�(KK��h�C8   !      <  }          	         !        �t�bhhK ��h��R�(KK	��h�C$:   T   X   �   Z   >   "        �t�bhhK ��h��R�(KK��h�C8      
   #     
   `   7         $  2         �t�bhhK ��h��R�(KK��h�C\D   9   %  �   t     �  &     "   !     !      v   V  s      '     (        �t�bhhK ��h��R�(KK��h�C         z        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C)     �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C*        �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C,+     �   �     �                 �t�bhhK ��h��R�(KK��h�C  �     �t�bhhK ��h��R�(KK��h�C`   !   )     �   m           �      F   k   	   t          �      r  �         �t�bhhK ��h��R�(KK��h�C0p     �     :   �   �  ,     �        �t�bhhK ��h��R�(KK��h�C H  �   -   �      C         �t�bhhK ��h��R�(KK
��h�C(      7         !   Q   2         �t�bhhK ��h��R�(KK��h�C         W   �        �t�bhhK ��h��R�(KK��h�C%   )        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C%   )        �t�bhhK ��h��R�(KK	��h�C$�      )         �      �      �t�bhhK ��h��R�(KK��h�C-        �t�bhhK ��h��R�(KK��h�C.     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CV           L      �t�bhhK ��h��R�(KK��h�Cz     �t�bhhK ��h��R�(KK��h�C  �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK
��h�C(   !      �  �     �   �         �t�bhhK ��h��R�(KK��h�C ]  6  D   &   �   &        �t�bhhK ��h��R�(KK��h�C8   !   V  �      )   	      	   E               �t�bhhK ��h��R�(KK��h�C0�   &  V  -   s      )      W   k         �t�bhhK ��h��R�(KK
��h�C(�   �   D   �   �        �        �t�bhhK ��h��R�(KK��h�CLB   6   i   
   �     v  $   w  �   n    z   6   f     &        �t�bhhK ��h��R�(KK��h�CD      i   
         &   �  &  M   �           7        �t�bhhK ��h��R�(KK��h�C8      '  `   5      �   �        '  [        �t�bhhK ��h��R�(KK��h�C,�     �     F      ^     U        �t�bhhK ��h��R�(KK��h�C �   �  �  .     T        �t�bhhK ��h��R�(KK��h�C\�   :  �      `   
   �        &     �          �  �     �     �        �t�bhhK ��h��R�(KK��h�C,�  �   B   
   �     &   �   ]        �t�bhhK ��h��R�(KK��h�CL
   K  �  �  �     9      *   	         D   g   �     �        �t�bhhK ��h��R�(KK��h�C4   6   c  �   �   J   `      &   �   ]        �t�bhhK ��h��R�(KK	��h�C$      7      M   q   �        �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�   �                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�   �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C `   
   d                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK	��h�C$'  x     �                 �t�bhhK ��h��R�(KK	��h�C$   
   &  )                  �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CL�      �     �      �  �     �   �   \      �     �  �        �t�bhhK ��h��R�(KK��h�C8   !      B   @   �      )   	                  �t�bhhK ��h��R�(KK	��h�C$   �   i   
                 �t�bhhK ��h��R�(KK��h�C4`      �  m  M   H   2            7        �t�bhhK ��h��R�(KK��h�Chf          	   5  `      -   �  �     \  	   
   K     F        !   '  ?   �        �t�bhhK ��h��R�(KK��h�CP�   s   8     �     4   "     k     )          D  a              �t�bhhK ��h��R�(KK��h�C8&   �        �     �     H  $      �        �t�bhhK ��h��R�(KK��h�C&   �      �  �        �t�bhhK ��h��R�(KK��h�C<T  8  z      &   �             �             �t�bhhK ��h��R�(KK��h�Cl   7         
     	   �          
   s      �     �      !   Q      �   9     2         �t�bhhK ��h��R�(KK��h�C,      -   �   
            U        �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C `                       �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
   &   �   �           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK	��h�C$'  x     g                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�      p              �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK��h�C0   !      �     �  �     �           �t�bhhK ��h��R�(KK��h�CD   !      -      �    	   v   B      �   �              �t�bhhK ��h��R�(KK��h�CH      
   �     !   7         !   Q      �   9     2         �t�bhhK ��h��R�(KK	��h�C$�     �  6   �     %        �t�bhhK ��h��R�(KK��h�C�     �             �t�bhhK ��h��R�(KK��h�C<   H   2   7      P     �           
   �        �t�bhhK ��h��R�(KK��h�C         [   X      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�  �      �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�   X   �  h     �t�bhhK ��h��R�(KK��h�Ct
   �   k     .   )   �   4      �  �     R     &   �  �  	      z   @   �   X      �  �           �t�bhhK ��h��R�(KK��h�C8   &   �      �  k  .   )   �      l  �        �t�bhhK ��h��R�(KK��h�C   s  �     '   I         �t�bhhK ��h��R�(KK��h�Cx
      "   �     1         �  }   `     "   $   ?   �   6      w   �      :     r   ;     <           �t�bhhK ��h��R�(KK��h�CD:  �  
   �    �      x   /      �      �  �   �        �t�bhhK ��h��R�(KK��h�C   
   &   �   �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C=     �t�bhhK ��h��R�(KK��h�C[   X      L   C      �t�bhhK ��h��R�(KK��h�CL   !   )     �   m        _     �     H  �  �   l  >        �t�bhhK ��h��R�(KK��h�CX
   B   "   �     �  	      B   �   l  �  D      �  
     �  �           �t�bhhK ��h��R�(KK��h�C[   X      �      �t�bhhK ��h��R�(KK��h�C�  
        �t�bhhK ��h��R�(KK��h�C�     ?     �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK*��h�C�      i      &   [   �  �  	   .   �   �        �  �     �     	   
      �  l  >    I      �    	   5  4   "   �     �      W   �        �t�bhhK ��h��R�(KK��h�CP   �  �        @    �  U   �        O      �     �  R        �t�bhhK ��h��R�(KK��h�CX�     !         �     �  !      �  !        �  �      A  n           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�CC      [   X      �t�bhhK ��h��R�(KK��h�C0   �     !   V  �     ^   >   k         �t�bhhK ��h��R�(KK+��h�C�   �  V  -   X      )      �     �  �  �             "   '   e   f  B  )   	         �  	      �  k     .   )   �   4         *     �        �t�bhhK ��h��R�(KK��h�CXN      �  /      @  	         �  �   /      �     s      J   �   �         �t�bhhK ��h��R�(KK��h�C\      -   �   /        2              �  	         O   U   J   �           �t�bhhK ��h��R�(KK
��h�C(&   �  �  �     &   �   @        �t�bhhK ��h��R�(KK��h�C@s      &   �   �     �   
   �  �     w             �t�bhhK ��h��R�(KK��h�C`      
   �     
   s        �   �   7         H   2      d   �     <           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�Cs      &   �   �     �t�bhhK ��h��R�(KK	��h�C$)      W   k      &   [   �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C=     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CT   !   �   �      �  �   �  �  	   �  �  \   �  B  C  �     !         �t�bhhK ��h��R�(KK��h�C<   �  �   -   �  s   \   �  �  .  N     C         �t�bhhK ��h��R�(KK��h�C�  �   �      �         �t�bhhK ��h��R�(KK��h�C<   !      -   �  �  �     p   X      >   �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�CD  �     !         �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C    B  C  �     !         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK	��h�C$X      '     �      �        �t�bhhK ��h��R�(KK��h�ChX      '     [   �                   �     �     #     �   �      [   �         �t�bhhK ��h��R�(KK��h�CL?   �        O           �     x   /        �    R        �t�bhhK ��h��R�(KK��h�C<      -   �  J              D   @    	        �t�bhhK ��h��R�(KK
��h�C(   !   �   �     X      �        �t�bhhK ��h��R�(KK��h�C@      
   �           j   �   P     '     �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   �     
     �t�bhhK ��h��R�(KK��h�CD  �     !         �t�bhhK ��h��R�(KK��h�CH   !         �      �     n        )   	                  �t�bhhK ��h��R�(KK��h�C8s                            n        �t�bhhK ��h��R�(KK��h�C    !      -   '   
        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   E           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�   |     �        �t�bhhK ��h��R�(KK��h�Ch
      �   �    k     )              �     '   �   	         g         �   |        �t�bhhK ��h��R�(KK��h�C&      �     C         �t�bhhK ��h��R�(KK��h�C,   !   �   �     X      A  n        �t�bhhK ��h��R�(KK��h�C4      
   �           j   �     |        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�   E     �t�bhhK ��h��R�(KK��h�CV           L      �t�bhhK ��h��R�(KK��h�CL
         ?     I   �        @   f        M        q         �t�bhhK ��h��R�(KK��h�C<    x   /   
      4   "   '   �         �         �t�bhhK ��h��R�(KK��h�CD      -   �   
   W   �  	         F   �      Q  �         �t�bhhK ��h��R�(KK��h�C        �t�bhhK ��h��R�(KK��h�C V           *           �t�bhhK ��h��R�(KK��h�C  o     �t�bhhK ��h��R�(KK��h�Cx
         ?     I   �  	   �     !      4   "   '   �         �   	         @   f           o        �t�bhhK ��h��R�(KK	��h�C$�      �      }      �        �t�bhhK ��h��R�(KK��h�CD�   b        �   o          F  y                   �t�bhhK ��h��R�(KK��h�C       7         =        �t�bhhK ��h��R�(KK��h�Co     �t�bhhK ��h��R�(KK��h�CG    	   �     �t�bhhK ��h��R�(KK��h�C(        �t�bhhK ��h��R�(KK��h�C      V      *           �t�bhhK ��h��R�(KK��h�Cz     �t�bhhK ��h��R�(KK��h�C8   !      <  }          	         !        �t�bhhK ��h��R�(KK	��h�C$:   T   X   �   Z   >   "        �t�bhhK ��h��R�(KK��h�C8      
   #     
   `   7         $  2         �t�bhhK ��h��R�(KK��h�C\D   9   %  �   t     �  &     "   !     !      v   V  s      '     (        �t�bhhK ��h��R�(KK��h�C         z        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C)     �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C*        �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C,+     �   �     �                 �t�bhhK ��h��R�(KK��h�C  �     �t�bhhK ��h��R�(KK��h�C`   !   )     �   m           �      F   k   	   t          �      r  �         �t�bhhK ��h��R�(KK��h�C0p     �     :   �   �  ,     �        �t�bhhK ��h��R�(KK��h�C H  �   -   �      C         �t�bhhK ��h��R�(KK
��h�C(      7         !   Q   2         �t�bhhK ��h��R�(KK��h�C         W   �        �t�bhhK ��h��R�(KK��h�C%   )        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C%   )        �t�bhhK ��h��R�(KK	��h�C$�      )         �      �      �t�bhhK ��h��R�(KK��h�C-        �t�bhhK ��h��R�(KK��h�C.     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CV           L      �t�bhhK ��h��R�(KK��h�Cz     �t�bhhK ��h��R�(KK��h�C  �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK
��h�C(   !      �  �     �   �         �t�bhhK ��h��R�(KK��h�C ]  6  D   &   �   &        �t�bhhK ��h��R�(KK��h�C8   !   V  �      )   	      	   E               �t�bhhK ��h��R�(KK��h�C0�   &  V  -   s      )      W   k         �t�bhhK ��h��R�(KK
��h�C(�   �   D   �   �        �        �t�bhhK ��h��R�(KK��h�CLB   6   i   
   �     v  $   w  �   n    z   6   f     &        �t�bhhK ��h��R�(KK��h�CD      i   
         &   �  &  M   �           7        �t�bhhK ��h��R�(KK��h�C8      '  `   5      �   �        '  [        �t�bhhK ��h��R�(KK��h�C,�     �     F      ^     U        �t�bhhK ��h��R�(KK��h�C �   �  �  .     T        �t�bhhK ��h��R�(KK��h�C\�   :  �      `   
   �        &     �          �  �     �     �        �t�bhhK ��h��R�(KK��h�C,�  �   B   
   �     &   �   ]        �t�bhhK ��h��R�(KK��h�CL
   K  �  �  �     9      *   	         D   g   �     �        �t�bhhK ��h��R�(KK��h�C4   6   c  �   �   J   `      &   �   ]        �t�bhhK ��h��R�(KK	��h�C$      7      M   q   �        �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�   �                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�   �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C `   
   d                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK	��h�C$'  x     �                 �t�bhhK ��h��R�(KK	��h�C$   
   &  )                  �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CL�      �     �      �  �     �   �   \      �     �  �        �t�bhhK ��h��R�(KK��h�C8   !      B   @   �      )   	                  �t�bhhK ��h��R�(KK	��h�C$   �   i   
                 �t�bhhK ��h��R�(KK��h�C4`      �  m  M   H   2            7        �t�bhhK ��h��R�(KK��h�Chf          	   5  `      -   �  �     \  	   
   K     F        !   '  ?   �        �t�bhhK ��h��R�(KK��h�CP�   s   8     �     4   "     k     )          D  a              �t�bhhK ��h��R�(KK��h�C8&   �        �     �     H  $      �        �t�bhhK ��h��R�(KK��h�C&   �      �  �        �t�bhhK ��h��R�(KK��h�C<T  8  z      &   �             �             �t�bhhK ��h��R�(KK��h�Cl   7         
     	   �          
   s      �     �      !   Q      �   9     2         �t�bhhK ��h��R�(KK��h�C,      -   �   
            U        �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C `                       �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C    
   &   �   �           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK	��h�C$'  x     g                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�      p              �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK��h�C0   !      �     �  �     �           �t�bhhK ��h��R�(KK��h�CD   !      -      �    	   v   B      �   �              �t�bhhK ��h��R�(KK��h�CH      
   �     !   7         !   Q      �   9     2         �t�bhhK ��h��R�(KK	��h�C$�     �  6   �     %        �t�bhhK ��h��R�(KK��h�C�     �             �t�bhhK ��h��R�(KK��h�C<   H   2   7      P     �           
   �        �t�bhhK ��h��R�(KK��h�C         [   X      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�  �      �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�   X   �  h     �t�bhhK ��h��R�(KK��h�Ct
   �   k     .   )   �   4      �  �     R     &   �  �  	      z   @   �   X      �  �           �t�bhhK ��h��R�(KK��h�C8   &   �      �  k  .   )   �      l  �        �t�bhhK ��h��R�(KK��h�C   s  �     '   I         �t�bhhK ��h��R�(KK��h�Cx
      "   �     1         �  }   `     "   $   ?   �   6      w   �      :     r   ;     <           �t�bhhK ��h��R�(KK��h�CD:  �  
   �    �      x   /      �      �  �   �        �t�bhhK ��h��R�(KK��h�C   
   &   �   �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C=     �t�bhhK ��h��R�(KK��h�C[   X      L   C      �t�bhhK ��h��R�(KK��h�CL   !   )     �   m        _     �     H  �  �   l  >        �t�bhhK ��h��R�(KK��h�CX
   B   "   �     �  	      B   �   l  �  D      �  
     �  �           �t�bhhK ��h��R�(KK��h�C[   X      �      �t�bhhK ��h��R�(KK��h�C�  
        �t�bhhK ��h��R�(KK��h�C�     ?     �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK*��h�C�      i      &   [   �  �  	   .   �   �        �  �     �     	   
      �  l  >    I      �    	   5  4   "   �     �      W   �        �t�bhhK ��h��R�(KK��h�CP   �  �        @    �  U   �        O      �     �  R        �t�bhhK ��h��R�(KK��h�CX�     !         �     �  !      �  !        �  �      A  n           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�CC      [   X      �t�bhhK ��h��R�(KK��h�C0   �     !   V  �     ^   >   k         �t�bhhK ��h��R�(KK+��h�C�   �  V  -   X      )      �     �  �  �             "   '   e   f  B  )   	         �  	      �  k     .   )   �   4         *     �        �t�bhhK ��h��R�(KK��h�CXN      �  /      @  	         �  �   /      �     s      J   �   �         �t�bhhK ��h��R�(KK��h�C\      -   �   /        2              �  	         O   U   J   �           �t�bhhK ��h��R�(KK
��h�C(&   �  �  �     &   �   @        �t�bhhK ��h��R�(KK��h�C@s      &   �   �     �   
   �  �     w             �t�bhhK ��h��R�(KK��h�C`      
   �     
   s        �   �   7         H   2      d   �     <           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�Cs      &   �   �     �t�bhhK ��h��R�(KK	��h�C$)      W   k      &   [   �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C=     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CT   !   �   �      �  �   �  �  	   �  �  \   �  B  C  �     !         �t�bhhK ��h��R�(KK��h�C<   �  �   -   �  s   \   �  �  .  N     C         �t�bhhK ��h��R�(KK��h�C�  �   �      �         �t�bhhK ��h��R�(KK��h�C<   !      -   �  �  �     p   X      >   �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�CD  �     !         �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C    B  C  �     !         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK	��h�C$X      '     �      �        �t�bhhK ��h��R�(KK��h�ChX      '     [   �                   �     �     #     �   �      [   �         �t�bhhK ��h��R�(KK��h�CL?   �        O           �     x   /        �    R        �t�bhhK ��h��R�(KK��h�C<      -   �  J              D   @    	        �t�bhhK ��h��R�(KK
��h�C(   !   �   �     X      �        �t�bhhK ��h��R�(KK��h�C@      
   �           j   �   P     '     �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   �     
     �t�bhhK ��h��R�(KK��h�CD  �     !         �t�bhhK ��h��R�(KK��h�CH   !         �      �     n        )   	                  �t�bhhK ��h��R�(KK��h�C8s                            n        �t�bhhK ��h��R�(KK��h�C    !      -   '   
        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   E           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�   |     �        �t�bhhK ��h��R�(KK��h�Ch
      �   �    k     )              �     '   �   	         g         �   |        �t�bhhK ��h��R�(KK��h�C&      �     C         �t�bhhK ��h��R�(KK��h�C,   !   �   �     X      A  n        �t�bhhK ��h��R�(KK��h�C4      
   �           j   �     |        �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�   E     �t�bhhK ��h��R�(KK��h�CV           L      �t�bhhK ��h��R�(KK��h�CL
         ?     I   �        @   f        M        q         �t�bhhK ��h��R�(KK��h�C<    x   /   
      4   "   '   �         �         �t�bhhK ��h��R�(KK��h�CD      -   �   
   W   �  	         F   �      Q  �         �t�bhhK ��h��R�(KK��h�C        �t�bhhK ��h��R�(KK��h�C V           *           �t�bhhK ��h��R�(KK��h�C  o     �t�bhhK ��h��R�(KK��h�Cx
         ?     I   �  	   �     !      4   "   '   �         �   	         @   f           o        �t�bhhK ��h��R�(KK	��h�C$�      �      }      �        �t�bhhK ��h��R�(KK��h�CD�   b        �   o          F  y                   �t�bhhK ��h��R�(KK��h�C       7         =        �t�bhhK ��h��R�(KK��h�Co     �t�bhhK ��h��R�(KK��h�CG    	   �     �t�bhhK ��h��R�(KK��h�C(        �t�bhhK ��h��R�(KK��h�C      V      *           �t�bhhK ��h��R�(KK��h�Cz     �t�bhhK ��h��R�(KK��h�C8   !      <  }          	         !        �t�bhhK ��h��R�(KK	��h�C$:   T   X   �   Z   >   "        �t�bhhK ��h��R�(KK��h�C8      
   #     
   `   7         $  2         �t�bhhK ��h��R�(KK��h�C\D   9   %  �   t     �  &     "   !     !      v   V  s      '     (        �t�bhhK ��h��R�(KK��h�C          }  	            �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C)     �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C*        �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C,+     �   �     �                 �t�bhhK ��h��R�(KK��h�C  �     �t�bhhK ��h��R�(KK��h�C`   !   )     �   m           �      F   k   	   t          �      r  �         �t�bhhK ��h��R�(KK��h�C0p     �     :   �   �  ,     �        �t�bhhK ��h��R�(KK��h�C H  �   -   �      C         �t�bhhK ��h��R�(KK
��h�C(      7         !   Q   2         �t�bhhK ��h��R�(KK��h�C          R     �        �t�bhhK ��h��R�(KK��h�C%   )        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C%   )        �t�bhhK ��h��R�(KK	��h�C$�      )         �      �      �t�bhhK ��h��R�(KK��h�C-        �t�bhhK ��h��R�(KK��h�C.     �t�bhhK ��h��R�(KK��h�C4�  �     4      .   k         "           �t�bhhK ��h��R�(KK��h�C  �   e   k         �t�bhhK ��h��R�(KK��h�C)      �t�bhhK ��h��R�(KK��h�C4�  �     4      .   k         "           �t�bhhK ��h��R�(KK��h�C  �   e   k         �t�bhhK ��h��R�(KK��h�C)      �t�bhhK ��h��R�(KK��h�C4�  �     4      .   k         "           �t�bhhK ��h��R�(KK��h�C  �   e   k         �t�bhhK ��h��R�(KK��h�C)      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�         �     �t�bhhK ��h��R�(KK��h�C7     �t�bhhK ��h��R�(KK��h�Cj          �t�bhhK ��h��R�(KK��h�CI  k     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C u     O  v     �         �t�bhhK ��h��R�(KK��h�C4      %  /         0  �   1  /   %        �t�bhhK ��h��R�(KK��h�C42  �      W   J  "   3      �  /   �         �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�CL   !      D   Z   W   J  	   @  :   P     4  	   5     6        �t�bhhK ��h��R�(KK��h�CD_    �      !      Z     	   7  8     9     :        �t�bhhK ��h��R�(KK��h�C4.        s      @   �   M      �   ;        �t�bhhK ��h��R�(KK��h�C`
                 i   
      �   M   X  x  y     �  �  <     =  y           �t�bhhK ��h��R�(KK��h�Cl
         ~  B    I   	         g   �   d   >     K     ?        @  L     L           �t�bhhK ��h��R�(KK��h�CA        �t�bhhK ��h��R�(KK��h�C!           �t�bhhK ��h��R�(KK��h�CB        �t�bhhK ��h��R�(KK��h�C!     �t�bhhK ��h��R�(KK��h�CC        �t�bhhK ��h��R�(KK��h�C!                 �t�bhhK ��h��R�(KK��h�C|     K        �t�bhhK ��h��R�(KK	��h�C$�      Y   ?     D           �t�bhhK ��h��R�(KK��h�C�      *           �t�bhhK ��h��R�(KK��h�Cy        �t�bhhK ��h��R�(KK��h�C �      z                 �t�bhhK ��h��R�(KK��h�CH   �      �t�bhhK ��h��R�(KK��h�CDH   �      �  "  B  :   �       �      �      w        �t�bhhK ��h��R�(KK��h�CTE     �  �     �  �  �     x     �       :   M  O      �         �t�bhhK ��h��R�(KK��h�C4!   Q   �          �      N    �        �t�bhhK ��h��R�(KK��h�CF  �     �t�bhhK ��h��R�(KK��h�C(   G     H        �t�bhhK ��h��R�(KK��h�C0      �      �     N      2         �t�bhhK ��h��R�(KK��h�C0`      I     �   n     �   `  J        �t�bhhK ��h��R�(KK��h�CD   K     |      H   �   L  :   M     "   '     M        �t�bhhK ��h��R�(KK��h�CDD   N  �  O  	     {  �     N     Y      �  �        �t�bhhK ��h��R�(KK��h�C   
   H   !           �t�bhhK ��h��R�(KK��h�C `   
   �      +           �t�bhhK ��h��R�(KK��h�C�         �     �t�bhhK ��h��R�(KK��h�C`
   J   �   "   �     F      �     �     �     �     �  �  �  :   �  �        �t�bhhK ��h��R�(KK
��h�C(=   r     .  N   �  "   �        �t�bhhK ��h��R�(KK��h�Cd   o  O   B   -   +      !   Q   0           )  }  *     	      "   �   �   �         �t�bhhK ��h��R�(KK��h�C,l     0      �         <      +     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C 0                       �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cd
        J   �  G  l   p  /      �  /      l   	         =   '   �      �           �t�bhhK ��h��R�(KK��h�C�  "   �  �   �         �t�bhhK ��h��R�(KK��h�C4#  �     '   �   �     �     �  $         �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�C0      -        !   �      �  �         �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�Cz  O     �t�bhhK ��h��R�(KK��h�C(      <      ]     �t�bhhK ��h��R�(KK��h�C�  �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C+      �     �     �t�bhhK ��h��R�(KK��h�CP+      V      I           E      �      �      �      �     �     �t�bhhK ��h��R�(KK��h�C:   _   (     �t�bhhK ��h��R�(KK��h�Cp�   	  
  !  _   (     �  �  �  �  �     p   V      +      o     J     %     H  �         �t�bhhK ��h��R�(KK��h�C<"  "   �   y      _     =  	   �  �   �   �         �t�bhhK ��h��R�(KK��h�C�  :     �  �        �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C�   	  
        �t�bhhK ��h��R�(KK��h�C :   _   #                 �t�bhhK ��h��R�(KK��h�C7     �t�bhhK ��h��R�(KK��h�CD
          6      =   P     Q        r   �   �        �t�bhhK ��h��R�(KK	��h�C$P  7         !   Q   2         �t�bhhK ��h��R�(KK��h�CH
   J   S     !   	         @      �   M   R  �     S        �t�bhhK ��h��R�(KK��h�C         7     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�CO                 �t�bhhK ��h��R�(KK��h�C�     T     �t�bhhK ��h��R�(KK	��h�C$U     Y      q  V          �t�bhhK ��h��R�(KK��h�Cj          �t�bhhK ��h��R�(KK��h�C\�   �   �     F      q     �   	      "   {      D     :   |  }  �   +         �t�bhhK ��h��R�(KK��h�Clq     �      4   �         �  W  	      �          X              Y     Z           �t�bhhK ��h��R�(KK��h�CT      
   �  ;   O      U   2     [  �      \  ]        r   ;        �t�bhhK ��h��R�(KK��h�C          j             �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
     �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   H   ^     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�   _     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�CO                 �t�bhhK ��h��R�(KK��h�CI  k     �t�bhhK ��h��R�(KK��h�CD   
   u   J   |  `     a     �   7         =  b        �t�bhhK ��h��R�(KK��h�C          k     &        �t�bhhK ��h��R�(KK��h�Cc        �t�bhhK ��h��R�(KK��h�CP     �t�bhhK ��h��R�(KK��h�Cd        �t�bhhK ��h��R�(KK��h�CP                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�         �     �t�bhhK ��h��R�(KK��h�C7     �t�bhhK ��h��R�(KK��h�Cj          �t�bhhK ��h��R�(KK��h�CI  k     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C u     O  v     �         �t�bhhK ��h��R�(KK��h�C4      %  /         0  �   1  /   %        �t�bhhK ��h��R�(KK��h�C42  �      W   J  "   3      �  /   �         �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�CL   !      D   Z   W   J  	   @  :   P     4  	   5     6        �t�bhhK ��h��R�(KK��h�CD_    �      !      Z     	   7  8     9     :        �t�bhhK ��h��R�(KK��h�C4.        s      @   �   M      �   ;        �t�bhhK ��h��R�(KK��h�C`
                 i   
      �   M   X  x  y     �  �  <     =  y           �t�bhhK ��h��R�(KK��h�Cl
         ~  B    I   	         g   �   d   >     K     ?        @  L     L           �t�bhhK ��h��R�(KK��h�CA        �t�bhhK ��h��R�(KK��h�C!           �t�bhhK ��h��R�(KK��h�CB        �t�bhhK ��h��R�(KK��h�C!     �t�bhhK ��h��R�(KK��h�CC        �t�bhhK ��h��R�(KK��h�C!                 �t�bhhK ��h��R�(KK��h�C|     K        �t�bhhK ��h��R�(KK	��h�C$�      Y   ?     D           �t�bhhK ��h��R�(KK��h�C�      *           �t�bhhK ��h��R�(KK��h�Cy        �t�bhhK ��h��R�(KK��h�C �      z                 �t�bhhK ��h��R�(KK��h�CH   �      �t�bhhK ��h��R�(KK��h�CDH   �      �  "  B  :   �       �      �      w        �t�bhhK ��h��R�(KK��h�CTE     �  �     �  �  �     x     �       :   M  O      �         �t�bhhK ��h��R�(KK��h�C4!   Q   �          �      N    �        �t�bhhK ��h��R�(KK��h�CF  �     �t�bhhK ��h��R�(KK��h�C(   G     H        �t�bhhK ��h��R�(KK��h�C0      �      �     N      2         �t�bhhK ��h��R�(KK��h�C0`      I     �   n     �   `  J        �t�bhhK ��h��R�(KK��h�CD   K     |      H   �   L  :   M     "   '     M        �t�bhhK ��h��R�(KK��h�CDD   N  �  O  	     {  �     N     Y      �  �        �t�bhhK ��h��R�(KK��h�C   
   H   !           �t�bhhK ��h��R�(KK��h�C `   
   �      +           �t�bhhK ��h��R�(KK��h�C�         �     �t�bhhK ��h��R�(KK��h�C`
   J   �   "   �     F      �     �     �     �     �  �  �  :   �  �        �t�bhhK ��h��R�(KK
��h�C(=   r     .  N   �  "   �        �t�bhhK ��h��R�(KK��h�Cd   o  O   B   -   +      !   Q   0           )  }  *     	      "   �   �   �         �t�bhhK ��h��R�(KK��h�C,l     0      �         <      +     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C 0                       �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cd
        J   �  G  l   p  /      �  /      l   	         =   '   �      �           �t�bhhK ��h��R�(KK��h�C�  "   �  �   �         �t�bhhK ��h��R�(KK��h�C4#  �     '   �   �     �     �  $         �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�C0      -        !   �      �  �         �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�Cz  O     �t�bhhK ��h��R�(KK��h�C(      <      ]     �t�bhhK ��h��R�(KK��h�C�  �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C+      �     �     �t�bhhK ��h��R�(KK��h�CP+      V      I           E      �      �      �      �     �     �t�bhhK ��h��R�(KK��h�C:   _   (     �t�bhhK ��h��R�(KK��h�Cp�   	  
  !  _   (     �  �  �  �  �     p   V      +      o     J     %     H  �         �t�bhhK ��h��R�(KK��h�C<"  "   �   y      _     =  	   �  �   �   �         �t�bhhK ��h��R�(KK��h�C�  :     �  �        �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C�   	  
        �t�bhhK ��h��R�(KK��h�C :   _   #                 �t�bhhK ��h��R�(KK��h�C7     �t�bhhK ��h��R�(KK��h�CD
          6      =   P     Q        r   �   �        �t�bhhK ��h��R�(KK	��h�C$P  7         !   Q   2         �t�bhhK ��h��R�(KK��h�CH
   J   S     !   	         @      �   M   R  �     S        �t�bhhK ��h��R�(KK��h�C         7     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�CO                 �t�bhhK ��h��R�(KK��h�C�     T     �t�bhhK ��h��R�(KK	��h�C$U     Y      q  V          �t�bhhK ��h��R�(KK��h�Cj          �t�bhhK ��h��R�(KK��h�C\�   �   �     F      q     �   	      "   {      D     :   |  }  �   +         �t�bhhK ��h��R�(KK��h�Clq     �      4   �         �  W  	      �          X              Y     Z           �t�bhhK ��h��R�(KK��h�CT      
   �  ;   O      U   2     [  �      \  ]        r   ;        �t�bhhK ��h��R�(KK��h�C          j             �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
     �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   H   ^     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�   _     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�CO                 �t�bhhK ��h��R�(KK��h�CI  k     �t�bhhK ��h��R�(KK��h�CD   
   u   J   |  `     a     �   7         =  b        �t�bhhK ��h��R�(KK��h�C          k     &        �t�bhhK ��h��R�(KK��h�Cc        �t�bhhK ��h��R�(KK��h�CP     �t�bhhK ��h��R�(KK��h�Cd        �t�bhhK ��h��R�(KK��h�CP                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�         �     �t�bhhK ��h��R�(KK��h�C7     �t�bhhK ��h��R�(KK��h�Cj          �t�bhhK ��h��R�(KK��h�CI  k     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C u     O  v     �         �t�bhhK ��h��R�(KK��h�C4      %  /         0  �   1  /   %        �t�bhhK ��h��R�(KK��h�C42  �      W   J  "   3      �  /   �         �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�CL   !      D   Z   W   J  	   @  :   P     4  	   5     6        �t�bhhK ��h��R�(KK��h�CD_    �      !      Z     	   7  8     9     :        �t�bhhK ��h��R�(KK��h�C4.        s      @   �   M      �   ;        �t�bhhK ��h��R�(KK��h�C`
                 i   
      �   M   X  x  y     �  �  <     =  y           �t�bhhK ��h��R�(KK��h�Cl
         ~  B    I   	         g   �   d   >     K     ?        @  L     L           �t�bhhK ��h��R�(KK��h�CA        �t�bhhK ��h��R�(KK��h�C!           �t�bhhK ��h��R�(KK��h�CB        �t�bhhK ��h��R�(KK��h�C!     �t�bhhK ��h��R�(KK��h�CC        �t�bhhK ��h��R�(KK��h�C!                 �t�bhhK ��h��R�(KK��h�C|     K        �t�bhhK ��h��R�(KK	��h�C$�      Y   ?     D           �t�bhhK ��h��R�(KK��h�C�      *           �t�bhhK ��h��R�(KK��h�Cy        �t�bhhK ��h��R�(KK��h�C �      z                 �t�bhhK ��h��R�(KK��h�CH   �      �t�bhhK ��h��R�(KK��h�CDH   �      �  "  B  :   �       �      �      w        �t�bhhK ��h��R�(KK��h�CTE     �  �     �  �  �     x     �       :   M  O      �         �t�bhhK ��h��R�(KK��h�C4!   Q   �          �      N    �        �t�bhhK ��h��R�(KK��h�CF  �     �t�bhhK ��h��R�(KK��h�C(   G     H        �t�bhhK ��h��R�(KK��h�C0      �      �     N      2         �t�bhhK ��h��R�(KK��h�C0`      I     �   n     �   `  J        �t�bhhK ��h��R�(KK��h�CD   K     |      H   �   L  :   M     "   '     M        �t�bhhK ��h��R�(KK��h�CDD   N  �  O  	     {  �     N     Y      �  �        �t�bhhK ���&      h��R�(KK��h�C   
   H   !           �t�bhhK ��h��R�(KK��h�C `   
   �      +           �t�bhhK ��h��R�(KK��h�C�         �     �t�bhhK ��h��R�(KK��h�C`
   J   �   "   �     F      �     �     �     �     �  �  �  :   �  �        �t�bhhK ��h��R�(KK
��h�C(=   r     .  N   �  "   �        �t�bhhK ��h��R�(KK��h�Cd   o  O   B   -   +      !   Q   0           )  }  *     	      "   �   �   �         �t�bhhK ��h��R�(KK��h�C,l     0      �         <      +     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C 0                       �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cd
        J   �  G  l   p  /      �  /      l   	         =   '   �      �           �t�bhhK ��h��R�(KK��h�C�  "   �  �   �         �t�bhhK ��h��R�(KK��h�C4#  �     '   �   �     �     �  $         �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�C0      -        !   �      �  �         �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�Cz  O     �t�bhhK ��h��R�(KK��h�C(      <      ]     �t�bhhK ��h��R�(KK��h�C�  �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C+      �     �     �t�bhhK ��h��R�(KK��h�CP+      V      I           E      �      �      �      �     �     �t�bhhK ��h��R�(KK��h�C:   _   (     �t�bhhK ��h��R�(KK��h�Cp�   	  
  !  _   (     �  �  �  �  �     p   V      +      o     J     %     H  �         �t�bhhK ��h��R�(KK��h�C<"  "   �   y      _     =  	   �  �   �   �         �t�bhhK ��h��R�(KK��h�C�  :     �  �        �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C�   	  
        �t�bhhK ��h��R�(KK��h�C :   _   #                 �t�bhhK ��h��R�(KK��h�C7     �t�bhhK ��h��R�(KK��h�CD
          6      =   P     Q        r   �   �        �t�bhhK ��h��R�(KK	��h�C$P  7         !   Q   2         �t�bhhK ��h��R�(KK��h�CH
   J   S     !   	         @      �   M   R  �     S        �t�bhhK ��h��R�(KK��h�C         7     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�CO                 �t�bhhK ��h��R�(KK��h�C�     T     �t�bhhK ��h��R�(KK	��h�C$U     Y      q  V          �t�bhhK ��h��R�(KK��h�Cj          �t�bhhK ��h��R�(KK��h�C\�   �   �     F      q     �   	      "   {      D     :   |  }  �   +         �t�bhhK ��h��R�(KK��h�Clq     �      4   �         �  W  	      �          X              Y     Z           �t�bhhK ��h��R�(KK��h�CT      
   �  ;   O      U   2     [  �      \  ]        r   ;        �t�bhhK ��h��R�(KK��h�C          j             �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
     �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   H   ^     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�   _     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�CO                 �t�bhhK ��h��R�(KK��h�CI  k     �t�bhhK ��h��R�(KK��h�CD   
   u   J   |  `     a     �   7         =  b        �t�bhhK ��h��R�(KK��h�C          k     &        �t�bhhK ��h��R�(KK��h�Cc        �t�bhhK ��h��R�(KK��h�CP     �t�bhhK ��h��R�(KK��h�Cd        �t�bhhK ��h��R�(KK��h�CP                 �t�bhhK ��h��R�(KK	��h�C$�      �   .   )         �      �t�bhhK ��h��R�(KK��h�C~     �t�bhhK ��h��R�(KK��h�C\   +      q           g      Y  �     )      9   	   !   	   *      8         �t�bhhK ��h��R�(KK��h�C<p        7      2      e     0     f  g        �t�bhhK ��h��R�(KK
��h�C(p     q        �               �t�bhhK ��h��R�(KK	��h�C$q   �  4   �        �         �t�bhhK ��h��R�(KK��h�Cl   !   �  �      )         �      C      !   )     �   m     h          �               �t�bhhK ��h��R�(KK��h�C4H  �      �  	   5  �   �   �     !         �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�Ci  �     �t�bhhK ��h��R�(KK��h�C(      <      j     �t�bhhK ��h��R�(KK��h�CD     
   �      �  7         !   k  2         Q        �t�bhhK ��h��R�(KK��h�CL   O   Q     F      �      ^  \      m  �     !   Q   2         �t�bhhK ��h��R�(KK��h�C@�        8  C      �      )   �      $     l        �t�bhhK ��h��R�(KK#��h�C�               m     n  o     /   	         D   @   D      �         p  q     D         r     s        �         �t�bhhK ��h��R�(KK
��h�C(      7         �              �t�bhhK ��h��R�(KK	��h�C$         R     )            �t�bhhK ��h��R�(KK��h�C,�      )         �           E      �t�bhhK ��h��R�(KK��h�C%   )        �t�bhhK ��h��R�(KK	��h�C$�      )         �      �      �t�bhhK ��h��R�(KK��h�C�      w        �t�bhhK ��h��R�(KK��h�C,X      )         �                 �t�bhhK ��h��R�(KK��h�C%   )        �t�bhhK ��h��R�(KK��h�C�     ?     �t�bhhK ��h��R�(KK��h�C�     )      �t�bhhK ��h��R�(KK��h�CL   !   �  �  �     t     	   v   B      u         L  )         �t�bhhK ��h��R�(KK��h�C4      �   R  a   �  )           v        �t�bhhK ��h��R�(KK��h�CH   �    w  )   	   i  .      �  
           x  )         �t�bhhK ��h��R�(KK��h�C�     v        �t�bhhK ��h��R�(KK
��h�C(      
   �  O      U   a        �t�bhhK ��h��R�(KK��h�Cl   !   �  y     )   D      z  �     �  �        {     |  }     ~  }    S           �t�bhhK ��h��R�(KK��h�Ch�  N     �     �  $      �   �     �     �           :   �   U     �             �t�bhhK ��h��R�(KK��h�C,         R  a   �  )      v        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CXT  7  �  ?     �  �     �     T   s      �     .   )   �      �        �t�bhhK ��h��R�(KK��h�C@^   >   7  �  ?     �     ?     >   �     !         �t�bhhK ��h��R�(KK	��h�C$.      �      �      �        �t�bhhK ��h��R�(KK��h�C�           E      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�CU           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�CU           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C,     |      �   r                 �t�bhhK ��h��R�(KK��h�C�  �  ?     T        �t�bhhK ��h��R�(KK
��h�C(7  �  ?     �                 �t�bhhK ��h��R�(KK��h�C'  �     �t�bhhK ��h��R�(KK��h�C0      �   '  �     )         �         �t�bhhK ��h��R�(KK��h�C\   �     �     2         �     ,        �  u      N         �   	        �t�bhhK ��h��R�(KK��h�C<   !   �   �     F      !   )     �   m           �t�bhhK ��h��R�(KK	��h�C$         �  �     �        �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C8    �   a         '  �     �                 �t�bhhK ��h��R�(KK��h�C%   )        �t�bhhK ��h��R�(KK��h�C'  �     �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK	��h�C$�      �   .   )         �      �t�bhhK ��h��R�(KK��h�C~     �t�bhhK ��h��R�(KK��h�C\   +      q           g      Y  �     )      9   	   !   	   *      8         �t�bhhK ��h��R�(KK��h�C<p        7      2      e     0     f  g        �t�bhhK ��h��R�(KK
��h�C(p     q        �               �t�bhhK ��h��R�(KK	��h�C$q   �  4   �        �         �t�bhhK ��h��R�(KK��h�Cl   !   �  �      )         �      C      !   )     �   m     h          �               �t�bhhK ��h��R�(KK��h�C4H  �      �  	   5  �   �   �     !         �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�Ci  �     �t�bhhK ��h��R�(KK��h�C(      <      j     �t�bhhK ��h��R�(KK��h�CD     
   �      �  7         !   k  2         Q        �t�bhhK ��h��R�(KK��h�CL   O   Q     F      �      ^  \      m  �     !   Q   2         �t�bhhK ��h��R�(KK��h�C@�        8  C      �      )   �      $     l        �t�bhhK ��h��R�(KK#��h�C�               m     n  o     /   	         D   @   D      �         p  q     D         r     s        �         �t�bhhK ��h��R�(KK
��h�C(      7         �              �t�bhhK ��h��R�(KK	��h�C$         R     )            �t�bhhK ��h��R�(KK��h�C,�      )         �           E      �t�bhhK ��h��R�(KK��h�C%   )        �t�bhhK ��h��R�(KK	��h�C$�      )         �      �      �t�bhhK ��h��R�(KK��h�C�      w        �t�bhhK ��h��R�(KK��h�C,X      )         �                 �t�bhhK ��h��R�(KK��h�C%   )        �t�bhhK ��h��R�(KK��h�C�     ?     �t�bhhK ��h��R�(KK��h�C�     )      �t�bhhK ��h��R�(KK��h�CL   !   �  �  �     t     	   v   B      u         L  )         �t�bhhK ��h��R�(KK��h�C4      �   R  a   �  )           v        �t�bhhK ��h��R�(KK��h�CH   �    w  )   	   i  .      �  
           x  )         �t�bhhK ��h��R�(KK��h�C�     v        �t�bhhK ��h��R�(KK
��h�C(      
   �  O      U   a        �t�bhhK ��h��R�(KK��h�Cl   !   �  y     )   D      z  �     �  �        {     |  }     ~  }    S           �t�bhhK ��h��R�(KK��h�Ch�  N     �     �  $      �   �     �     �           :   �   U     �             �t�bhhK ��h��R�(KK��h�C,         R  a   �  )      v        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CXT  7  �  ?     �  �     �     T   s      �     .   )   �      �        �t�bhhK ��h��R�(KK��h�C@^   >   7  �  ?     �     ?     >   �     !         �t�bhhK ��h��R�(KK	��h�C$.      �      �      �        �t�bhhK ��h��R�(KK��h�C�           E      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�CU           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�CU           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C,     |      �   r                 �t�bhhK ��h��R�(KK��h�C�  �  ?     T        �t�bhhK ��h��R�(KK
��h�C(7  �  ?     �                 �t�bhhK ��h��R�(KK��h�C'  �     �t�bhhK ��h��R�(KK��h�C0      �   '  �     )         �         �t�bhhK ��h��R�(KK��h�C\   �     �     2         �     ,        �  u      N         �   	        �t�bhhK ��h��R�(KK��h�C<   !   �   �     F      !   )     �   m           �t�bhhK ��h��R�(KK	��h�C$         �  �     �        �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C8    �   a         '  �     �                 �t�bhhK ��h��R�(KK��h�C%   )        �t�bhhK ��h��R�(KK��h�C'  �     �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK	��h�C$�      �   .   )         �      �t�bhhK ��h��R�(KK��h�C~     �t�bhhK ��h��R�(KK��h�C\   +      q           g      Y  �     )      9   	   !   	   *      8         �t�bhhK ��h��R�(KK��h�C<p        7      2      e     0     f  g        �t�bhhK ��h��R�(KK
��h�C(p     q        �               �t�bhhK ��h��R�(KK	��h�C$q   �  4   �        �         �t�bhhK ��h��R�(KK��h�Cl   !   �  �      )         �      C      !   )     �   m     h          �               �t�bhhK ��h��R�(KK��h�C4H  �      �  	   5  �   �   �     !         �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�Ci  �     �t�bhhK ��h��R�(KK��h�C(      <      j     �t�bhhK ��h��R�(KK��h�CD     
   �      �  7         !   k  2         Q        �t�bhhK ��h��R�(KK��h�CL   O   Q     F      �      ^  \      m  �     !   Q   2         �t�bhhK ��h��R�(KK��h�C@�        8  C      �      )   �      $     l        �t�bhhK ��h��R�(KK#��h�C�               m     n  o     /   	         D   @   D      �         p  q     D         r     s        �         �t�bhhK ��h��R�(KK
��h�C(      7         �              �t�bhhK ��h��R�(KK	��h�C$         R     )            �t�bhhK ��h��R�(KK��h�C,�      )         �           E      �t�bhhK ��h��R�(KK��h�C%   )        �t�bhhK ��h��R�(KK	��h�C$�      )         �      �      �t�bhhK ��h��R�(KK��h�C�      w        �t�bhhK ��h��R�(KK��h�C,X      )         �                 �t�bhhK ��h��R�(KK��h�C%   )        �t�bhhK ��h��R�(KK��h�C�     ?     �t�bhhK ��h��R�(KK��h�C�     )      �t�bhhK ��h��R�(KK��h�CL   !   �  �  �     t     	   v   B      u         L  )         �t�bhhK ��h��R�(KK��h�C4      �   R  a   �  )           v        �t�bhhK ��h��R�(KK��h�CH   �    w  )   	   i  .      �  
           x  )         �t�bhhK ��h��R�(KK��h�C�     v        �t�bhhK ��h��R�(KK
��h�C(      
   �  O      U   a        �t�bhhK ��h��R�(KK��h�Cl   !   �  y     )   D      z  �     �  �        {     |  }     ~  }    S           �t�bhhK ��h��R�(KK��h�Ch�  N     �     �  $      �   �     �     �           :   �   U     �             �t�bhhK ��h��R�(KK��h�C,         R  a   �  )      v        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CXT  7  �  ?     �  �     �     T   s      �     .   )   �      �        �t�bhhK ��h��R�(KK��h�C@^   >   7  �  ?     �     ?     >   �     !         �t�bhhK ��h��R�(KK	��h�C$.      �      �      �        �t�bhhK ��h��R�(KK��h�C�           E      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�CU           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�CU           �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C,     |      �   r                 �t�bhhK ��h��R�(KK��h�C�  �  ?     T        �t�bhhK ��h��R�(KK
��h�C(7  �  ?     �                 �t�bhhK ��h��R�(KK��h�C'  �     �t�bhhK ��h��R�(KK��h�C0      �   '  �     )         �         �t�bhhK ��h��R�(KK��h�C\   �     �     2         �     ,        �  u      N         �   	        �t�bhhK ��h��R�(KK��h�C<   !   �   �     F      !   )     �   m           �t�bhhK ��h��R�(KK	��h�C$         �  �     �        �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C8    �   a         '  �     �                 �t�bhhK ��h��R�(KK��h�C%   )        �t�bhhK ��h��R�(KK��h�C'  �     �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�Cu   7   F  �   h      �t�bhhK ��h��R�(KK��h�C+      �     �t�bhhK ��h��R�(KK��h�C    H  '   �      �t�bhhK ��h��R�(KK��h�CG     �t�bhhK ��h��R�(KK��h�Cu   7   F  �   h      �t�bhhK ��h��R�(KK��h�C<S      �      S      V     x   /       g   �         �t�bhhK ��h��R�(KK��h�CT
         �     �  g  �   	   6      �   /        d   S      �         �t�bhhK ��h��R�(KK��h�C<      �   /   w  M        1  d   S      �         �t�bhhK ��h��R�(KK��h�C\�     m     �  	   �  	   �     �     �   a        M   S      �           �t�bhhK ��h��R�(KK��h�C4  �  �  �   �   a   1  d   S      �         �t�bhhK ��h��R�(KK
��h�C(w      /   J   [     r   {         �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�CD   
   S      �  ;   7         j   �   �       �        �t�bhhK ��h��R�(KK��h�CL   
       g   �      1   7         j   �      u   7   F  �   h      �t�bhhK ��h��R�(KK��h�C%   �      +        �t�bhhK ��h��R�(KK��h�C�      �           �t�bhhK ��h��R�(KK��h�C�      w        �t�be(hhK ��h��R�(KK��h�C*  �           �t�bhhK ��h��R�(KK��h�C�      �        �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK
��h�C(V          E  �                 �t�bhhK ��h��R�(KK��h�C+      �     �t�bhhK ��h��R�(KK��h�CH   ;           �t�bhhK ��h��R�(KK��h�CP!      u  >   ;      "     x   #      @   �      W     E  �         �t�bhhK ��h��R�(KK��h�C0   !   �   -   Z   �  v   �  �  �        �t�bhhK ��h��R�(KK��h�C4   7         
   H   ;      !   Q   2         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK	��h�C$H   ;      �                 �t�bhhK ��h��R�(KK��h�Cd
      5   +      �            E     �         =   �     �  ~  X  �     %        �t�bhhK ��h��R�(KK
��h�C(   7   P     �  ~  X  2         �t�bhhK ��h��R�(KK��h�C,�  �  H  x   "  �      E  �         �t�bhhK ��h��R�(KK��h�CP      @   +          �  J   �        �  	   �   �     �  �        �t�bhhK ��h��R�(KK��h�CY  $     �t�bhhK ��h��R�(KK��h�C`Y  Z        �  	      T     c      C      �  �   e   �      {  �     �        �t�bhhK ��h��R�(KK	��h�C$�      [     �              �t�bhhK ��h��R�(KK
��h�C(f   
   �                 /     �t�bhhK ��h��R�(KK	��h�C$�  �     �     \  C         �t�bhhK ��h��R�(KK��h�CdM   �        @      �  	        /      �  g  �      �            H  �   �         �t�bhhK ��h��R�(KK��h�C�  y     )         �t�bhhK ��h��R�(KK��h�C �     �   
   �           �t�bhhK ��h��R�(KK��h�CH
         ?     I   	         @   f        M   q   d        �t�bhhK ��h��R�(KK��h�C@�     d  x   /   
      4   "   �   �         �         �t�bhhK ��h��R�(KK��h�CX�     L   C   ]     ]  �  �  ^     x   �      �      �  X      �        �t�bhhK ��h��R�(KK	��h�C$      7         _  2         �t�bhhK ��h��R�(KK��h�CV      L   �      �t�bhhK ��h��R�(KK��h�C    H  '   �      �t�bhhK ��h��R�(KK��h�CD
      "   '   �      !   	         �  �     !   `        �t�bhhK ��h��R�(KK��h�CD!   `  �     �  �     T   �  �     F   X      c         �t�bhhK ��h��R�(KK	��h�C$      7         _  2         �t�bhhK ��h��R�(KK��h�Ctr  0  T   c      +          H  �   �      )   	      	      	   E   	   �   	   s  	   }             �t�bhhK ��h��R�(KK��h�C\   r  0  �   �  
       H  �      C      )   	      	   E   	   �      s        �t�bhhK ��h��R�(KK��h�C�     v        �t�bhhK ��h��R�(KK��h�C0r  0  �   �     )   	         E         �t�bhhK ��h��R�(KK��h�Cd        p     N     Y      6   H  �   �              #       "   �   �         �t�bhhK ��h��R�(KK
��h�C(�   a     )   	         E         �t�bhhK ��h��R�(KK��h�C,         �        r  0  2         �t�bhhK ��h��R�(KK��h�C|~   S      �     S      V     T   �  ;      Y      �         H  �      #           �      H  �         �t�bhhK ��h��R�(KK��h�CX   ~   S      �           F   �      �     g   �         H  �   �         �t�bhhK ��h��R�(KK��h�C              �  '   �      �t�bhhK ��h��R�(KK��h�C ;      �     �           �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�Cb                 �t�bhhK ��h��R�(KK��h�Cb           �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�CG     �t�bhhK ��h��R�(KK	��h�C$�  !  �   Q       9         �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C�  �     �        �t�bhhK ��h��R�(KK��h�C(      �     �t�bhhK ��h��R�(KK��h�C0C      -   9  �        <  =  0        �t�bhhK ��h��R�(KK��h�C`     x   2     �  �  C      U     1          0     �      �  G     (  Z     �t�bhhK ��h��R�(KK��h�C �        <  =  0        �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C         G     �t�bhhK ��h��R�(KK��h�C5        �t�bhhK ��h��R�(KK��h�C�                  �t�bhhK ��h��R�(KK��h�C,c   
   (  Z     �                 �t�bhhK ��h��R�(KK��h�C,4  �   �     /           1         �t�bhhK ��h��R�(KK��h�Cu   7   F  �   h      �t�bhhK ��h��R�(KK��h�C+      �     �t�bhhK ��h��R�(KK��h�C    H  '   �      �t�bhhK ��h��R�(KK��h�CG     �t�bhhK ��h��R�(KK��h�Cu   7   F  �   h      �t�bhhK ��h��R�(KK��h�C<S      �      S      V     x   /       g   �         �t�bhhK ��h��R�(KK��h�CT
         �     �  g  �   	   6      �   /        d   S      �         �t�bhhK ��h��R�(KK��h�C<      �   /   w  M        1  d   S      �         �t�bhhK ��h��R�(KK��h�C\�     m     �  	   �  	   �     �     �   a        M   S      �           �t�bhhK ��h��R�(KK��h�C4  �  �  �   �   a   1  d   S      �         �t�bhhK ��h��R�(KK
��h�C(w      /   J   [     r   {         �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�CD   
   S      �  ;   7         j   �   �       �        �t�bhhK ��h��R�(KK��h�CL   
       g   �      1   7         j   �      u   7   F  �   h      �t�bhhK ��h��R�(KK��h�C%   �      +        �t�bhhK ��h��R�(KK��h�C�      �           �t�bhhK ��h��R�(KK��h�C�      w        �t�bhhK ��h��R�(KK��h�C*  �           �t�bhhK ��h��R�(KK��h�C�      �        �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK
��h�C(V          E  �                 �t�bhhK ��h��R�(KK��h�C+      �     �t�bhhK ��h��R�(KK��h�CH   ;           �t�bhhK ��h��R�(KK��h�CP!      u  >   ;      "     x   #      @   �      W     E  �         �t�bhhK ��h��R�(KK��h�C0   !   �   -   Z   �  v   �  �  �        �t�bhhK ��h��R�(KK��h�C4   7         
   H   ;      !   Q   2         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK	��h�C$H   ;      �                 �t�bhhK ��h��R�(KK��h�Cd
      5   +      �            E     �         =   �     �  ~  X  �     %        �t�bhhK ��h��R�(KK
��h�C(   7   P     �  ~  X  2         �t�bhhK ��h��R�(KK��h�C,�  �  H  x   "  �      E  �         �t�bhhK ��h��R�(KK��h�CP      @   +          �  J   �        �  	   �   �     �  �        �t�bhhK ��h��R�(KK��h�CY  $     �t�bhhK ��h��R�(KK��h�C`Y  Z        �  	      T     c      C      �  �   e   �      {  �     �        �t�bhhK ��h��R�(KK	��h�C$�      [     �              �t�bhhK ��h��R�(KK
��h�C(f   
   �                 /     �t�bhhK ��h��R�(KK	��h�C$�  �     �     \  C         �t�bhhK ��h��R�(KK��h�CdM   �        @      �  	        /      �  g  �      �            H  �   �         �t�bhhK ��h��R�(KK��h�C�  y     )         �t�bhhK ��h��R�(KK��h�C �     �   
   �           �t�bhhK ��h��R�(KK��h�CH
         ?     I   	         @   f        M   q   d        �t�bhhK ��h��R�(KK��h�C@�     d  x   /   
      4   "   �   �         �         �t�bhhK ��h��R�(KK��h�CX�     L   C   ]     ]  �  �  ^     x   �      �      �  X      �        �t�bhhK ��h��R�(KK	��h�C$      7         _  2         �t�bhhK ��h��R�(KK��h�CV      L   �      �t�bhhK ��h��R�(KK��h�C    H  '   �      �t�bhhK ��h��R�(KK��h�CD
      "   '   �      !   	         �  �     !   `        �t�bhhK ��h��R�(KK��h�CD!   `  �     �  �     T   �  �     F   X      c         �t�bhhK ��h��R�(KK	��h�C$      7         _  2         �t�bhhK ��h��R�(KK��h�Ctr  0  T   c      +          H  �   �      )   	      	      	   E   	   �   	   s  	   }             �t�bhhK ��h��R�(KK��h�C\   r  0  �   �  
       H  �      C      )   	      	   E   	   �      s        �t�bhhK ��h��R�(KK��h�C�     v        �t�bhhK ��h��R�(KK��h�C0r  0  �   �     )   	         E         �t�bhhK ��h��R�(KK��h�Cd        p     N     Y      6   H  �   �              #       "   �   �         �t�bhhK ��h��R�(KK
��h�C(�   a     )   	         E         �t�bhhK ��h��R�(KK��h�C,         �        r  0  2         �t�bhhK ��h��R�(KK��h�C|~   S      �     S      V     T   �  ;      Y      �         H  �      #           �      H  �         �t�bhhK ��h��R�(KK��h�CX   ~   S      �           F   �      �     g   �         H  �   �         �t�bhhK ��h��R�(KK��h�C              �  '   �      �t�bhhK ��h��R�(KK��h�C ;      �     �           �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�Cb                 �t�bhhK ��h��R�(KK��h�Cb           �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�CG     �t�bhhK ��h��R�(KK	��h�C$�  !  �   Q       9         �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C�  �     �        �t�bhhK ��h��R�(KK��h�C(      �     �t�bhhK ��h��R�(KK��h�C0C      -   9  �        <  =  0        �t�bhhK ��h��R�(KK��h�C`     x   2     �  �  C      U     1          0     �      �  G     (  Z     �t�bhhK ��h��R�(KK��h�C �        <  =  0        �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C         G     �t�bhhK ��h��R�(KK��h�C5        �t�bhhK ��h��R�(KK��h�C�                  �t�bhhK ��h��R�(KK��h�C,c   
   (  Z     �                 �t�bhhK ��h��R�(KK��h�C,4  �   �     /           1         �t�bhhK ��h��R�(KK��h�Cu   7   F  �   h      �t�bhhK ��h��R�(KK��h�C+      �     �t�bhhK ��h��R�(KK��h�C    H  '   �      �t�bhhK ��h��R�(KK��h�CG     �t�bhhK ��h��R�(KK��h�Cu   7   F  �   h      �t�bhhK ��h��R�(KK��h�C<S      �      S      V     x   /       g   �         �t�bhhK ��h��R�(KK��h�CT
         �     �  g  �   	   6      �   /        d   S      �         �t�bhhK ��h��R�(KK��h�C<      �   /   w  M        1  d   S      �         �t�bhhK ��h��R�(KK��h�C\�     m     �  	   �  	   �     �     �   a        M   S      �           �t�bhhK ��h��R�(KK��h�C4  �  �  �   �   a   1  d   S      �         �t�bhhK ��h��R�(KK
��h�C(w      /   J   [     r   {         �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�CD   
   S      �  ;   7         j   �   �       �        �t�bhhK ��h��R�(KK��h�CL   
       g   �      1   7         j   �      u   7   F  �   h      �t�bhhK ��h��R�(KK��h�C%   �      +        �t�bhhK ��h��R�(KK��h�C�      �           �t�bhhK ��h��R�(KK��h�C�      w        �t�bhhK ��h��R�(KK��h�C*  �           �t�bhhK ��h��R�(KK��h�C�      �        �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK
��h�C(V          E  �                 �t�bhhK ��h��R�(KK��h�C+      �     �t�bhhK ��h��R�(KK��h�CH   ;           �t�bhhK ��h��R�(KK��h�CP!      u  >   ;      "     x   #      @   �      W     E  �         �t�bhhK ��h��R�(KK��h�C0   !   �   -   Z   �  v   �  �  �        �t�bhhK ��h��R�(KK��h�C4   7         
   H   ;      !   Q   2         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK	��h�C$H   ;      �                 �t�bhhK ��h��R�(KK��h�Cd
      5   +      �            E     �         =   �     �  ~  X  �     %        �t�bhhK ��h��R�(KK
��h�C(   7   P     �  ~  X  2         �t�bhhK ��h��R�(KK��h�C,�  �  H  x   "  �      E  �         �t�bhhK ��h��R�(KK��h�CP      @   +          �  J   �        �  	   �   �     �  �        �t�bhhK ��h��R�(KK��h�CY  $     �t�bhhK ��h��R�(KK��h�C`Y  Z        �  	      T     c      C      �  �   e   �      {  �     �        �t�bhhK ��h��R�(KK	��h�C$�      [     �              �t�bhhK ��h��R�(KK
��h�C(f   
   �                 /     �t�bhhK ��h��R�(KK	��h�C$�  �     �     \  C         �t�bhhK ��h��R�(KK��h�CdM   �        @      �  	        /      �  g  �      �            H  �   �         �t�bhhK ��h��R�(KK��h�C�  y     )         �t�bhhK ��h��R�(KK��h�C �     �   
   �           �t�bhhK ��h��R�(KK��h�CH
         ?     I   	         @   f        M   q   d        �t�bhhK ��h��R�(KK��h�C@�     d  x   /   
      4   "   �   �         �         �t�bhhK ��h��R�(KK��h�CX�     L   C   ]     ]  �  �  ^     x   �      �      �  X      �        �t�bhhK ��h��R�(KK	��h�C$      7         _  2         �t�bhhK ��h��R�(KK��h�CV      L   �      �t�bhhK ��h��R�(KK��h�C    H  '   �      �t�bhhK ��h��R�(KK��h�CD
      "   '   �      !   	         �  �     !   `        �t�bhhK ��h��R�(KK��h�CD!   `  �     �  �     T   �  �     F   X      c         �t�bhhK ��h��R�(KK	��h�C$      7         _  2         �t�bhhK ��h��R�(KK��h�Ctr  0  T   c      +          H  �   �      )   	      	      	   E   	   �   	   s  	   }             �t�bhhK ��h��R�(KK��h�C\   r  0  �   �  
       H  �      C      )   	      	   E   	   �      s        �t�bhhK ��h��R�(KK��h�C�     v        �t�bhhK ��h��R�(KK��h�C0r  0  �   �     )   	         E         �t�bhhK ��h��R�(KK��h�Cd        p     N     Y      6   H  �   �              #       "   �   �         �t�bhhK ��h��R�(KK
��h�C(�   a     )   	         E         �t�bhhK ��h��R�(KK��h�C,         �        r  0  2         �t�bhhK ��h��R�(KK��h�C|~   S      �     S      V     T   �  ;      Y      �         H  �      #           �      H  �         �t�bhhK ��h��R�(KK��h�CX   ~   S      �           F   �      �     g   �         H  �   �         �t�bhhK ��h��R�(KK��h�C              �  '   �      �t�bhhK ��h��R�(KK��h�C ;      �     �           �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�Cb                 �t�bhhK ��h��R�(KK��h�Cb           �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�CG     �t�bhhK ��h��R�(KK	��h�C$�  !  �   Q       9         �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C�  �     �        �t�bhhK ��h��R�(KK��h�C(      �     �t�bhhK ��h��R�(KK��h�C0C      -   9  �        <  =  0        �t�bhhK ��h��R�(KK��h�C`     x   2     �  �  C      U     1          0     �      �  G     (  Z     �t�bhhK ��h��R�(KK��h�C �        <  =  0        �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C         G     �t�bhhK ��h��R�(KK��h�C5        �t�bhhK ��h��R�(KK��h�C�                  �t�bhhK ��h��R�(KK��h�C,c   
   (  Z     �                 �t�bhhK ��h��R�(KK��h�C,4  �   �     /           1         �t�bhhK ��h��R�(KK��h�Cc         $     C      �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C5         �   h      �t�bhhK ��h��R�(KK��h�Cc         $     C      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C!   Q   ;      C   �     �t�bhhK ��h��R�(KK��h�C�     C      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�Cl!   Q   ;      C      �   �     p   /      
   $  	   0      �      
   H      >   �  ;         �t�bhhK ��h��R�(KK��h�Ct      �  �  
      �     1      �     �  	        	   �     �     "   �         �   �         �t�bhhK ��h��R�(KK��h�C,(      <      �        <      �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�CH         �  �     p   c      C      v   �   Z   �  �        �t�bhhK ��h��R�(KK��h�C         	   �        �t�bhhK ��h��R�(KK��h�C(      <            �t�bhhK ��h��R�(KK��h�C   �        �t�bhhK ��h��R�(KK��h�C c      +     �            �t�bhhK ��h��R�(KK��h�C4^  p   /      
   
  �  Q      �  ;         �t�bhhK ��h��R�(KK
��h�C(�        �  	   �     �        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK	��h�C$�  	   G  �  	   �  �        �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C,P     �  7         !   Q   2         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK/��h�C�&   ~  �     �     �  �  �     "      �     �   C      �  	   �     W   p     !   	      �   �     
      F   R  	   ~  	   �   	   �  	   o     M  �         �t�bhhK ��h��R�(KK��h�C,�    �  	   �     :     �        �t�bhhK ��h��R�(KK	��h�C$(      <      �     �        �t�bhhK ��h��R�(KK��h�C�  �     �        �t�bhhK ��h��R�(KK��h�C0c      �            E      �      �      �t�bhhK ��h��R�(KK#��h�C�   �     �  �   c  ^     �   c  �  �  �           �   
   �     �     F   W  	   (  Z  	   G   	   X      {         �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�CS  �     �t�bhhK ��h��R�(KK
��h�C(�  C     �  =  e  	   �        �t�bhhK ��h��R�(KK	��h�C$!   �     <      �     �     �t�bhhK ��h��R�(KK��h�C�  :     �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�Cc      �      �t�bhhK ��h��R�(KK��h�Cp
      "   �     �   �  	            <  =  0     4     @   c      �     '                �t�bhhK ��h��R�(KK��h�C,4  �   �     /           1         �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�CD&   �   �     �     x   /       E  �  ;      J   �        �t�bhhK ��h��R�(KK��h�CL!         ~   S      �  �      �   �      d    C      !         �t�bhhK ��h��R�(KK
��h�C(   "   �       @      �   �   
      �t�bhhK ��h��R�(KK��h�CJ   S     !      �t�bhhK ��h��R�(KK��h�C@   "   �     !   U   '   e   #        z       1      �t�bhhK ��h��R�(KK
��h�C(  �   �   4   "   �     /         �t�bhhK ��h��R�(KK��h�C0   "   �  S     1           I         �t�bhhK ��h��R�(KK��h�C\   &   �   �  O         
   X      )         	   �  	   X      ;      !         �t�bhhK ��h��R�(KK��h�C4   &   �   �  [  B         +      �         �t�bhhK ��h��R�(KK��h�C&   �   �     �        �t�bhhK ��h��R�(KK��h�C�  
   �   �      �t�bhhK ��h��R�(KK��h�CT      $     �   �   M             i        �      }   �   ]         �t�bhhK ��h��R�(KK��h�C(   �  	   �     �     �t�bhhK ��h��R�(KK��h�C<
      �  �   	   �     �   /      S      �         �t�bhhK ��h��R�(KK	��h�C$S      �   �  &   �   �        �t�bhhK ��h��R�(KK��h�C<      
   &   �   �     )     j   2   Z     1      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�C5         �   h      �t�bhhK ��h��R�(KK$��h�C�
      �   9  �      {  	   5  4      )            .   4        �   e   k      �            	         �      �        �t�bhhK ��h��R�(KK��h�C0         �  
      5      �         �t�bhhK ��h��R�(KK��h�C,  �       �   O      �  �        �t�bhhK ��h��R�(KK��h�CL
      %  �       �  �  	         �     �   N      a        �t�bhhK ��h��R�(KK	��h�C$         5         �   h      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   �     �t�bhhK ��h��R�(KK��h�C�   �     �        �t�bhhK ��h��R�(KK	��h�C$�  �      �                 �t�bhhK ��h��R�(KK��h�Cc         $     C      �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C5         �   h      �t�bhhK ��h��R�(KK��h�Cc         $     C      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C!   Q   ;      C   �     �t�bhhK ��h��R�(KK��h�C�     C      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�Cl!   Q   ;      C      �   �     p   /      
   $  	   0      �      
   H      >   �  ;         �t�bhhK ��h��R�(KK��h�Ct      �  �  
      �     1      �     �  	        	   �     �     "   �         �   �         �t�bhhK ��h��R�(KK��h�C,(      <      �        <      �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�CH         �  �     p   c      C      v   �   Z   �  �        �t�bhhK ��h��R�(KK��h�C         	   �        �t�bhhK ��h��R�(KK��h�C(      <            �t�bhhK ��h��R�(KK��h�C   �        �t�bhhK ��h��R�(KK��h�C c      +     �            �t�bhhK ��h��R�(KK��h�C4^  p   /      
   
  �  Q      �  ;         �t�bhhK ��h��R�(KK
��h�C(�        �  	   �     �        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK	��h�C$�  	   G  �  	   �  �        �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C,P     �  7         !   Q   2         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK/��h�C�&   ~  �     �     �  �  �     "      �     �   C      �  	   �     W   p     !   	      �   �     
      F   R  	   ~  	   �   	   �  	   o     M  �         �t�bhhK ��h��R�(KK��h�C,�    �  	   �     :     �        �t�bhhK ��h��R�(KK	��h�C$(      <      �     �        �t�bhhK ��h��R�(KK��h�C�  �     �        �t�bhhK ��h��R�(KK��h�C0c      �            E      �      �      �t�bhhK ��h��R�(KK#��h�C�   �     �  �   c  ^     �   c  �  �  �           �   
   �     �     F   W  	   (  Z  	   G   	   X      {         �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�CS  �     �t�bhhK ��h��R�(KK
��h�C(�  C     �  =  e  	   �        �t�bhhK ��h��R�(KK	��h�C$!   �     <      �     �     �t�bhhK ��h��R�(KK��h�C�  :     �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�Cc      �      �t�bhhK ��h��R�(KK��h�Cp
      "   �     �   �  	            <  =  0     4     @   c      �     '                �t�bhhK ��h��R�(KK��h�C,4  �   �     /           1         �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�CD&   �   �     �     x   /       E  �  ;      J   �        �t�bhhK ��h��R�(KK��h�CL!         ~   S      �  �      �   �      d    C      !         �t�bhhK ��h��R�(KK
��h�C(   "   �       @      �   �   
      �t�bhhK ��h��R�(KK��h�CJ   S     !      �t�bhhK ��h��R�(KK��h�C@   "   �     !   U   '   e   #        z       1      �t�bhhK ��h��R�(KK
��h�C(  �   �   4   "   �     /         �t�bhhK ��h��R�(KK��h�C0   "   �  S     1           I         �t�bhhK ��h��R�(KK��h�C\   &   �   �  O         
   X      )         	   �  	   X      ;      !         �t�bhhK ��h��R�(KK��h�C4   &   �   �  [  B         +      �         �t�bhhK ��h��R�(KK��h�C&   �   �     �        �t�bhhK ��h��R�(KK��h�C�  
   �   �      �t�bhhK ��h��R�(KK��h�CT      $     �   �   M             i        �      }   �   ]         �t�bhhK ��h��R�(KK��h�C(   �  	   �     �     �t�bhhK ��h��R�(KK��h�C<
      �  �   	   �     �   /      S      �         �t�bhhK ��h��R�(KK	��h�C$S      �   �  &   �   �        �t�bhhK ��h��R�(KK��h�C<      
   &   �   �     )     j   2   Z     1      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�C5         �   h      �t�bhhK ��h��R�(KK$��h�C�
      �   9  �      {  	   5  4      )            .   4        �   e   k      �            	         �      �        �t�bhhK ��h��R�(KK��h�C0         �  
      5      �         �t�bhhK ��h��R�(KK��h�C,  �       �   O      �  �        �t�bhhK ��h��R�(KK��h�CL
      %  �       �  �  	         �     �   N      a        �t�bhhK ��h��R�(KK	��h�C$         5         �   h      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   �     �t�bhhK ��h��R�(KK��h�C�   �     �        �t�bhhK ��h��R�(KK	��h�C$�  �      �                 �t�bhhK ��h��R�(KK��h�Cc         $     C      �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C5         �   h      �t�bhhK ��h��R�(KK��h�Cc         $     C      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C!   Q   ;      C   �     �t�bhhK ��h��R�(KK��h�C�     C      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�Cl!   Q   ;      C      �   �     p   /      
   $  	   0      �      
   H      >   �  ;         �t�bhhK ��h��R�(KK��h�Ct      �  �  
      �     1      �     �  	        	   �     �     "   �         �   �         �t�bhhK ��h��R�(KK��h�C,(      <      �        <      �     �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C4^  p   /      
   
  �  Q      �  ;         �t�bhhK ��h��R�(KK
��h�C(�        �  	   �     �        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK	��h�C$�  	   G  �  	   �  �        �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C,P     �  7         !   Q   2         �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK/��h�C�&   ~  �     �     �  �  �     "      �     �   C      �  	   �     W   p     !   	      �   �     
      F   R  	   ~  	   �   	   �  	   o     M  �         �t�bhhK ��h��R�(KK��h�C,�    �  	   �     :     �        �t�bhhK ��h��R�(KK	��h�C$(      <      �     �        �t�bhhK ��h��R�(KK��h�C�  �     �        �t�bhhK ��h��R�(KK��h�C0c      �            E      �      �      �t�bhhK ��h��R�(KK#��h�C�   �     �  �   c  ^     �   c  �  �  �           �   
   �     �     F   W  	   (  Z  	   G   	   X      {         �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�CS  �     �t�bhhK ��h��R�(KK
��h�C(�  C     �  =  e  	   �        �t�bhhK ��h��R�(KK	��h�C$!   �     <      �     �     �t�bhhK ��h��R�(KK��h�C�  :     �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�Cc      �      �t�bhhK ��h��R�(KK��h�Cp
      "   �     �   �  	            <  =  0     4     @   c      �     '                �t�bhhK ��h��R�(KK��h�C,4  �   �     /           1         �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�CD&   �   �     �     x   /       E  �  ;      J   �        �t�bhhK ��h��R�(KK��h�CL!         ~   S      �  �      �   �      d    C      !         �t�bhhK ��h��R�(KK
��h�C(   "   �       @      �   �   
      �t�bhhK ��h��R�(KK��h�CJ   S     !      �t�bhhK ��h��R�(KK��h�C@   "   �     !   U   '   e   #        z       1      �t�bhhK ��h��R�(KK
��h�C(  �   �   4   "   �     /         �t�bhhK ��h��R�(KK��h�C0   "   �  S     1           I         �t�bhhK ��h��R�(KK��h�C\   &   �   �  O         
   X      )         	   �  	   X      ;      !         �t�bhhK ��h��R�(KK��h�C4   &   �   �  [  B         +      �         �t�bhhK ��h��R�(KK��h�C&   �   �     �        �t�bhhK ��h��R�(KK��h�C�  
   �   �      �t�bhhK ��h��R�(KK��h�CT      $     �   �   M             i        �      }   �   ]         �t�bhhK ��h��R�(KK��h�C(   �  	   �     �     �t�bhhK ��h��R�(KK��h�C<
      �  �   	   �     �   /      S      �         �t�bhhK ��h��R�(KK	��h�C$S      �   �  &   �   �        �t�bhhK ��h��R�(KK��h�C<      
   &   �   �     )     j   2   Z     1      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�C5         �   h      �t�bhhK ��h��R�(KK$��h�C�
      �   9  �      {  	   5  4      )            .   4        �   e   k      �            	         �      �        �t�bhhK ��h��R�(KK��h�C0         �  
      5      �         �t�bhhK ��h��R�(KK��h�C,  �       �   O      �  �        �t�bhhK ��h��R�(KK��h�CL
      %  �       �  �  	         �     �   N      a        �t�bhhK ��h��R�(KK	��h�C$         5         �   h      �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C   
   �     �t�bhhK ��h��R�(KK��h�C�   �     �        �t�bhhK ��h��R�(KK	��h�C$�  �      �                 �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CH   �  �     9         i   
   {      I  m     �  ,        �t�bhhK ��h��R�(KK��h�C�  �     9         �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�CP      D   i   
   Z   �  {      m          "     q   �  1         �t�bhhK ��h��R�(KK��h�Ch
      4      �         �      B  	   �        `      �     �   �   &      �  �        �t�bhhK ��h��R�(KK��h�C8�       �      �      }      �     d        �t�bhhK ��h��R�(KK
��h�C(      �      }      �  �        �t�bhhK ��h��R�(KK��h�C,3      d  4      e  c   
   �        �t�bhhK ��h��R�(KK��h�C          �     1         �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C'  �                 �t�bhhK ��h��R�(KK��h�C'  �                 �t�bhhK ��h��R�(KK��h�C     |      �t�bhhK ��h��R�(KK��h�CL
        r   �  �      !   	   6      I  /      |      ]        �t�bhhK ��h��R�(KK��h�C       I  /      �         �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�Ck  �     �t�bhhK ��h��R�(KK��h�C     �  �     �t�bhhK ��h��R�(KK��h�C,N      �     �   6      w      /      �t�bhhK ��h��R�(KK��h�C[        F   �        �t�bhhK ��h��R�(KK��h�C0{      *     
      5   {      1         �t�bhhK ��h��R�(KK��h�C<+  ;  �     �  �     
         m     �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C  n   -        �t�bhhK ��h��R�(KK	��h�C$3      4  �  6   �  .        �t�bhhK ��h��R�(KK��h�CT   O         
       �    �     �      �     r   �   #     1         �t�bhhK ��h��R�(KK��h�C               |         �t�bhhK ��h��R�(KK��h�C      �                 �t�bhhK ��h��R�(KK��h�Cp
      "   �     �   �  	            <  =  0     4     @   c      �     '                �t�bhhK ��h��R�(KK��h�C      @         �t�bhhK ��h��R�(KK��h�C0�  c         :      �     ^   >   k      �t�bhhK ��h��R�(KK��h�C4   4  �  	   I  /      |      �   J   �      �t�bhhK ��h��R�(KK��h�C �     �  \   c   
   �     �t�bhhK ��h��R�(KK	��h�C$   
   &   �  �     �  �     �t�bhhK ��h��R�(KK��h�C4c   
   �      �     
       �  �     �     �t�bhhK ��h��R�(KK	��h�C$c   
   �     
              �t�bhhK ��h��R�(KK��h�Cc   
        �t�bhhK ��h��R�(KK��h�Cc      �              �t�bhhK ��h��R�(KK��h�Cpf  4  �  g  h  x   /       E  �   {        &   7         
   _       6   w                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C,4  �   �     /           1         �t�bhhK ��h��R�(KK��h�Cf  4  �  g  h        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CH   �  �     9         i   
   {      I  m     �  ,        �t�bhhK ��h��R�(KK��h�C�  �     9         �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�CP      D   i   
   Z   �  {      m          "     q   �  1         �t�bhhK ��h��R�(KK��h�Ch
      4      �         �      B  	   �        `      �     �   �   &      �  �        �t�bhhK ��h��R�(KK��h�C8�       �      �      }      �     d        �t�bhhK ��h��R�(KK
��h�C(      �      }      �  �        �t�bhhK ��h��R�(KK��h�C,3      d  4      e  c   
   �        �t�bhhK ��h��R�(KK��h�C          �     1         �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C'  �                 �t�bhhK ��h��R�(KK��h�C'  �                 �t�bhhK ��h��R�(KK��h�C     |      �t�bhhK ��h��R�(KK��h�CL
        r   �  �      !   	   6      I  /      |      ]        �t�bhhK ��h��R�(KK��h�C       I  /      �         �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�Ck  �     �t�bhhK ��h��R�(KK��h�C     �  �     �t�bhhK ��h��R�(KK��h�C,N      �     �   6      w      /      �t�bhhK ��h��R�(KK��h�C[        F   �        �t�bhhK ��h��R�(KK��h�C0{      *     
      5   {      1         �t�bhhK ��h��R�(KK��h�C<+  ;  �     �  �     
         m     �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C  n   -        �t�bhhK ��h��R�(KK	��h�C$3      4  �  6   �  .        �t�bhhK ��h��R�(KK��h�CT   O         
       �    �     �      �     r   �   #     1         �t�bhhK ��h��R�(KK��h�C               |         �t�bhhK ��h��R�(KK��h�C      �                 �t�bhhK ��h��R�(KK��h�Cp
      "   �     �   �  	            <  =  0     4     @   c      �     '                �t�bhhK ��h��R�(KK��h�C      @         �t�bhhK ��h��R�(KK��h�C0�  c         :      �     ^   >   k      �t�bhhK ��h��R�(KK��h�C4   4  �  	   I  /      |      �   J   �      �t�bhhK ��h��R�(KK��h�C �     �  \   c   
   �     �t�bhhK ��h��R�(KK	��h�C$   
   &   �  �     �  �     �t�bhhK ��h��R�(KK��h�C4c   
   �      �     
       �  �     �     �t�bhhK ��h��R�(KK	��h�C$c   
   �     
              �t�bhhK ��h��R�(KK��h�Cc   
        �t�bhhK ��h��R�(KK��h�Cc      �              �t�bhhK ��h��R�(KK��h�Cpf  4  �  g  h  x   /       E  �   {        &   7         
   _       6   w                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C,4  �   �     /           1         �t�bhhK ��h��R�(KK��h�Cf  4  �  g  h        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CH   �  �     9         i   
   {      I  m     �  ,        �t�bhhK ��h��R�(KK��h�C�  �     9         �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�CP      D   i   
   Z   �  {      m          "     q   �  1         �t�bhhK ��h��R�(KK��h�Ch
      4      �         �      B  	   �        `      �     �   �   &      �  �        �t�bhhK ��h��R�(KK��h�C8�       �      �      }      �     d        �t�bhhK ��h��R�(KK
��h�C(      �      }      �  �        �t�bhhK ��h��R�(KK��h�C,3      d  4      e  c   
   �        �t�bhhK ��h��R�(KK��h�C          �     1         �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C'  �                 �t�bhhK ��h��R�(KK��h�C'  �                 �t�bhhK ��h��R�(KK��h�C     |      �t�bhhK ��h��R�(KK��h�CL
        r   �  �      !   	   6      I  /      |      ]        �t�bhhK ��h��R�(KK��h�C       I  /      �         �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�Ck  �     �t�bhhK ��h��R�(KK��h�C     �  �     �t�bhhK ��h��R�(KK��h�C,N      �     �   6      w      /      �t�bhhK ��h��R�(KK��h�C[        F   �        �t�bhhK ��h��R�(KK��h�C0{      *     
      5   {      1         �t�bhhK ��h��R�(KK��h�C<+  ;  �     �  �     
         m     �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C  n   -        �t�bhhK ��h��R�(KK	��h�C$3      4  �  6   �  .        �t�bhhK ��h��R�(KK��h�CT   O         
       �    �     �      �     r   �   #     1         �t�bhhK ��h��R�(KK��h�C               |         �t�bhhK ��h��R�(KK��h�C      �                 �t�bhhK ��h��R�(KK��h�Cp
      "   �     �   �  	            <  =  0     4     @   c      �     '                �t�bhhK ��h��R�(KK��h�C      @         �t�bhhK ��h��R�(KK��h�C0�  c         :      �     ^   >   k      �t�bhhK ��h��R�(KK��h�C4   4  �  	   I  /      |      �   J   �      �t�bhhK ��h��R�(KK��h�C �     �  \   c   
   �     �t�bhhK ��h��R�(KK	��h�C$   
   &   �  �     �  �     �t�bhhK ��h��R�(KK��h�C4c   
   �      �     
       �  �     �     �t�bhhK ��h��R�(KK	��h�C$c   
   �     
              �t�bhhK ��h��R�(KK��h�Cc   
        �t�bhhK ��h��R�(KK��h�Cc      �              �t�bhhK ��h��R�(KK��h�Cpf  4  �  g  h  x   /       E  �   {        &   7         
   _       6   w                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C,4  �   �     /           1         �t�bhhK ��h��R�(KK��h�Cf  4  �  g  h        �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CJ     �t�bhhK ��h��R�(KK	��h�C$*      �  �   "   R          �t�bhhK ��h��R�(KK	��h�C$   *      ^                �t�bhhK ��h��R�(KK��h�C   �      ^   >        �t�bhhK ��h��R�(KK
��h�C(      f      �                 �t�bhhK ��h��R�(KK��h�CD*   �  �  X  �   �     �     	      �   J     �         �t�bhhK ��h��R�(KK��h�C4      g      
   �          �           �t�bhhK ��h��R�(KK��h�C<q   p   /   f   
   >     U   '   x     '   e         �t�bhhK ��h��R�(KK��h�C ?                 E      �t�bhhK ��h��R�(KK��h�C,   J        �     9     &        �t�bhhK ��h��R�(KK
��h�C(   :  �      �   @     �        �t�bhhK ��h��R�(KK��h�C@      
   	     �  �     *   7         �  2         �t�bhhK ��h��R�(KK��h�C@      -   �      B     <        C        �        �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK��h�C         ]     �t�bhhK ��h��R�(KK��h�CX
      �        ]     *         g      Y  �     �     �     �        �t�bhhK ��h��R�(KK��h�C0
                           E      �t�bhhK ��h��R�(KK��h�C@      9   	   !      *      �               �        �t�bhhK ��h��R�(KK��h�C�     R        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�C8      �  �     Z   �     �  �     J        �t�bhhK ��h��R�(KK
��h�C(9      !   >  �   �    !         �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C
                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C    *   E  �      �        �t�bhhK ��h��R�(KK��h�C0   �  F    G     H  >   �  {        �t�bhhK ��h��R�(KK	��h�C$I  �  u   �  I   2  �        �t�bhhK ��h��R�(KK��h�C@     *      �  �     �     �      Z   >   �        �t�bhhK ��h��R�(KK��h�C@      e  %               F   M   .   &          �t�bhhK ��h��R�(KK��h�C0      �             w   '           �t�bhhK ��h��R�(KK��h�C4      
   �        �     *   Q   2         �t�bhhK ��h��R�(KK��h�C<   *         �     �  �        H   �          �t�bhhK ��h��R�(KK��h�CP   *      Z   �  �   	   �     W   �   M   _     D      �  �        �t�bhhK ��h��R�(KK��h�C              Y     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C    
                    �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cm                   �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                   �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C,Z     S     ?     *      9         �t�bhhK ��h��R�(KK��h�C@M   q   �  �        g      g  .     K     L        �t�bhhK ��h��R�(KK
��h�C(         T     �     1         �t�bhhK ��h��R�(KK��h�C  M           �t�bhhK ��h��R�(KK��h�CA   �   �        �t�bhhK ��h��R�(KK	��h�C$�      �   O                 �t�bhhK ��h��R�(KK��h�C�   �   �        �t�bhhK ��h��R�(KK��h�C�   N     E      �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK	��h�C$*            �  �   6        �t�bhhK ��h��R�(KK
��h�C(.   �     9   	     
   �         �t�bhhK ��h��R�(KK��h�C<7  �     .   ^     �  	             *         �t�bhhK ��h��R�(KK��h�C*   "       |         �t�bhhK ��h��R�(KK��h�C:   �       �        �t�bhhK ��h��R�(KK��h�C<i  �  �          �     /  �  "   W   f        �t�bhhK ��h��R�(KK��h�C<�  *         �  	   @       �     �        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C,!  u   �       i  "  I   `        �t�bhhK ��h��R�(KK��h�C �   u   #  *   $  %        �t�bhhK ��h��R�(KK��h�C4   &     Z  '  Z   (  U   )     *         �t�bhhK ��h��R�(KK��h�C8   *     Z  �   *      +  �     Z   ,        �t�bhhK ��h��R�(KK��h�C8   *   -  �  .     A    /     j  �        �t�bhhK ��h��R�(KK��h�C8N   1   �           0  �   9   1  I   2        �t�bhhK ��h��R�(KK��h�C<-   
   9   3  s  	   u   *   4  �     5  6        �t�bhhK ��h��R�(KK��h�C47     *   �   8  U         9     Z        �t�bhhK ��h��R�(KK��h�C<I   :  A  *   ;  |      h  I   �    <  |         �t�bhhK ��h��R�(KK��h�C *   �         I   P        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CJ     �t�bhhK ��h��R�(KK	��h�C$*      �  �   "   R          �t�bhhK ��h��R�(KK	��h�C$   *      ^                �t�bhhK ��h��R�(KK��h�C   �      ^   >        �t�bhhK ��h��R�(KK
��h�C(      f      �                 �t�bhhK ��h��R�(KK��h�CD*   �  �  X  �   �     �     	      �   J     �         �t�bhhK ��h��R�(KK��h�C4      g      
   �          �           �t�bhhK ��h��R�(KK��h�C<q   p   /   f   
   >     U   '   x     '   e         �t�bhhK ��h��R�(KK��h�C ?                 E      �t�bhhK ��h��R�(KK��h�C,   J        �     9     &        �t�bhhK ��h��R�(KK
��h�C(   :  �      �   @     �        �t�bhhK ��h��R�(KK��h�C@      
   	     �  �     *   7         �  2         �t�bhhK ��h��R�(KK��h�C@      -   �      B     <        C        �        �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK��h�C         ]     �t�bhhK ��h��R�(KK��h�CX
      �        ]     *         g      Y  �     �     �     �        �t�bhhK ��h��R�(KK��h�C0
                           E      �t�bhhK ��h��R�(KK��h�C@      9   	   !      *      �               �        �t�bhhK ��h��R�(KK��h�C�     R        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�C8      �  �     Z   �     �  �     J        �t�b�
      hhK ��h��R�(KK
��h�C(9      !   >  �   �    !         �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C
                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C    *   E  �      �        �t�bhhK ��h��R�(KK��h�C0   �  F    G     H  >   �  {        �t�bhhK ��h��R�(KK	��h�C$I  �  u   �  I   2  �        �t�bhhK ��h��R�(KK��h�C@     *      �  �     �     �      Z   >   �        �t�bhhK ��h��R�(KK��h�C@      e  %               F   M   .   &          �t�bhhK ��h��R�(KK��h�C0      �             w   '           �t�bhhK ��h��R�(KK��h�C4      
   �        �     *   Q   2         �t�bhhK ��h��R�(KK��h�C<   *         �     �  �        H   �          �t�bhhK ��h��R�(KK��h�CP   *      Z   �  �   	   �     W   �   M   _     D      �  �        �t�bhhK ��h��R�(KK��h�C              Y     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C    
                    �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cm                   �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                   �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C,Z     S     ?     *      9         �t�bhhK ��h��R�(KK��h�C@M   q   �  �        g      g  .     K     L        �t�bhhK ��h��R�(KK
��h�C(         T     �     1         �t�bhhK ��h��R�(KK��h�C  M           �t�bhhK ��h��R�(KK��h�CA   �   �        �t�bhhK ��h��R�(KK	��h�C$�      �   O                 �t�bhhK ��h��R�(KK��h�C�   �   �        �t�bhhK ��h��R�(KK��h�C�   N     E      �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK	��h�C$*            �  �   6        �t�bhhK ��h��R�(KK
��h�C(.   �     9   	     
   �         �t�bhhK ��h��R�(KK��h�C<7  �     .   ^     �  	             *         �t�bhhK ��h��R�(KK��h�C*   "       |         �t�bhhK ��h��R�(KK��h�C:   �       �        �t�bhhK ��h��R�(KK��h�C<i  �  �          �     /  �  "   W   f        �t�bhhK ��h��R�(KK��h�C<�  *         �  	   @       �     �        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C,!  u   �       i  "  I   `        �t�bhhK ��h��R�(KK��h�C �   u   #  *   $  %        �t�bhhK ��h��R�(KK��h�C4   &     Z  '  Z   (  U   )     *         �t�bhhK ��h��R�(KK��h�C8   *     Z  �   *      +  �     Z   ,        �t�bhhK ��h��R�(KK��h�C8   *   -  �  .     A    /     j  �        �t�bhhK ��h��R�(KK��h�C8N   1   �           0  �   9   1  I   2        �t�bhhK ��h��R�(KK��h�C<-   
   9   3  s  	   u   *   4  �     5  6        �t�bhhK ��h��R�(KK��h�C47     *   �   8  U         9     Z        �t�bhhK ��h��R�(KK��h�C<I   :  A  *   ;  |      h  I   �    <  |         �t�bhhK ��h��R�(KK��h�C *   �         I   P        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CJ     �t�bhhK ��h��R�(KK	��h�C$*      �  �   "   R          �t�bhhK ��h��R�(KK	��h�C$   *      ^                �t�bhhK ��h��R�(KK��h�C   �      ^   >        �t�bhhK ��h��R�(KK
��h�C(      f      �                 �t�bhhK ��h��R�(KK��h�CD*   �  �  X  �   �     �     	      �   J     �         �t�bhhK ��h��R�(KK��h�C4      g      
   �          �           �t�bhhK ��h��R�(KK��h�C<q   p   /   f   
   >     U   '   x     '   e         �t�bhhK ��h��R�(KK��h�C?                 �t�bhhK ��h��R�(KK��h�C,   J        �     9     &        �t�bhhK ��h��R�(KK
��h�C(   :  �      �   @     �        �t�bhhK ��h��R�(KK��h�C@      
   	     �  �     *   7         �  2         �t�bhhK ��h��R�(KK��h�C@      -   �      B     <        C        �        �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK��h�C         ]     �t�bhhK ��h��R�(KK��h�CX
      �        ]     *         g      Y  �     �     �     �        �t�bhhK ��h��R�(KK��h�C0
                           E      �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�C8      �  �     Z   �     �  �     J        �t�bhhK ��h��R�(KK
��h�C(9      !   >  �   �    !         �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C
                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C    *   E  �      �        �t�bhhK ��h��R�(KK��h�C0   �  F    G     H  >   �  {        �t�bhhK ��h��R�(KK	��h�C$I  �  u   �  I   2  �        �t�bhhK ��h��R�(KK��h�C@     *      �  �     �     �      Z   >   �        �t�bhhK ��h��R�(KK��h�C@      e  %               F   M   .   &          �t�bhhK ��h��R�(KK��h�C0      �             w   '           �t�bhhK ��h��R�(KK��h�C4      
   �        �     *   Q   2         �t�bhhK ��h��R�(KK��h�C<   *         �     �  �        H   �          �t�bhhK ��h��R�(KK��h�CP   *      Z   �  �   	   �     W   �   M   _     D      �  �        �t�bhhK ��h��R�(KK��h�C              Y     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C    
                    �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cm                   �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                   �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C,Z     S     ?     *      9         �t�bhhK ��h��R�(KK��h�C@M   q   �  �        g      g  .     K     L        �t�bhhK ��h��R�(KK
��h�C(         T     �     1         �t�bhhK ��h��R�(KK��h�C  M           �t�bhhK ��h��R�(KK��h�CA   �   �        �t�bhhK ��h��R�(KK	��h�C$�      �   O                 �t�bhhK ��h��R�(KK��h�C�   �   �        �t�bhhK ��h��R�(KK��h�C�   N     E      �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK	��h�C$*            �  �   6        �t�bhhK ��h��R�(KK
��h�C(.   �     9   	     
   �         �t�bhhK ��h��R�(KK��h�C<7  �     .   ^     �  	             *         �t�bhhK ��h��R�(KK��h�C*   "       |         �t�bhhK ��h��R�(KK��h�C:   �       �        �t�bhhK ��h��R�(KK��h�C<i  �  �          �     /  �  "   W   f        �t�bhhK ��h��R�(KK��h�C<�  *         �  	   @       �     �        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C,!  u   �       i  "  I   `        �t�bhhK ��h��R�(KK��h�C �   u   #  *   $  %        �t�bhhK ��h��R�(KK��h�C4   &     Z  '  Z   (  U   )     *         �t�bhhK ��h��R�(KK��h�C8   *     Z  �   *      +  �     Z   ,        �t�bhhK ��h��R�(KK��h�C8   *   -  �  .     A    /     j  �        �t�bhhK ��h��R�(KK��h�C8N   1   �           0  �   9   1  I   2        �t�bhhK ��h��R�(KK��h�C<-   
   9   3  s  	   u   *   4  �     5  6        �t�bhhK ��h��R�(KK��h�C47     *   �   8  U         9     Z        �t�bhhK ��h��R�(KK��h�C<I   :  A  *   ;  |      h  I   �    <  |         �t�bhhK ��h��R�(KK��h�C *   �         I   P        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C    �   a      �      �t�bhhK ��h��R�(KK��h�C�      7     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cn     $      L      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C   *      Z   �        �t�bhhK ��h��R�(KK
��h�C(k  �     l     �               �t�bhhK ��h��R�(KK��h�C<   k     j  |   �     =  \   @   �     f         �t�bhhK ��h��R�(KK��h�Cm  �     �t�bhhK ��h��R�(KK��h�C>  C  �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�  ?                 �t�bhhK ��h��R�(KK��h�Cm  l     �t�bhhK ��h��R�(KK��h�C@  �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�CA  B     �t�bhhK ��h��R�(KK��h�Cd   *   C     D  E        B      F   8  ^  	   Q  	   R  S  	   T     F  �         �t�bhhK ��h��R�(KK��h�C,v      B   -   �   )      W   k         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�CG                 �t�bhhK ��h��R�(KK��h�CD   *      ^   �     p   �     �  �     $      L         �t�bhhK ��h��R�(KK��h�C8>   �     �   	   �  	   �  	   �      H        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�              �t�bhhK ��h��R�(KK	��h�C$�  I  J  �   �     $         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK��h�C         X        �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK
��h�C(�                 E      �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C0   *      ^   �      >   �     �         �t�bhhK ��h��R�(KK��h�CL           [  9  	   �  	   �   	   W  	   X     [  e         �t�bhhK ��h��R�(KK��h�C0a  "   9     e   Z     ^   >   k         �t�bhhK ��h��R�(KK	��h�C$           D   �   B        �t�bhhK ��h��R�(KK
��h�C(O  a  D   �     �      a        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�CK                 �t�bhhK ��h��R�(KK��h�C�       �t�bhhK ��h��R�(KK��h�C �    �           9      �t�bhhK ��h��R�(KK��h�CD�     9  	   �   	   �     0  \   1     ^   >   k         �t�bhhK ��h��R�(KK��h�C8                �  Z     r   �   2        �t�bhhK ��h��R�(KK��h�C�   �        �t�bhhK ��h��R�(KK��h�C�  Y                 �t�bhhK ��h��R�(KK��h�C8�  �  /                 �      �     �      �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CD   *      �  	   ^   �  	   �     W   �     >   �        �t�bhhK ��h��R�(KK��h�C8   �     B   �     �       �     �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C    
   L                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C    �   a      �      �t�bhhK ��h��R�(KK��h�C4   *      ^   M  v   B      N     �         �t�bhhK ��h��R�(KK��h�C,   F   O  P  �   N     �  �        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C Q     �                 �t�bhhK ��h��R�(KK
��h�C(6                 E      �     �t�bhhK ��h��R�(KK��h�CR                 �t�bhhK ��h��R�(KK��h�C0   n  S  o  �     	   �      �        �t�bhhK ��h��R�(KK��h�C8n     �            �      �     T  U        �t�bhhK ��h��R�(KK��h�CV  o        �t�bhhK ��h��R�(KK��h�CW  X                 �t�bhhK ��h��R�(KK��h�C4   *      �     Y     >   �     �         �t�bhhK ��h��R�(KK��h�C    Z     Z   �          �t�bhhK ��h��R�(KK��h�C     '     [        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C\                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK
��h�C(   ]        ^     Z           �t�bhhK ��h��R�(KK��h�C,   p  O   ,  �     _     `        �t�bhhK ��h��R�(KK��h�C0
      �  W   a  6      �  '   b        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C L     c                 �t�bhhK ��h��R�(KK
��h�C(             �   a      �         �t�bhhK ��h��R�(KK��h�C�      7     �t�bhhK ��h��R�(KK	��h�C$   *      ^   �     �        �t�bhhK ��h��R�(KK��h�C   *         �        �t�bhhK ��h��R�(KK��h�C,      
   �  7         �  �        �t�bhhK ��h��R�(KK��h�C_  �   *      �        �t�bhhK ��h��R�(KK��h�C          �      7        �t�bhhK ��h��R�(KK��h�Cd        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C e     �                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C   *      ^   �         �t�bhhK ��h��R�(KK��h�C0*   f  �  g     '      �   P  h        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C0�     �  ^  i                 E      �t�bhhK ��h��R�(KK��h�Cn     $      L      �t�bhhK ��h��R�(KK��h�CD   *      ^   �     p   �     �  �     $      L         �t�bhhK ��h��R�(KK��h�C8>   �     �   	   �  	   �  	   �      �        �t�bhhK ��h��R�(KK��h�C0   *      �     \  j     6  �        �t�bhhK ��h��R�(KK��h�C4q     �         �      �  �     _        �t�bhhK ��h��R�(KK
��h�C(   q     :   L   �     k        �t�bhhK ��h��R�(KK��h�C0v   �  .   -   l     �   �      �         �t�bhhK ��h��R�(KK��h�C,D   �        �   [  +     �         �t�bhhK ��h��R�(KK
��h�C(         n     $      L         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C +     *                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C c      *                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8   *      Z   >   �   	      F   Z             �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�Cm     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�      n           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C    �   a      �      �t�bhhK ��h��R�(KK��h�C�      7     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cn     $      L      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C   *      Z   �        �t�bhhK ��h��R�(KK
��h�C(k  �     l     �               �t�bhhK ��h��R�(KK��h�C<   k     j  |   �     =  \   @   �     f         �t�bhhK ��h��R�(KK��h�Cm  �     �t�bhhK ��h��R�(KK��h�C>  C  �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�  ?                 �t�bhhK ��h��R�(KK��h�Cm  l     �t�bhhK ��h��R�(KK��h�C@  �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�CA  B     �t�bhhK ��h��R�(KK��h�Cd   *   C     D  E        B      F   8  ^  	   Q  	   R  S  	   T     F  �         �t�bhhK ��h��R�(KK��h�C,v      B   -   �   )      W   k         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�CG                 �t�bhhK ��h��R�(KK��h�CD   *      ^   �     p   �     �  �     $      L         �t�bhhK ��h��R�(KK��h�C8>   �     �   	   �  	   �  	   �      H        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�              �t�bhhK ��h��R�(KK	��h�C$�  I  J  �   �     $         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK��h�C         X        �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C �                 E      �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C0   *      ^   �      >   �     �         �t�bhhK ��h��R�(KK��h�CL           [  9  	   �  	   �   	   W  	   X     [  e         �t�bhhK ��h��R�(KK��h�C0a  "   9     e   Z     ^   >   k         �t�bhhK ��h��R�(KK	��h�C$           D   �   B        �t�bhhK ��h��R�(KK
��h�C(O  a  D   �     �      a        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�CK                 �t�bhhK ��h��R�(KK��h�C�       �t�bhhK ��h��R�(KK��h�C �    �           9      �t�bhhK ��h��R�(KK��h�CD�     9  	   �   	   �     0  \   1     ^   >   k         �t�bhhK ��h��R�(KK��h�C8                �  Z     r   �   2        �t�be(hhK ��h��R�(KK��h�C�   �        �t�bhhK ��h��R�(KK��h�C�  Y                 �t�bhhK ��h��R�(KK��h�C8�  �  /                 �      �     �      �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CD   *      �  	   ^   �  	   �     W   �     >   �        �t�bhhK ��h��R�(KK��h�C8   �     B   �     �       �     �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C    
   L                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C    �   a      �      �t�bhhK ��h��R�(KK��h�C4   *      ^   M  v   B      N     �         �t�bhhK ��h��R�(KK��h�C,   F   O  P  �   N     �  �        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C Q     �                 �t�bhhK ��h��R�(KK
��h�C(6                 E      �     �t�bhhK ��h��R�(KK��h�CR                 �t�bhhK ��h��R�(KK��h�C0   n  S  o  �     	   �      �        �t�bhhK ��h��R�(KK��h�C8n     �            �      �     T  U        �t�bhhK ��h��R�(KK��h�CV  o        �t�bhhK ��h��R�(KK��h�CW  X                 �t�bhhK ��h��R�(KK��h�C4   *      �     Y     >   �     �         �t�bhhK ��h��R�(KK��h�C    Z     Z   �          �t�bhhK ��h��R�(KK��h�C     '     [        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C\                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK
��h�C(   ]        ^     Z           �t�bhhK ��h��R�(KK��h�C,   p  O   ,  �     _     `        �t�bhhK ��h��R�(KK��h�C0
      �  W   a  6      �  '   b        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C L     c                 �t�bhhK ��h��R�(KK
��h�C(             �   a      �         �t�bhhK ��h��R�(KK��h�C�      7     �t�bhhK ��h��R�(KK	��h�C$   *      ^   �     �        �t�bhhK ��h��R�(KK��h�C   *         �        �t�bhhK ��h��R�(KK��h�C,      
   �  7         �  �        �t�bhhK ��h��R�(KK��h�C_  �   *      �        �t�bhhK ��h��R�(KK��h�C          �      7        �t�bhhK ��h��R�(KK��h�Cd        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C e     �                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C   *      ^   �         �t�bhhK ��h��R�(KK��h�C0*   f  �  g     '      �   P  h        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C0�     �  ^  i                 E      �t�bhhK ��h��R�(KK��h�Cn     $      L      �t�bhhK ��h��R�(KK��h�CD   *      ^   �     p   �     �  �     $      L         �t�bhhK ��h��R�(KK��h�C8>   �     �   	   �  	   �  	   �      �        �t�bhhK ��h��R�(KK��h�C0   *      �     \  j     6  �        �t�bhhK ��h��R�(KK��h�C4q     �         �      �  �     _        �t�bhhK ��h��R�(KK
��h�C(   q     :   L   �     k        �t�bhhK ��h��R�(KK��h�C0v   �  .   -   l     �   �      �         �t�bhhK ��h��R�(KK��h�C,D   �        �   [  +     �         �t�bhhK ��h��R�(KK
��h�C(         n     $      L         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C +     *                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C c      *                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8   *      Z   >   �   	      F   Z             �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�Cm     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�      n           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C    �   a      �      �t�bhhK ��h��R�(KK��h�C�      7     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cn     $      L      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C   *      Z   �        �t�bhhK ��h��R�(KK
��h�C(k  �     l     �               �t�bhhK ��h��R�(KK��h�C<   k     j  |   �     =  \   @   �     f         �t�bhhK ��h��R�(KK��h�Cm  �     �t�bhhK ��h��R�(KK��h�C>  C  �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�  ?                 �t�bhhK ��h��R�(KK��h�Cm  l     �t�bhhK ��h��R�(KK��h�C@  �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�CA  B     �t�bhhK ��h��R�(KK��h�Cd   *   C     D  E        B      F   8  ^  	   Q  	   R  S  	   T     F  �         �t�bhhK ��h��R�(KK��h�C,v      B   -   �   )      W   k         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�CG                 �t�bhhK ��h��R�(KK��h�CD   *      ^   �     p   �     �  �     $      L         �t�bhhK ��h��R�(KK��h�C8>   �     �   	   �  	   �  	   �      H        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�              �t�bhhK ��h��R�(KK	��h�C$�  I  J  �   �     $         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK��h�C         X        �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C �                 E      �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C0   *      ^   �      >   �     �         �t�bhhK ��h��R�(KK��h�CL           [  9  	   �  	   �   	   W  	   X     [  e         �t�bhhK ��h��R�(KK��h�C0a  "   9     e   Z     ^   >   k         �t�bhhK ��h��R�(KK	��h�C$           D   �   B        �t�bhhK ��h��R�(KK
��h�C(O  a  D   �     �      a        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�CK                 �t�bhhK ��h��R�(KK��h�C�       �t�bhhK ��h��R�(KK��h�C �    �           9      �t�bhhK ��h��R�(KK��h�CD�     9  	   �   	   �     0  \   1     ^   >   k         �t�bhhK ��h��R�(KK��h�C8                �  Z     r   �   2        �t�bhhK ��h��R�(KK��h�C�   �        �t�bhhK ��h��R�(KK��h�C�  Y                 �t�bhhK ��h��R�(KK��h�C8�  �  /                 �      �     �      �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CD   *      �  	   ^   �  	   �     W   �     >   �        �t�bhhK ��h��R�(KK��h�C8   �     B   �     �       �     �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C    
   L                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C    �   a      �      �t�bhhK ��h��R�(KK��h�C4   *      ^   M  v   B      N     �         �t�bhhK ��h��R�(KK��h�C,   F   O  P  �   N     �  �        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C Q     �                 �t�bhhK ��h��R�(KK
��h�C(6                 E      �     �t�bhhK ��h��R�(KK��h�CR                 �t�bhhK ��h��R�(KK��h�C0   n  S  o  �     	   �      �        �t�bhhK ��h��R�(KK��h�C8n     �            �      �     T  U        �t�bhhK ��h��R�(KK��h�CV  o        �t�bhhK ��h��R�(KK��h�CW  X                 �t�bhhK ��h��R�(KK��h�C4   *      �     Y     >   �     �         �t�bhhK ��h��R�(KK��h�C    Z     Z   �          �t�bhhK ��h��R�(KK��h�C     '     [        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C\                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK
��h�C(   ]        ^     Z           �t�bhhK ��h��R�(KK��h�C,   p  O   ,  �     _     `        �t�bhhK ��h��R�(KK��h�C0
      �  W   a  6      �  '   b        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C L     c                 �t�bhhK ��h��R�(KK
��h�C(             �   a      �         �t�bhhK ��h��R�(KK��h�C�      7     �t�bhhK ��h��R�(KK	��h�C$   *      ^   �     �        �t�bhhK ��h��R�(KK��h�C   *         �        �t�bhhK ��h��R�(KK��h�C,      
   �  7         �  �        �t�bhhK ��h��R�(KK��h�C_  �   *      �        �t�bhhK ��h��R�(KK��h�C          �      7        �t�bhhK ��h��R�(KK��h�Cd        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C e     �                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C   *      ^   �         �t�bhhK ��h��R�(KK��h�C0*   f  �  g     '      �   P  h        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C0�     �  ^  i                 E      �t�bhhK ��h��R�(KK��h�Cn     $      L      �t�bhhK ��h��R�(KK��h�CD   *      ^   �     p   �     �  �     $      L         �t�bhhK ��h��R�(KK��h�C8>   �     �   	   �  	   �  	   �      �        �t�bhhK ��h��R�(KK��h�C0   *      �     \  j     6  �        �t�bhhK ��h��R�(KK��h�C4q     �         �      �  �     _        �t�bhhK ��h��R�(KK
��h�C(   q     :   L   �     k        �t�bhhK ��h��R�(KK��h�C0v   �  .   -   l     �   �      �         �t�bhhK ��h��R�(KK��h�C,D   �        �   [  +     �         �t�bhhK ��h��R�(KK
��h�C(         n     $      L         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C +     *                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C c      *                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8   *      Z   >   �   	      F   Z             �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�Cm     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�      n           �t�bhhK ��h��R�(KK��h�C,      �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�Cl   �     m      �      �t�bhhK ��h��R�(KK��h�Cn      _   ,      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C0�   �   �   
   .      �   
      M        �t�bhhK ��h��R�(KK��h�C0M   �         5  6  	   7     8        �t�bhhK ��h��R�(KK��h�C,�   4   �   
   .   4         M        �t�bhhK ��h��R�(KK��h�C         �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C`0      �      )  }  *     x   �   �   
         J   �  5   +           �        �t�bhhK ��h��R�(KK��h�C@o        F   �     l   	   b     �  ,       �         �t�bhhK ��h��R�(KK��h�Cx      -   =   0      �   
      "   ,      J   `  G   	   �      
      p  �         q  r     3        �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�Cs  �      �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C(      <      D     �t�bhhK ��h��R�(KK��h�C�   d  E  �   �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C 0                       �t�bhhK ��h��R�(KK��h�CD�     �   G      1      �  t     "      u     C         �t�bhhK ��h��R�(KK��h�C r  �           9         �t�bhhK ��h��R�(KK��h�C,v  p   /   +      V      w          �t�bhhK ��h��R�(KK��h�C4�      }   �   ]      �     <      x        �t�bhhK ��h��R�(KK��h�C 9     �   G      1         �t�bhhK ��h��R�(KK��h�C@�     �                  E      �      �      �     �t�bhhK ��h��R�(KK��h�C,      �     �t�bhhK ��h��R�(KK��h�CD
      "   ,      �     �  	   6      w   �      y        �t�bhhK ��h��R�(KK��h�C         ,      {      �t�bhhK ��h��R�(KK��h�C�  z                 �t�bhhK ��h��R�(KK��h�Cl
           	   {     �     1        z  |        >  
   s  +      c      :  �        �t�bhhK ��h��R�(KK��h�Cr  �      9         �t�bhhK ��h��R�(KK��h�C�      }  1  �     �t�bhhK ��h��R�(KK��h�C(   ~     �t�bhhK ��h��R�(KK��h�C<  =        �t�bhhK ��h��R�(KK��h�C �     >                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C<
        b     '   �   	   �        d   �        �t�bhhK ��h��R�(KK��h�C       �         "        �t�bhhK ��h��R�(KK��h�C<      -           �     �   &      *   E        �t�bhhK ��h��R�(KK��h�C*   E     �t�bhhK ��h��R�(KK��h�C  1     �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C�                  �t�bhhK ��h��R�(KK��h�C'  \                 �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�C8
      5   s  +   	         =   �   ~           �t�bhhK ��h��R�(KK��h�C�  �  e     �t�bhhK ��h��R�(KK��h�C(   @     �t�bhhK ��h��R�(KK	��h�C$         5           h      �t�bhhK ��h��R�(KK��h�CF  ~           �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�CL�     �     x   /   
      "   �  b     �     l   �   K        �t�bhhK ��h��R�(KK��h�C0�  �      �  �      /        $         �t�bhhK ��h��R�(KK��h�CP      �   �     q   �   �         5   4     r   �  N      �        �t�bhhK ��h��R�(KK��h�Cx      D   �  �   b         L  
   J   �  	   �     �  y      �     �     F  y      /     O        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C2     t     �t�bhhK ��h��R�(KK��h�C�  �  �     �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�C         l      �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK
��h�C(+      �     �                 �t�bhhK ��h��R�(KK��h�Cp�  u     �  u                x   G  	      "   b  �  �     l      q      �     _        �t�bhhK ��h��R�(KK��h�C�  :  e     �t�bhhK ��h��R�(KK��h�C(      <      a     �t�bhhK ��h��R�(KK��h�C+      B           �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK��h�C<
      "   ,      r   m      �         =   �         �t�bhhK ��h��R�(KK��h�C,�        �  N          $         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cc                 �t�bhhK ��h��R�(KK��h�C4i  T   c      �     �     )               �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C8c      C   �     M        �                 �t�bhhK ��h��R�(KK��h�CD�  �  %  �  T   v     �  U   <  T     )               �t�bhhK ��h��R�(KK��h�CL             �t�bhhK ��h��R�(KK	��h�C$v     �  U   <  �           �t�bhhK ��h��R�(KK��h�C,D   �  Y  T   �     ,      b        �t�bhhK ��h��R�(KK��h�C�  �                 �t�bhhK ��h��R�(KK	��h�C$         ,      m      �      �t�bhhK ��h��R�(KK��h�Cn      _   ,      �t�bhhK ��h��R�(KK��h�CH?     J  p   f      �      �  a     �     $   ?   �         �t�bhhK ��h��R�(KK
��h�C(   *      ^   Q  �     �         �t�bhhK ��h��R�(KK��h�Cj  b     c      �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cj  �                  �t�bhhK ��h��R�(KK��h�C8   ,      �  $      �   x      F   j  0        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK
��h�C(   
   �     �                 �t�bhhK ��h��R�(KK��h�CP
      5   f      �   :  n   C  �  	         �      }   d   �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cc                 �t�bhhK ��h��R�(KK��h�C8i  p   f      �     �   w  �     A  �        �t�bhhK ��h��R�(KK��h�CL     >   k         �t�bhhK ��h��R�(KK��h�C (   �     E   	            �t�bhhK ��h��R�(KK��h�C@L      L  
   �  ,      ?     &   �   @     �        �t�bhhK ��h��R�(KK��h�C0.      -   W     v   B      @   +         �t�bhhK ��h��R�(KK ��h�C�        �  r     �  I      @   +      x  -  
   �  "   ,      F      &   `  a  	   �  	   �     �        �t�bhhK ��h��R�(KK��h�C B      �      �   -        �t�bhhK ��h��R�(KK	��h�C$     -     R     �        �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C -  �   +      *           �t�bhhK ��h��R�(KK��h�CX
   &   L   4           v  �   M  	      �  =   �   	  
  !  _   (        �t�bhhK ��h��R�(KK��h�C"        �        �t�bhhK ��h��R�(KK��h�C:   _   (     �t�bhhK ��h��R�(KK��h�C(      <      C     �t�bhhK ��h��R�(KK��h�C�   	  
        �t�bhhK ��h��R�(KK��h�C:   _   #     �t�bhhK ��h��R�(KK��h�C          n      _   ,      �t�bhhK ��h��R�(KK��h�C<
      "   Q  ,         �   
   f   d   t  %        �t�bhhK ��h��R�(KK��h�Cd
         J   �  4   "     �     �     &   �  |  �        g   [   �  d           �t�bhhK ��h��R�(KK��h�C0   
                    E      s     �t�bhhK ��h��R�(KK��h�C8
      "   ,      �  	   =   �  �     �        �t�bhhK ��h��R�(KK��h�Cq      �        �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C �                      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CT     �     �  T   �   p  +      o      ,      &   `  a     �        �t�bhhK ��h��R�(KK��h�C}  �        �t�bhhK ��h��R�(KK��h�C]      �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C    
   4                 �t�bhhK ��h��R�(KK��h�C@L      �  r     �     �      @   +      x  -        �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C -  �   +      *           �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C,�  x      :   �           	        �t�bhhK ��h��R�(KK��h�C4      g   �     F      �         2         �t�bhhK ��h��R�(KK��h�C�             �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK��h�C    *      �     �        �t�bhhK ��h��R�(KK
��h�C(      c     '                  �t�bhhK ��h��R�(KK��h�CHv      :   �  R     A     z        4         �           �t�bhhK ��h��R�(KK��h�CA   �        �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK��h�Cd
      �  S  D        5   V         =   0      �      *   	   ]      <      D        �t�bhhK ��h��R�(KK��h�C         �     �t�bhhK ��h��R�(KK��h�C,      �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�Cl   �     m      �      �t�bhhK ��h��R�(KK��h�Cn      _   ,      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C0�   �   �   
   .      �   
      M        �t�bhhK ��h��R�(KK��h�C0M   �         5  6  	   7     8        �t�bhhK ��h��R�(KK��h�C,�   4   �   
   .   4         M        �t�bhhK ��h��R�(KK��h�C         �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C`0      �      )  }  *     x   �   �   
         J   �  5   +           �        �t�bhhK ��h��R�(KK��h�C@o        F   �     l   	   b     �  ,       �         �t�bhhK ��h��R�(KK��h�Cx      -   =   0      �   
      "   ,      J   `  G   	   �      
      p  �         q  r     3        �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�Cs  �      �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C(      <      D     �t�bhhK ��h��R�(KK��h�C�   d  E  �   �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C 0                       �t�bhhK ��h��R�(KK��h�CD�     �   G      1      �  t     "      u     C         �t�bhhK ��h��R�(KK��h�C r  �           9         �t�bhhK ��h��R�(KK��h�C,v  p   /   +      V      w          �t�bhhK ��h��R�(KK��h�C4�      }   �   ]      �     <      x        �t�bhhK ��h��R�(KK��h�C 9     �   G      1         �t�bhhK ��h��R�(KK��h�C@�     �                  E      �      �      �     �t�bhhK ��h��R�(KK��h�C,      �     �t�bhhK ��h��R�(KK��h�CD
      "   ,      �     �  	   6      w   �      y        �t�bhhK ��h��R�(KK��h�C         ,      {      �t�bhhK ��h��R�(KK��h�C�  z                 �t�bhhK ��h��R�(KK��h�Cl
           	   {     �     1        z  |        >  
   s  +      c      :  �        �t�bhhK ��h��R�(KK��h�Cr  �      9         �t�bhhK ��h��R�(KK��h�C�      }  1  �     �t�bhhK ��h��R�(KK��h�C(   ~     �t�bhhK ��h��R�(KK��h�C<  =        �t�bhhK ��h��R�(KK��h�C �     >                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C<
        b     '   �   	   �        d   �        �t�bhhK ��h��R�(KK��h�C       �         "        �t�bhhK ��h��R�(KK��h�C<      -           �     �   &      *   E        �t�bhhK ��h��R�(KK��h�C*   E     �t�bhhK ��h��R�(KK��h�C  1     �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C�                  �t�bhhK ��h��R�(KK��h�C'  \                 �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�C8
      5   s  +   	         =   �   ~           �t�bhhK ��h��R�(KK��h�C�  �  e     �t�bhhK ��h��R�(KK��h�C(   @     �t�bhhK ��h��R�(KK	��h�C$         5           h      �t�bhhK ��h��R�(KK��h�CF  ~           �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�CL�     �     x   /   
      "   �  b     �     l   �   K        �t�bhhK ��h��R�(KK��h�C0�  �      �  �      /        $         �t�bhhK ��h��R�(KK��h�CP      �   �     q   �   �         5   4     r   �  N      �        �t�bhhK ��h��R�(KK��h�Cx      D   �  �   b         L  
   J   �  	   �     �  y      �     �     F  y      /     O        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C2     t     �t�bhhK ��h��R�(KK��h�C�  �  �     �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�C         l      �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK
��h�C(+      �     �                 �t�bhhK ��h��R�(KK��h�Cp�  u     �  u                x   G  	      "   b  �  �     l      q      �     _        �t�bhhK ��h��R�(KK��h�C�  :  e     �t�bhhK ��h��R�(KK��h�C(      <      a     �t�bhhK ��h��R�(KK��h�C+      B           �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK��h�C<
      "   ,      r   m      �         =   �         �t�bhhK ��h��R�(KK��h�C,�        �  N          $         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cc                 �t�bhhK ��h��R�(KK��h�C4i  T   c      �     �     )               �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C8c      C   �     M        �                 �t�bhhK ��h��R�(KK��h�CD�  �  %  �  T   v     �  U   <  T     )               �t�bhhK ��h��R�(KK��h�CL             �t�bhhK ��h��R�(KK	��h�C$v     �  U   <  �           �t�bhhK ��h��R�(KK��h�C,D   �  Y  T   �     ,      b        �t�bhhK ��h��R�(KK��h�C�  �                 �t�bhhK ��h��R�(KK	��h�C$         ,      m      �      �t�bhhK ��h��R�(KK��h�Cn      _   ,      �t�bhhK ��h��R�(KK��h�CH?     J  p   f      �      �  a     �     $   ?   �         �t�bhhK ��h��R�(KK
��h�C(   *      ^   Q  �     �         �t�bhhK ��h��R�(KK��h�Cj  b     c      �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cj  �                  �t�bhhK ��h��R�(KK��h�C8   ,      �  $      �   x      F   j  0        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK
��h�C(   
   �     �                 �t�bhhK ��h��R�(KK��h�CP
      5   f      �   :  n   C  �  	         �      }   d   �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cc                 �t�bhhK ��h��R�(KK��h�C8i  p   f      �     �   w  �     A  �        �t�bhhK ��h��R�(KK��h�CL     >   k         �t�bhhK ��h��R�(KK��h�C (   �     E   	            �t�bhhK ��h��R�(KK��h�C@L      L  
   �  ,      ?     &   �   @     �        �t�bhhK ��h��R�(KK��h�C0.      -   W     v   B      @   +         �t�bhhK ��h��R�(KK ��h�C�        �  r     �  I      @   +      x  -  
   �  "   ,      F      &   `  a  	   �  	   �     �        �t�bhhK ��h��R�(KK��h�C B      �      �   -        �t�bhhK ��h��R�(KK	��h�C$     -     R     �        �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C -  �   +      *           �t�bhhK ��h��R�(KK��h�CX
   &   L   4           v  �   M  	      �  =   �   	  
  !  _   (        �t�bhhK ��h��R�(KK��h�C"        �        �t�bhhK ��h��R�(KK��h�C:   _   (     �t�bhhK ��h��R�(KK��h�C(      <      C     �t�bhhK ��h��R�(KK��h�C�   	  
        �t�bhhK ��h��R�(KK��h�C:   _   #     �t�bhhK ��h��R�(KK��h�C          n      _   ,      �t�bhhK ��h��R�(KK��h�C<
      "   Q  ,         �   
   f   d   t  %        �t�bhhK ��h��R�(KK��h�Cd
         J   �  4   "     �     �     &   �  |  �        g   [   �  d           �t�bhhK ��h��R�(KK��h�C0   
                    E      s     �t�bhhK ��h��R�(KK��h�C8
      "   ,      �  	   =   �  �     �        �t�bhhK ��h��R�(KK��h�Cq      �        �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C �                      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CT     �     �  T   �   p  +      o      ,      &   `  a     �        �t�bhhK ��h��R�(KK��h�C}  �        �t�bhhK ��h��R�(KK��h�C]      �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C    
   4                 �t�bhhK ��h��R�(KK��h�C@L      �  r     �     �      @   +      x  -        �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C -  �   +      *           �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C,�  x      :   �           	        �t�bhhK ��h��R�(KK��h�C4      g   �     F      �         2         �t�bhhK ��h��R�(KK��h�C�             �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C    *      �     �        �t�bhhK ��h��R�(KK
��h�C(      c     '                  �t�bhhK ��h��R�(KK��h�CHv      :   �  R     A     z        4         �           �t�bhhK ��h��R�(KK��h�CA   �        �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK��h�Cd
      �  S  D        5   V         =   0      �      *   	   ]      <      D        �t�bhhK ��h��R�(KK��h�C         �     �t�bhhK ��h��R�(KK��h�C,      �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�Cl   �     m      �      �t�bhhK ��h��R�(KK��h�Cn      _   ,      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C0�   �   �   
   .      �   
      M        �t�bhhK ��h��R�(KK��h�C0M   �         5  6  	   7     8        �t�bhhK ��h��R�(KK��h�C,�   4   �   
   .   4         M        �t�bhhK ��h��R�(KK��h�C         �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�C`0      �      )  }  *     x   �   �   
         J   �  5   +           �        �t�bhhK ��h��R�(KK��h�C@o        F   �     l   	   b     �  ,       �         �t�bhhK ��h��R�(KK��h�Cx      -   =   0      �   
      "   ,      J   `  G   	   �      
      p  �         q  r     3        �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�Cs  �      �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C(      <      D     �t�bhhK ��h��R�(KK��h�C�   d  E  �   �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C 0                       �t�bhhK ��h��R�(KK��h�CD�     �   G      1      �  t     "      u     C         �t�bhhK ��h��R�(KK��h�C r  �           9         �t�bhhK ��h��R�(KK��h�C,v  p   /   +      V      w          �t�bhhK ��h��R�(KK��h�C4�      }   �   ]      �     <      x        �t�bhhK ��h��R�(KK��h�C 9     �   G      1         �t�bhhK ��h��R�(KK��h�C@�     �                  E      �      �      �     �t�bhhK ��h��R�(KK��h�C,      �     �t�bhhK ��h��R�(KK��h�CD
      "   ,      �     �  	   6      w   �      y        �t�bhhK ��h��R�(KK��h�C         ,      {      �t�bhhK ��h��R�(KK��h�C�  z                 �t�bhhK ��h��R�(KK��h�Cl
           	   {     �     1        z  |        >  
   s  +      c      :  �        �t�bhhK ��h��R�(KK��h�Cr  �      9         �t�bhhK ��h��R�(KK��h�C�      }  1  �     �t�bhhK ��h��R�(KK��h�C(   ~     �t�bhhK ��h��R�(KK��h�C<  =        �t�bhhK ��h��R�(KK��h�C �     >                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C<
        b     '   �   	   �        d   �        �t�bhhK ��h��R�(KK��h�C       �         "        �t�bhhK ��h��R�(KK��h�C<      -           �     �   &      *   E        �t�bhhK ��h��R�(KK��h�C*   E     �t�bhhK ��h��R�(KK��h�C  1     �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C�                  �t�bhhK ��h��R�(KK��h�C'  \                 �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�C8
      5   s  +   	         =   �   ~           �t�bhhK ��h��R�(KK��h�C�  �  e     �t�bhhK ��h��R�(KK��h�C(   @     �t�bhhK ��h��R�(KK	��h�C$         5           h      �t�bhhK ��h��R�(KK��h�CF  ~           �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�CL�     �     x   /   
      "   �  b     �     l   �   K        �t�bhhK ��h��R�(KK��h�C0�  �      �  �      /        $         �t�bhhK ��h��R�(KK��h�CP      �   �     q   �   �         5   4     r   �  N      �        �t�bhhK ��h��R�(KK��h�Cx      D   �  �   b         L  
   J   �  	   �     �  y      �     �     F  y      /     O        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C2     t     �t�bhhK ��h��R�(KK��h�C�  �  �     �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�C         l      �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK
��h�C(+      �     �                 �t�bhhK ��h��R�(KK��h�Cp�  u     �  u                x   G  	      "   b  �  �     l      q      �     _        �t�bhhK ��h��R�(KK��h�C�  :  e     �t�bhhK ��h��R�(KK��h�C(      <      a     �t�bhhK ��h��R�(KK��h�C+      B           �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK��h�C<
      "   ,      r   m      �         =   �         �t�bhhK ��h��R�(KK��h�C,�        �  N          $         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cc                 �t�bhhK ��h��R�(KK��h�C4i  T   c      �     �     )               �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C8c      C   �     M        �                 �t�bhhK ��h��R�(KK��h�CD�  �  %  �  T   v     �  U   <  T     )               �t�bhhK ��h��R�(KK��h�CL             �t�bhhK ��h��R�(KK	��h�C$v     �  U   <  �           �t�bhhK ��h��R�(KK��h�C,D   �  Y  T   �     ,      b        �t�bhhK ��h��R�(KK��h�C�  �                 �t�bhhK ��h��R�(KK	��h�C$         ,      m      �      �t�bhhK ��h��R�(KK��h�Cn      _   ,      �t�bhhK ��h��R�(KK��h�CH?     J  p   f      �      �  a     �     $   ?   �         �t�bhhK ��h��R�(KK
��h�C(   *      ^   Q  �     �         �t�bhhK ��h��R�(KK��h�Cj  b     c      �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cj  �                  �t�bhhK ��h��R�(KK��h�C8   ,      �  $      �   x      F   j  0        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK
��h�C(   
   �     �                 �t�bhhK ��h��R�(KK��h�CP
      5   f      �   :  n   C  �  	         �      }   d   �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cc                 �t�bhhK ��h��R�(KK��h�C8i  p   f      �     �   w  �     A  �        �t�bhhK ��h��R�(KK��h�CL     >   k         �t�bhhK ��h��R�(KK��h�C (   �     E   	            �t�bhhK ��h��R�(KK��h�C@L      L  
   �  ,      ?     &   �   @     �        �t�bhhK ��h��R�(KK��h�C0.      -   W     v   B      @   +         �t�bhhK ��h��R�(KK ��h�C�        �  r     �  I      @   +      x  -  
   �  "   ,      F      &   `  a  	   �  	   �     �        �t�bhhK ��h��R�(KK��h�C B      �      �   -        �t�bhhK ��h��R�(KK	��h�C$     -     R     �        �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C -  �   +      *           �t�bhhK ��h��R�(KK��h�CX
   &   L   4           v  �   M  	      �  =   �   	  
  !  _   (        �t�bhhK ��h��R�(KK��h�C"        �        �t�bhhK ��h��R�(KK��h�C:   _   (     �t�bhhK ��h��R�(KK��h�C(      <      C     �t�bhhK ��h��R�(KK��h�C�   	  
        �t�bhhK ��h��R�(KK��h�C:   _   #     �t�bhhK ��h��R�(KK��h�C          n      _   ,      �t�bhhK ��h��R�(KK��h�C<
      "   Q  ,         �   
   f   d   t  %        �t�bhhK ��h��R�(KK��h�Cd
         J   �  4   "     �     �     &   �  |  �        g   [   �  d           �t�bhhK ��h��R�(KK��h�C0   
                    E      s     �t�bhhK ��h��R�(KK��h�C8
      "   ,      �  	   =   �  �     �        �t�bhhK ��h��R�(KK��h�Cq      �        �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C �                      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CT     �     �  T   �   p  +      o      ,      &   `  a     �        �t�bhhK ��h��R�(KK��h�C}  �        �t�bhhK ��h��R�(KK��h�C]      �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C    
   4                 �t�bhhK ��h��R�(KK��h�C@L      �  r     �     �      @   +      x  -        �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C -  �   +      *           �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C,�  x      :   �           	        �t�bhhK ��h��R�(KK��h�C4      g   �     F      �         2         �t�bhhK ��h��R�(KK��h�C�             �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C    *      �     �        �t�bhhK ��h��R�(KK
��h�C(      c     '                  �t�bhhK ��h��R�(KK��h�CHv      :   �  R     A     z        4         �           �t�bhhK ��h��R�(KK��h�CA   �        �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK��h�Cd
      �  S  D        5   V         =   0      �      *   	   ]      <      D        �t�bhhK ��h��R�(KK��h�C         �     �t�bhhK ��h��R�(KK��h�Cm      �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C   �      �t�bhhK ��h��R�(KK��h�Co      $         �     �t�bhhK ��h��R�(KK��h�C,      K     �t�bhhK ��h��R�(KK��h�Cm      �t�bhhK ��h��R�(KK��h�C8�  �  6      d  $  g                    �t�bhhK ��h��R�(KK	��h�C$e  �     �                 �t�bhhK ��h��R�(KK��h�C,      $  g     ,  �     a        �t�bhhK ��h��R�(KK��h�C�      �  	   *   �     �t�bhhK ��h��R�(KK��h�C   :     �t�bhhK ��h��R�(KK��h�C(         �t�bhhK ��h��R�(KK��h�C         m         �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK
��h�C(  
   �     O  p  �           �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C8d     e     �   �   g     �   ~   f  �        �t�bhhK ��h��R�(KK��h�C<      D   g   b   g  	   �   J   E     F  G        �t�bhhK ��h��R�(KK��h�CL        �   `      h  �  �     	   i     M                �t�bhhK ��h��R�(KK��h�C(         �t�bhhK ��h��R�(KK��h�C         b         �t�bhhK ��h��R�(KK��h�CF  ~   h        �t�bhhK ��h��R�(KK��h�C�            �t�bhhK ��h��R�(KK��h�C$      b      �t�bhhK ��h��R�(KK��h�CX
      "   $   ?   r  I      �      j  /   	   w   �      �      �           �t�bhhK ��h��R�(KK��h�C0   �         �  A  �     :           �t�bhhK ��h��R�(KK	��h�C$   �         *   Q   2         �t�bhhK ��h��R�(KK��h�CP
      1  b         D   w   �      �             2     t        �t�bhhK ��h��R�(KK��h�C,   �        �        �           �t�bhhK ��h��R�(KK��h�C8�  6      '   k  
   �  �   	   �     �        �t�bhhK ��h��R�(KK��h�C�  �  8        �t�bhhK ��h��R�(KK
��h�C(P     �        *   Q   2         �t�bhhK ��h��R�(KK��h�CT*      "         v   B      �   
   f      �   w  k  N         a         �t�bhhK ��h��R�(KK��h�C(         �t�bhhK ��h��R�(KK��h�C          $      b         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cb                     �t�bhhK ��h��R�(KK��h�Co      $      �t�bhhK ��h��R�(KK��h�C@   
   �      $      *         j   �   P     *         �t�bhhK ��h��R�(KK��h�C  o      $      �t�bhhK ��h��R�(KK��h�C0         z                 o         �t�bhhK ��h��R�(KK��h�CP.   �             :     �   �     o                           �t�bhhK ��h��R�(KK
��h�C(   O   �          �   ]         �t�bhhK ��h��R�(KK	��h�C$   7   �     *   Q   2         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CD
      5           M  	         =   #  �     i        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C$  �        �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�Co     �t�bhhK ��h��R�(KK��h�Cp
   A  }  $      ?      I   	      �   �  @   o       �     N          �  z      �         �t�bhhK ��h��R�(KK��h�C<
      "   �      h        i   
   .   d           �t�bhhK ��h��R�(KK��h�C8           `      �        &              �t�bhhK ��h��R�(KK��h�C       D   �   2          �t�bhhK ��h��R�(KK��h�CH*      �  '        :        �  '   ?     $      �         �t�bhhK ��h��R�(KK��h�CPB      i   
      
      �  �   �   
   A     $   ?   �      �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK
��h�C(o      $                        �t�bhhK ��h��R�(KK��h�C    
   �                 �t�b��K      hhK ��h��R�(KK	��h�C$9  �      �                 �t�bhhK ��h��R�(KK��h�C �                        �t�bhhK ��h��R�(KK��h�C,     �     �t�bhhK ��h��R�(KK��h�Ch*      �   [  +     :   �     �  $      �      .         F   ,  	   �   �      �        �t�bhhK ��h��R�(KK��h�C,         V      o      $      �      �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C,                 �t�bhhK ��h��R�(KK��h�C,      K     �t�bhhK ��h��R�(KK!��h�C�   j   �   &       *   7        
   �        y  /      *          @   +      n      _   ,      ,      K        �t�bhhK ��h��R�(KK��h�Ct   7     
   n      _   ,   D      j   �   '     _   ,      �  7   F  +   N   $      L   "   ,   h      �t�bhhK ��h��R�(KK��h�Ch   j   �   �     m      �        
   �        y  /          @   +      ,      b        �t�bhhK ��h��R�(KK��h�Cm      �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C   �      �t�bhhK ��h��R�(KK��h�Co      $         �     �t�bhhK ��h��R�(KK��h�C,      K     �t�bhhK ��h��R�(KK��h�Cm      �t�bhhK ��h��R�(KK��h�C8�  �  6      d  $  g                    �t�bhhK ��h��R�(KK	��h�C$e  �     �                 �t�bhhK ��h��R�(KK��h�C,      $  g     ,  �     a        �t�bhhK ��h��R�(KK��h�C�      �  	   *   �     �t�bhhK ��h��R�(KK��h�C   :     �t�bhhK ��h��R�(KK��h�C(         �t�bhhK ��h��R�(KK��h�C         m         �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK
��h�C(  
   �     O  p  �           �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C8d     e     �   �   g     �   ~   f  �        �t�bhhK ��h��R�(KK��h�C<      D   g   b   g  	   �   J   E     F  G        �t�bhhK ��h��R�(KK��h�CL        �   `      h  �  �     	   i     M                �t�bhhK ��h��R�(KK��h�C(         �t�bhhK ��h��R�(KK��h�C         b         �t�bhhK ��h��R�(KK��h�CF  ~   h        �t�bhhK ��h��R�(KK��h�C�            �t�bhhK ��h��R�(KK��h�C$      b      �t�bhhK ��h��R�(KK��h�CX
      "   $   ?   r  I      �      j  /   	   w   �      �      �           �t�bhhK ��h��R�(KK��h�C0   �         �  A  �     :           �t�bhhK ��h��R�(KK	��h�C$   �         *   Q   2         �t�bhhK ��h��R�(KK��h�CP
      1  b         D   w   �      �             2     t        �t�bhhK ��h��R�(KK��h�C,   �        �        �           �t�bhhK ��h��R�(KK��h�C8�  6      '   k  
   �  �   	   �     �        �t�bhhK ��h��R�(KK��h�C�  �  8        �t�bhhK ��h��R�(KK
��h�C(P     �        *   Q   2         �t�bhhK ��h��R�(KK��h�CT*      "         v   B      �   
   f      �   w  k  N         a         �t�bhhK ��h��R�(KK��h�C(         �t�bhhK ��h��R�(KK��h�C          $      b         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cb                     �t�bhhK ��h��R�(KK��h�Co      $      �t�bhhK ��h��R�(KK��h�C@   
   �      $      *         j   �   P     *         �t�bhhK ��h��R�(KK��h�C  o      $      �t�bhhK ��h��R�(KK��h�C0         z                 o         �t�bhhK ��h��R�(KK��h�CP.   �             :     �   �     o                           �t�bhhK ��h��R�(KK
��h�C(   O   �          �   ]         �t�bhhK ��h��R�(KK	��h�C$   7   �     *   Q   2         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CD
      5           M  	         =   #  �     i        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C$  �        �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�Co     �t�bhhK ��h��R�(KK��h�Cp
   A  }  $      ?      I   	      �   �  @   o       �     N          �  z      �         �t�bhhK ��h��R�(KK��h�C<
      "   �      h        i   
   .   d           �t�bhhK ��h��R�(KK��h�C8           `      �        &              �t�bhhK ��h��R�(KK��h�C       D   �   2          �t�bhhK ��h��R�(KK��h�CH*      �  '        :        �  '   ?     $      �         �t�bhhK ��h��R�(KK��h�CPB      i   
      
      �  �   �   
   A     $   ?   �      �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK
��h�C(o      $                        �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK	��h�C$9  �      �                 �t�bhhK ��h��R�(KK��h�C �                        �t�bhhK ��h��R�(KK��h�C,     �     �t�bhhK ��h��R�(KK��h�Ch*      �   [  +     :   �     �  $      �      .         F   ,  	   �   �      �        �t�bhhK ��h��R�(KK��h�C,         V      o      $      �      �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C,                 �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK
��h�C(q     �   �      :   �  �        �t�bhhK ��h��R�(KK��h�C8�     q     *   �   ;   	      F     ;         �t�bhhK ��h��R�(KK��h�CL
      �   �        
   ;      �         =   ;     �           �t�bhhK ��h��R�(KK��h�C(      <            �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK
��h�C(N      �   �   
      N     �      �t�bhhK ��h��R�(KK��h�C|
      �   �   
      �   	   /     �  N  �  i      �  6   �  �  �  	         �  �      V      |        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�CV      �           �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C,      K     �t�bhhK ��h��R�(KK!��h�C�   j   �   &       *   7        
   �        y  /      *          @   +      n      _   ,      ,      K        �t�bhhK ��h��R�(KK��h�Ct   7     
   n      _   ,   D      j   �   '     _   ,      �  7   F  +   N   $      L   "   ,   h      �t�bhhK ��h��R�(KK��h�Ch   j   �   �     m      �        
   �        y  /          @   +      ,      b        �t�bhhK ��h��R�(KK��h�Cm      �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C   �      �t�bhhK ��h��R�(KK��h�Co      $         �     �t�bhhK ��h��R�(KK��h�C,      K     �t�bhhK ��h��R�(KK��h�Cm      �t�bhhK ��h��R�(KK��h�C8�  �  6      d  $  g                    �t�bhhK ��h��R�(KK	��h�C$e  �     �                 �t�bhhK ��h��R�(KK��h�C,      $  g     ,  �     a        �t�bhhK ��h��R�(KK��h�C�      �  	   *   �     �t�bhhK ��h��R�(KK��h�C   :     �t�bhhK ��h��R�(KK��h�C(         �t�bhhK ��h��R�(KK��h�C         m         �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK
��h�C(  
   �     O  p  �           �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C8d     e     �   �   g     �   ~   f  �        �t�bhhK ��h��R�(KK��h�C<      D   g   b   g  	   �   J   E     F  G        �t�bhhK ��h��R�(KK��h�CL        �   `      h  �  �     	   i     M                �t�bhhK ��h��R�(KK��h�C(         �t�bhhK ��h��R�(KK��h�C         b         �t�bhhK ��h��R�(KK��h�CF  ~   h        �t�bhhK ��h��R�(KK��h�C�            �t�bhhK ��h��R�(KK��h�C$      b      �t�bhhK ��h��R�(KK��h�CX
      "   $   ?   r  I      �      j  /   	   w   �      �      �           �t�bhhK ��h��R�(KK��h�C0   �         �  A  �     :           �t�bhhK ��h��R�(KK	��h�C$   �         *   Q   2         �t�bhhK ��h��R�(KK��h�CP
      1  b         D   w   �      �             2     t        �t�bhhK ��h��R�(KK��h�C,   �        �        �           �t�bhhK ��h��R�(KK��h�C8�  6      '   k  
   �  �   	   �     �        �t�bhhK ��h��R�(KK��h�C�  �  8        �t�bhhK ��h��R�(KK
��h�C(P     �        *   Q   2         �t�bhhK ��h��R�(KK��h�CT*      "         v   B      �   
   f      �   w  k  N         a         �t�bhhK ��h��R�(KK��h�C(         �t�bhhK ��h��R�(KK��h�C          $      b         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cb                     �t�bhhK ��h��R�(KK��h�Co      $      �t�bhhK ��h��R�(KK��h�C@   
   �      $      *         j   �   P     *         �t�bhhK ��h��R�(KK��h�C  o      $      �t�bhhK ��h��R�(KK��h�C0         z                 o         �t�bhhK ��h��R�(KK��h�CP.   �             :     �   �     o                           �t�bhhK ��h��R�(KK
��h�C(   O   �          �   ]         �t�bhhK ��h��R�(KK	��h�C$   7   �     *   Q   2         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�CD
      5           M  	         =   #  �     i        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C$  �        �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�Co     �t�bhhK ��h��R�(KK��h�Cp
   A  }  $      ?      I   	      �   �  @   o       �     N          �  z      �         �t�bhhK ��h��R�(KK��h�C<
      "   �      h        i   
   .   d           �t�bhhK ��h��R�(KK��h�C8           `      �        &              �t�bhhK ��h��R�(KK��h�C       D   �   2          �t�bhhK ��h��R�(KK��h�CH*      �  '        :        �  '   ?     $      �         �t�bhhK ��h��R�(KK��h�CPB      i   
      
      �  �   �   
   A     $   ?   �      �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK
��h�C(o      $                        �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK	��h�C$9  �      �                 �t�bhhK ��h��R�(KK��h�C �                        �t�bhhK ��h��R�(KK��h�C,     �     �t�bhhK ��h��R�(KK��h�Ch*      �   [  +     :   �     �  $      �      .         F   ,  	   �   �      �        �t�bhhK ��h��R�(KK��h�C,         V      o      $      �      �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C,                 �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK
��h�C(q     �   �      :   �  �        �t�bhhK ��h��R�(KK��h�C8�     q     *   �   ;   	      F     ;         �t�bhhK ��h��R�(KK��h�CL
      �   �        
   ;      �         =   ;     �           �t�bhhK ��h��R�(KK��h�C(      <            �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK
��h�C(N      �   �   
      N     �      �t�bhhK ��h��R�(KK��h�C|
      �   �   
      �   	   /     �  N  �  i      �  6   �  �  �  	         �  �      V      |        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�CV      �           �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C,      K     �t�bhhK ��h��R�(KK!��h�C�   j   �   &       *   7        
   �        y  /      *          @   +      n      _   ,      ,      K        �t�bhhK ��h��R�(KK��h�Ct   7     
   n      _   ,   D      j   �   '     _   ,      �  7   F  +   N   $      L   "   ,   h      �t�bhhK ��h��R�(KK��h�Ch   j   �   �     m      �        
   �        y  /          @   +      ,      b        �t�bhhK ��h��R�(KK��h�C�     *      �t�bhhK ��h��R�(KK��h�C�   �  G      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�   G      �t�bhhK ��h��R�(KK��h�C4  G      �t�bhhK ��h��R�(KK��h�CN      u  $      �t�bhhK ��h��R�(KK��h�C�   Y      �t�bhhK ��h��R�(KK��h�C4�   �   �   
   .      �   
      �   M        �t�bhhK ��h��R�(KK��h�CD�   �      F         �  �     N     �        L        �t�bhhK ��h��R�(KK��h�C,�   4   �   
   .   4         M        �t�bhhK ��h��R�(KK��h�C<
      "   J   S     *         �  :   �   �        �t�bhhK ��h��R�(KK��h�C4�   �   8     5  	   �  	   Q     �         �t�bhhK ��h��R�(KK��h�CP
      4   "   �      :   �   �  	         g   +         �   �        �t�bhhK ��h��R�(KK��h�C0      �   �  �      �  3  ~  %        �t�bhhK ��h��R�(KK��h�C         G         �t�bhhK ��h��R�(KK��h�C�     *      �t�bhhK ��h��R�(KK
��h�C(�   �   8     �     )           �t�bhhK ��h��R�(KK
��h�C(�  "   �   \     �     /        �t�bhhK ��h��R�(KK��h�C0   �     �  N  	   O     P  Q        �t�bhhK ��h��R�(KK
��h�C(      �   }      �   �   ]         �t�bhhK ��h��R�(KK��h�C0   *   Q   2      P     �     �        �t�bhhK ��h��R�(KK��h�C4N      �  �   	   �  r   �  4               �t�bhhK ��h��R�(KK��h�C4r   �     �        �                   �t�bhhK ��h��R�(KK��h�C      }      �        �t�bhhK ��h��R�(KK��h�CX
      4      �     �  	             �  J   }            �     p        �t�bhhK ��h��R�(KK��h�C@
      5   �  �  s  	         �     �   �            �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Ct                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C,      a             �   �         �t�bhhK ��h��R�(KK��h�CLD   :   Y      4   "   �      &   �   �     1      �   �   5        �t�bhhK ��h��R�(KK��h�C0      �   �   �      %  �  3  ~        �t�bhhK ��h��R�(KK��h�C    *      ^   �   *        �t�bhhK ��h��R�(KK��h�C0�      �   @  7         F      �        �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C�   �                 �t�bhhK ��h��R�(KK��h�C�   �                 �t�bhhK ��h��R�(KK��h�C-     �t�bhhK ��h��R�(KK��h�C4   
   �     -  7         j   �   �        �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�CL   9      3  X  	   v   Y      �     1   �   >     @   �        �t�bhhK ��h��R�(KK
��h�C(�      3  X     v     Q        �t�bhhK ��h��R�(KK��h�C03  X  �  4   Q     �     W   {        �t�bhhK ��h��R�(KK��h�C4       �  Q  �  4   �  �      �  �        �t�bhhK ��h��R�(KK
��h�C(l     3  X     9      �        �t�bhhK ��h��R�(KK
��h�C(�  �        �        @        �t�bhhK ��h��R�(KK��h�C@�     �           E      �      �      �     �     �t�bhhK ��h��R�(KK��h�C         �      1      �t�bhhK ��h��R�(KK	��h�C$�     ?   B  "   �   �        �t�bhhK ��h��R�(KK��h�C4�     z        �     �      �           �t�bhhK ��h��R�(KK��h�C,&   |  �      �         W  �         �t�bhhK ��h��R�(KK��h�C8�   &   R  �     (          U     �         �t�bhhK ��h��R�(KK��h�C�      W  �      �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C(      <      �     �t�bhhK ��h��R�(KK��h�C@      $   ?   /  I         W        �     9         �t�bhhK ��h��R�(KK	��h�C$   5   4   �   }      �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C         �      1      �t�bhhK ��h��R�(KK��h�Cn   G      �t�bhhK ��h��R�(KK��h�CX   �     C     �     H  $   O   B   +            �     0     @        �t�bhhK ��h��R�(KK��h�C<#        �   
   f      @   +      �     $         �t�bhhK ��h��R�(KK��h�C8   �  6      z                  .   6         �t�bhhK ��h��R�(KK��h�C0   *      ^   Q     >   �     �         �t�bhhK ��h��R�(KK	��h�C$j  �         *   Q   2         �t�bhhK ��h��R�(KK��h�C0      �   }         Q       �        �t�bhhK ��h��R�(KK��h�CL
   '   $     �     5   s  o   	   w   �      �      )           �t�bhhK ��h��R�(KK��h�C �  "   �   
   �  G         �t�bhhK ��h��R�(KK��h�CT?   �     B     �      $   ?   /  I      W  �         �     9         �t�bhhK ��h��R�(KK��h�C0      D   w   r   $         �   �        �t�bhhK ��h��R�(KK��h�C         n   G         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C   �                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cj  �                  �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Ct                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK
��h�C(   
   �     �                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�   �  G      �t�bhhK ��h��R�(KK
��h�C(q     �   �      :   �  �        �t�bhhK ��h��R�(KK��h�C8�     q     *   �   ;   	      F     ;         �t�bhhK ��h��R�(KK��h�CL
      �   �        
   ;      �         =   ;     �           �t�bhhK ��h��R�(KK��h�C(      <            �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK
��h�C(N      �   �   
      N     �      �t�bhhK ��h��R�(KK��h�C|
      �   �   
      �   	   /     �  N  �  i      �  6   �  �  �  	         �  �      V      |        �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�CV      �           �t�bhhK ��h��R�(KK��h�C�   �  G   	           �t�bhhK ��h��R�(KK��h�C�     �t�be.