grundläggande information
historia
trafik
religion
beslutsfattande och påverkan
grundläggande information
Karleby finns i Mellersta Österbotten invid Bottniska viken .
Karleby stad är grundad 1620 och hette då Gamlakarleby .
senare blev Kokkola stadens finska namn .
vid Karleby centrum finns en av landets mest omfattande historiska trästadshelheter .
Stadsplanen är från 1650 @-@ talet .
den omfattar 12 kvarter med hundratals trähus och gårdsbyggnader .
de äldsta av dessa är från 1600 @-@ talet .
Karleby är en kulturstad med mycket att se och uppleva .
Karleby hamn ligger i stadsdelen Yxpila och är en av Finlands mest trafikerade godshamnar .
Grunden för näringslivet i Karleby är den internationella storindustrin .
i Karleby är den kemiska industrin och industri i anslutning till denna särskilt viktig .
Karleby är även en betydande handelsstad .
information om Karlebyfinska _ svenska _ engelska
historia
redan under medeltiden fanns det hamn , båtbygge och handelsplats i Karleby .
Landhöjningen har varit en central faktor i Karlebys historia .
den har format omgivningen i hög grad och bland annat påverkat utvecklingen av hamnverksamheten och handeln .
Handel bedrevs längs med Bottniska vikens kust och jordbruk , jakt , fiske och sälfångst var även viktiga näringar .
Exporten av tjära , som blev mycket viktig för Karlebys historia , inleddes redan på 1500 @-@ talet .
den sjunde september 1620 undertecknade Sveriges kung Gustav II Adolf en handling som gav den lilla jordbruks- och fiskebyn vid Ristrand status som stad .
Dagens stadssund var då en smal havsvik som sträckte sig ända till Kyrkbacken .
Sakta men säkert blev Karleby en viktig stad för sjöfart och skeppsbygge .
Skeppsvarv fanns bland annat i Kaustarviken , Svartskär och Soldatskär .
Inledningsvis seglade man endast till Åbo och Stockholm , eftersom Karleby som s.k. uppstad inte fick bedriva utrikeshandel .
år 1765 erhöll staden stapelrättigheter , dvs. rätt till fri utrikeshandel , främst tack vare den aktiva kyrkoherden och lantdagsmannen Anders Chydenius .
Karleby blev snabbt en förmögen stad i början av 1800 @-@ talet tack vare just handeln med tjära och rederiverksamheten .
stadens borgare köpte tjära av bönder och exporterade den , ofta till hamnar vid Medelhavet och i England .
Karleby handelsflotta var under perioder Finlands största .
den snabba ekonomiska utvecklingen avtog i mitten av 1800 @-@ talet , men tog ny fart i slutet av århundradet tack vare industrialiseringen .
Karleby blev en viktig industristad främst tack vare läder- och metallindustrin .
Karlebys historiafinska _ svenska _ engelska
trafik
Karleby har goda trafikförbindelser .
via Karleby löper riksväg 8 och 13 .
Järnvägsstationen finns i stadens centrum .
Restiden med tåg till Helsingfors är cirka fyra timmar .
Flygplatsen finns i Kronoby på endast 22 kilometers avstånd från Karleby centrum .
Stadsborna erbjuds även ett tryggt , omfattande , fungerande och trivsamt nätverk för den lätta trafiken .
Karleby har satsat på att förbättra förhållandena för cyklister .
Lokalbussarna trafikerar de olika delarna av staden på vardagar .
Läs mer : trafik .
Gator och trafikfinska _ svenska
Kollektivtrafikfinska _ svenska
linkkiVR :
Tågtidtabellerfinska _ svenska _ engelska _ ryska
Busstidtabellerfinska _ svenska _ engelska
flyg från Karleby @-@ Jakobstad flygplatsfinska _ svenska _ engelska
religion
i Karleby finns flera olika religiösa samfund .
i tjänsten Uskonnot Suomessa ( Religioner i Finland ) finns information om religiösa samfund enligt ort .
den evangelisk @-@ lutherska kyrkan har fyra finskspråkiga församlingar och en svenskspråkig församling i Karleby .
Läs mer på Karleby kyrkliga samfällighets webbplats .
i Karleby finns en ortodox kyrka .
mer information om den ortodoxa församlingens verksamhet i Karleby finns på Vasa ortodoxa församlings webbplats .
Läs mer : kulturer och religioner i Finland .
linkkiKarleby kyrkliga samfällighet :
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiVasa ortodoxa församling :
Vasa ortodoxa församlingfinska _ engelska _ ryska
beslutsfattande och påverkan
den högsta beslutsfattande makten i Karleby stad innehas av stadsfullmäktige .
Fullmäktigeledamöterna och deras suppleanter väljs vid kommunalval vart fjärde år .
på stadens webbplats finns information om stadsfullmäktige och dess beslut .
invånarna kan påverka stadens beslutsfattande redan då beslut bereds .
information om olika sätt att delta och påverka finns på stadens webbplats .
kommunens invånare har enligt kommunallagen rätt att lämna in motioner till kommunen i ärenden som gäller dess verksamhet .
i Karleby finns ungdomsfullmäktige , äldre- och handikappråd samt ett råd för kulturell mångfald .
Läs mer : Finlands förvaltning , Val och röstning i Finland
beslutsfattandefinska _ svenska _ engelska
grundläggande information
historia
trafik
religion
beslutsfattande och påverkan
grundläggande information
Karleby finns i Mellersta Österbotten invid Bottniska viken .
Karleby stad är grundad 1620 och hette då Gamlakarleby .
senare blev Kokkola stadens finska namn .
vid Karleby centrum finns en av landets mest omfattande historiska trästadshelheter .
Stadsplanen är från 1650 @-@ talet .
den omfattar 12 kvarter med hundratals trähus och gårdsbyggnader .
de äldsta av dessa är från 1600 @-@ talet .
Karleby är en kulturstad med mycket att se och uppleva .
Karleby hamn ligger i stadsdelen Yxpila och är en av Finlands mest trafikerade godshamnar .
Grunden för näringslivet i Karleby är den internationella storindustrin .
i Karleby är den kemiska industrin och industri i anslutning till denna särskilt viktig .
Karleby är även en betydande handelsstad .
information om Karlebyfinska _ svenska _ engelska
historia
redan under medeltiden fanns det hamn , båtbygge och handelsplats i Karleby .
Landhöjningen har varit en central faktor i Karlebys historia .
den har format omgivningen i hög grad och bland annat påverkat utvecklingen av hamnverksamheten och handeln .
Handel bedrevs längs med Bottniska vikens kust och jordbruk , jakt , fiske och sälfångst var även viktiga näringar .
Exporten av tjära , som blev mycket viktig för Karlebys historia , inleddes redan på 1500 @-@ talet .
den sjunde september 1620 undertecknade Sveriges kung Gustav II Adolf en handling som gav den lilla jordbruks- och fiskebyn vid Ristrand status som stad .
Dagens stadssund var då en smal havsvik som sträckte sig ända till Kyrkbacken .
Sakta men säkert blev Karleby en viktig stad för sjöfart och skeppsbygge .
Skeppsvarv fanns bland annat i Kaustarviken , Svartskär och Soldatskär .
Inledningsvis seglade man endast till Åbo och Stockholm , eftersom Karleby som s.k. uppstad inte fick bedriva utrikeshandel .
år 1765 erhöll staden stapelrättigheter , dvs. rätt till fri utrikeshandel , främst tack vare den aktiva kyrkoherden och lantdagsmannen Anders Chydenius .
Karleby blev snabbt en förmögen stad i början av 1800 @-@ talet tack vare just handeln med tjära och rederiverksamheten .
stadens borgare köpte tjära av bönder och exporterade den , ofta till hamnar vid Medelhavet och i England .
Karleby handelsflotta var under perioder Finlands största .
den snabba ekonomiska utvecklingen avtog i mitten av 1800 @-@ talet , men tog ny fart i slutet av århundradet tack vare industrialiseringen .
Karleby blev en viktig industristad främst tack vare läder- och metallindustrin .
Karlebys historiafinska _ svenska _ engelska
trafik
Karleby har goda trafikförbindelser .
via Karleby löper riksväg 8 och 13 .
Järnvägsstationen finns i stadens centrum .
Restiden med tåg till Helsingfors är cirka fyra timmar .
Flygplatsen finns i Kronoby på endast 22 kilometers avstånd från Karleby centrum .
Stadsborna erbjuds även ett tryggt , omfattande , fungerande och trivsamt nätverk för den lätta trafiken .
Karleby har satsat på att förbättra förhållandena för cyklister .
Lokalbussarna trafikerar de olika delarna av staden på vardagar .
Läs mer : trafik .
Gator och trafikfinska _ svenska
Kollektivtrafikfinska _ svenska
linkkiVR :
Tågtidtabellerfinska _ svenska _ engelska _ ryska
Busstidtabellerfinska _ svenska _ engelska
flyg från Karleby @-@ Jakobstad flygplatsfinska _ svenska _ engelska
religion
i Karleby finns flera olika religiösa samfund .
i tjänsten Uskonnot Suomessa ( Religioner i Finland ) finns information om religiösa samfund enligt ort .
den evangelisk @-@ lutherska kyrkan har fyra finskspråkiga församlingar och en svenskspråkig församling i Karleby .
Läs mer på Karleby kyrkliga samfällighets webbplats .
i Karleby finns en ortodox kyrka .
mer information om den ortodoxa församlingens verksamhet i Karleby finns på Vasa ortodoxa församlings webbplats .
Läs mer : kulturer och religioner i Finland .
linkkiKarleby kyrkliga samfällighet :
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiVasa ortodoxa församling :
Vasa ortodoxa församlingfinska _ engelska _ ryska
beslutsfattande och påverkan
den högsta beslutsfattande makten i Karleby stad innehas av stadsfullmäktige .
Fullmäktigeledamöterna och deras suppleanter väljs vid kommunalval vart fjärde år .
på stadens webbplats finns information om stadsfullmäktige och dess beslut .
invånarna kan påverka stadens beslutsfattande redan då beslut bereds .
information om olika sätt att delta och påverka finns på stadens webbplats .
kommunens invånare har enligt kommunallagen rätt att lämna in motioner till kommunen i ärenden som gäller dess verksamhet .
i Karleby finns ungdomsfullmäktige , äldre- och handikappråd samt ett råd för kulturell mångfald .
Läs mer : Finlands förvaltning , Val och röstning i Finland
beslutsfattandefinska _ svenska _ engelska
grundläggande information
historia
trafik
religion
beslutsfattande och påverkan
grundläggande information
Karleby finns i Mellersta Österbotten invid Bottniska viken .
Karleby stad är grundad 1620 och hette då Gamlakarleby .
senare blev Kokkola stadens finska namn .
vid Karleby centrum finns en av landets mest omfattande historiska trästadshelheter .
Stadsplanen är från 1650 @-@ talet .
den omfattar 12 kvarter med hundratals trähus och gårdsbyggnader .
de äldsta av dessa är från 1600 @-@ talet .
Karleby är en kulturstad med mycket att se och uppleva .
Karleby hamn ligger i stadsdelen Yxpila och är en av Finlands mest trafikerade godshamnar .
Grunden för näringslivet i Karleby är den internationella storindustrin .
i Karleby är den kemiska industrin och industri i anslutning till denna särskilt viktig .
Karleby är även en betydande handelsstad .
information om Karlebyfinska _ svenska _ engelska
historia
redan under medeltiden fanns det hamn , båtbygge och handelsplats i Karleby .
Landhöjningen har varit en central faktor i Karlebys historia .
den har format omgivningen i hög grad och bland annat påverkat utvecklingen av hamnverksamheten och handeln .
Handel bedrevs längs med Bottniska vikens kust och jordbruk , jakt , fiske och sälfångst var även viktiga näringar .
Exporten av tjära , som blev mycket viktig för Karlebys historia , inleddes redan på 1500 @-@ talet .
den sjunde september 1620 undertecknade Sveriges kung Gustav II Adolf en handling som gav den lilla jordbruks- och fiskebyn vid Ristrand status som stad .
Dagens stadssund var då en smal havsvik som sträckte sig ända till Kyrkbacken .
Sakta men säkert blev Karleby en viktig stad för sjöfart och skeppsbygge .
Skeppsvarv fanns bland annat i Kaustarviken , Svartskär och Soldatskär .
Inledningsvis seglade man endast till Åbo och Stockholm , eftersom Karleby som s.k. uppstad inte fick bedriva utrikeshandel .
år 1765 erhöll staden stapelrättigheter , dvs. rätt till fri utrikeshandel , främst tack vare den aktiva kyrkoherden och lantdagsmannen Anders Chydenius .
Karleby blev snabbt en förmögen stad i början av 1800 @-@ talet tack vare just handeln med tjära och rederiverksamheten .
stadens borgare köpte tjära av bönder och exporterade den , ofta till hamnar vid Medelhavet och i England .
Karleby handelsflotta var under perioder Finlands största .
den snabba ekonomiska utvecklingen avtog i mitten av 1800 @-@ talet , men tog ny fart i slutet av århundradet tack vare industrialiseringen .
Karleby blev en viktig industristad främst tack vare läder- och metallindustrin .
Karlebys historiafinska _ svenska _ engelska
trafik
Karleby har goda trafikförbindelser .
via Karleby löper riksväg 8 och 13 .
Järnvägsstationen finns i stadens centrum .
Restiden med tåg till Helsingfors är cirka fyra timmar .
Flygplatsen finns i Kronoby på endast 22 kilometers avstånd från Karleby centrum .
Stadsborna erbjuds även ett tryggt , omfattande , fungerande och trivsamt nätverk för den lätta trafiken .
Karleby har satsat på att förbättra förhållandena för cyklister .
Lokalbussarna trafikerar de olika delarna av staden på vardagar .
Läs mer : trafik .
Gator och trafikfinska _ svenska
Kollektivtrafikfinska _ svenska
linkkiVR :
Tågtidtabellerfinska _ svenska _ engelska _ ryska
Busstidtabellerfinska _ svenska _ engelska
flyg från Karleby @-@ Jakobstad flygplatsfinska _ svenska _ engelska
religion
i Karleby finns flera olika religiösa samfund .
i tjänsten Uskonnot Suomessa ( Religioner i Finland ) finns information om religiösa samfund enligt ort .
den evangelisk @-@ lutherska kyrkan har fyra finskspråkiga församlingar och en svenskspråkig församling i Karleby .
Läs mer på Karleby kyrkliga samfällighets webbplats .
i Karleby finns en ortodox kyrka .
mer information om den ortodoxa församlingens verksamhet i Karleby finns på Vasa ortodoxa församlings webbplats .
Läs mer : kulturer och religioner i Finland .
linkkiKarleby kyrkliga samfällighet :
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiVasa ortodoxa församling :
Vasa ortodoxa församlingfinska _ engelska _ ryska
beslutsfattande och påverkan
den högsta beslutsfattande makten i Karleby stad innehas av stadsfullmäktige .
Fullmäktigeledamöterna och deras suppleanter väljs vid kommunalval vart fjärde år .
på stadens webbplats finns information om stadsfullmäktige och dess beslut .
invånarna kan påverka stadens beslutsfattande redan då beslut bereds .
information om olika sätt att delta och påverka finns på stadens webbplats .
kommunens invånare har enligt kommunallagen rätt att lämna in motioner till kommunen i ärenden som gäller dess verksamhet .
i Karleby finns ungdomsfullmäktige , äldre- och handikappråd samt ett råd för kulturell mångfald .
Läs mer : Finlands förvaltning , Val och röstning i Finland
beslutsfattandefinska _ svenska _ engelska
detta innehåll finns inte på det språk som du har valt .
Välj något annat språk .
finska
detta innehåll finns inte på det språk som du har valt .
Välj något annat språk .
finska
detta innehåll finns inte på det språk som du har valt .
Välj något annat språk .
finska
bibliotek
motion
att röra sig i naturen
teater och film
museer
hobbyer för barn och unga
föreningar
Karleby är en gammal sjöstad som erbjuder mångsidiga möjligheter för utfärder och friluftsliv .
personer ntresserad av friluftsliv bör läsa mer om allemansrätten under rubriken &quot; Att röra sig i naturen &quot; i denna tjänst .
flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet .
föreningar och organisationer samt hobbygrupper och kommunala institut erbjuder kurser i idrott och kultur samt bl.a. språk och hantverk .
i Snellman @-@ salen och i stadens övriga kulturlokaler erbjuds kulturevenemang av varierande slag .
Årliga evenemang i Karleby är bland annat Veneziansk afton i slutet av sommaren , Kokkola Cup för fotbollsjuniorer , Stadsfestivalen Karleby sommarveckor , Lochteå kyrkomusikfest samt Vinterdans i Karleby och festivalen Karleby Vinterharmonika .
mer information om fritidstjänsterna i Karleby finns på Karleby stads webbplats .
på stadens webbplats finns även en länk till Evenemangskalendern med daglig information om stadens kultur- och motionsevenemang .
Läs mer : Fritid .
Evenemangskalenderfinska
Kulturtjänsterfinska _ svenska _ engelska
Idrottstjänsterfinska _ svenska _ engelska
bibliotek
Karleby stadsbibliotek finns i stadens centrum .
Närbiblioteken finns i Björkhagen , Kelviå , Lochteå samt Ullava kyrkby och Rahkonen .
information om bibliotekets öppettider och tjänster finns på dess webbplats .
biblioteket finns även på nätet .
där kan kunderna bläddra i bibliotekets samlingar , reservera material , förnya sina lån , beställa fjärrlån och låna e @-@ böcker under alla tider på dygnet .
tack vare det effektiva biblioteksnätverket i Finland är nästan alla finländska biblioteks samlingar tillgängliga för bibliotekskunderna i Karleby .
Karleby stadsbibliotek / huvudbiblioteket
Storgatan 3 , 67100 Karleby
telefon : 040.806.5124 , 040.806.5133
Läs mer : bibliotek .
Bibliotekstjänsterfinska _ svenska _ engelska
motion
i Karleby finns mångsidiga motionsmöjligheter året runt .
staden anordnar ledda aktiviteter i Simcentret VesiVeijari och motionshallarna .
dessutom finns det gym av flera olika slag .
gym anpassade för äldre finns i Furuåsens aktivitetscenter och Kuusikumpu servicehus .
staden underhåller cykelvägar , motionsrutter , joggingbanor , skidspår , badstränder , bollplaner och skridskobanor samt platser för närmotion .
i Karlebynejdens instituts nättjänst finns information om institutets mångsidiga motionsutbud .
i Karleby finns nära på hundra idrottsföreningar för olika grenar samt föreningar som arrangerar övrig motion .
mer information om motionsmöjligheter i Karleby finns på Karleby stads webbplats .
Läs mer :
motion .
Idrottstjänsterfinska _ svenska _ engelska
Motionsplatserfinska _ svenska
gym för äldrefinska
Karlebynejdens institutfinska _ svenska
att röra sig i naturen
att röra sig i naturen är en traditionell och populär form av avkoppling för finländarna under alla årstider .
i Finland kan man med stöd av allemansrätten plocka bär och svamp i skogen och röra sig till fots , med cykel eller skidor vintertid .
det är inte tillåtet att beträda folks gårdar utan lov .
för fiske krävs fiskelov , med undantag för mete och pilkning .
även jakt fordrar jakttillstånd .
allemansrätten ger inte rätt att skräpa ner i naturen , skada träd eller växter , störa eller skada fågelbon eller fågelungar , köra motorfordon utan markägarens tillstånd eller bygga ens tillfälliga byggen .
mer information om motionsrutterna , rastplatser , möjligheter till fiske och båtliv samt exempelvis fågeltorn i Karleby finns på stadens webbplats .
rutterna för camping , paddling , vandring , cykling och övriga rutter i Karleby finns i karttjänsten på nätet .
i karttjänsten visas även var största delen av motionsplatserna finns .
du kan köpa friluftskartor över Karleby hos Karleby Turism : Salutorget 5 , 67100 Karleby .
Läs mer : att röra sig i naturen .
linkkiMiljöförvaltningen :
Allemansrättenfinska _ svenska _ engelska _ ryska
Motionskarta över Karlebyfinska _ svenska
motionsrutter i Karlebyfinska _ svenska
teater och film
Karleby är en teaterstad med långa anor , som erbjuder scenkonst på hög nivå framförd av både proffs och amatörer .
Karleby stadsteater finns i det stämningsfulla Vartiolinna ( Torggatan 48 ) .
du kan läsa mer om amatörteatrarnas verksamhet på deras webbplats och i evenemangskalendern .
i Karleby finns biografen Bio Rex , vars två salar använder digital- och 3D @-@ teknik .
Bio Rex program finns under länken här intill .
Läs mer : teater och film .
Stadsteaternfinska
Biograffinska
teater och danskonst i Karlebyfinska _ svenska _ engelska
Evenemangskalenderfinska
museer
i hjärtat av staden , i det anrika Rooska gården , finns K.H.Renlunds museum .
Karleby stad grundade museet 1909 utgående från en testamentsgåva av affärsmannen Karl Herman Renlund ( 1850 @-@ 1908 ) .
på museet finns Renlunds samling av finländsk konst från guldåldern och tillfälliga utställningar i en kulturhistorisk miljö .
även i museikvarterens övriga byggnader finns utställningar om stadens kulturhistoria och utställningar med ITE @-@ konst .
på K.H.Renlunds museums webbplats finns mer information om museets tjänster , utställningar samt aktuell verksamhet .
Utöver K.H.Renlunds museum lönar det sig att besöka det naturhistoriska museet Kieppi ( Kieppi är stängt tills vidare på grund av brand ) samt de många hembygdsmuseerna och övriga de historiska resmålen i regionen .
exempelvis i Konst @-@ Vionoja @-@ centret presenteras konstnären Veikko Vionojas verk .
i Kelviå , ca 10 km norrut från Karleby , finns Toivonen djurpark och drängmuseum .
mer information om dessa museer finns under länkarna här intill .
Läs mer : museer .
museer och traditionsarbetefinska _ svenska _ engelska
K.H. Renlunds museum - Mellersta Österbottens landskapsmuseumfinska _ svenska _ engelska
Kieppi , Karleby naturvetenskapliga museumfinska _ svenska _ engelska
linkkiToivonens djurpark och drängmuseum :
Toivonens djurpark och drängmuseum finska _ svenska _ engelska
konst Vionojafinska
hobbyer för barn och unga
flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet .
flera olika föreningar samt kommunala institut ger unga möjlighet att studera idrott och kultur samt bl.a. språk och hantverk .
barn och unga kan delta i grundläggande undervisning i musik , dans , bildkonst och hantverk .
dessutom erbjuder stadens ungdomstjänster en rockskola .
stadens ungdomstjänster driver sju ungdomsgårdar runt om i Karleby .
de rusmedels- och rökfria ungdomslokalerna erbjuder handledd verksamhet för barn i årskurserna 3 @-@ 6 och unga i åldern 13 @-@ 17 år i olika delar av Karleby .
information om hobbyverksamheter för barn och unga finns på stadens webbplats .
rådgivningen vid Ungdomsgården Vinge ger aktuell information om bl.a. internationalisering , studier , arbetsliv , hälsa , hobbyverksamhet och boende .
Karlebynejdens institut erbjuder barn och unga olika former av hobbyverksamhet , exempelvis i konstämnen och musik .
kontrollera vilka kurser som är aktuella i institutets webbtjänst .
Karleby evangelisk @-@ lutherska församlingar erbjuder även hobbyverksamhet för barn och unga , såsom lekparksträffar , klubbar , musikverksamhet och läger .
mer information om verksamheten finns på Karleby församlingssammanslutnings webbplats .
ungdomsgården Vinge
67100 Karleby
Läs mer : hobbyer för barn och unga .
övrig undervisning i Karlebyfinska _ svenska
Ungdomstjänsterfinska _ svenska _ engelska
Karlebynejdens institutfinska _ svenska
linkkiKarleby kyrkliga samfällighet :
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
föreningar
Karleby har ett aktivt och mångsidigt föreningsliv för invånare i alla åldrar .
Läs mer : föreningar .
bibliotek
motion
att röra sig i naturen
teater och film
museer
hobbyer för barn och unga
föreningar
Karleby är en gammal sjöstad som erbjuder mångsidiga möjligheter för utfärder och friluftsliv .
personer ntresserad av friluftsliv bör läsa mer om allemansrätten under rubriken &quot; Att röra sig i naturen &quot; i denna tjänst .
flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet .
föreningar och organisationer samt hobbygrupper och kommunala institut erbjuder kurser i idrott och kultur samt bl.a. språk och hantverk .
i Snellman @-@ salen och i stadens övriga kulturlokaler erbjuds kulturevenemang av varierande slag .
Årliga evenemang i Karleby är bland annat Veneziansk afton i slutet av sommaren , Kokkola Cup för fotbollsjuniorer , Stadsfestivalen Karleby sommarveckor , Lochteå kyrkomusikfest samt Vinterdans i Karleby och festivalen Karleby Vinterharmonika .
mer information om fritidstjänsterna i Karleby finns på Karleby stads webbplats .
på stadens webbplats finns även en länk till Evenemangskalendern med daglig information om stadens kultur- och motionsevenemang .
Läs mer : Fritid .
Evenemangskalenderfinska
Kulturtjänsterfinska _ svenska _ engelska
Idrottstjänsterfinska _ svenska _ engelska
bibliotek
Karleby stadsbibliotek finns i stadens centrum .
Närbiblioteken finns i Björkhagen , Kelviå , Lochteå samt Ullava kyrkby och Rahkonen .
information om bibliotekets öppettider och tjänster finns på dess webbplats .
biblioteket finns även på nätet .
där kan kunderna bläddra i bibliotekets samlingar , reservera material , förnya sina lån , beställa fjärrlån och låna e @-@ böcker under alla tider på dygnet .
tack vare det effektiva biblioteksnätverket i Finland är nästan alla finländska biblioteks samlingar tillgängliga för bibliotekskunderna i Karleby .
Karleby stadsbibliotek / huvudbiblioteket
Storgatan 3 , 67100 Karleby
telefon : 040.806.5124 , 040.806.5133
Läs mer : bibliotek .
Bibliotekstjänsterfinska _ svenska _ engelska
motion
i Karleby finns mångsidiga motionsmöjligheter året runt .
staden anordnar ledda aktiviteter i Simcentret VesiVeijari och motionshallarna .
dessutom finns det gym av flera olika slag .
gym anpassade för äldre finns i Furuåsens aktivitetscenter och Kuusikumpu servicehus .
staden underhåller cykelvägar , motionsrutter , joggingbanor , skidspår , badstränder , bollplaner och skridskobanor samt platser för närmotion .
i Karlebynejdens instituts nättjänst finns information om institutets mångsidiga motionsutbud .
i Karleby finns nära på hundra idrottsföreningar för olika grenar samt föreningar som arrangerar övrig motion .
mer information om motionsmöjligheter i Karleby finns på Karleby stads webbplats .
Läs mer :
motion .
Idrottstjänsterfinska _ svenska _ engelska
Motionsplatserfinska _ svenska
gym för äldrefinska
Karlebynejdens institutfinska _ svenska
att röra sig i naturen
att röra sig i naturen är en traditionell och populär form av avkoppling för finländarna under alla årstider .
i Finland kan man med stöd av allemansrätten plocka bär och svamp i skogen och röra sig till fots , med cykel eller skidor vintertid .
det är inte tillåtet att beträda folks gårdar utan lov .
för fiske krävs fiskelov , med undantag för mete och pilkning .
även jakt fordrar jakttillstånd .
allemansrätten ger inte rätt att skräpa ner i naturen , skada träd eller växter , störa eller skada fågelbon eller fågelungar , köra motorfordon utan markägarens tillstånd eller bygga ens tillfälliga byggen .
mer information om motionsrutterna , rastplatser , möjligheter till fiske och båtliv samt exempelvis fågeltorn i Karleby finns på stadens webbplats .
rutterna för camping , paddling , vandring , cykling och övriga rutter i Karleby finns i karttjänsten på nätet .
i karttjänsten visas även var största delen av motionsplatserna finns .
du kan köpa friluftskartor över Karleby hos Karleby Turism : Salutorget 5 , 67100 Karleby .
Läs mer : att röra sig i naturen .
linkkiMiljöförvaltningen :
Allemansrättenfinska _ svenska _ engelska _ ryska
Motionskarta över Karlebyfinska _ svenska
motionsrutter i Karlebyfinska _ svenska
teater och film
Karleby är en teaterstad med långa anor , som erbjuder scenkonst på hög nivå framförd av både proffs och amatörer .
Karleby stadsteater finns i det stämningsfulla Vartiolinna ( Torggatan 48 ) .
du kan läsa mer om amatörteatrarnas verksamhet på deras webbplats och i evenemangskalendern .
i Karleby finns biografen Bio Rex , vars två salar använder digital- och 3D @-@ teknik .
Bio Rex program finns under länken här intill .
Läs mer : teater och film .
Stadsteaternfinska
Biograffinska
teater och danskonst i Karlebyfinska _ svenska _ engelska
Evenemangskalenderfinska
museer
i hjärtat av staden , i det anrika Rooska gården , finns K.H.Renlunds museum .
Karleby stad grundade museet 1909 utgående från en testamentsgåva av affärsmannen Karl Herman Renlund ( 1850 @-@ 1908 ) .
på museet finns Renlunds samling av finländsk konst från guldåldern och tillfälliga utställningar i en kulturhistorisk miljö .
även i museikvarterens övriga byggnader finns utställningar om stadens kulturhistoria och utställningar med ITE @-@ konst .
på K.H.Renlunds museums webbplats finns mer information om museets tjänster , utställningar samt aktuell verksamhet .
Utöver K.H.Renlunds museum lönar det sig att besöka det naturhistoriska museet Kieppi ( Kieppi är stängt tills vidare på grund av brand ) samt de många hembygdsmuseerna och övriga de historiska resmålen i regionen .
exempelvis i Konst @-@ Vionoja @-@ centret presenteras konstnären Veikko Vionojas verk .
i Kelviå , ca 10 km norrut från Karleby , finns Toivonen djurpark och drängmuseum .
mer information om dessa museer finns under länkarna här intill .
Läs mer : museer .
museer och traditionsarbetefinska _ svenska _ engelska
K.H. Renlunds museum - Mellersta Österbottens landskapsmuseumfinska _ svenska _ engelska
Kieppi , Karleby naturvetenskapliga museumfinska _ svenska _ engelska
linkkiToivonens djurpark och drängmuseum :
Toivonens djurpark och drängmuseum finska _ svenska _ engelska
konst Vionojafinska
hobbyer för barn och unga
flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet .
flera olika föreningar samt kommunala institut ger unga möjlighet att studera idrott och kultur samt bl.a. språk och hantverk .
barn och unga kan delta i grundläggande undervisning i musik , dans , bildkonst och hantverk .
dessutom erbjuder stadens ungdomstjänster en rockskola .
stadens ungdomstjänster driver sju ungdomsgårdar runt om i Karleby .
de rusmedels- och rökfria ungdomslokalerna erbjuder handledd verksamhet för barn i årskurserna 3 @-@ 6 och unga i åldern 13 @-@ 17 år i olika delar av Karleby .
information om hobbyverksamheter för barn och unga finns på stadens webbplats .
rådgivningen vid Ungdomsgården Vinge ger aktuell information om bl.a. internationalisering , studier , arbetsliv , hälsa , hobbyverksamhet och boende .
Karlebynejdens institut erbjuder barn och unga olika former av hobbyverksamhet , exempelvis i konstämnen och musik .
kontrollera vilka kurser som är aktuella i institutets webbtjänst .
Karleby evangelisk @-@ lutherska församlingar erbjuder även hobbyverksamhet för barn och unga , såsom lekparksträffar , klubbar , musikverksamhet och läger .
mer information om verksamheten finns på Karleby församlingssammanslutnings webbplats .
ungdomsgården Vinge
67100 Karleby
Läs mer : hobbyer för barn och unga .
övrig undervisning i Karlebyfinska _ svenska
Ungdomstjänsterfinska _ svenska _ engelska
Karlebynejdens institutfinska _ svenska
linkkiKarleby kyrkliga samfällighet :
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
föreningar
Karleby har ett aktivt och mångsidigt föreningsliv för invånare i alla åldrar .
Läs mer : föreningar .
bibliotek
motion
att röra sig i naturen
teater och film
museer
hobbyer för barn och unga
föreningar
Karleby är en gammal sjöstad som erbjuder mångsidiga möjligheter för utfärder och friluftsliv .
personer ntresserad av friluftsliv bör läsa mer om allemansrätten under rubriken &quot; Att röra sig i naturen &quot; i denna tjänst .
flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet .
föreningar och organisationer samt hobbygrupper och kommunala institut erbjuder kurser i idrott och kultur samt bl.a. språk och hantverk .
i Snellman @-@ salen och i stadens övriga kulturlokaler erbjuds kulturevenemang av varierande slag .
Årliga evenemang i Karleby är bland annat Veneziansk afton i slutet av sommaren , Kokkola Cup för fotbollsjuniorer , Stadsfestivalen Karleby sommarveckor , Lochteå kyrkomusikfest samt Vinterdans i Karleby och festivalen Karleby Vinterharmonika .
mer information om fritidstjänsterna i Karleby finns på Karleby stads webbplats .
på stadens webbplats finns även en länk till Evenemangskalendern med daglig information om stadens kultur- och motionsevenemang .
Läs mer : Fritid .
Evenemangskalenderfinska
Kulturtjänsterfinska _ svenska _ engelska
Idrottstjänsterfinska _ svenska _ engelska
bibliotek
Karleby stadsbibliotek finns i stadens centrum .
Närbiblioteken finns i Björkhagen , Kelviå , Lochteå samt Ullava kyrkby och Rahkonen .
information om bibliotekets öppettider och tjänster finns på dess webbplats .
biblioteket finns även på nätet .
där kan kunderna bläddra i bibliotekets samlingar , reservera material , förnya sina lån , beställa fjärrlån och låna e @-@ böcker under alla tider på dygnet .
tack vare det effektiva biblioteksnätverket i Finland är nästan alla finländska biblioteks samlingar tillgängliga för bibliotekskunderna i Karleby .
Karleby stadsbibliotek / huvudbiblioteket
Storgatan 3 , 67100 Karleby
telefon : 040.806.5124 , 040.806.5133
Läs mer : bibliotek .
Bibliotekstjänsterfinska _ svenska _ engelska
motion
i Karleby finns mångsidiga motionsmöjligheter året runt .
staden anordnar ledda aktiviteter i Simcentret VesiVeijari och motionshallarna .
dessutom finns det gym av flera olika slag .
gym anpassade för äldre finns i Furuåsens aktivitetscenter och Kuusikumpu servicehus .
staden underhåller cykelvägar , motionsrutter , joggingbanor , skidspår , badstränder , bollplaner och skridskobanor samt platser för närmotion .
i Karlebynejdens instituts nättjänst finns information om institutets mångsidiga motionsutbud .
i Karleby finns nära på hundra idrottsföreningar för olika grenar samt föreningar som arrangerar övrig motion .
mer information om motionsmöjligheter i Karleby finns på Karleby stads webbplats .
Läs mer :
motion .
Idrottstjänsterfinska _ svenska _ engelska
Motionsplatserfinska _ svenska
gym för äldrefinska
Karlebynejdens institutfinska _ svenska
att röra sig i naturen
att röra sig i naturen är en traditionell och populär form av avkoppling för finländarna under alla årstider .
i Finland kan man med stöd av allemansrätten plocka bär och svamp i skogen och röra sig till fots , med cykel eller skidor vintertid .
det är inte tillåtet att beträda folks gårdar utan lov .
för fiske krävs fiskelov , med undantag för mete och pilkning .
även jakt fordrar jakttillstånd .
allemansrätten ger inte rätt att skräpa ner i naturen , skada träd eller växter , störa eller skada fågelbon eller fågelungar , köra motorfordon utan markägarens tillstånd eller bygga ens tillfälliga byggen .
mer information om motionsrutterna , rastplatser , möjligheter till fiske och båtliv samt exempelvis fågeltorn i Karleby finns på stadens webbplats .
rutterna för camping , paddling , vandring , cykling och övriga rutter i Karleby finns i karttjänsten på nätet .
i karttjänsten visas även var största delen av motionsplatserna finns .
du kan köpa friluftskartor över Karleby hos Karleby Turism : Salutorget 5 , 67100 Karleby .
Läs mer : att röra sig i naturen .
linkkiMiljöförvaltningen :
Allemansrättenfinska _ svenska _ engelska _ ryska
Motionskarta över Karlebyfinska _ svenska
motionsrutter i Karlebyfinska _ svenska
teater och film
Karleby är en teaterstad med långa anor , som erbjuder scenkonst på hög nivå framförd av både proffs och amatörer .
Karleby stadsteater finns i det stämningsfulla Vartiolinna ( Torggatan 48 ) .
du kan läsa mer om amatörteatrarnas verksamhet på deras webbplats och i evenemangskalendern .
i Karleby finns biografen Bio Rex , vars två salar använder digital- och 3D @-@ teknik .
Bio Rex program finns under länken här intill .
Läs mer : teater och film .
Stadsteaternfinska
Biograffinska
teater och danskonst i Karlebyfinska _ svenska _ engelska
Evenemangskalenderfinska
museer
i hjärtat av staden , i det anrika Rooska gården , finns K.H.Renlunds museum .
Karleby stad grundade museet 1909 utgående från en testamentsgåva av affärsmannen Karl Herman Renlund ( 1850 @-@ 1908 ) .
på museet finns Renlunds samling av finländsk konst från guldåldern och tillfälliga utställningar i en kulturhistorisk miljö .
även i museikvarterens övriga byggnader finns utställningar om stadens kulturhistoria och utställningar med ITE @-@ konst .
på K.H.Renlunds museums webbplats finns mer information om museets tjänster , utställningar samt aktuell verksamhet .
Utöver K.H.Renlunds museum lönar det sig att besöka det naturhistoriska museet Kieppi ( Kieppi är stängt tills vidare på grund av brand ) samt de många hembygdsmuseerna och övriga de historiska resmålen i regionen .
exempelvis i Konst @-@ Vionoja @-@ centret presenteras konstnären Veikko Vionojas verk .
i Kelviå , ca 10 km norrut från Karleby , finns Toivonen djurpark och drängmuseum .
mer information om dessa museer finns under länkarna här intill .
Läs mer : museer .
museer och traditionsarbetefinska _ svenska _ engelska
K.H. Renlunds museum - Mellersta Österbottens landskapsmuseumfinska _ svenska _ engelska
Kieppi , Karleby naturvetenskapliga museumfinska _ svenska _ engelska
linkkiToivonens djurpark och drängmuseum :
Toivonens djurpark och drängmuseum finska _ svenska _ engelska
konst Vionojafinska
hobbyer för barn och unga
flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet .
flera olika föreningar samt kommunala institut ger unga möjlighet att studera idrott och kultur samt bl.a. språk och hantverk .
barn och unga kan delta i grundläggande undervisning i musik , dans , bildkonst och hantverk .
dessutom erbjuder stadens ungdomstjänster en rockskola .
stadens ungdomstjänster driver sju ungdomsgårdar runt om i Karleby .
de rusmedels- och rökfria ungdomslokalerna erbjuder handledd verksamhet för barn i årskurserna 3 @-@ 6 och unga i åldern 13 @-@ 17 år i olika delar av Karleby .
information om hobbyverksamheter för barn och unga finns på stadens webbplats .
rådgivningen vid Ungdomsgården Vinge ger aktuell information om bl.a. internationalisering , studier , arbetsliv , hälsa , hobbyverksamhet och boende .
Karlebynejdens institut erbjuder barn och unga olika former av hobbyverksamhet , exempelvis i konstämnen och musik .
kontrollera vilka kurser som är aktuella i institutets webbtjänst .
Karleby evangelisk @-@ lutherska församlingar erbjuder även hobbyverksamhet för barn och unga , såsom lekparksträffar , klubbar , musikverksamhet och läger .
mer information om verksamheten finns på Karleby församlingssammanslutnings webbplats .
ungdomsgården Vinge
67100 Karleby
Läs mer : hobbyer för barn och unga .
övrig undervisning i Karlebyfinska _ svenska
Ungdomstjänsterfinska _ svenska _ engelska
Karlebynejdens institutfinska _ svenska
linkkiKarleby kyrkliga samfällighet :
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
föreningar
Karleby har ett aktivt och mångsidigt föreningsliv för invånare i alla åldrar .
Läs mer : föreningar .
problem med uppehållstillstånd
brott
våld
diskriminering och rasism
behöver du en jurist ?
Död
problem i äktenskap eller parförhållande
skilsmässa
problem med den mentala hälsan
missbruksproblem
i en krissituation kan du ringa nödcentralen på numret 112 .
de slussar vid behov dig vidare till socialjouren .
du ska endast ringa nödcentralen i brådskande nödsituationer , där liv , egendom eller miljön är i fara .
problem med uppehållstillstånd
om du har problem eller oklarheter med ditt uppehållstillstånd kan du kontakta Migrationsverket .
Migrationsverket
Korsholmsesplanaden 45
Vasa
Läs mer : problem med uppehållstillstånd .
brott
om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112 .
ring inte nödnumret om det inte är fråga om en nödsituation .
du kan göra en polisanmälan på nätet .
mer information finns på Polisens webbplats .
du kan även skriva ut anmälningsblanketten på nätet och lämna in den till polisstationen .
Karleby polisstation
Karlebygatan 74
67100 Karleby
Läs mer : brott .
tidsbokningfinska _ svenska _ engelska
Polisamälanfinska _ svenska _ engelska
våld
om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112 .
Läs mer : våld .
diskriminering och rasism
om du misstänker att du blivit utsatt för diskriminering då du sökt arbete eller på arbetsplatsen ska du först ta upp detta på din arbetsplats .
om saken inte kan lösas på arbetsplatsen ska du kontakta arbetarskyddet vid Regionförvaltningsverket i Västra och Inre Finland .
Besöksadress :
Regionförvaltningsverket i Västra och Inre Finland
Wollfskavägen 35
65101 Vasa
telefon : 0295.018.450
om du utsätts för diskriminering kan du be om hjälp av Diskrimineringsombudsmannen .
om du fallit offer för ett rasistiskt motiverat brott kan du göra en polisanmälan på nätet eller polisstationen .
Läs mer : diskriminering och rasism .
linkkiRegionförvaltningsverket i Västra och Inre Finland :
Regionförvaltningsverket i Västra och Inre Finlandfinska _ svenska _ engelska
hjälp och information för personer som drabbats av etnisk diskrimineringfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
behöver du en jurist ?
juridiska tjänster är avgiftsbelagda men om du har små eller medelstora inkomster , kan du få helt eller delvis avgiftsfri rättshjälp från statens rättshjälpsbyrå .
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
Besöksadress : Ämbetshuset , Torggatan 40 , 67100 Karleby
telefon : 029.566.1270
information om enskilda jurister finns bland annat på Finlands Advokatförbunds webbplats .
Läs mer :
behöver du en jurist ?
linkkiFinlands advokatförbund :
Finlands advokatförbundfinska _ svenska _ engelska
Död
den evangelisk @-@ lutherska kyrkans församlingars begravningsplatser fungerar som allmänna begravningsplatser .
där kan även avlidna som inte är medlemmar i kyrkan begravas .
de är alltså avsedda för alla invånare i staden .
mer information finns på Karleby kyrkliga samfällighets webbplats .
om en närstående plötsligt dör kan du söka krishjälp vid din egen hälsostation , eller utanför tjänstetid vid samjouren för Mellersta Österbottens centralsjukhus .
de evangelisk @-@ lutherska församlingarna i Karlebynejden erbjuder även sorggrupper .
även församlingarnas diakonimottagningar erbjuder samtalshjälp för sorgearbetet .
Läs mer : Död .
linkkiKarleby kyrkliga samfällighet :
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Hälsostationernafinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
problem i äktenskap eller parförhållande
vid problem i äktenskap eller parförhållande får du hjälp av Mellersta Österbottens familjerådgivningscentral som underhålls av Karleby kyrkliga samfällighets och Mellersta Österbottens social- och hälsovårdssamkommun Soites familjerådgivning .
Familjerågivningscentralen
telefon : 050.3147.464 .
Karleby familjerådgivning
67100 Karleby
tel . 044.730.7640
Läs mer : problem i äktenskap eller parförhållande .
linkkiMellersta Österbottens Familjerådgivningscentral :
familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
familjerådgivningfinska _ svenska
skilsmässa
skilsmässa kan sökas av kvinnan , av mannen eller av båda makarna tillsammans .
man ansöker om skilsmässa i tingsrätten .
till att börja med görs en skriftlig skilsmässoansökan .
Österbottens tingsrätt Karleby kansli
Besöksadress : Karlebygatan 27 , 67100 Karleby
telefon : 029.56.49294
Läs mer : skilsmässa .
hälsovårdaren på barnrådgivningsbyrån ger råd i frågor som gäller små barns hälsa , tillväxt och utveckling .
barnrådgivningsbyrån ger information om platser som erbjuder hjälp vid behov .
vid problem hos unga i skolåldern hjälper exempelvis skolans hälsovårdare eller skolkuratorn .
Läs mer : barns och ungas problem .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Skolhälsovårdfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Barnrådgivningarfinska _ svenska
du kan ta upp problem med hälsovårdaren på skolan eller studieplatsen eller vuxna på ungdomsgården .
mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats .
föräldrar eller unga själva kan kontakta familjerådgivningen .
där kan man tala om problem och få hjälp och stöd .
mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats .
Familjerådgivningens telefonnummer : 044.730.7640 .
Läs mer : barns och ungas problem .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Studerandehälsovårdfinska _ svenska
ungdomsgårdar och -lokaler finska _ svenska
problem med den mentala hälsan
om du behöver hjälp och stöd för din mentala hälsa kan du boka en läkartid vid hälsostationen .
läkaren bedömer situationen .
vid behov skriver läkaren en remiss till psykiatrisk specialsjukvård .
Läs mer : mental hälsa .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Mentalvårdstjänsterfinska _ svenska
om du har ekonomiska problem kan du be om råd hos Mellersta Österbottens social- och hälsovårdssamkommun Soites enheter för socialarbete eller utkomststöd , tfn 040.806.5095 eller tjänstestyrningen , tfn 040.806.5093 .
om du har problem med skulder , kontakta rättshjälpsbyrån .
du kan anlita vilken som helst rättshjälpsbyrå oberoende av din hemkommun .
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
telefon : 029.566.1270
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Servicehandledningfinska _ svenska
missbruksproblem
om du har problem med alkohol , droger , läkemedel eller hasardspel kan du få vård och rehabilitering vid Porten , Mellersta Österbottens social- och hälsovårdssamkommun Soites center för missbruksproblem .
du kan ta upp problemet med proffs inom hälsovården eller företagshälsovården , som kan slussa dig vidare i vårdsystemet , eller direkt kontakta Soites missbrukstjänster , tfn 040.8068.101 .
för tillnyktrings- och avgiftningsvård debiteras en patientavgift liksom även för korttidsrehabilitering , öppen rehabilitering är gratis .
även Karleby evangelisk @-@ lutherska församlingssammanslutnings specialdiakoner erbjuder samtalshjälp vid missbruksproblem .
kontaktuppgifter
Hälsovägen 4
67200 Karleby
telefon : 040.806.8101
Läs mer : missbruksproblem .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Service för missbrukarefinska _ svenska
linkkiKarleby evangelisk @-@ lutherska församlingssammansutning :
Karleby evangelisk @-@ lutherska församlings arbete bland missbrukarefinska _ svenska
problem med uppehållstillstånd
brott
våld
diskriminering och rasism
behöver du en jurist ?
Död
problem i äktenskap eller parförhållande
skilsmässa
problem med den mentala hälsan
missbruksproblem
i en krissituation kan du ringa nödcentralen på numret 112 .
de slussar vid behov dig vidare till socialjouren .
du ska endast ringa nödcentralen i brådskande nödsituationer , där liv , egendom eller miljön är i fara .
problem med uppehållstillstånd
om du har problem eller oklarheter med ditt uppehållstillstånd kan du kontakta Migrationsverket .
Migrationsverket
Korsholmsesplanaden 45
Vasa
Läs mer : problem med uppehållstillstånd .
brott
om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112 .
ring inte nödnumret om det inte är fråga om en nödsituation .
du kan göra en polisanmälan på nätet .
mer information finns på Polisens webbplats .
du kan även skriva ut anmälningsblanketten på nätet och lämna in den till polisstationen .
Karleby polisstation
Karlebygatan 74
67100 Karleby
Läs mer : brott .
tidsbokningfinska _ svenska _ engelska
Polisamälanfinska _ svenska _ engelska
våld
om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112 .
Läs mer : våld .
diskriminering och rasism
om du misstänker att du blivit utsatt för diskriminering då du sökt arbete eller på arbetsplatsen ska du först ta upp detta på din arbetsplats .
om saken inte kan lösas på arbetsplatsen ska du kontakta arbetarskyddet vid Regionförvaltningsverket i Västra och Inre Finland .
Besöksadress :
Regionförvaltningsverket i Västra och Inre Finland
Wollfskavägen 35
65101 Vasa
telefon : 0295.018.450
om du utsätts för diskriminering kan du be om hjälp av Diskrimineringsombudsmannen .
om du fallit offer för ett rasistiskt motiverat brott kan du göra en polisanmälan på nätet eller polisstationen .
Läs mer : diskriminering och rasism .
linkkiRegionförvaltningsverket i Västra och Inre Finland :
Regionförvaltningsverket i Västra och Inre Finlandfinska _ svenska _ engelska
hjälp och information för personer som drabbats av etnisk diskrimineringfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
behöver du en jurist ?
juridiska tjänster är avgiftsbelagda men om du har små eller medelstora inkomster , kan du få helt eller delvis avgiftsfri rättshjälp från statens rättshjälpsbyrå .
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
Besöksadress : Ämbetshuset , Torggatan 40 , 67100 Karleby
telefon : 029.566.1270
information om enskilda jurister finns bland annat på Finlands Advokatförbunds webbplats .
Läs mer :
behöver du en jurist ?
linkkiFinlands advokatförbund :
Finlands advokatförbundfinska _ svenska _ engelska
Död
den evangelisk @-@ lutherska kyrkans församlingars begravningsplatser fungerar som allmänna begravningsplatser .
där kan även avlidna som inte är medlemmar i kyrkan begravas .
de är alltså avsedda för alla invånare i staden .
mer information finns på Karleby kyrkliga samfällighets webbplats .
om en närstående plötsligt dör kan du söka krishjälp vid din egen hälsostation , eller utanför tjänstetid vid samjouren för Mellersta Österbottens centralsjukhus .
de evangelisk @-@ lutherska församlingarna i Karlebynejden erbjuder även sorggrupper .
även församlingarnas diakonimottagningar erbjuder samtalshjälp för sorgearbetet .
Läs mer : Död .
linkkiKarleby kyrkliga samfällighet :
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Hälsostationernafinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
problem i äktenskap eller parförhållande
vid problem i äktenskap eller parförhållande får du hjälp av Mellersta Österbottens familjerådgivningscentral som underhålls av Karleby kyrkliga samfällighets och Mellersta Österbottens social- och hälsovårdssamkommun Soites familjerådgivning .
Familjerågivningscentralen
telefon : 050.3147.464 .
Karleby familjerådgivning
67100 Karleby
tel . 044.730.7640
Läs mer : problem i äktenskap eller parförhållande .
linkkiMellersta Österbottens Familjerådgivningscentral :
familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
familjerådgivningfinska _ svenska
skilsmässa
skilsmässa kan sökas av kvinnan , av mannen eller av båda makarna tillsammans .
man ansöker om skilsmässa i tingsrätten .
till att börja med görs en skriftlig skilsmässoansökan .
Österbottens tingsrätt Karleby kansli
Besöksadress : Karlebygatan 27 , 67100 Karleby
telefon : 029.56.49294
Läs mer : skilsmässa .
hälsovårdaren på barnrådgivningsbyrån ger råd i frågor som gäller små barns hälsa , tillväxt och utveckling .
barnrådgivningsbyrån ger information om platser som erbjuder hjälp vid behov .
vid problem hos unga i skolåldern hjälper exempelvis skolans hälsovårdare eller skolkuratorn .
Läs mer : barns och ungas problem .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Skolhälsovårdfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Barnrådgivningarfinska _ svenska
du kan ta upp problem med hälsovårdaren på skolan eller studieplatsen eller vuxna på ungdomsgården .
mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats .
föräldrar eller unga själva kan kontakta familjerådgivningen .
där kan man tala om problem och få hjälp och stöd .
mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats .
Familjerådgivningens telefonnummer : 044.730.7640 .
Läs mer : barns och ungas problem .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Studerandehälsovårdfinska _ svenska
ungdomsgårdar och -lokaler finska _ svenska
problem med den mentala hälsan
om du behöver hjälp och stöd för din mentala hälsa kan du boka en läkartid vid hälsostationen .
läkaren bedömer situationen .
vid behov skriver läkaren en remiss till psykiatrisk specialsjukvård .
Läs mer : mental hälsa .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Mentalvårdstjänsterfinska _ svenska
om du har ekonomiska problem kan du be om råd hos Mellersta Österbottens social- och hälsovårdssamkommun Soites enheter för socialarbete eller utkomststöd , tfn 040.806.5095 eller tjänstestyrningen , tfn 040.806.5093 .
om du har problem med skulder , kontakta rättshjälpsbyrån .
du kan anlita vilken som helst rättshjälpsbyrå oberoende av din hemkommun .
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
telefon : 029.566.1270
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Servicehandledningfinska _ svenska
missbruksproblem
om du har problem med alkohol , droger , läkemedel eller hasardspel kan du få vård och rehabilitering vid Porten , Mellersta Österbottens social- och hälsovårdssamkommun Soites center för missbruksproblem .
du kan ta upp problemet med proffs inom hälsovården eller företagshälsovården , som kan slussa dig vidare i vårdsystemet , eller direkt kontakta Soites missbrukstjänster , tfn 040.8068.101 .
för tillnyktrings- och avgiftningsvård debiteras en patientavgift liksom även för korttidsrehabilitering , öppen rehabilitering är gratis .
även Karleby evangelisk @-@ lutherska församlingssammanslutnings specialdiakoner erbjuder samtalshjälp vid missbruksproblem .
kontaktuppgifter
Hälsovägen 4
67200 Karleby
telefon : 040.806.8101
Läs mer : missbruksproblem .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Service för missbrukarefinska _ svenska
linkkiKarleby evangelisk @-@ lutherska församlingssammansutning :
Karleby evangelisk @-@ lutherska församlings arbete bland missbrukarefinska _ svenska
problem med uppehållstillstånd
brott
våld
diskriminering och rasism
behöver du en jurist ?
Död
problem i äktenskap eller parförhållande
skilsmässa
problem med den mentala hälsan
missbruksproblem
i en krissituation kan du ringa nödcentralen på numret 112 .
de slussar vid behov dig vidare till socialjouren .
du ska endast ringa nödcentralen i brådskande nödsituationer , där liv , egendom eller miljön är i fara .
problem med uppehållstillstånd
om du har problem eller oklarheter med ditt uppehållstillstånd kan du kontakta Migrationsverket .
Migrationsverket
Korsholmsesplanaden 45
Vasa
Läs mer : problem med uppehållstillstånd .
brott
om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112 .
ring inte nödnumret om det inte är fråga om en nödsituation .
du kan göra en polisanmälan på nätet .
mer information finns på Polisens webbplats .
du kan även skriva ut anmälningsblanketten på nätet och lämna in den till polisstationen .
Karleby polisstation
Karlebygatan 74
67100 Karleby
Läs mer : brott .
tidsbokningfinska _ svenska _ engelska
Polisamälanfinska _ svenska _ engelska
våld
om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112 .
Läs mer : våld .
diskriminering och rasism
om du misstänker att du blivit utsatt för diskriminering då du sökt arbete eller på arbetsplatsen ska du först ta upp detta på din arbetsplats .
om saken inte kan lösas på arbetsplatsen ska du kontakta arbetarskyddet vid Regionförvaltningsverket i Västra och Inre Finland .
Besöksadress :
Regionförvaltningsverket i Västra och Inre Finland
Wollfskavägen 35
65101 Vasa
telefon : 0295.018.450
om du utsätts för diskriminering kan du be om hjälp av Diskrimineringsombudsmannen .
om du fallit offer för ett rasistiskt motiverat brott kan du göra en polisanmälan på nätet eller polisstationen .
Läs mer : diskriminering och rasism .
linkkiRegionförvaltningsverket i Västra och Inre Finland :
Regionförvaltningsverket i Västra och Inre Finlandfinska _ svenska _ engelska
hjälp och information för personer som drabbats av etnisk diskrimineringfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
behöver du en jurist ?
juridiska tjänster är avgiftsbelagda men om du har små eller medelstora inkomster , kan du få helt eller delvis avgiftsfri rättshjälp från statens rättshjälpsbyrå .
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
Besöksadress : Ämbetshuset , Torggatan 40 , 67100 Karleby
telefon : 029.566.1270
information om enskilda jurister finns bland annat på Finlands Advokatförbunds webbplats .
Läs mer :
behöver du en jurist ?
linkkiFinlands advokatförbund :
Finlands advokatförbundfinska _ svenska _ engelska
Död
den evangelisk @-@ lutherska kyrkans församlingars begravningsplatser fungerar som allmänna begravningsplatser .
där kan även avlidna som inte är medlemmar i kyrkan begravas .
de är alltså avsedda för alla invånare i staden .
mer information finns på Karleby kyrkliga samfällighets webbplats .
om en närstående plötsligt dör kan du söka krishjälp vid din egen hälsostation , eller utanför tjänstetid vid samjouren för Mellersta Österbottens centralsjukhus .
de evangelisk @-@ lutherska församlingarna i Karlebynejden erbjuder även sorggrupper .
även församlingarnas diakonimottagningar erbjuder samtalshjälp för sorgearbetet .
Läs mer : Död .
linkkiKarleby kyrkliga samfällighet :
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Hälsostationernafinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
problem i äktenskap eller parförhållande
vid problem i äktenskap eller parförhållande får du hjälp av Mellersta Österbottens familjerådgivningscentral som underhålls av Karleby kyrkliga samfällighets och Mellersta Österbottens social- och hälsovårdssamkommun Soites familjerådgivning .
Familjerågivningscentralen
telefon : 050.3147.464 .
Karleby familjerådgivning
67100 Karleby
tel . 044.730.7640
Läs mer : problem i äktenskap eller parförhållande .
linkkiMellersta Österbottens Familjerådgivningscentral :
familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
familjerådgivningfinska _ svenska
skilsmässa
skilsmässa kan sökas av kvinnan , av mannen eller av båda makarna tillsammans .
man ansöker om skilsmässa i tingsrätten .
till att börja med görs en skriftlig skilsmässoansökan .
Österbottens tingsrätt Karleby kansli
Besöksadress : Karlebygatan 27 , 67100 Karleby
telefon : 029.56.49294
Läs mer : skilsmässa .
hälsovårdaren på barnrådgivningsbyrån ger råd i frågor som gäller små barns hälsa , tillväxt och utveckling .
barnrådgivningsbyrån ger information om platser som erbjuder hjälp vid behov .
vid problem hos unga i skolåldern hjälper exempelvis skolans hälsovårdare eller skolkuratorn .
Läs mer : barns och ungas problem .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Skolhälsovårdfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Barnrådgivningarfinska _ svenska
du kan ta upp problem med hälsovårdaren på skolan eller studieplatsen eller vuxna på ungdomsgården .
mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats .
föräldrar eller unga själva kan kontakta familjerådgivningen .
där kan man tala om problem och få hjälp och stöd .
mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats .
Familjerådgivningens telefonnummer : 044.730.7640 .
Läs mer : barns och ungas problem .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Studerandehälsovårdfinska _ svenska
ungdomsgårdar och -lokaler finska _ svenska
problem med den mentala hälsan
om du behöver hjälp och stöd för din mentala hälsa kan du boka en läkartid vid hälsostationen .
läkaren bedömer situationen .
vid behov skriver läkaren en remiss till psykiatrisk specialsjukvård .
Läs mer : mental hälsa .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Mentalvårdstjänsterfinska _ svenska
om du har ekonomiska problem kan du be om råd hos Mellersta Österbottens social- och hälsovårdssamkommun Soites enheter för socialarbete eller utkomststöd , tfn 040.806.5095 eller tjänstestyrningen , tfn 040.806.5093 .
om du har problem med skulder , kontakta rättshjälpsbyrån .
du kan anlita vilken som helst rättshjälpsbyrå oberoende av din hemkommun .
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
telefon : 029.566.1270
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Servicehandledningfinska _ svenska
missbruksproblem
om du har problem med alkohol , droger , läkemedel eller hasardspel kan du få vård och rehabilitering vid Porten , Mellersta Österbottens social- och hälsovårdssamkommun Soites center för missbruksproblem .
du kan ta upp problemet med proffs inom hälsovården eller företagshälsovården , som kan slussa dig vidare i vårdsystemet , eller direkt kontakta Soites missbrukstjänster , tfn 040.8068.101 .
för tillnyktrings- och avgiftningsvård debiteras en patientavgift liksom även för korttidsrehabilitering , öppen rehabilitering är gratis .
även Karleby evangelisk @-@ lutherska församlingssammanslutnings specialdiakoner erbjuder samtalshjälp vid missbruksproblem .
kontaktuppgifter
Hälsovägen 4
67200 Karleby
telefon : 040.806.8101
Läs mer : missbruksproblem .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Service för missbrukarefinska _ svenska
linkkiKarleby evangelisk @-@ lutherska församlingssammansutning :
Karleby evangelisk @-@ lutherska församlings arbete bland missbrukarefinska _ svenska
äktenskap
skilsmässa
barn vid skilsmässa
när du väntar barn
vård av barnet
vård av barnet i hemmet
äktenskap
innan äktenskapet ingås ska du skriftligen be om prövning av äktenskapshinder .
Prövningen görs vid magistraten . du kan lämna in ansökan om prövning vid vilken magistrat som helst .
Civilvigsel äger rum vid magistraten .
magistraten i Västra Finland
Karleby enhet
Karlebygatan 27 , PB 581
67701 Karleby
telefon : 029.553.9451
Läs mer :
äktenskap .
skilsmässa
skilsmässa kan sökas av kvinnan , av mannen eller av båda makarna tillsammans .
man ansöker om skilsmässa i tingsrätten .
till att börja med görs en skriftlig skilsmässoansökan .
Österbottens tingsrätt Karleby kansli
Besöksadress : Karlebygatan 27 , 67100 Karleby
telefon : 029.56.49294
Läs mer : skilsmässa .
barn vid skilsmässa
om du har barn och går igenom en skilsmässa ska du ta kontakt med barnatillsyningsmannen .
barnatillsyningsmannen bekräftar överenskommelsen om var barnen ska bo , vården av barnen , umgängesrätt och underhållsbidrag .
barnatillsyningsmannen
67100 Karleby
Telefontid och tidsbokning
tel . 06.826.4111
Läs mer : barn vid skilsmässa .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Barnatillsyningsmannenfinska _ svenska
när du väntar barn
ta kontakt med rådgivningen då du märker att du är gravid .
på rådgivningen följer man med moderns , barnets och hela familjens välmående under graviditeten .
du kan be om råd per telefon ( 06 ) 826.4477 .
Läs mer :
när du väntar barn .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Mödrarådgivningfinska _ svenska
vård av barnet
i Karleby finns stadens daghem , gruppfamiljedaghem , familjedagvårdare samt barnklubbar .
dessutom finns det daghem som köptjänst ( svenskspråkiga ) , ett privat daghem och privata familjedagvårdare i Karleby .
du kan ansöka om plats inom småbarnspedagogiken för ditt barn elektroniskt via tjänsten suomi.fi eller med en blankett på stadens webbplats ( ansökan om småbarnspedagogik ) .
ansökan ska lämnas in fyra månader innan du behöver plats inom småbarnspedagogiken .
det är möjligt att få en plats snabbare om den behövs för att du exempelvis erhållit arbete eller studieplats .
ansökan kan returneras till platsen för småbarnspedagogik , kontorstjänster för småbarnspedagogik eller lämnas i brevlådan i den nedre aulan i Bildningscentralen .
du kan ansöka om en plats i stadens barnklubbar med blanketten som finns på stadens webbplats .
ansökan kan även skickas per post till följande adress :
Bildningscentralen
tjänster för småbarnspedagogik
Strandgatan16
67100 Karleby
Läs mer :
daghem och andra dagvårdsplatserfinska _ svenska
Gruppfamiljedaghemfinska _ svenska
Dagvårdsblanketterfinska _ svenska
att ansöka om kommunal dagvårdfinska _ svenska
vård av barnet i hemmet
om familjens yngsta barn är yngre än tre år kan föräldern få hemvårdsstöd för vård av barnet i hemmet .
om du har rätt till stödet kan du ansöka om stödet hos FPA .
du kan fylla i ansökan på nätet eller skicka den per post till FPA .
du kan även besöka FPA:s kontor .
Karleby stad betalar extra Karlebystöd för de familjer som tar hand om barn under tre år i hemmet .
du kan ansöka om Karlebystödet om den ena av föräldrarna vårdar samtliga av familjens barn under skolåldern i hemmet .
om din familj fyller villkoren , beviljas Karlebystödet i samband med beviljandet av vårdnadsbidraget .
Läs mer :
stöd för vård av barn i hemmet .
Karlebystödfinska _ svenska
information om FPA:s hemvårdsstödfinska _ svenska _ engelska
FPA kontaktuppgifterfinska _ svenska _ engelska
äktenskap
skilsmässa
barn vid skilsmässa
när du väntar barn
vård av barnet
vård av barnet i hemmet
äktenskap
innan äktenskapet ingås ska du skriftligen be om prövning av äktenskapshinder .
Prövningen görs vid magistraten . du kan lämna in ansökan om prövning vid vilken magistrat som helst .
Civilvigsel äger rum vid magistraten .
magistraten i Västra Finland
Karleby enhet
Karlebygatan 27 , PB 581
67701 Karleby
telefon : 029.553.9451
Läs mer :
äktenskap .
skilsmässa
skilsmässa kan sökas av kvinnan , av mannen eller av båda makarna tillsammans .
man ansöker om skilsmässa i tingsrätten .
till att börja med görs en skriftlig skilsmässoansökan .
Österbottens tingsrätt Karleby kansli
Besöksadress : Karlebygatan 27 , 67100 Karleby
telefon : 029.56.49294
Läs mer : skilsmässa .
barn vid skilsmässa
om du har barn och går igenom en skilsmässa ska du ta kontakt med barnatillsyningsmannen .
barnatillsyningsmannen bekräftar överenskommelsen om var barnen ska bo , vården av barnen , umgängesrätt och underhållsbidrag .
barnatillsyningsmannen
67100 Karleby
Telefontid och tidsbokning
tel . 06.826.4111
Läs mer : barn vid skilsmässa .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Barnatillsyningsmannenfinska _ svenska
när du väntar barn
ta kontakt med rådgivningen då du märker att du är gravid .
på rådgivningen följer man med moderns , barnets och hela familjens välmående under graviditeten .
du kan be om råd per telefon ( 06 ) 826.4477 .
Läs mer :
när du väntar barn .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Mödrarådgivningfinska _ svenska
vård av barnet
i Karleby finns stadens daghem , gruppfamiljedaghem , familjedagvårdare samt barnklubbar .
dessutom finns det daghem som köptjänst ( svenskspråkiga ) , ett privat daghem och privata familjedagvårdare i Karleby .
du kan ansöka om plats inom småbarnspedagogiken för ditt barn elektroniskt via tjänsten suomi.fi eller med en blankett på stadens webbplats ( ansökan om småbarnspedagogik ) .
ansökan ska lämnas in fyra månader innan du behöver plats inom småbarnspedagogiken .
det är möjligt att få en plats snabbare om den behövs för att du exempelvis erhållit arbete eller studieplats .
ansökan kan returneras till platsen för småbarnspedagogik , kontorstjänster för småbarnspedagogik eller lämnas i brevlådan i den nedre aulan i Bildningscentralen .
du kan ansöka om en plats i stadens barnklubbar med blanketten som finns på stadens webbplats .
ansökan kan även skickas per post till följande adress :
Bildningscentralen
tjänster för småbarnspedagogik
Strandgatan16
67100 Karleby
Läs mer :
daghem och andra dagvårdsplatserfinska _ svenska
Gruppfamiljedaghemfinska _ svenska
Dagvårdsblanketterfinska _ svenska
att ansöka om kommunal dagvårdfinska _ svenska
vård av barnet i hemmet
om familjens yngsta barn är yngre än tre år kan föräldern få hemvårdsstöd för vård av barnet i hemmet .
om du har rätt till stödet kan du ansöka om stödet hos FPA .
du kan fylla i ansökan på nätet eller skicka den per post till FPA .
du kan även besöka FPA:s kontor .
Karleby stad betalar extra Karlebystöd för de familjer som tar hand om barn under tre år i hemmet .
du kan ansöka om Karlebystödet om den ena av föräldrarna vårdar samtliga av familjens barn under skolåldern i hemmet .
om din familj fyller villkoren , beviljas Karlebystödet i samband med beviljandet av vårdnadsbidraget .
Läs mer :
stöd för vård av barn i hemmet .
Karlebystödfinska _ svenska
information om FPA:s hemvårdsstödfinska _ svenska _ engelska
FPA kontaktuppgifterfinska _ svenska _ engelska
äktenskap
skilsmässa
barn vid skilsmässa
när du väntar barn
vård av barnet
vård av barnet i hemmet
äktenskap
innan äktenskapet ingås ska du skriftligen be om prövning av äktenskapshinder .
Prövningen görs vid magistraten . du kan lämna in ansökan om prövning vid vilken magistrat som helst .
Civilvigsel äger rum vid magistraten .
magistraten i Västra Finland
Karleby enhet
Karlebygatan 27 , PB 581
67701 Karleby
telefon : 029.553.9451
Läs mer :
äktenskap .
skilsmässa
skilsmässa kan sökas av kvinnan , av mannen eller av båda makarna tillsammans .
man ansöker om skilsmässa i tingsrätten .
till att börja med görs en skriftlig skilsmässoansökan .
Österbottens tingsrätt Karleby kansli
Besöksadress : Karlebygatan 27 , 67100 Karleby
telefon : 029.56.49294
Läs mer : skilsmässa .
barn vid skilsmässa
om du har barn och går igenom en skilsmässa ska du ta kontakt med barnatillsyningsmannen .
barnatillsyningsmannen bekräftar överenskommelsen om var barnen ska bo , vården av barnen , umgängesrätt och underhållsbidrag .
barnatillsyningsmannen
67100 Karleby
Telefontid och tidsbokning
tel . 06.826.4111
Läs mer : barn vid skilsmässa .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Barnatillsyningsmannenfinska _ svenska
när du väntar barn
ta kontakt med rådgivningen då du märker att du är gravid .
på rådgivningen följer man med moderns , barnets och hela familjens välmående under graviditeten .
du kan be om råd per telefon ( 06 ) 826.4477 .
Läs mer : graviditet och förlossning .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Mödrarådgivningfinska _ svenska
vård av barnet
i Karleby finns stadens daghem , gruppfamiljedaghem , familjedagvårdare samt barnklubbar .
dessutom finns det daghem som köptjänst ( svenskspråkiga ) , ett privat daghem och privata familjedagvårdare i Karleby .
du kan ansöka om plats inom småbarnspedagogiken för ditt barn elektroniskt via tjänsten suomi.fi eller med en blankett på stadens webbplats ( ansökan om småbarnspedagogik ) .
ansökan ska lämnas in fyra månader innan du behöver plats inom småbarnspedagogiken .
det är möjligt att få en plats snabbare om den behövs för att du exempelvis erhållit arbete eller studieplats .
ansökan kan returneras till platsen för småbarnspedagogik , kontorstjänster för småbarnspedagogik eller lämnas i brevlådan i den nedre aulan i Bildningscentralen .
du kan ansöka om en plats i stadens barnklubbar med blanketten som finns på stadens webbplats .
ansökan kan även skickas per post till följande adress :
Bildningscentralen
tjänster för småbarnspedagogik
Strandgatan16
67100 Karleby
Läs mer :
vård av barnet .
daghem och andra dagvårdsplatserfinska _ svenska
Gruppfamiljedaghemfinska _ svenska
Dagvårdsblanketterfinska _ svenska
att ansöka om kommunal dagvårdfinska _ svenska
vård av barnet i hemmet
om familjens yngsta barn är yngre än tre år kan föräldern få hemvårdsstöd för vård av barnet i hemmet .
om du har rätt till stödet kan du ansöka om stödet hos FPA .
du kan fylla i ansökan på nätet eller skicka den per post till FPA .
du kan även besöka FPA:s kontor .
Karleby stad betalar extra Karlebystöd för de familjer som tar hand om barn under tre år i hemmet .
du kan ansöka om Karlebystödet om den ena av föräldrarna vårdar samtliga av familjens barn under skolåldern i hemmet .
om din familj fyller villkoren , beviljas Karlebystödet i samband med beviljandet av vårdnadsbidraget .
Läs mer :
stöd för vård av barn i hemmet .
Karlebystödfinska _ svenska
information om FPA:s hemvårdsstödfinska _ svenska _ engelska
FPA kontaktuppgifterfinska _ svenska _ engelska
hälsovårdstjänster i Karleby
äldre människors hälsa
tandvård
mental hälsa
sexuell hälsa
när du väntar barn
förlossning
läkemedel
handikappade personer
ett handikappat barn
hälsovårdstjänster i Karleby
i Karleby finns hälsostationer i olika delar av staden .
varje hälsostation har ett eget telefonnummer för tidsbokning , som man kan ringa för att boka tid till sjukskötare eller läkare .
kontaktuppgifter :
Karleby huvudhälsostation
Mariegatan 28
67200 Karleby
telefon : ( 06 ) 8287.580
på Karleby huvudhälsostationen styrs patienterna till mottagningen på basis av hur akuta deras symptom är .
Klienten får en tid till akutvården , mottagningen eller Min Soite @-@ mottagningen .
samtal till huvudhälsostationen styrs till ett och samma telefonnummer , ( 06 ) 8287.310 .
67800 Karleby
telefon : ( 06 ) 8287.580
mottagning / Kelviå
Ellfolkgatan 5
68300 Kelviå
telefon : ( 06 ) 8287.701
mottagning / Lochteå
telefon : ( 06 ) 8287.750
mottagning / Ullava
Ullavavägen 701
68370 Ullava
telefon : ( 06 ) 8287.639
om du kommer som flykting till Finland ska du komma överens om en hälsokontroll med Utlänningsbyrån .
Läs mer : hälsa .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Hälsostationernafinska _ svenska
under kvällar och helger är hälsostationerna stängda .
då hanteras plötsliga sjukdomar och olyckor vid jouren .
jouren är avsedd för patienter vars sjukdom kräver brådskande bedömning och vård .
i livshotande situationer ska du ringa nödnumret 112 .
om du besöker jouren kvällstid eller under helger ska du först ringa jourens telefonrådgivning ( 06 ) 826.4500 .
Samjourens adress :
Mellersta Österbottens centralsjukhus
Mariegatan 16 @-@ 20 ( l @-@ flygeln , ingång B1 )
67200 Karleby
Läs mer : hälsovårdstjänster i Finland
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
barns hälsa
om ditt barn insjuknar ska du kontakta hälsostationen vid behov .
ådgivningarna erbjuder tjänster för gravida och barn under skolåldern .
vid rådgivningarna utförs vaccinationer av barn och vuxna .
du kan kontakta rådgivningen via den centraliserade telefontjänsten ( 06 ) 826.4477 .
genom regelbundna besök på barnrådgivningsbyrån följs barnets hälsa , tillväxt och utveckling upp .
på rådgivningen vårdas inte barn som insjuknar plötsligt , men du kan be om råd via den centraliserade telefontjänsten ( 06 ) 826.4477 .
Skolhälsovårdaren har hand om skolelevers hälsa .
mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats .
Läs mer : barns hälsa .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Barnrådgivningarfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Rådgivningarfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Skolhälsovårdfinska _ svenska
äldre människors hälsa
vid hälsopunkten Daalia ges vägledning och rådgivning för personer över 65 år om diet , motion och livsstil .
Vaccinering av personer över 65 år utförs vid seniorrådgivning .
Läs mer :
äldre människors hälsa .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Seniorernas hälsopunkterfinska _ svenska
tandvård
om du behöver icke @-@ brådskande tandvård ska du ringa munhälsans centraliserade tidsbokningen .
Centraliserad tidsbokning per telefon : ( 06 ) 8287.400
Huvudhälsostationens tandklinik
Mariegatan 28 , 67200 Karleby
Björkhagens tandklinik
Storkisbackens tandklinik
Korpvägen 11 , 67100 Karleby
Kelviå tandklinik
Ellfolkgatan 5 , 68300 , Kelviå
Lochteå tandklinik
Ullava tandklinik
Ullavavägen 701 , 68370 Ullava
vardagar kan tider till smärtjouren bokas enligt överenskommelse vid samtliga tandkliniker .
brådskande tandvård / första hjälpen ( kvälls- , vardags- , helg- och nattjour ) :
vid smärtjouren får du första hjälpen vid plötslig tandvärk och tandolyckor .
Tandläkarjouren ( kvälls- , vardags- och helgjour ) ordnas vid polikliniken för tand- och munsjukdomar vid Mellersta Österbottens social- och hälsovårdssamkommun Soite , Mariegatan 16 @-@ 20 , 67200 Karleby ( vån 1 , del D ) , vardagkvällar kl . 16.00 @-@ 21.00 samt veckoslut och helgdagar kl . 8.00 @-@ 21.00 .
du kan i regel komma till jourmottagningen genom att först kontakta jouren via telefon .
för frågor gällande jouren ring tel . ( 06 ) 828.7450 .
när du kommer till jourmottagningen ska du ta en kölapp , såvida du inte har en bokad tid .
brådskande tandvård / första hjälpen ( nattjour ) :
Allvarliga fall i samjour Uleåborgs universitetssjukhus ( Oulun yliopistollinen sairaala OYS ) kl . 21.00 − 8.00 , tel . ( 08 ) 315.2655
Läs mer : tandvård .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Munhälsovårdenfinska _ svenska
mental hälsa
vid problem med din mentala hälsa ska du i första hand kontakta din egen hälsostation eller företagshälsovårdens mottagning .
vid brådskande problem , kontakta hälsovårdcentralens jour .
Läs mer : mental hälsa .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Hälsostationernafinska _ svenska
sexuell hälsa
om du känner att du behöver information om familjeplanering och prevention kan du kontakta din egen hälsostation .
boka tid till hälsostationen om du behöver preventivmedel , överväger att göra en abort eller misstänker att du lider av en könssjukdom .
du kan även boka en tid hos en allmänläkare för en gynekologisk eller urologisk undersökning .
i preventionsfrågor kan du kontakta den centraliserade telefontjänsten ( 06 ) 826.4477 .
Läs mer :
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Hälsostationernafinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Preventivrådgivningfinska _ svenska
när du väntar barn
ta kontakt med rådgivningen då du märker att du är gravid .
på rådgivningen följer man med moderns , barnets och hela familjens välmående under graviditeten .
Läs mer :
när du väntar barn .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Mödrarådgivningfinska _ svenska
förlossning
förlossningsavdelningen är öppen dygnet runt .
om du önskar kan du ringa förlossningsavdelning då din förlossning satt igång eller om du vill fråga om råd .
då du kommer till sjukhuset ska du använda centralsjukhusets huvudingång kl . 7 @-@ 20 och övriga tider bör du använda den gemensamma jourens / poliklinikens dörr .
kontaktuppgifter för förlossningsavdelningen :
Mariegatan 16 @-@ 20 ,
67200 Karleby
telefon : ( 06 ) 8264355 .
Läs mer : förlossning .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Förlossningarfinska _ svenska
läkemedel
du kan köpa läkemedel på apoteket .
du kan besöka vilket apotek som helst .
du kan även besöka apotek som inte finns i din egen kommun .
Läs mer : läkemedel .
handikappade personer
en handikappad person bosatt i Karleby har rätt att erhålla de tjänster han eller hon behöver på samma grunder som de övriga invånarna i kommunen .
Personen kan dock på grund av sitt handikapp eller sin sjukdom även behöva särskilda tjänster för handikappade för att klara vardagen .
för tjänsterna för handikappade i Karleby svarar Mellersta Österbottens social- och hälsovårdssamkommun Soite , där man kan ansöka om tjänster och stödfunktioner .
tjänster av flera olika slag erbjuds även för personer med gravt handikapp .
dessa tjänster inkluderar bland annat :
transporttjänster
ombyggnad och nödvändig utrustning för hemmet
maskiner och utrustning
personlig hjälp och dagverksamhet
stödboende
stöd för närståendevård av personer under 65 och arbetsverksamhet .
dessutom är det möjligt att ansöka om specialboende , korttidsvård eller tillfällig vård samt handledning hos den öppna vården .
mer information om tjänster för handikappade får du från Mellersta Österbottens social- och hälsovårdssamkommun Soites handikapptjänster per telefon : 040.804.2122 .
Läs mer : handikappade personer .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
tjänster för handikappadefinska _ svenska
Specialpedagogik i förskolanfinska _ svenska
kontaktuppgifter för den grundläggande utbildningenfinska
ett handikappat barn
särskilt stöd erbjuds barn med handikapp inom småbarnspedagogiken och skolan .
kontakta Karleby stads förskoleundervisning för information om specialsmåbarnspedagogiken .
du kan be undervisningsväsendet om mer information om tjänster som skolan erbjuder .
Bildningscentralen
Strandgatan 16 ( våning 5 och 6 )
67100 Karleby
telefon : 040.8065.149
Läs mer : ett handikappat barn .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
tjänster för handikappadefinska _ svenska
Specialpedagogik i förskolanfinska _ svenska
kontaktuppgifter för den grundläggande utbildningenfinska
hälsovårdstjänster i Karleby
äldre människors hälsa
tandvård
mental hälsa
sexuell hälsa
när du väntar barn
förlossning
läkemedel
handikappade personer
ett handikappat barn
hälsovårdstjänster i Karleby
i Karleby finns hälsostationer i olika delar av staden .
varje hälsostation har ett eget telefonnummer för tidsbokning , som man kan ringa för att boka tid till sjukskötare eller läkare .
kontaktuppgifter :
Karleby huvudhälsostation
Mariegatan 28
67200 Karleby
telefon : ( 06 ) 8287.580
på Karleby huvudhälsostationen styrs patienterna till mottagningen på basis av hur akuta deras symptom är .
Klienten får en tid till akutvården , mottagningen eller Min Soite @-@ mottagningen .
samtal till huvudhälsostationen styrs till ett och samma telefonnummer , ( 06 ) 8287.310 .
67800 Karleby
telefon : ( 06 ) 8287.580
mottagning / Kelviå
Ellfolkgatan 5
68300 Kelviå
telefon : ( 06 ) 8287.701
mottagning / Lochteå
telefon : ( 06 ) 8287.750
mottagning / Ullava
Ullavavägen 701
68370 Ullava
telefon : ( 06 ) 8287.639
om du kommer som flykting till Finland ska du komma överens om en hälsokontroll med Utlänningsbyrån .
Läs mer : hälsa .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Hälsostationernafinska _ svenska
under kvällar och helger är hälsostationerna stängda .
då hanteras plötsliga sjukdomar och olyckor vid jouren .
jouren är avsedd för patienter vars sjukdom kräver brådskande bedömning och vård .
i livshotande situationer ska du ringa nödnumret 112 .
om du besöker jouren kvällstid eller under helger ska du först ringa jourens telefonrådgivning ( 06 ) 826.4500 .
Samjourens adress :
Mellersta Österbottens centralsjukhus
Mariegatan 16 @-@ 20 ( l @-@ flygeln , ingång B1 )
67200 Karleby
Läs mer : hälsovårdstjänster i Finland
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
barns hälsa
om ditt barn insjuknar ska du kontakta hälsostationen vid behov .
ådgivningarna erbjuder tjänster för gravida och barn under skolåldern .
vid rådgivningarna utförs vaccinationer av barn och vuxna .
du kan kontakta rådgivningen via den centraliserade telefontjänsten ( 06 ) 826.4477 .
genom regelbundna besök på barnrådgivningsbyrån följs barnets hälsa , tillväxt och utveckling upp .
på rådgivningen vårdas inte barn som insjuknar plötsligt , men du kan be om råd via den centraliserade telefontjänsten ( 06 ) 826.4477 .
Skolhälsovårdaren har hand om skolelevers hälsa .
mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats .
Läs mer : barns hälsa .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Barnrådgivningarfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Rådgivningarfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Skolhälsovårdfinska _ svenska
äldre människors hälsa
vid hälsopunkten Daalia ges vägledning och rådgivning för personer över 65 år om diet , motion och livsstil .
Vaccinering av personer över 65 år utförs vid seniorrådgivning .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Seniorernas hälsopunkterfinska _ svenska
tandvård
om du behöver icke @-@ brådskande tandvård ska du ringa munhälsans centraliserade tidsbokningen .
Centraliserad tidsbokning per telefon : ( 06 ) 8287.400
Huvudhälsostationens tandklinik
Mariegatan 28 , 67200 Karleby
Björkhagens tandklinik
Storkisbackens tandklinik
Korpvägen 11 , 67100 Karleby
Kelviå tandklinik
Ellfolkgatan 5 , 68300 , Kelviå
Lochteå tandklinik
Ullava tandklinik
Ullavavägen 701 , 68370 Ullava
vardagar kan tider till smärtjouren bokas enligt överenskommelse vid samtliga tandkliniker .
brådskande tandvård / första hjälpen ( kvälls- , vardags- , helg- och nattjour ) :
vid smärtjouren får du första hjälpen vid plötslig tandvärk och tandolyckor .
Tandläkarjouren ( kvälls- , vardags- och helgjour ) ordnas vid polikliniken för tand- och munsjukdomar vid Mellersta Österbottens social- och hälsovårdssamkommun Soite , Mariegatan 16 @-@ 20 , 67200 Karleby ( vån 1 , del D ) , vardagkvällar kl . 16.00 @-@ 21.00 samt veckoslut och helgdagar kl . 8.00 @-@ 21.00 .
du kan i regel komma till jourmottagningen genom att först kontakta jouren via telefon .
för frågor gällande jouren ring tel . ( 06 ) 828.7450 .
när du kommer till jourmottagningen ska du ta en kölapp , såvida du inte har en bokad tid .
brådskande tandvård / första hjälpen ( nattjour ) :
Allvarliga fall i samjour Uleåborgs universitetssjukhus ( Oulun yliopistollinen sairaala OYS ) kl . 21.00 − 8.00 , tel . ( 08 ) 315.2655
Läs mer : tandvård .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Munhälsovårdenfinska _ svenska
mental hälsa
vid problem med din mentala hälsa ska du i första hand kontakta din egen hälsostation eller företagshälsovårdens mottagning .
vid brådskande problem , kontakta hälsovårdcentralens jour .
Läs mer : mental hälsa .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Hälsostationernafinska _ svenska
sexuell hälsa
om du känner att du behöver information om familjeplanering och prevention kan du kontakta din egen hälsostation .
boka tid till hälsostationen om du behöver preventivmedel , överväger att göra en abort eller misstänker att du lider av en könssjukdom .
du kan även boka en tid hos en allmänläkare för en gynekologisk eller urologisk undersökning .
i preventionsfrågor kan du kontakta den centraliserade telefontjänsten ( 06 ) 826.4477 .
Läs mer :
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Hälsostationernafinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Preventivrådgivningfinska _ svenska
när du väntar barn
ta kontakt med rådgivningen då du märker att du är gravid .
på rådgivningen följer man med moderns , barnets och hela familjens välmående under graviditeten .
Läs mer :
när du väntar barn .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Mödrarådgivningfinska _ svenska
förlossning
förlossningsavdelningen är öppen dygnet runt .
om du önskar kan du ringa förlossningsavdelning då din förlossning satt igång eller om du vill fråga om råd .
då du kommer till sjukhuset ska du använda centralsjukhusets huvudingång kl . 7 @-@ 20 och övriga tider bör du använda den gemensamma jourens / poliklinikens dörr .
kontaktuppgifter för förlossningsavdelningen :
Mariegatan 16 @-@ 20 ,
67200 Karleby
telefon : ( 06 ) 8264355 .
Läs mer : förlossning .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Förlossningarfinska _ svenska
läkemedel
du kan köpa läkemedel på apoteket .
du kan besöka vilket apotek som helst .
du kan även besöka apotek som inte finns i din egen kommun .
Läs mer : läkemedel .
handikappade personer
en handikappad person bosatt i Karleby har rätt att erhålla de tjänster han eller hon behöver på samma grunder som de övriga invånarna i kommunen .
Personen kan dock på grund av sitt handikapp eller sin sjukdom även behöva särskilda tjänster för handikappade för att klara vardagen .
för tjänsterna för handikappade i Karleby svarar Mellersta Österbottens social- och hälsovårdssamkommun Soite , där man kan ansöka om tjänster och stödfunktioner .
tjänster av flera olika slag erbjuds även för personer med gravt handikapp .
dessa tjänster inkluderar bland annat :
transporttjänster
ombyggnad och nödvändig utrustning för hemmet
maskiner och utrustning
personlig hjälp och dagverksamhet
stödboende
stöd för närståendevård av personer under 65 och arbetsverksamhet .
dessutom är det möjligt att ansöka om specialboende , korttidsvård eller tillfällig vård samt handledning hos den öppna vården .
mer information om tjänster för handikappade får du från Mellersta Österbottens social- och hälsovårdssamkommun Soites handikapptjänster per telefon : 040.804.2122 .
Läs mer : handikappade personer .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
tjänster för handikappadefinska _ svenska
Specialpedagogik i förskolanfinska _ svenska
kontaktuppgifter för den grundläggande utbildningenfinska
ett handikappat barn
särskilt stöd erbjuds barn med handikapp inom småbarnspedagogiken och skolan .
kontakta Karleby stads förskoleundervisning för information om specialsmåbarnspedagogiken .
du kan be undervisningsväsendet om mer information om tjänster som skolan erbjuder .
Bildningscentralen
Strandgatan 16 ( våning 5 och 6 )
67100 Karleby
telefon : 040.8065.149
Läs mer : ett handikappat barn .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
tjänster för handikappadefinska _ svenska
Specialpedagogik i förskolanfinska _ svenska
kontaktuppgifter för den grundläggande utbildningenfinska
hälsovårdstjänster i Karleby
äldre människors hälsa
tandvård
mental hälsa
sexuell hälsa
när du väntar barn
förlossning
läkemedel
handikappade personer
ett handikappat barn
hälsovårdstjänster i Karleby
i Karleby finns hälsostationer i olika delar av staden .
varje hälsostation har ett eget telefonnummer för tidsbokning , som man kan ringa för att boka tid till sjukskötare eller läkare .
kontaktuppgifter :
Karleby huvudhälsostation
Mariegatan 28
67200 Karleby
telefon : ( 06 ) 8287.580
på Karleby huvudhälsostationen styrs patienterna till mottagningen på basis av hur akuta deras symptom är .
Klienten får en tid till akutvården , mottagningen eller Min Soite @-@ mottagningen .
samtal till huvudhälsostationen styrs till ett och samma telefonnummer , ( 06 ) 8287.310 .
67800 Karleby
telefon : ( 06 ) 8287.580
mottagning / Kelviå
Ellfolkgatan 5
68300 Kelviå
telefon : ( 06 ) 8287.701
mottagning / Lochteå
telefon : ( 06 ) 8287.750
mottagning / Ullava
Ullavavägen 701
68370 Ullava
telefon : ( 06 ) 8287.639
om du kommer som flykting till Finland ska du komma överens om en hälsokontroll med Utlänningsbyrån .
Läs mer : hälsa .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Hälsostationernafinska _ svenska
under kvällar och helger är hälsostationerna stängda .
då hanteras plötsliga sjukdomar och olyckor vid jouren .
jouren är avsedd för patienter vars sjukdom kräver brådskande bedömning och vård .
i livshotande situationer ska du ringa nödnumret 112 .
om du besöker jouren kvällstid eller under helger ska du först ringa jourens telefonrådgivning ( 06 ) 826.4500 .
Samjourens adress :
Mellersta Österbottens centralsjukhus
Mariegatan 16 @-@ 20 ( l @-@ flygeln , ingång B1 )
67200 Karleby
Läs mer : hälsovårdstjänster i Finland
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
barns hälsa
om ditt barn insjuknar ska du kontakta hälsostationen vid behov .
ådgivningarna erbjuder tjänster för gravida och barn under skolåldern .
vid rådgivningarna utförs vaccinationer av barn och vuxna .
du kan kontakta rådgivningen via den centraliserade telefontjänsten ( 06 ) 826.4477 .
genom regelbundna besök på barnrådgivningsbyrån följs barnets hälsa , tillväxt och utveckling upp .
på rådgivningen vårdas inte barn som insjuknar plötsligt , men du kan be om råd via den centraliserade telefontjänsten ( 06 ) 826.4477 .
Skolhälsovårdaren har hand om skolelevers hälsa .
mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats .
Läs mer : barns hälsa .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Barnrådgivningarfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Rådgivningarfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Skolhälsovårdfinska _ svenska
äldre människors hälsa
vid hälsopunkten Daalia ges vägledning och rådgivning för personer över 65 år om diet , motion och livsstil .
Vaccinering av personer över 65 år utförs vid seniorrådgivning .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Seniorernas hälsopunkterfinska _ svenska
tandvård
om du behöver icke @-@ brådskande tandvård ska du ringa munhälsans centraliserade tidsbokningen .
Centraliserad tidsbokning per telefon : ( 06 ) 8287.400
Huvudhälsostationens tandklinik
Mariegatan 28 , 67200 Karleby
Björkhagens tandklinik
Storkisbackens tandklinik
Korpvägen 11 , 67100 Karleby
Kelviå tandklinik
Ellfolkgatan 5 , 68300 , Kelviå
Lochteå tandklinik
Ullava tandklinik
Ullavavägen 701 , 68370 Ullava
vardagar kan tider till smärtjouren bokas enligt överenskommelse vid samtliga tandkliniker .
brådskande tandvård / första hjälpen ( kvälls- , vardags- , helg- och nattjour ) :
vid smärtjouren får du första hjälpen vid plötslig tandvärk och tandolyckor .
Tandläkarjouren ( kvälls- , vardags- och helgjour ) ordnas vid polikliniken för tand- och munsjukdomar vid Mellersta Österbottens social- och hälsovårdssamkommun Soite , Mariegatan 16 @-@ 20 , 67200 Karleby ( vån 1 , del D ) , vardagkvällar kl . 16.00 @-@ 21.00 samt veckoslut och helgdagar kl . 8.00 @-@ 21.00 .
du kan i regel komma till jourmottagningen genom att först kontakta jouren via telefon .
för frågor gällande jouren ring tel . ( 06 ) 828.7450 .
när du kommer till jourmottagningen ska du ta en kölapp , såvida du inte har en bokad tid .
brådskande tandvård / första hjälpen ( nattjour ) :
Allvarliga fall i samjour Uleåborgs universitetssjukhus ( Oulun yliopistollinen sairaala OYS ) kl . 21.00 − 8.00 , tel . ( 08 ) 315.2655
Läs mer : tandvård .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Munhälsovårdenfinska _ svenska
mental hälsa
vid problem med din mentala hälsa ska du i första hand kontakta din egen hälsostation eller företagshälsovårdens mottagning .
vid brådskande problem , kontakta hälsovårdcentralens jour .
Läs mer : mental hälsa .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Hälsostationernafinska _ svenska
sexuell hälsa
om du känner att du behöver information om familjeplanering och prevention kan du kontakta din egen hälsostation .
boka tid till hälsostationen om du behöver preventivmedel , överväger att göra en abort eller misstänker att du lider av en könssjukdom .
du kan även boka en tid hos en allmänläkare för en gynekologisk eller urologisk undersökning .
i preventionsfrågor kan du kontakta den centraliserade telefontjänsten ( 06 ) 826.4477 .
Läs mer :
sexuell hälsa och prevention .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Hälsostationernafinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Preventivrådgivningfinska _ svenska
när du väntar barn
ta kontakt med rådgivningen då du märker att du är gravid .
på rådgivningen följer man med moderns , barnets och hela familjens välmående under graviditeten .
Läs mer : graviditet och förlossning .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Mödrarådgivningfinska _ svenska
förlossning
förlossningsavdelningen är öppen dygnet runt .
om du önskar kan du ringa förlossningsavdelning då din förlossning satt igång eller om du vill fråga om råd .
då du kommer till sjukhuset ska du använda centralsjukhusets huvudingång kl . 7 @-@ 20 och övriga tider bör du använda den gemensamma jourens / poliklinikens dörr .
kontaktuppgifter för förlossningsavdelningen :
Mariegatan 16 @-@ 20 ,
67200 Karleby
telefon : ( 06 ) 8264355 .
Läs mer : graviditet och förlossning .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Förlossningarfinska _ svenska
läkemedel
du kan köpa läkemedel på apoteket .
du kan besöka vilket apotek som helst .
du kan även besöka apotek som inte finns i din egen kommun .
Läs mer : läkemedel .
handikappade personer
en handikappad person bosatt i Karleby har rätt att erhålla de tjänster han eller hon behöver på samma grunder som de övriga invånarna i kommunen .
Personen kan dock på grund av sitt handikapp eller sin sjukdom även behöva särskilda tjänster för handikappade för att klara vardagen .
för tjänsterna för handikappade i Karleby svarar Mellersta Österbottens social- och hälsovårdssamkommun Soite , där man kan ansöka om tjänster och stödfunktioner .
tjänster av flera olika slag erbjuds även för personer med gravt handikapp .
dessa tjänster inkluderar bland annat :
transporttjänster
ombyggnad och nödvändig utrustning för hemmet
maskiner och utrustning
personlig hjälp och dagverksamhet
stödboende
stöd för närståendevård av personer under 65 och arbetsverksamhet .
dessutom är det möjligt att ansöka om specialboende , korttidsvård eller tillfällig vård samt handledning hos den öppna vården .
mer information om tjänster för handikappade får du från Mellersta Österbottens social- och hälsovårdssamkommun Soites handikapptjänster per telefon : 040.804.2122 .
Läs mer : handikappade personer .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
tjänster för handikappadefinska _ svenska
Specialpedagogik i förskolanfinska _ svenska
kontaktuppgifter för den grundläggande utbildningenfinska
ett handikappat barn
särskilt stöd erbjuds barn med handikapp inom småbarnspedagogiken och skolan .
kontakta Karleby stads förskoleundervisning för information om specialsmåbarnspedagogiken .
du kan be undervisningsväsendet om mer information om tjänster som skolan erbjuder .
Bildningscentralen
Strandgatan 16 ( våning 5 och 6 )
67100 Karleby
telefon : 040.8065.149
Läs mer : ett handikappat barn .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
tjänster för handikappadefinska _ svenska
Specialpedagogik i förskolanfinska _ svenska
kontaktuppgifter för den grundläggande utbildningenfinska
småbarnspedagogik
förskoleundervisning
grundläggande utbildning
undervisning i det egna modersmålet för invandrare
yrkesutbildning
gymnasium
unga utan studieplats
Högskoleutbildning
andra studiemöjligheter
småbarnspedagogik
i Karleby finns stadens egna daghem , gruppfamiljedaghem , familjedagvårdare samt barnklubbar .
dessutom finns det daghem som köptjänst ( svenskspråkiga ) , ett privat daghem och privata familjedagvårdare i Karleby .
du kan ansöka om plats inom småbarnspedagogiken för ditt barn elektroniskt via tjänsten Suomi.fi eller med en blankett på stadens webbplats ( ansökan till småbarnspedagogiken ) .
ansökan ska lämnas in fyra månader innan du behöver plats inom småbarnspedagogiken .
det är möjligt att få en plats snabbare om den behövs för att du exempelvis erhållit arbete eller studieplats .
ansökan kan returneras till platsen för småbarnspedagogik , kontorstjänster för småbarnspedagogik eller lämnas i brevlådan i den nedre aulan i Bildningscentralen .
du kan ansöka om en plats i stadens barnklubbar med blanketten som finns på stadens webbplats .
ansökan kan även skickas per post till följande adress :
Bildningscentralen
tjänster för småbarnspedagogik
Strandgatan16
67100 Karleby
Läs mer :
daghem och andra dagvårdsplatserfinska _ svenska
Gruppfamiljedaghemfinska _ svenska
Dagvårdsblanketterfinska _ svenska
att ansöka om kommunal dagvårdfinska _ svenska
förskoleundervisning
Karleby stad erbjuder gratis förskoleundervisning för alla 6 år fyllda barn .
förskoleundervisningen ges av lärare med utbildning i pedagogik i minst 700 timmar om året , dvs. cirka fyra timmar om dagen , enligt skolans arbetstider .
förskoleundervisningen är gratis .
om barnet dessutom behöver avgiftsbelagd småbarnspedagogisk verksamhet arrangeras denna på samma ställe som förskoleundervisningen , dock med undantag för skiftesvård .
Anmälningar till förskoleundervisningen sker i januari @-@ februari .
detta meddelas i lokaltidningarna och på stadens webbplats .
om du inte fått ett brev om förskoleplats eller ansöker om förskoleplats under annan tid på året , ta kontakt med kontorstjänster för småbarnspedagogik per telefon på numret 040.806.5089 .
Läs mer : förskoleundervisning .
förskoleundervisningfinska _ svenska
grundläggande utbildning
i Finland har alla barn som fyllt 7 år läroplikt , vilket innebär att de måste delta i den grundläggande utbildningen .
Läroplikten upphör i slutet av det läsår då barnet fyller 17 .
det är föräldrarna som har ansvaret för att barnet går i skolan .
anmälan till grundskolan sker i början av året .
på stadens webbplats finns skolornas kontaktuppgifter och mer information om anmälan .
om du har frågor om den grundläggande utbildningen kan du även kontakta stadens undervisningstjänster .
varje barn och ung person har rätt att gå i skola .
om barnet flyttar till Karleby under läsåret kan han eller hon genast börja i skolan .
om barnet saknar tillräckliga färdigheter i finska eller svenska för att delta i undervisningen i klassen inleder han eller hon studierna i förberedande undervisning i en egen grupp eller i klassen enligt det egna studieprogrammet .
i Karleby finns grupper för den förberedande utbildningen i lågstadiet i Hollihaan koulu och Koivuhaan koulu och i högstadiet i Stenängens skola .
Övergången till den vanliga undervisningen sker steg för steg enligt elevens förutsättningar .
undervisning i enlighet med lärokursen finska som andra språk och litteratur stödjer en helhetsmässig utveckling av språket .
stöd för lärande arrangeras i mån av möjlighet på elevens eget modersmål i skolan .
mer information om den förberedande undervisningen för invandrare får du av stadens undervisningstjänster .
Läs mer : grundläggande utbildning .
kontaktuppgifter för den grundläggande utbildningenfinska
undervisning i det egna modersmålet för invandrare
undervisning i elevens eget modersmål arrangeras i Karleby på flera olika språk , till exempel under läsåret 2017 @-@ 2018 arrangerades undervisning på nio olika språk .
Undervisningsgruppen ska ha minst fyra elever .
undervisningen sker vanligtvis i de skolor där det finns flest elever som talar språket i fråga .
som elevens egen religion undervisas bland annat islam , buddhism och ortodox religion , beroende på antalet elever .
information om undervisning i elevens eget modersmål och religion får du av koordinatoren för undervisningen för olika språk- och kulturgrupper :
tfn 040.489.2129
utbildning för invandrarefinska
yrkesutbildning
Mellersta Österbottens yrkesinstitut erbjuder yrkesutbildning i Karleby , Kelviå , Kannus , Kaustby , Perho och Jakobstad .
yrkesinstitutet anordnar även handledande utbildning för grundläggande yrkesutbildning , dvs . VALMA @-@ utbildning samt förberedande utbildningar för vuxna invandrare vid Mellersta Österbottens folkhögskola i Kelviå .
Läs mer : yrkesutbildning .
linkkiMellersta Österbottens utbildningskoncern :
Mellersta Österbottens utbildningskoncernfinska _ engelska
linkkiMellersta Österbottens utbildningskoncern :
utbildning för invandrarefinska _ engelska
linkkiMellersta Österbottens folkhögskola :
Folkhögskolans invandrarlinjefinska
gymnasium
i Karleby ges gymnasieutbildning för ungdomar vid Karleby finska gymnasium och Karleby svenska gymnasium , samt för vuxna vid Karleby vuxengymnasium .
till gymnasieutbildning för ungdomar ansöker man under våren via gemensam ansökning för gymnasierna och man kan bli antagen om man i slutbetyget från grundskolan har tillräckligt högt snittbetyg i läsämnena .
du kan ansöka till vuxenutbildningen direkt hos vuxengymnasiet året runt .
Karleby finska gymnasium erbjuder förberedande undervisning för gymnasiet även för invandrare .
den förberedande undervisningen för gymnasiet är ett läsår och målet med den är att förbättra möjligheterna för elever med ett annat modersmål att klara av gymnasiestudierna .
varje år fattas ett skilt beslut om undervisningens start .
för varje studerande utarbetas ett eget studieprogram .
man ansöker till förberedande undervisning för gymnasiet under sommaren på webbsidan Opintopolku.fi .
Undervisningsspråket i vid Karleby finska gymnasium och Karleby vuxengymnasium är finska och svenska vid Karleby svenska gymnasium .
vid Karleby finska gymnasium anordnas undervisning i finska som andraspråk för invandrare invandrare .
målet är att invandrarna ska klara av gymnasiestudierna och efter gymnasiet kunna söka sig till fortsatta studier .
mer information om gymnasieskolorna och den förberedande undervisningen för gymnasiet fås av stadens undervisningstjänster .
kontaktuppgifterna för gymnasierna finns på stadens undervisningstjänsters webbplats .
Bildningscentralen
Strandgatan 16 ( våning 5 och 6 )
67100 Karleby
telefon : 044.756.7673
Läs mer :
gymnasium .
Gymnasie- och yrkesutbildningfinska _ svenska
unga utan studieplats
unga som saknar studieplats eller arbete kan få hjälp av det uppsökande ungdomsarbetet .
det uppsökande ungdomsarbetet hjälper unga i åldern 15 @-@ 28 år hitta rätt tjänster till stöd för utbildning , arbete och utkomst .
de anställda inom uppsökande ungdomsarbete hjälper med att klara upp den ungas livssituation , hantera praktiska ärenden , såsom besök hos olika myndigheter , och ger personlig handledning enligt den ungas önskemål .
uppsökande ungdomsarbetefinska _ svenska
Högskoleutbildning
vid Centria yrkeshögskola kan man avlägga högskoleexamen i teknik , företagsekonomi , social- och hälsovård .
man kan även avlägga en examen inom musikpedagogik och samhällspedagogik .
det är dessutom möjligt att studera vid den öppna yrkeshögskolan .
vid Karleby universitetscenter Chydenius kan man avlägga såväl högre högskoleexamen som doktorsexamen .
vid Chydenius anordnas även vuxenutbildning och vetenskaplig forskning bedrivs .
Läs mer : Högskoleutbildning .
Högskole- och universitetsutbildningfinska
linkkiCentria yrkeshögskola :
Centria yrkeshögskolafinska _ svenska _ engelska
Universitetscentret Chydeniusfinska _ svenska _ engelska
andra studiemöjligheter
Karlebynejdens institut , som ägs och drivs av Karleby stad , är ett tvåspråkigt ( finska och svenska ) medborgarinstitut .
institutet erbjuder undervisning i datateknik , musik , idrott och dans , konstämnen , hantverk , matlagning och första hjälpen .
institutet erbjuder även undervisning i flera olika språk , bland annat finska , svenska , engelska , tyska , franska , ryska , spanska och italienska .
Undervisningsutbudet varierar från år till år , så det lönar sig att kontrollera aktuella kurser på institutets webbplats .
invandrare ges rabatt på vissa kurser .
i kursuppgifterna anges om det är möjligt att få rabatt på kursen .
kontrollera på institutets webbplats vilka kurser som är aktuella .
Vasavägen 7
67100 Karleby
telefon : 040.8065.169 , 040.8065.168
vid Mellersta Österbottens sommaruniversitet kan du läsa kurser på universitetsnivå vid det öppna universitetet , delta i kompletterande yrkesutbildning samt läsa språk- och kulturkurser .
under sommaren är det möjligt att repetera gymnasiestudier vid sommaruniversitetet .
dessutom är det även möjligt att läsa normala gymnasiekurser vid sommaruniversitetets sommargymnasium .
Sommaruniversitets kurser är avgiftsbelagda för deltagarna .
Läs mer :
studier som hobby , Arbetskraftsutbildning
Karlebynejdens institutfinska _ svenska
linkkiArbets- och näringsbyråns tjänster :
offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiMellersta Österbottens sommaruniversitet :
Mellersta Österbottens sommaruniversitetfinska
övrig undervisning i Karlebyfinska _ svenska
småbarnspedagogik
förskoleundervisning
grundläggande utbildning
undervisning i det egna modersmålet för invandrare
yrkesutbildning
gymnasium
unga utan studieplats
Högskoleutbildning
andra studiemöjligheter
småbarnspedagogik
i Karleby finns stadens egna daghem , gruppfamiljedaghem , familjedagvårdare samt barnklubbar .
dessutom finns det daghem som köptjänst ( svenskspråkiga ) , ett privat daghem och privata familjedagvårdare i Karleby .
du kan ansöka om plats inom småbarnspedagogiken för ditt barn elektroniskt via tjänsten Suomi.fi eller med en blankett på stadens webbplats ( ansökan till småbarnspedagogiken ) .
ansökan ska lämnas in fyra månader innan du behöver plats inom småbarnspedagogiken .
det är möjligt att få en plats snabbare om den behövs för att du exempelvis erhållit arbete eller studieplats .
ansökan kan returneras till platsen för småbarnspedagogik , kontorstjänster för småbarnspedagogik eller lämnas i brevlådan i den nedre aulan i Bildningscentralen .
du kan ansöka om en plats i stadens barnklubbar med blanketten som finns på stadens webbplats .
ansökan kan även skickas per post till följande adress :
Bildningscentralen
tjänster för småbarnspedagogik
Strandgatan16
67100 Karleby
Läs mer :
daghem och andra dagvårdsplatserfinska _ svenska
Gruppfamiljedaghemfinska _ svenska
Dagvårdsblanketterfinska _ svenska
att ansöka om kommunal dagvårdfinska _ svenska
förskoleundervisning
Karleby stad erbjuder gratis förskoleundervisning för alla 6 år fyllda barn .
förskoleundervisningen ges av lärare med utbildning i pedagogik i minst 700 timmar om året , dvs. cirka fyra timmar om dagen , enligt skolans arbetstider .
förskoleundervisningen är gratis .
om barnet dessutom behöver avgiftsbelagd småbarnspedagogisk verksamhet arrangeras denna på samma ställe som förskoleundervisningen , dock med undantag för skiftesvård .
Anmälningar till förskoleundervisningen sker i januari @-@ februari .
detta meddelas i lokaltidningarna och på stadens webbplats .
om du inte fått ett brev om förskoleplats eller ansöker om förskoleplats under annan tid på året , ta kontakt med kontorstjänster för småbarnspedagogik per telefon på numret 040.806.5089 .
Läs mer : förskoleundervisning .
förskoleundervisningfinska _ svenska
grundläggande utbildning
i Finland har alla barn som fyllt 7 år läroplikt , vilket innebär att de måste delta i den grundläggande utbildningen .
Läroplikten upphör i slutet av det läsår då barnet fyller 17 .
det är föräldrarna som har ansvaret för att barnet går i skolan .
anmälan till grundskolan sker i början av året .
på stadens webbplats finns skolornas kontaktuppgifter och mer information om anmälan .
om du har frågor om den grundläggande utbildningen kan du även kontakta stadens undervisningstjänster .
varje barn och ung person har rätt att gå i skola .
om barnet flyttar till Karleby under läsåret kan han eller hon genast börja i skolan .
om barnet saknar tillräckliga färdigheter i finska eller svenska för att delta i undervisningen i klassen inleder han eller hon studierna i förberedande undervisning i en egen grupp eller i klassen enligt det egna studieprogrammet .
i Karleby finns grupper för den förberedande utbildningen i lågstadiet i Hollihaan koulu och Koivuhaan koulu och i högstadiet i Stenängens skola .
Övergången till den vanliga undervisningen sker steg för steg enligt elevens förutsättningar .
undervisning i enlighet med lärokursen finska som andra språk och litteratur stödjer en helhetsmässig utveckling av språket .
stöd för lärande arrangeras i mån av möjlighet på elevens eget modersmål i skolan .
mer information om den förberedande undervisningen för invandrare får du av stadens undervisningstjänster .
Läs mer : grundläggande utbildning .
kontaktuppgifter för den grundläggande utbildningenfinska
undervisning i det egna modersmålet för invandrare
undervisning i elevens eget modersmål arrangeras i Karleby på flera olika språk , till exempel under läsåret 2017 @-@ 2018 arrangerades undervisning på nio olika språk .
Undervisningsgruppen ska ha minst fyra elever .
undervisningen sker vanligtvis i de skolor där det finns flest elever som talar språket i fråga .
som elevens egen religion undervisas bland annat islam , buddhism och ortodox religion , beroende på antalet elever .
information om undervisning i elevens eget modersmål och religion får du av koordinatoren för undervisningen för olika språk- och kulturgrupper :
tfn 040.489.2129
utbildning för invandrarefinska
yrkesutbildning
Mellersta Österbottens yrkesinstitut erbjuder yrkesutbildning i Karleby , Kelviå , Kannus , Kaustby , Perho och Jakobstad .
yrkesinstitutet anordnar även handledande utbildning för grundläggande yrkesutbildning , dvs . VALMA @-@ utbildning samt förberedande utbildningar för vuxna invandrare vid Mellersta Österbottens folkhögskola i Kelviå .
Läs mer : yrkesutbildning .
linkkiMellersta Österbottens utbildningskoncern :
Mellersta Österbottens utbildningskoncernfinska _ engelska
linkkiMellersta Österbottens utbildningskoncern :
utbildning för invandrarefinska _ engelska
linkkiMellersta Österbottens folkhögskola :
Folkhögskolans invandrarlinjefinska
gymnasium
i Karleby ges gymnasieutbildning för ungdomar vid Karleby finska gymnasium och Karleby svenska gymnasium , samt för vuxna vid Karleby vuxengymnasium .
till gymnasieutbildning för ungdomar ansöker man under våren via gemensam ansökning för gymnasierna och man kan bli antagen om man i slutbetyget från grundskolan har tillräckligt högt snittbetyg i läsämnena .
du kan ansöka till vuxenutbildningen direkt hos vuxengymnasiet året runt .
Karleby finska gymnasium erbjuder förberedande undervisning för gymnasiet även för invandrare .
den förberedande undervisningen för gymnasiet är ett läsår och målet med den är att förbättra möjligheterna för elever med ett annat modersmål att klara av gymnasiestudierna .
varje år fattas ett skilt beslut om undervisningens start .
för varje studerande utarbetas ett eget studieprogram .
man ansöker till förberedande undervisning för gymnasiet under sommaren på webbsidan Opintopolku.fi .
Undervisningsspråket i vid Karleby finska gymnasium och Karleby vuxengymnasium är finska och svenska vid Karleby svenska gymnasium .
vid Karleby finska gymnasium anordnas undervisning i finska som andraspråk för invandrare invandrare .
målet är att invandrarna ska klara av gymnasiestudierna och efter gymnasiet kunna söka sig till fortsatta studier .
mer information om gymnasieskolorna och den förberedande undervisningen för gymnasiet fås av stadens undervisningstjänster .
kontaktuppgifterna för gymnasierna finns på stadens undervisningstjänsters webbplats .
Bildningscentralen
Strandgatan 16 ( våning 5 och 6 )
67100 Karleby
telefon : 044.756.7673
Läs mer :
gymnasium .
Gymnasie- och yrkesutbildningfinska _ svenska
unga utan studieplats
unga som saknar studieplats eller arbete kan få hjälp av det uppsökande ungdomsarbetet .
det uppsökande ungdomsarbetet hjälper unga i åldern 15 @-@ 28 år hitta rätt tjänster till stöd för utbildning , arbete och utkomst .
de anställda inom uppsökande ungdomsarbete hjälper med att klara upp den ungas livssituation , hantera praktiska ärenden , såsom besök hos olika myndigheter , och ger personlig handledning enligt den ungas önskemål .
uppsökande ungdomsarbetefinska _ svenska
Högskoleutbildning
vid Centria yrkeshögskola kan man avlägga högskoleexamen i teknik , företagsekonomi , social- och hälsovård .
man kan även avlägga en examen inom musikpedagogik och samhällspedagogik .
det är dessutom möjligt att studera vid den öppna yrkeshögskolan .
vid Karleby universitetscenter Chydenius kan man avlägga såväl högre högskoleexamen som doktorsexamen .
vid Chydenius anordnas även vuxenutbildning och vetenskaplig forskning bedrivs .
Läs mer : Högskoleutbildning .
Högskole- och universitetsutbildningfinska
linkkiCentria yrkeshögskola :
Centria yrkeshögskolafinska _ svenska _ engelska
Universitetscentret Chydeniusfinska _ svenska _ engelska
andra studiemöjligheter
Karlebynejdens institut , som ägs och drivs av Karleby stad , är ett tvåspråkigt ( finska och svenska ) medborgarinstitut .
institutet erbjuder undervisning i datateknik , musik , idrott och dans , konstämnen , hantverk , matlagning och första hjälpen .
institutet erbjuder även undervisning i flera olika språk , bland annat finska , svenska , engelska , tyska , franska , ryska , spanska och italienska .
Undervisningsutbudet varierar från år till år , så det lönar sig att kontrollera aktuella kurser på institutets webbplats .
invandrare ges rabatt på vissa kurser .
i kursuppgifterna anges om det är möjligt att få rabatt på kursen .
kontrollera på institutets webbplats vilka kurser som är aktuella .
Vasavägen 7
67100 Karleby
telefon : 040.8065.169 , 040.8065.168
vid Mellersta Österbottens sommaruniversitet kan du läsa kurser på universitetsnivå vid det öppna universitetet , delta i kompletterande yrkesutbildning samt läsa språk- och kulturkurser .
under sommaren är det möjligt att repetera gymnasiestudier vid sommaruniversitetet .
dessutom är det även möjligt att läsa normala gymnasiekurser vid sommaruniversitetets sommargymnasium .
Sommaruniversitets kurser är avgiftsbelagda för deltagarna .
Läs mer :
studier som hobby , Arbetskraftsutbildning
Karlebynejdens institutfinska _ svenska
linkkiArbets- och näringsbyråns tjänster :
offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiMellersta Österbottens sommaruniversitet :
Mellersta Österbottens sommaruniversitetfinska
övrig undervisning i Karlebyfinska _ svenska
småbarnspedagogik
förskoleundervisning
grundläggande utbildning
undervisning i det egna modersmålet för invandrare
yrkesutbildning
gymnasium
unga utan studieplats
Högskoleutbildning
andra studiemöjligheter
småbarnspedagogik
i Karleby finns stadens egna daghem , gruppfamiljedaghem , familjedagvårdare samt barnklubbar .
dessutom finns det daghem som köptjänst ( svenskspråkiga ) , ett privat daghem och privata familjedagvårdare i Karleby .
du kan ansöka om plats inom småbarnspedagogiken för ditt barn elektroniskt via tjänsten Suomi.fi eller med en blankett på stadens webbplats ( ansökan till småbarnspedagogiken ) .
ansökan ska lämnas in fyra månader innan du behöver plats inom småbarnspedagogiken .
det är möjligt att få en plats snabbare om den behövs för att du exempelvis erhållit arbete eller studieplats .
ansökan kan returneras till platsen för småbarnspedagogik , kontorstjänster för småbarnspedagogik eller lämnas i brevlådan i den nedre aulan i Bildningscentralen .
du kan ansöka om en plats i stadens barnklubbar med blanketten som finns på stadens webbplats .
ansökan kan även skickas per post till följande adress :
Bildningscentralen
tjänster för småbarnspedagogik
Strandgatan16
67100 Karleby
Läs mer :
småbarnspedagogik .
daghem och andra dagvårdsplatserfinska _ svenska
Gruppfamiljedaghemfinska _ svenska
Dagvårdsblanketterfinska _ svenska
att ansöka om kommunal dagvårdfinska _ svenska
förskoleundervisning
Karleby stad erbjuder gratis förskoleundervisning för alla 6 år fyllda barn .
förskoleundervisningen ges av lärare med utbildning i pedagogik i minst 700 timmar om året , dvs. cirka fyra timmar om dagen , enligt skolans arbetstider .
förskoleundervisningen är gratis .
om barnet dessutom behöver avgiftsbelagd småbarnspedagogisk verksamhet arrangeras denna på samma ställe som förskoleundervisningen , dock med undantag för skiftesvård .
Anmälningar till förskoleundervisningen sker i januari @-@ februari .
detta meddelas i lokaltidningarna och på stadens webbplats .
om du inte fått ett brev om förskoleplats eller ansöker om förskoleplats under annan tid på året , ta kontakt med kontorstjänster för småbarnspedagogik per telefon på numret 040.806.5089 .
Läs mer : förskoleundervisning .
förskoleundervisningfinska _ svenska
grundläggande utbildning
i Finland har alla barn som fyllt 7 år läroplikt , vilket innebär att de måste delta i den grundläggande utbildningen .
Läroplikten upphör i slutet av det läsår då barnet fyller 17 .
det är föräldrarna som har ansvaret för att barnet går i skolan .
anmälan till grundskolan sker i början av året .
på stadens webbplats finns skolornas kontaktuppgifter och mer information om anmälan .
om du har frågor om den grundläggande utbildningen kan du även kontakta stadens undervisningstjänster .
varje barn och ung person har rätt att gå i skola .
om barnet flyttar till Karleby under läsåret kan han eller hon genast börja i skolan .
om barnet saknar tillräckliga färdigheter i finska eller svenska för att delta i undervisningen i klassen inleder han eller hon studierna i förberedande undervisning i en egen grupp eller i klassen enligt det egna studieprogrammet .
i Karleby finns grupper för den förberedande utbildningen i lågstadiet i Hollihaan koulu och Koivuhaan koulu och i högstadiet i Stenängens skola .
Övergången till den vanliga undervisningen sker steg för steg enligt elevens förutsättningar .
undervisning i enlighet med lärokursen finska som andra språk och litteratur stödjer en helhetsmässig utveckling av språket .
stöd för lärande arrangeras i mån av möjlighet på elevens eget modersmål i skolan .
mer information om den förberedande undervisningen för invandrare får du av stadens undervisningstjänster .
Läs mer : grundläggande utbildning .
kontaktuppgifter för den grundläggande utbildningenfinska
undervisning i det egna modersmålet för invandrare
undervisning i elevens eget modersmål arrangeras i Karleby på flera olika språk , till exempel under läsåret 2017 @-@ 2018 arrangerades undervisning på nio olika språk .
Undervisningsgruppen ska ha minst fyra elever .
undervisningen sker vanligtvis i de skolor där det finns flest elever som talar språket i fråga .
som elevens egen religion undervisas bland annat islam , buddhism och ortodox religion , beroende på antalet elever .
information om undervisning i elevens eget modersmål och religion får du av koordinatoren för undervisningen för olika språk- och kulturgrupper :
tfn 040.489.2129
utbildning för invandrarefinska
yrkesutbildning
Mellersta Österbottens yrkesinstitut erbjuder yrkesutbildning i Karleby , Kelviå , Kannus , Kaustby , Perho och Jakobstad .
yrkesinstitutet anordnar även handledande utbildning för grundläggande yrkesutbildning , dvs . VALMA @-@ utbildning samt förberedande utbildningar för vuxna invandrare vid Mellersta Österbottens folkhögskola i Kelviå .
Läs mer : yrkesutbildning .
linkkiMellersta Österbottens utbildningskoncern :
Mellersta Österbottens utbildningskoncernfinska _ engelska
linkkiMellersta Österbottens utbildningskoncern :
utbildning för invandrarefinska _ engelska
linkkiMellersta Österbottens folkhögskola :
Folkhögskolans invandrarlinjefinska
gymnasium
i Karleby ges gymnasieutbildning för ungdomar vid Karleby finska gymnasium och Karleby svenska gymnasium , samt för vuxna vid Karleby vuxengymnasium .
till gymnasieutbildning för ungdomar ansöker man under våren via gemensam ansökning för gymnasierna och man kan bli antagen om man i slutbetyget från grundskolan har tillräckligt högt snittbetyg i läsämnena .
du kan ansöka till vuxenutbildningen direkt hos vuxengymnasiet året runt .
Karleby finska gymnasium erbjuder förberedande undervisning för gymnasiet även för invandrare .
den förberedande undervisningen för gymnasiet är ett läsår och målet med den är att förbättra möjligheterna för elever med ett annat modersmål att klara av gymnasiestudierna .
varje år fattas ett skilt beslut om undervisningens start .
för varje studerande utarbetas ett eget studieprogram .
man ansöker till förberedande undervisning för gymnasiet under sommaren på webbsidan Opintopolku.fi .
Undervisningsspråket i vid Karleby finska gymnasium och Karleby vuxengymnasium är finska och svenska vid Karleby svenska gymnasium .
vid Karleby finska gymnasium anordnas undervisning i finska som andraspråk för invandrare invandrare .
målet är att invandrarna ska klara av gymnasiestudierna och efter gymnasiet kunna söka sig till fortsatta studier .
mer information om gymnasieskolorna och den förberedande undervisningen för gymnasiet fås av stadens undervisningstjänster .
kontaktuppgifterna för gymnasierna finns på stadens undervisningstjänsters webbplats .
Bildningscentralen
Strandgatan 16 ( våning 5 och 6 )
67100 Karleby
telefon : 044.756.7673
Läs mer :
gymnasium .
Gymnasie- och yrkesutbildningfinska _ svenska
unga utan studieplats
unga som saknar studieplats eller arbete kan få hjälp av det uppsökande ungdomsarbetet .
det uppsökande ungdomsarbetet hjälper unga i åldern 15 @-@ 28 år hitta rätt tjänster till stöd för utbildning , arbete och utkomst .
de anställda inom uppsökande ungdomsarbete hjälper med att klara upp den ungas livssituation , hantera praktiska ärenden , såsom besök hos olika myndigheter , och ger personlig handledning enligt den ungas önskemål .
uppsökande ungdomsarbetefinska _ svenska
Högskoleutbildning
vid Centria yrkeshögskola kan man avlägga högskoleexamen i teknik , företagsekonomi , social- och hälsovård .
man kan även avlägga en examen inom musikpedagogik och samhällspedagogik .
det är dessutom möjligt att studera vid den öppna yrkeshögskolan .
vid Karleby universitetscenter Chydenius kan man avlägga såväl högre högskoleexamen som doktorsexamen .
vid Chydenius anordnas även vuxenutbildning och vetenskaplig forskning bedrivs .
Läs mer :
yrkeshögskolor , Universitet .
Högskole- och universitetsutbildningfinska
linkkiCentria yrkeshögskola :
Centria yrkeshögskolafinska _ svenska _ engelska
Universitetscentret Chydeniusfinska _ svenska _ engelska
andra studiemöjligheter
Karlebynejdens institut , som ägs och drivs av Karleby stad , är ett tvåspråkigt ( finska och svenska ) medborgarinstitut .
institutet erbjuder undervisning i datateknik , musik , idrott och dans , konstämnen , hantverk , matlagning och första hjälpen .
institutet erbjuder även undervisning i flera olika språk , bland annat finska , svenska , engelska , tyska , franska , ryska , spanska och italienska .
Undervisningsutbudet varierar från år till år , så det lönar sig att kontrollera aktuella kurser på institutets webbplats .
invandrare ges rabatt på vissa kurser .
i kursuppgifterna anges om det är möjligt att få rabatt på kursen .
kontrollera på institutets webbplats vilka kurser som är aktuella .
Vasavägen 7
67100 Karleby
telefon : 040.8065.169 , 040.8065.168
vid Mellersta Österbottens sommaruniversitet kan du läsa kurser på universitetsnivå vid det öppna universitetet , delta i kompletterande yrkesutbildning samt läsa språk- och kulturkurser .
under sommaren är det möjligt att repetera gymnasiestudier vid sommaruniversitetet .
dessutom är det även möjligt att läsa normala gymnasiekurser vid sommaruniversitetets sommargymnasium .
Sommaruniversitets kurser är avgiftsbelagda för deltagarna .
Läs mer :
studier som hobby , Arbetskraftsutbildning
Karlebynejdens institutfinska _ svenska
linkkiArbets- och näringsbyråns tjänster :
offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiMellersta Österbottens sommaruniversitet :
Mellersta Österbottens sommaruniversitetfinska
övrig undervisning i Karlebyfinska _ svenska
hyresbostad
Ägarbostad
tillfälligt boende
Stöd- och serviceboende
Bostadslöshet
avfallshantering för bostaden
hyresbostad
Karleby stads blankett för ansökan om hyresbostad kan fyllas i och skickas in på nätet .
Bilagor till ansökningen ska tillhandahållas då bostad erbjuds , men kan även lämnas in tidigare .
man kan även lämna in bostadsansökan på papper .
Ansökningsblanketterna kan hämtas från och lämnas in till Kokkolan Vuokra Asunnot Oy:s verksamhetsställen .
67800 Karleby
telefon : 040.1817.400
Studiebostäder hyrs ut av Kiinteistöyhtiö Tankkari , som erbjuder möblerade kollektivbostäder samt familjebostäder i olika storlek .
en familjebostad är en omöblerad lägenhet som endast hyrs ut till personer i samma hushåll .
såväl individer som sambor / gifta par kan ansöka om en hyresetta .
Bondegatan 2
67100 Karleby
telefon : 040.193.6468
Läs mer :
hyresbostad .
hyresbostäderfinska _ svenska
ansökan om Karleby stads hyresbostadfinska _ svenska _ engelska
hyresbostäder enligt stadsdelfinska _ svenska
Studiebostäderfinska _ engelska
privata hyresbostäderfinska _ svenska
Ägarbostad
de flesta finländarna bor i en ägarbostad , alltså i en bostad som de själva äger .
på lång sikt är det ofta förmånligare att köpa sin egen bostad än att hyra .
bland annat hos bostadsförmedlingen , på internet och i lokala tidningar finns annonser om bostäder som är till salu .
Läs mer :
Ägarbostad .
tillfälligt boende
i Karlebynejden erbjuds olika inkvarteringsalternativ .
kontaktuppgifterna finns under länkarna nedan .
Läs mer :
tillfälligt boende .
Övernattningsalternativ i Karlebyfinska _ svenska _ engelska
om du saknar boende på grund av kris eller olycka ska du kontakta Kokkolan Vuokra Asunnot Oy eller bostadsbyrån .
om din bostad har skadats , till exempel till följd av brand eller vattenskada , kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna .
kontakta ditt försäkringsbolag direkt när skadan har inträffat .
om en familjemedlem är våldsam eller hotar med våld , ta kontakt med Karleby mödra- och skyddshem .
du kan ringa skyddshemmet under alla tider på dygnet .
du behöver inte uppge ditt namn då du ringer .
Karleby mödra- och skyddshem
telefon : 044.336.0056
hyresbostäderfinska _ svenska
Karleby mödra- och skyddshemfinska
Stöd- och serviceboende
äldre människor erbjuds boendeservice anordnad av Mellersta Österbottens social- och hälsovårdssamkommun Soite samt privata servicebostäder .
serviceboende för äldre är avsett för personer över 65 år som behöver vård och omsorg dygnet runt .
serviceboende är lämpat för personer som inte längre klarar sig på egen hand med tjänster som tillhandahålls i hemmet .
mer information om boendeservice anordnad av Mellersta Österbottens social- och hälsovårdssamkommun Soite får du av bland annat samkommunens servicestyrcentral , tfn 040.806.5093 .
för handikappade och personer som återhämtar sig från mentala problem erbjuds bostäder som beaktar invånarnas särskilda behov .
hemvårdens stödtjänster erbjuds personer som har svårigheter med att klara vardagen utan hjälp , såsom äldre och handikappade personer .
tjänster av detta slag är bland annat måltidstjänst och transporttjänst .
målet med hemvården är att erbjuda trygg vård och omsorg samt främja invånarnas ork , handlingskraft och företagsamhet .
Läs mer :
Stöd- och serviceboende .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Servicehandledningscentretfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Seniorernas tjänster , hemvårdfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Seniorernas tjänster , serviceboendet och anstaltsvårdenfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
boendetjänster för utvecklingsstörda och handikappadefinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Socialrådgivningfinska _ svenska
Bostadslöshet
om du blir bostadslös bör du kontakta Kokkolan Vuokra Asunnot Oy eller bostadsbyrån .
hyresbostäderfinska _ svenska
avfallshantering för bostaden
med bioavfall avses bl.a. :
matrester
skämda och torra livsmedel
skal från frukt och grönsaker
separat insamlat bioavfall packas i en papperspåse , en påse vikt av en dagstidning eller en plastkasse . Kassen eller påsen får vara högst 30l stor .
en full sopsäck ska tillslutas noggrant .
med energiavfall avses bl.a. :
bakplåtspapper , hushållspapper och våtservetter
kläder ( inte skor , regnställ eller läderplagg )
små plastleksaker och bruksföremål i plast såsom disk- och tandborstar .
separat insamlat energiavfall ska packas i plastkasse eller papperspåsar .
Kassen eller påsen får vara högst 30 l stor .
påsen tillsluts noga .
avfall som inte får läggas i det egna husets sopbehållare kan föras till återvinningsstationer .
kontrollera på förhand vilken typ av avfall stationen tar emot .
mer information om avfallshanteringen i Karlebynejden finns på Karleby stads och på Ab Ekorosk Oy:s ( kommunalt avfallshanteringsbolag ) webbplats .
Läs mer : avfallshantering och återvinning .
avfallshantering för bostaden finska _ svenska
ett kommunalt avfallshanteringsbolagfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ vietnamesiska _ polska _ kroatiska
hyresbostad
köpa bostad
tillfälligt boende
Stöd- och serviceboende
Bostadslöshet
avfallshantering för bostaden
hyresbostad
Karleby stads blankett för ansökan om hyresbostad kan fyllas i och skickas in på nätet .
Bilagor till ansökningen ska tillhandahållas då bostad erbjuds , men kan även lämnas in tidigare .
man kan även lämna in bostadsansökan på papper .
Ansökningsblanketterna kan hämtas från och lämnas in till Kokkolan Vuokra Asunnot Oy:s verksamhetsställen .
67800 Karleby
telefon : 040.1817.400
Studiebostäder hyrs ut av Kiinteistöyhtiö Tankkari , som erbjuder möblerade kollektivbostäder samt familjebostäder i olika storlek .
en familjebostad är en omöblerad lägenhet som endast hyrs ut till personer i samma hushåll .
såväl individer som sambor / gifta par kan ansöka om en hyresetta .
Bondegatan 2
67100 Karleby
telefon : 040.193.6468
Läs mer : hyresbostad .
hyresbostäderfinska _ svenska
ansökan om Karleby stads hyresbostadfinska _ svenska _ engelska
hyresbostäder enligt stadsdelfinska _ svenska
Studiebostäderfinska _ engelska
privata hyresbostäderfinska _ svenska
köpa bostad
de flesta finländarna bor i en ägarbostad , alltså i en bostad som de själva äger .
på lång sikt är det ofta förmånligare att köpa sin egen bostad än att hyra .
bland annat hos bostadsförmedlingen , på internet och i lokala tidningar finns annonser om bostäder som är till salu .
Läs mer : köpa bostad .
tillfälligt boende
i Karlebynejden erbjuds olika inkvarteringsalternativ .
kontaktuppgifterna finns under länkarna nedan .
Läs mer :
tillfälligt boende .
Övernattningsalternativ i Karlebyfinska _ svenska _ engelska
om du saknar boende på grund av kris eller olycka ska du kontakta Kokkolan Vuokra Asunnot Oy eller bostadsbyrån .
om din bostad har skadats , till exempel till följd av brand eller vattenskada , kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna .
kontakta ditt försäkringsbolag direkt när skadan har inträffat .
om en familjemedlem är våldsam eller hotar med våld , ta kontakt med Karleby mödra- och skyddshem .
du kan ringa skyddshemmet under alla tider på dygnet .
du behöver inte uppge ditt namn då du ringer .
Karleby mödra- och skyddshem
telefon : 044.336.0056
Läs mer : boende .
hyresbostäderfinska _ svenska
Karleby mödra- och skyddshemfinska
Stöd- och serviceboende
äldre människor erbjuds boendeservice anordnad av Mellersta Österbottens social- och hälsovårdssamkommun Soite samt privata servicebostäder .
serviceboende för äldre är avsett för personer över 65 år som behöver vård och omsorg dygnet runt .
serviceboende är lämpat för personer som inte längre klarar sig på egen hand med tjänster som tillhandahålls i hemmet .
mer information om boendeservice anordnad av Mellersta Österbottens social- och hälsovårdssamkommun Soite får du av bland annat samkommunens servicestyrcentral , tfn 040.806.5093 .
för handikappade och personer som återhämtar sig från mentala problem erbjuds bostäder som beaktar invånarnas särskilda behov .
hemvårdens stödtjänster erbjuds personer som har svårigheter med att klara vardagen utan hjälp , såsom äldre och handikappade personer .
tjänster av detta slag är bland annat måltidstjänst och transporttjänst .
målet med hemvården är att erbjuda trygg vård och omsorg samt främja invånarnas ork , handlingskraft och företagsamhet .
Läs mer :
Stöd- och serviceboende .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Servicehandledningscentretfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Seniorernas tjänster , hemvårdfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Seniorernas tjänster , serviceboendet och anstaltsvårdenfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
boendetjänster för utvecklingsstörda och handikappadefinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Socialrådgivningfinska _ svenska
Bostadslöshet
om du blir bostadslös bör du kontakta Kokkolan Vuokra Asunnot Oy eller bostadsbyrån .
Läs mer : Bostadslöshet .
hyresbostäderfinska _ svenska
avfallshantering för bostaden
med bioavfall avses bl.a. :
matrester
skämda och torra livsmedel
skal från frukt och grönsaker
separat insamlat bioavfall packas i en papperspåse , en påse vikt av en dagstidning eller en plastkasse . Kassen eller påsen får vara högst 30l stor .
en full sopsäck ska tillslutas noggrant .
med energiavfall avses bl.a. :
bakplåtspapper , hushållspapper och våtservetter
kläder ( inte skor , regnställ eller läderplagg )
små plastleksaker och bruksföremål i plast såsom disk- och tandborstar .
separat insamlat energiavfall ska packas i plastkasse eller papperspåsar .
Kassen eller påsen får vara högst 30 l stor .
påsen tillsluts noga .
avfall som inte får läggas i det egna husets sopbehållare kan föras till återvinningsstationer .
kontrollera på förhand vilken typ av avfall stationen tar emot .
mer information om avfallshanteringen i Karlebynejden finns på Karleby stads och på Ab Ekorosk Oy:s ( kommunalt avfallshanteringsbolag ) webbplats .
Läs mer : avfallshantering och återvinning .
avfallshantering för bostaden finska _ svenska
ett kommunalt avfallshanteringsbolagfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ vietnamesiska _ polska _ kroatiska
hyresbostad
köpa bostad
tillfälligt boende
Stöd- och serviceboende
Bostadslöshet
avfallshantering för bostaden
hyresbostad
Karleby stads blankett för ansökan om hyresbostad kan fyllas i och skickas in på nätet .
Bilagor till ansökningen ska tillhandahållas då bostad erbjuds , men kan även lämnas in tidigare .
man kan även lämna in bostadsansökan på papper .
Ansökningsblanketterna kan hämtas från och lämnas in till Kokkolan Vuokra Asunnot Oy:s verksamhetsställen .
67800 Karleby
telefon : 040.1817.400
Studiebostäder hyrs ut av Kiinteistöyhtiö Tankkari , som erbjuder möblerade kollektivbostäder samt familjebostäder i olika storlek .
en familjebostad är en omöblerad lägenhet som endast hyrs ut till personer i samma hushåll .
såväl individer som sambor / gifta par kan ansöka om en hyresetta .
Bondegatan 2
67100 Karleby
telefon : 040.193.6468
Läs mer : hyresbostad .
hyresbostäderfinska _ svenska
ansökan om Karleby stads hyresbostadfinska _ svenska _ engelska
hyresbostäder enligt stadsdelfinska _ svenska
Studiebostäderfinska _ engelska
privata hyresbostäderfinska _ svenska
köpa bostad
de flesta finländarna bor i en ägarbostad , alltså i en bostad som de själva äger .
på lång sikt är det ofta förmånligare att köpa sin egen bostad än att hyra .
bland annat hos bostadsförmedlingen , på internet och i lokala tidningar finns annonser om bostäder som är till salu .
Läs mer : köpa bostad .
tillfälligt boende
i Karlebynejden erbjuds olika inkvarteringsalternativ .
kontaktuppgifterna finns under länkarna nedan .
Läs mer :
tillfälligt boende .
Övernattningsalternativ i Karlebyfinska _ svenska _ engelska
om du saknar boende på grund av kris eller olycka ska du kontakta Kokkolan Vuokra Asunnot Oy eller bostadsbyrån .
om din bostad har skadats , till exempel till följd av brand eller vattenskada , kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna .
kontakta ditt försäkringsbolag direkt när skadan har inträffat .
om en familjemedlem är våldsam eller hotar med våld , ta kontakt med Karleby mödra- och skyddshem .
du kan ringa skyddshemmet under alla tider på dygnet .
du behöver inte uppge ditt namn då du ringer .
Karleby mödra- och skyddshem
telefon : 044.336.0056
Läs mer : boende .
hyresbostäderfinska _ svenska
Karleby mödra- och skyddshemfinska
Stöd- och serviceboende
äldre människor erbjuds boendeservice anordnad av Mellersta Österbottens social- och hälsovårdssamkommun Soite samt privata servicebostäder .
serviceboende för äldre är avsett för personer över 65 år som behöver vård och omsorg dygnet runt .
serviceboende är lämpat för personer som inte längre klarar sig på egen hand med tjänster som tillhandahålls i hemmet .
mer information om boendeservice anordnad av Mellersta Österbottens social- och hälsovårdssamkommun Soite får du av bland annat samkommunens servicestyrcentral , tfn 040.806.5093 .
för handikappade och personer som återhämtar sig från mentala problem erbjuds bostäder som beaktar invånarnas särskilda behov .
hemvårdens stödtjänster erbjuds personer som har svårigheter med att klara vardagen utan hjälp , såsom äldre och handikappade personer .
tjänster av detta slag är bland annat måltidstjänst och transporttjänst .
målet med hemvården är att erbjuda trygg vård och omsorg samt främja invånarnas ork , handlingskraft och företagsamhet .
Läs mer :
Stöd- och serviceboende .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Servicehandledningscentretfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Seniorernas tjänster , hemvårdfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Seniorernas tjänster , serviceboendet och anstaltsvårdenfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
boendetjänster för utvecklingsstörda och handikappadefinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Socialrådgivningfinska _ svenska
Bostadslöshet
om du blir bostadslös bör du kontakta Kokkolan Vuokra Asunnot Oy eller bostadsbyrån .
Läs mer : Bostadslöshet .
hyresbostäderfinska _ svenska
avfallshantering för bostaden
med bioavfall avses bl.a. :
matrester
skämda och torra livsmedel
skal från frukt och grönsaker
separat insamlat bioavfall packas i en papperspåse , en påse vikt av en dagstidning eller en plastkasse . Kassen eller påsen får vara högst 30l stor .
en full sopsäck ska tillslutas noggrant .
med energiavfall avses bl.a. :
bakplåtspapper , hushållspapper och våtservetter
kläder ( inte skor , regnställ eller läderplagg )
små plastleksaker och bruksföremål i plast såsom disk- och tandborstar .
separat insamlat energiavfall ska packas i plastkasse eller papperspåsar .
Kassen eller påsen får vara högst 30 l stor .
påsen tillsluts noga .
avfall som inte får läggas i det egna husets sopbehållare kan föras till återvinningsstationer .
kontrollera på förhand vilken typ av avfall stationen tar emot .
mer information om avfallshanteringen i Karlebynejden finns på Karleby stads och på Ab Ekorosk Oy:s ( kommunalt avfallshanteringsbolag ) webbplats .
Läs mer : avfallshantering och återvinning .
avfallshantering för bostaden finska _ svenska
ett kommunalt avfallshanteringsbolagfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ vietnamesiska _ polska _ kroatiska
möjligheter att studera finska eller svenska
Karlebynejdens institut erbjuder undervisning i finska och svenska från grundnivå .
Mellersta Österbottens utbildningskoncern erbjuder kurser i finska vid Mellersta Österbottens folkhögskola i Kelviå inom utbildningen i läs- och skrivfärdigheter och den förberedande utbildningen för vuxna invandrare . det går också att studera finska inom utbildningen som handleder för yrkesutbildning ( VALMA ) vid Mellersta Österbottens Vuxeninstitut .
vuxenutbildningen anordnar även förberedande utbildning för vuxna invandrare vid Mellersta Österbottens folkhögskola i Kelviå .
vid Kronoby folkhögskola kan du studera finska och svenska på grund- och påbyggnadsnivå .
om du är berättigad till integrationsstöd ska du kontakta TE @-@ byrån innan du ansöker .
du kan be om information om undervisning i finska och svenska för invandrare hos utlänningsbyrån .
Läs mer : finska och svenska språket
Karlebynejdens institutfinska _ svenska
linkkiMellersta Österbottens utbildningskoncern :
utbildning för invandrarefinska _ engelska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Utlänningsbyrånfinska _ svenska
linkkiKronoby folkhögskola :
Kronoby folkhögskolafinska _ svenska _ engelska
möjligheter att studera finska eller svenska
Karlebynejdens institut erbjuder undervisning i finska och svenska från grundnivå .
Mellersta Österbottens utbildningskoncern erbjuder kurser i finska vid Mellersta Österbottens folkhögskola i Kelviå inom utbildningen i läs- och skrivfärdigheter och den förberedande utbildningen för vuxna invandrare . det går också att studera finska inom utbildningen som handleder för yrkesutbildning ( VALMA ) vid Mellersta Österbottens Vuxeninstitut .
vuxenutbildningen anordnar även förberedande utbildning för vuxna invandrare vid Mellersta Österbottens folkhögskola i Kelviå .
vid Kronoby folkhögskola kan du studera finska och svenska på grund- och påbyggnadsnivå .
om du är berättigad till integrationsstöd ska du kontakta TE @-@ byrån innan du ansöker .
du kan be om information om undervisning i finska och svenska för invandrare hos utlänningsbyrån .
Läs mer : finska och svenska språket
Karlebynejdens institutfinska _ svenska
linkkiMellersta Österbottens utbildningskoncern :
utbildning för invandrarefinska _ engelska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Utlänningsbyrånfinska _ svenska
linkkiKronoby folkhögskola :
Kronoby folkhögskolafinska _ svenska _ engelska
möjligheter att studera finska eller svenska
Karlebynejdens institut erbjuder undervisning i finska och svenska från grundnivå .
Mellersta Österbottens utbildningskoncern erbjuder kurser i finska vid Mellersta Österbottens folkhögskola i Kelviå inom utbildningen i läs- och skrivfärdigheter och den förberedande utbildningen för vuxna invandrare . det går också att studera finska inom utbildningen som handleder för yrkesutbildning ( VALMA ) vid Mellersta Österbottens Vuxeninstitut .
vuxenutbildningen anordnar även förberedande utbildning för vuxna invandrare vid Mellersta Österbottens folkhögskola i Kelviå .
vid Kronoby folkhögskola kan du studera finska och svenska på grund- och påbyggnadsnivå .
om du är berättigad till integrationsstöd ska du kontakta TE @-@ byrån innan du ansöker .
du kan be om information om undervisning i finska och svenska för invandrare hos utlänningsbyrån .
Läs mer : finska och svenska språket
Karlebynejdens institutfinska _ svenska
linkkiMellersta Österbottens utbildningskoncern :
utbildning för invandrarefinska _ engelska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Utlänningsbyrånfinska _ svenska
linkkiKronoby folkhögskola :
Kronoby folkhögskolafinska _ svenska _ engelska
var hittar jag jobb ?
att grunda ett företag
beskattning
om du blir arbetslös
var hittar jag jobb ?
du kan söka arbetsplatser på internet och i tidningar .
på internet hittar du jobbsajter när du skriver &quot; avoimet työpaikat &quot; ( lediga jobb ) i sökmotorns textfält .
på många jobbsajter kan du spara din jobbansökan och meritförteckning ( CV ) så att arbetsgivaren kan läsa dem .
vid Österbottens TE @-@ byrå ( arbets- och näringsbyrå ) får du hjälp med att hitta en arbetsplats .
du behöver inte alltid boka tid för att besöka TE @-@ byrån .
i Mina e @-@ tjänster på nätet kan du bl.a. ändra dina uppgifter som arbetssökande och kontrollera giltighetstiden för jobbsökningen och utlåtandet om arbetslöshetsförsäkring .
om du behöver boka en tid till TE @-@ byrån ska du kontakta TE @-@ byrån direkt per telefon eller boka en tid på plats .
var även direkt i kontakt med TE @-@ byrån om du önskar ändra en tidsbokning .
du kan ringa TE @-@ telefonservice då du behöver information om TE @-@ byråns tjänster eller vägledning i tjänsterna på nätet .
telefonnumret till TE @-@ telefonservice är 0295.025.500 på finska , 0295.025.510 på svenska , 0295.020.713 på engelska och 0295.020.715 på ryska .
TE @-@ byrån i Österbotten betjänar i Karleby , Kaustby , Jakobstad , Närpes , Kristinestad och Vasa .
du kan fritt välja vilken TE @-@ byrå du besöker .
adressen för TE @-@ byrån i Karleby är
67100 Karleby .
på TE @-@ byråns jobbsajt finns tusentals arbetsplatser runt om i Finland .
du hittar lediga arbetsplatser i din kommun genom att skriva kommunens namn i sökfältet &quot; Region &quot; .
Läs mer :
var hittar jag jobb ?
linkkiArbets- och näringsbyråns tjänster :
offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiArbets- och näringsbyråns tjänster :
Österbottens TE @-@ byråfinska _ svenska
linkkiArbets- och näringsbyråns tjänster :
TE @-@ telefonservicefinska _ svenska _ engelska _ ryska
linkkiArbets- och näringsbyråns tjänster :
arbets- och näringsbyråns arbetsplatssajtfinska _ svenska
att grunda ett företag
KOSEK ( Karlebynejdens Utveckling Ab ) erbjuder tjänster som nyttar företaget under hela dess livscykel , från och med att starta företagsverksamhet .
KOSEKs experter hjälper bland annat med att utarbeta en affärsverksamhetsplan och att ansöka startpeng .
tjänsterna är avgiftsfria .
verksamheten av Mellersta Österbottens Nyföretagarcentral FIRMAXI fortsätter som en del av KOSEKs tjänster .
du kan besöka Karlebynejdens Utveckling Ab om du behöver information om att grunda ett företag .
detta kan exempelvis inkludera
företagsfinansiering
rekrytering av anställda
samarbetsnätverk
verksamhetslokaler
Läs mer :
att grunda ett företag .
linkkiNyföretagarcentralen Firmaxi :
Nyföretagarcentralen Firmaxifinska
Karlebynejdens Utveckling Abfinska _ svenska _ engelska
beskattning
om du behöver ett skattekort eller skattenummer kan du besöka Västra Finlands skattebyrå .
Skattebyråns kontaktuppgifter :
PB 1002 , 67101 Karleby
Besöksadress : Karlebygatan 27 , Karleby
Skatteförvaltningens riksomfattande telefontjänst : 029.497.050
Läs mer : beskattning .
om du blir arbetslös
medborgare i EU- och EES @-@ länderna kan anmäla sig som arbetslösa på nätet i TE @-@ byråns &quot; Mina e @-@ tjänster &quot; .
du kan besöka TE @-@ byrån om du inte kan anmäla dig som arbetssökande på nätet eller om du är medborgare i något annat land .
du kan ringa till riksomfattande servicenummer om du behöver hjälp med att använda e @-@ tjänsterna eller mer information om TE @-@ byråns tjänster .
det riksomfattande servicenumret är 0295.025.500 på finska , 0295.025.510 på svenska , 0295.020.713 på engelska och 0295.020.715 på ryska .
TE @-@ byrån i Österbotten betjänar i Karleby , Kaustby , Jakobstad , Närpes , Kristinestad och Vasa .
du kan fritt välja vilken TE @-@ byrå du besöker .
TE @-@ byråns adress i Karleby
Läs mer : Arbetslöshetsförsäkring .
linkkiArbets- och näringsbyråns tjänster :
offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiArbets- och näringsbyråns tjänster :
Österbottens TE @-@ byråfinska _ svenska
linkkiArbets- och näringsbyråns tjänster :
TE @-@ telefonservicefinska _ svenska _ engelska _ ryska
Fennovoima bygger kärnkraftverksenheten Hanhikivi 1 i Pyhäjoki .
kärnkraftverket levereras av RAOS Project Oy , ett bolag som ingår i den ryska Rosatom @-@ koncernen .
enligt den överenskomna tidtabellen kommer kärnkraftverket att producera el år 2024 .
Planeringen och konstruktionen av kärnkraftverket är ett omfattande projekt som tar cirka 10 år att slutföra .
under tiden kärnkraftverket uppförs kommer som mest upp till 3.000 @-@ 4.000 personer att arbeta på området .
arbetsgivaren arrangerar logi för merparten av arbetstagarna , och man strävar efter att ordna inkvartering så nära bygget som möjligt .
i kärnkraftverkets omedelbara närhet byggs ett inkvarteringsområde för 1.000 personer .
i Pyhäjoki och det omgivande området har man förberett sig på kärnkraftverksprojektet redan i flera års tid .
information om området har sammanställts bl.a. i Hanhikivi @-@ guiden som publicerats på finska , engelska , svenska och ryska .
elektroniska versioner av guiden finns på storprojektets webbplats .
den tryckta guiden finns i företagsservicecentralerna i kommunerna på området .
som en del av förberedelserna för kärnkraftverksprojektet finns information samlad om tjänsterna på området på dessa lokala InfoFinland @-@ sidor .
mer information om Fennovoimas kärnkraftverksprojekt i Pyhäjoki :
Fennovoima Oyfinska _ engelska
linkkiBrahestadsregionens företagstjänster :
information om storprojekt som förverkligas i regionen och förberedelserna för dessafinska _ engelska _ ryska
Karlebynejdens Utveckling Abfinska _ svenska _ engelska
linkkiPyhäjoki kommun :
Pyhäjoki kommunfinska _ svenska _ engelska
information om verksamhetsmiljön för kärnkraftverksprojektetfinska _ svenska _ engelska _ ryska
var hittar jag jobb ?
att grunda ett företag
beskattning
om du blir arbetslös
var hittar jag jobb ?
du kan söka arbetsplatser på internet och i tidningar .
på internet hittar du jobbsajter när du skriver &quot; avoimet työpaikat &quot; ( lediga jobb ) i sökmotorns textfält .
på många jobbsajter kan du spara din jobbansökan och meritförteckning ( CV ) så att arbetsgivaren kan läsa dem .
vid Österbottens TE @-@ byrå ( arbets- och näringsbyrå ) får du hjälp med att hitta en arbetsplats .
du behöver inte alltid boka tid för att besöka TE @-@ byrån .
i Mina e @-@ tjänster på nätet kan du bl.a. ändra dina uppgifter som arbetssökande och kontrollera giltighetstiden för jobbsökningen och utlåtandet om arbetslöshetsförsäkring .
om du behöver boka en tid till TE @-@ byrån ska du kontakta TE @-@ byrån direkt per telefon eller boka en tid på plats .
var även direkt i kontakt med TE @-@ byrån om du önskar ändra en tidsbokning .
du kan ringa TE @-@ telefonservice då du behöver information om TE @-@ byråns tjänster eller vägledning i tjänsterna på nätet .
telefonnumret till TE @-@ telefonservice är 0295.025.500 på finska , 0295.025.510 på svenska , 0295.020.713 på engelska och 0295.020.715 på ryska .
TE @-@ byrån i Österbotten betjänar i Karleby , Kaustby , Jakobstad , Närpes , Kristinestad och Vasa .
du kan fritt välja vilken TE @-@ byrå du besöker .
adressen för TE @-@ byrån i Karleby är
67100 Karleby .
på TE @-@ byråns jobbsajt finns tusentals arbetsplatser runt om i Finland .
du hittar lediga arbetsplatser i din kommun genom att skriva kommunens namn i sökfältet &quot; Region &quot; .
Läs mer :
var hittar jag jobb ?
linkkiArbets- och näringsbyråns tjänster :
offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiArbets- och näringsbyråns tjänster :
Österbottens TE @-@ byråfinska _ svenska
linkkiArbets- och näringsbyråns tjänster :
TE @-@ telefonservicefinska _ svenska _ engelska _ ryska
linkkiArbets- och näringsbyråns tjänster :
arbets- och näringsbyråns arbetsplatssajtfinska _ svenska
att grunda ett företag
KOSEK ( Karlebynejdens Utveckling Ab ) erbjuder tjänster som nyttar företaget under hela dess livscykel , från och med att starta företagsverksamhet .
KOSEKs experter hjälper bland annat med att utarbeta en affärsverksamhetsplan och att ansöka startpeng .
tjänsterna är avgiftsfria .
verksamheten av Mellersta Österbottens Nyföretagarcentral FIRMAXI fortsätter som en del av KOSEKs tjänster .
du kan besöka Karlebynejdens Utveckling Ab om du behöver information om att grunda ett företag .
detta kan exempelvis inkludera
företagsfinansiering
rekrytering av anställda
samarbetsnätverk
verksamhetslokaler
Läs mer :
att grunda ett företag .
linkkiNyföretagarcentralen Firmaxi :
Nyföretagarcentralen Firmaxifinska
Karlebynejdens Utveckling Abfinska _ svenska _ engelska
beskattning
om du behöver ett skattekort eller skattenummer kan du besöka Västra Finlands skattebyrå .
Skattebyråns kontaktuppgifter :
PB 1002 , 67101 Karleby
Besöksadress : Karlebygatan 27 , Karleby
Skatteförvaltningens riksomfattande telefontjänst : 029.497.050
Läs mer : beskattning .
om du blir arbetslös
medborgare i EU- och EES @-@ länderna kan anmäla sig som arbetslösa på nätet i TE @-@ byråns &quot; Mina e @-@ tjänster &quot; .
du kan besöka TE @-@ byrån om du inte kan anmäla dig som arbetssökande på nätet eller om du är medborgare i något annat land .
du kan ringa till riksomfattande servicenummer om du behöver hjälp med att använda e @-@ tjänsterna eller mer information om TE @-@ byråns tjänster .
det riksomfattande servicenumret är 0295.025.500 på finska , 0295.025.510 på svenska , 0295.020.713 på engelska och 0295.020.715 på ryska .
TE @-@ byrån i Österbotten betjänar i Karleby , Kaustby , Jakobstad , Närpes , Kristinestad och Vasa .
du kan fritt välja vilken TE @-@ byrå du besöker .
TE @-@ byråns adress i Karleby
Läs mer : Arbetslöshetsförsäkring .
linkkiArbets- och näringsbyråns tjänster :
offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiArbets- och näringsbyråns tjänster :
Österbottens TE @-@ byråfinska _ svenska
linkkiArbets- och näringsbyråns tjänster :
TE @-@ telefonservicefinska _ svenska _ engelska _ ryska
Fennovoima bygger kärnkraftverksenheten Hanhikivi 1 i Pyhäjoki .
kärnkraftverket levereras av RAOS Project Oy , ett bolag som ingår i den ryska Rosatom @-@ koncernen .
enligt den överenskomna tidtabellen kommer kärnkraftverket att producera el år 2024 .
Planeringen och konstruktionen av kärnkraftverket är ett omfattande projekt som tar cirka 10 år att slutföra .
under tiden kärnkraftverket uppförs kommer som mest upp till 3.000 @-@ 4.000 personer att arbeta på området .
arbetsgivaren arrangerar logi för merparten av arbetstagarna , och man strävar efter att ordna inkvartering så nära bygget som möjligt .
i kärnkraftverkets omedelbara närhet byggs ett inkvarteringsområde för 1.000 personer .
i Pyhäjoki och det omgivande området har man förberett sig på kärnkraftverksprojektet redan i flera års tid .
information om området har sammanställts bl.a. i Hanhikivi @-@ guiden som publicerats på finska , engelska , svenska och ryska .
elektroniska versioner av guiden finns på storprojektets webbplats .
den tryckta guiden finns i företagsservicecentralerna i kommunerna på området .
som en del av förberedelserna för kärnkraftverksprojektet finns information samlad om tjänsterna på området på dessa lokala InfoFinland @-@ sidor .
mer information om Fennovoimas kärnkraftverksprojekt i Pyhäjoki :
Fennovoima Oyfinska _ engelska
linkkiBrahestadsregionens företagstjänster :
information om storprojekt som förverkligas i regionen och förberedelserna för dessafinska _ engelska _ ryska
Karlebynejdens Utveckling Abfinska _ svenska _ engelska
linkkiPyhäjoki kommun :
Pyhäjoki kommunfinska _ svenska _ engelska
information om verksamhetsmiljön för kärnkraftverksprojektetfinska _ svenska _ engelska _ ryska
var hittar jag jobb ?
att grunda ett företag
beskattning
om du blir arbetslös
var hittar jag jobb ?
du kan söka arbetsplatser på internet och i tidningar .
på internet hittar du jobbsajter när du skriver &quot; avoimet työpaikat &quot; ( lediga jobb ) i sökmotorns textfält .
på många jobbsajter kan du spara din jobbansökan och meritförteckning ( CV ) så att arbetsgivaren kan läsa dem .
vid Österbottens TE @-@ byrå ( arbets- och näringsbyrå ) får du hjälp med att hitta en arbetsplats .
du behöver inte alltid boka tid för att besöka TE @-@ byrån .
i Mina e @-@ tjänster på nätet kan du bl.a. ändra dina uppgifter som arbetssökande och kontrollera giltighetstiden för jobbsökningen och utlåtandet om arbetslöshetsförsäkring .
om du behöver boka en tid till TE @-@ byrån ska du kontakta TE @-@ byrån direkt per telefon eller boka en tid på plats .
var även direkt i kontakt med TE @-@ byrån om du önskar ändra en tidsbokning .
du kan ringa TE @-@ telefonservice då du behöver information om TE @-@ byråns tjänster eller vägledning i tjänsterna på nätet .
telefonnumret till TE @-@ telefonservice är 0295.025.500 på finska , 0295.025.510 på svenska , 0295.020.713 på engelska och 0295.020.715 på ryska .
TE @-@ byrån i Österbotten betjänar i Karleby , Kaustby , Jakobstad , Närpes , Kristinestad och Vasa .
du kan fritt välja vilken TE @-@ byrå du besöker .
adressen för TE @-@ byrån i Karleby är
67100 Karleby .
på TE @-@ byråns jobbsajt finns tusentals arbetsplatser runt om i Finland .
du hittar lediga arbetsplatser i din kommun genom att skriva kommunens namn i sökfältet &quot; Region &quot; .
Läs mer :
var hittar jag jobb ?
linkkiArbets- och näringsbyråns tjänster :
offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiArbets- och näringsbyråns tjänster :
Österbottens TE @-@ byråfinska _ svenska
linkkiArbets- och näringsbyråns tjänster :
TE @-@ telefonservicefinska _ svenska _ engelska _ ryska
linkkiArbets- och näringsbyråns tjänster :
arbets- och näringsbyråns arbetsplatssajtfinska _ svenska
att grunda ett företag
KOSEK ( Karlebynejdens Utveckling Ab ) erbjuder tjänster som nyttar företaget under hela dess livscykel , från och med att starta företagsverksamhet .
KOSEKs experter hjälper bland annat med att utarbeta en affärsverksamhetsplan och att ansöka startpeng .
tjänsterna är avgiftsfria .
verksamheten av Mellersta Österbottens Nyföretagarcentral FIRMAXI fortsätter som en del av KOSEKs tjänster .
du kan besöka Karlebynejdens Utveckling Ab om du behöver information om att grunda ett företag .
detta kan exempelvis inkludera
företagsfinansiering
rekrytering av anställda
samarbetsnätverk
verksamhetslokaler
Läs mer :
att grunda ett företag .
linkkiNyföretagarcentralen Firmaxi :
Nyföretagarcentralen Firmaxifinska
Karlebynejdens Utveckling Abfinska _ svenska _ engelska
beskattning
om du behöver ett skattekort eller skattenummer kan du besöka Västra Finlands skattebyrå .
Skattebyråns kontaktuppgifter :
PB 1002 , 67101 Karleby
Besöksadress : Karlebygatan 27 , Karleby
Skatteförvaltningens riksomfattande telefontjänst : 029.497.050
Läs mer : beskattning .
om du blir arbetslös
medborgare i EU- och EES @-@ länderna kan anmäla sig som arbetslösa på nätet i TE @-@ byråns &quot; Mina e @-@ tjänster &quot; .
du kan besöka TE @-@ byrån om du inte kan anmäla dig som arbetssökande på nätet eller om du är medborgare i något annat land .
du kan ringa till riksomfattande servicenummer om du behöver hjälp med att använda e @-@ tjänsterna eller mer information om TE @-@ byråns tjänster .
det riksomfattande servicenumret är 0295.025.500 på finska , 0295.025.510 på svenska , 0295.020.713 på engelska och 0295.020.715 på ryska .
TE @-@ byrån i Österbotten betjänar i Karleby , Kaustby , Jakobstad , Närpes , Kristinestad och Vasa .
du kan fritt välja vilken TE @-@ byrå du besöker .
TE @-@ byråns adress i Karleby
Läs mer : Arbetslöshetsförsäkring .
linkkiArbets- och näringsbyråns tjänster :
offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiArbets- och näringsbyråns tjänster :
Österbottens TE @-@ byråfinska _ svenska
linkkiArbets- och näringsbyråns tjänster :
TE @-@ telefonservicefinska _ svenska _ engelska _ ryska
Fennovoima bygger kärnkraftverksenheten Hanhikivi 1 i Pyhäjoki .
kärnkraftverket levereras av RAOS Project Oy , ett bolag som ingår i den ryska Rosatom @-@ koncernen .
enligt den överenskomna tidtabellen kommer kärnkraftverket att producera el år 2024 .
Planeringen och konstruktionen av kärnkraftverket är ett omfattande projekt som tar cirka 10 år att slutföra .
under tiden kärnkraftverket uppförs kommer som mest upp till 3.000 @-@ 4.000 personer att arbeta på området .
arbetsgivaren arrangerar logi för merparten av arbetstagarna , och man strävar efter att ordna inkvartering så nära bygget som möjligt .
i kärnkraftverkets omedelbara närhet byggs ett inkvarteringsområde för 1.000 personer .
i Pyhäjoki och det omgivande området har man förberett sig på kärnkraftverksprojektet redan i flera års tid .
information om området har sammanställts bl.a. i Hanhikivi @-@ guiden som publicerats på finska , engelska , svenska och ryska .
elektroniska versioner av guiden finns på storprojektets webbplats .
den tryckta guiden finns i företagsservicecentralerna i kommunerna på området .
som en del av förberedelserna för kärnkraftverksprojektet finns information samlad om tjänsterna på området på dessa lokala InfoFinland @-@ sidor .
mer information om Fennovoimas kärnkraftverksprojekt i Pyhäjoki :
Fennovoima Oyfinska _ engelska
linkkiBrahestadsregionens företagstjänster :
information om storprojekt som förverkligas i regionen och förberedelserna för dessafinska _ engelska _ ryska
Karlebynejdens Utveckling Abfinska _ svenska _ engelska
linkkiPyhäjoki kommun :
Pyhäjoki kommunfinska _ svenska _ engelska
information om verksamhetsmiljön för kärnkraftverksprojektetfinska _ svenska _ engelska _ ryska
rådgivning och integration för invandrare
inledande kartläggning och integrationsplan
behöver du en tolk ?
rådgivning och integration för invandrare
då du flyttar till Finland kan du använda dig av TE @-@ byråns ( arbets- och näringsbyrån ) tjänster som hjälper dig att göra dig hemmastadd i Finland och hitta en arbetsplats .
tjänster särskilt avsedda för invandrare är :
handledning och rådgivning för invandrare
inledande kartläggning
integrationsutbildning
Österbottens TE @-@ byrå
67100 Karleby
Telefonväxel : 0295.025.500
Karleby evangelisk @-@ lutherska församlingssammanslutnings invandrararbete stöder invandrares integrering i det finländska samhället .
linkkiArbets- och näringsbyråns tjänster :
offentliga arbets- och näringstjänsterfinska _ svenska
linkkiArbets- och näringsministeriet :
guiden Välkommen till Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
linkkiKarleby evangelisk @-@ lutherska församlingssammansutning :
Karleby evangelisk @-@ lutherska församlings invandrararbetefinska _ svenska _ engelska _ ryska
inledande kartläggning och integrationsplan
en inledande kartläggning och integrationsplan utarbetas för dig i arbets- och näringsbyrån . om du kommit till
Finland som flykting utarbetas en inledande kartläggning och integrationsplan för dig vid utlänningsbyrån .
du kan fråga mer om kartläggningen och integrationsplanen vid utlänningsbyrån eller TE @-@ byrån .
utlänningsbyrån
Vasavägen 6 C
67100 Karleby
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Utlänningsbyrånfinska _ svenska
behöver du en tolk ?
om du måste sköta ärenden med finländska myndigheter , men inte kan finska eller svenska och det inte heller finns något annat språk som både du och myndigheten talar , kan du i vissa fall ha rätt till tolkning .
myndigheten beställer tolken om du på förhand uppgett att du behöver en tolk .
i detta fall är det gratis för dig att använda dig av tolk .
du kan använda tolken när du själv önskar om du betalar kostnaderna och beställer tolken själv .
Läs mer :
behöver du en tolk ?
rådgivning och integration för invandrare
inledande kartläggning och integrationsplan
behöver du en tolk ?
rådgivning och integration för invandrare
då du flyttar till Finland kan du använda dig av TE @-@ byråns ( arbets- och näringsbyrån ) tjänster som hjälper dig att göra dig hemmastadd i Finland och hitta en arbetsplats .
tjänster särskilt avsedda för invandrare är :
handledning och rådgivning för invandrare
inledande kartläggning
integrationsutbildning
Österbottens TE @-@ byrå
67100 Karleby
Telefonväxel : 0295.025.500
Karleby evangelisk @-@ lutherska församlingssammanslutnings invandrararbete stöder invandrares integrering i det finländska samhället .
linkkiArbets- och näringsbyråns tjänster :
offentliga arbets- och näringstjänsterfinska _ svenska
linkkiArbets- och näringsministeriet :
guiden Välkommen till Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
linkkiKarleby evangelisk @-@ lutherska församlingssammansutning :
Karleby evangelisk @-@ lutherska församlings invandrararbetefinska _ svenska _ engelska _ ryska
inledande kartläggning och integrationsplan
en inledande kartläggning och integrationsplan utarbetas för dig i arbets- och näringsbyrån . om du kommit till
Finland som flykting utarbetas en inledande kartläggning och integrationsplan för dig vid utlänningsbyrån .
du kan fråga mer om kartläggningen och integrationsplanen vid utlänningsbyrån eller TE @-@ byrån .
utlänningsbyrån
Vasavägen 6 C
67100 Karleby
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Utlänningsbyrånfinska _ svenska
behöver du en tolk ?
om du måste sköta ärenden med finländska myndigheter , men inte kan finska eller svenska och det inte heller finns något annat språk som både du och myndigheten talar , kan du i vissa fall ha rätt till tolkning .
myndigheten beställer tolken om du på förhand uppgett att du behöver en tolk .
i detta fall är det gratis för dig att använda dig av tolk .
du kan använda tolken när du själv önskar om du betalar kostnaderna och beställer tolken själv .
Läs mer :
behöver du en tolk ?
rådgivning och integration för invandrare
inledande kartläggning och integrationsplan
behöver du en tolk ?
rådgivning och integration för invandrare
då du flyttar till Finland kan du använda dig av TE @-@ byråns ( arbets- och näringsbyrån ) tjänster som hjälper dig att göra dig hemmastadd i Finland och hitta en arbetsplats .
tjänster särskilt avsedda för invandrare är :
handledning och rådgivning för invandrare
inledande kartläggning
integrationsutbildning
Österbottens TE @-@ byrå
67100 Karleby
Telefonväxel : 0295.025.500
Karleby evangelisk @-@ lutherska församlingssammanslutnings invandrararbete stöder invandrares integrering i det finländska samhället .
linkkiArbets- och näringsbyråns tjänster :
offentliga arbets- och näringstjänsterfinska _ svenska
linkkiArbets- och näringsministeriet :
guiden Välkommen till Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
linkkiKarleby evangelisk @-@ lutherska församlingssammansutning :
Karleby evangelisk @-@ lutherska församlings invandrararbetefinska _ svenska _ engelska _ ryska
inledande kartläggning och integrationsplan
en inledande kartläggning och integrationsplan utarbetas för dig i arbets- och näringsbyrån . om du kommit till
Finland som flykting utarbetas en inledande kartläggning och integrationsplan för dig vid utlänningsbyrån .
du kan fråga mer om kartläggningen och integrationsplanen vid utlänningsbyrån eller TE @-@ byrån .
utlänningsbyrån
Vasavägen 6 C
67100 Karleby
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Utlänningsbyrånfinska _ svenska
behöver du en tolk ?
om du måste sköta ärenden med finländska myndigheter , men inte kan finska eller svenska och det inte heller finns något annat språk som både du och myndigheten talar , kan du i vissa fall ha rätt till tolkning .
myndigheten beställer tolken om du på förhand uppgett att du behöver en tolk .
i detta fall är det gratis för dig att använda dig av tolk .
du kan använda tolken när du själv önskar om du betalar kostnaderna och beställer tolken själv .
Läs mer :
behöver du en tolk ?
registrering som invånare
om du vill flytta till Finland behöver du vanligtvis ett uppehållstillstånd .
Uppehållstillståndsärenden hanteras av Finlands beskickningar i utlandet och Migrationsverket .
Läs mer : flytta till Finland .
då du flyttar till Karleby ( Kokkola ) ska du registrera dig som invånare i kommunen .
du kan personligen registrera dig på Karleby enheten för Magistraten i Västra Finland :
magistraten i Västra Finland
Karleby enhet
Karlebygatan 27
67701 Karleby
telefon : 029.553.9451
när du går till magistraten ska du ta med dig
uppehållstillstånd och uppehållskort ( om du behöver ett uppehållstillstånd i Finland )
registreringsintyget över uppehållsrätt för EU @-@ medborgare ( om du är EU @-@ medborgare )
äktenskapsbevis
födelseattester för dina barn
Observera att officiella handlingar som tagits med från utlandet ska vara legaliserade och i original samt översatta till finska , svenska eller engelska .
mer information om legalisering av handlingar får du hos magistraten eller hos ditt lands beskickning i Finland .
Läs mer :
registrering som invånare .
magistratens kontaktuppgifterfinska _ svenska _ engelska
fortsatt uppehållstillstånd
du ska ansöka om fortsatt uppehållstillstånd innan ditt tidigare uppehållstillstånd går ut .
du ansöker om tillståndet vid Migrationsverkets servicesställen .
du kan endast ansöka om fortsatt uppehållstillstånd i Finland .
Migrationsverket
Korsholmsesplanaden 45
Vasa
Läs mer : fortsatt uppehållstillstånd .
registrering som invånare
om du vill flytta till Finland behöver du vanligtvis ett uppehållstillstånd .
Uppehållstillståndsärenden hanteras av Finlands beskickningar i utlandet och Migrationsverket .
Läs mer : flytta till Finland .
då du flyttar till Karleby ( Kokkola ) ska du registrera dig som invånare i kommunen .
du kan personligen registrera dig på Karleby enheten för Magistraten i Västra Finland :
magistraten i Västra Finland
Karleby enhet
Karlebygatan 27
67701 Karleby
telefon : 029.553.9451
när du går till magistraten ska du ta med dig
uppehållstillstånd och uppehållskort ( om du behöver ett uppehållstillstånd i Finland )
registreringsintyget över uppehållsrätt för EU @-@ medborgare ( om du är EU @-@ medborgare )
äktenskapsbevis
födelseattester för dina barn
Observera att officiella handlingar som tagits med från utlandet ska vara legaliserade och i original samt översatta till finska , svenska eller engelska .
mer information om legalisering av handlingar får du hos magistraten eller hos ditt lands beskickning i Finland .
Läs mer :
registrering som invånare .
magistratens kontaktuppgifterfinska _ svenska _ engelska
fortsatt uppehållstillstånd
du ska ansöka om fortsatt uppehållstillstånd innan ditt tidigare uppehållstillstånd går ut .
du ansöker om tillståndet vid Migrationsverkets servicesställen .
du kan endast ansöka om fortsatt uppehållstillstånd i Finland .
Migrationsverket
Korsholmsesplanaden 45
Vasa
Läs mer : fortsatt uppehållstillstånd .
registrering som invånare
om du vill flytta till Finland behöver du vanligtvis ett uppehållstillstånd .
Uppehållstillståndsärenden hanteras av Finlands beskickningar i utlandet och Migrationsverket .
Läs mer : flytta till Finland .
då du flyttar till Karleby ( Kokkola ) ska du registrera dig som invånare i kommunen .
du kan personligen registrera dig på Karleby enheten för Magistraten i Västra Finland :
magistraten i Västra Finland
Karleby enhet
Karlebygatan 27
67701 Karleby
telefon : 029.553.9451
när du går till magistraten ska du ta med dig
uppehållstillstånd och uppehållskort ( om du behöver ett uppehållstillstånd i Finland )
registreringsintyget över uppehållsrätt för EU @-@ medborgare ( om du är EU @-@ medborgare )
äktenskapsbevis
födelseattester för dina barn
Observera att officiella handlingar som tagits med från utlandet ska vara legaliserade och i original samt översatta till finska , svenska eller engelska .
mer information om legalisering av handlingar får du hos magistraten eller hos ditt lands beskickning i Finland .
Läs mer :
registrering som invånare .
magistratens kontaktuppgifterfinska _ svenska _ engelska
fortsatt uppehållstillstånd
du ska ansöka om fortsatt uppehållstillstånd innan ditt tidigare uppehållstillstånd går ut .
du ansöker om tillståndet vid Migrationsverkets servicesställen .
du kan endast ansöka om fortsatt uppehållstillstånd i Finland .
Migrationsverket
Korsholmsesplanaden 45
Vasa
Läs mer : fortsatt uppehållstillstånd .
InfoFinland finansieras av Samarbetskommunerna och staten .
åren 2017 @-@ 2020 var statens finansiärer arbets- och näringsministeriet , undervisnings- och kulturministeriet , miljöministeriet , FPA och Skatteförvaltningen .
InfoFinland utvecklas i samarbete med finansiärerna .
den som planerar att flytta till Finland med hjälp av Infobanken hittar lätt information om att leva , bo , arbeta och studera i Finland på många olika språk .
staten
arbets- och näringsministeriet
arbets- och näringsministeriet svarar för beredningen av ärenden i anslutning till integrationen av invandrare i Finland .
Kompetenscentret för integration av invandrare stöder arbete som främjar integrationen av invandrare lokalt , regionalt och riksomfattande .
linkkiArbets- och näringsministeriet :
integration av invandrarefinska _ svenska _ engelska
undervisnings- och kulturministeriet
undervisnings- och kulturministeriet svarar för utvecklingen av och det internationella samarbetet inom utbildnings- , vetenskaps- , kultur- , motions- och ungdomspolitiken .
linkkiUndervisnings- och kulturministeriet :
Webbsidorfinska _ svenska _ engelska
miljöministeriet
linkkiMiljöministeriet :
Webbsidorfinska _ svenska _ engelska
FPA
FPA sköter grundtryggheten i olika skeden av livet för dem som bor i Finland .
FPA:s kunder är alla personer som bor i Finland och utomlands och som omfattas av socialskyddet i Finland .
FPA och Skatteförvaltningen erbjuder information till utländska anställda på servicestället In To Finland i Helsingfors .
Flyttning till eller från Finlandfinska _ svenska _ engelska
Skatteförvaltningen
linkkiSkatteförvaltningen :
Webbsidorfinska _ svenska _ engelska
kommunerna
Helsingfors stad
Publicerar och administrerar InfoFinland .
kommuner som är med i samarbetsavtalet
InfoFinlands samarbetsavtal
InfoFinlands finansiärer har ingått ett samarbetsavtal med vilket man överenskommit om principerna för genomförandet och finansieringen av nättjänsten InfoFinland ( tidigare Infobanken ) för åren 2017 @-@ 2020 .
samarbetet möjliggör riksomfattande webbinformation för invandrare och personer som planerar att flytta till Finland och för myndigheter inom invandrarsektorn på ett sätt som också stöder behovet av information i kommunerna .
det är lätt att på ett pålitligt sätt hitta väsentlig information om integration av invandrare och om att bo i Finland på ett ställe , www.infofinland.fi .
Avtalsparterna driver och utvecklar tjänsten tillsammans .
de vill dessutom stärka InfoFinlands riksomfattande ställning , så att det är möjligt för nya kommuner och andra organisationer att ansluta sig till tjänsten också i fortsättningen .
Kommunernas finansieringsandelar fastställs utgående från antalet invånare .
genomförandet av avtalet följs upp av en styrgrupp .
nya aktörer är välkomna att utveckla den flerspråkiga informationen till invandrare och ansluta sig till InfoFinlands samarbetsavtal .
närmare information om hur man ansluter sig till avtalet ger InfoFinlands chefredaktör Eija Kyllönen @-@ Saarnio , eija.kyllonen @-@ saarnio ( snabel @-@ a ) hel.fi , tfn 050.363.3285 .
InfoFinland finansieras av Samarbetskommunerna och staten .
åren 2017 @-@ 2020 var statens finansiärer arbets- och näringsministeriet , undervisnings- och kulturministeriet , miljöministeriet , FPA och Skatteförvaltningen .
InfoFinland utvecklas i samarbete med finansiärerna .
den som planerar att flytta till Finland med hjälp av Infobanken hittar lätt information om att leva , bo , arbeta och studera i Finland på många olika språk .
staten
arbets- och näringsministeriet
arbets- och näringsministeriet svarar för beredningen av ärenden i anslutning till integrationen av invandrare i Finland .
Kompetenscentret för integration av invandrare stöder arbete som främjar integrationen av invandrare lokalt , regionalt och riksomfattande .
linkkiArbets- och näringsministeriet :
integration av invandrarefinska _ svenska _ engelska
undervisnings- och kulturministeriet
undervisnings- och kulturministeriet svarar för utvecklingen av och det internationella samarbetet inom utbildnings- , vetenskaps- , kultur- , motions- och ungdomspolitiken .
linkkiUndervisnings- och kulturministeriet :
Webbsidorfinska _ svenska _ engelska
miljöministeriet
linkkiMiljöministeriet :
Webbsidorfinska _ svenska _ engelska
FPA
FPA sköter grundtryggheten i olika skeden av livet för dem som bor i Finland .
FPA:s kunder är alla personer som bor i Finland och utomlands och som omfattas av socialskyddet i Finland .
FPA och Skatteförvaltningen erbjuder information till utländska anställda på servicestället In To Finland i Helsingfors .
Flyttning till eller från Finlandfinska _ svenska _ engelska
Skatteförvaltningen
linkkiSkatteförvaltningen :
Webbsidorfinska _ svenska _ engelska
kommunerna
Helsingfors stad
Publicerar och administrerar InfoFinland .
kommuner som är med i samarbetsavtalet
InfoFinlands samarbetsavtal
InfoFinlands finansiärer har ingått ett samarbetsavtal med vilket man överenskommit om principerna för genomförandet och finansieringen av nättjänsten InfoFinland ( tidigare Infobanken ) för åren 2017 @-@ 2020 .
samarbetet möjliggör riksomfattande webbinformation för invandrare och personer som planerar att flytta till Finland och för myndigheter inom invandrarsektorn på ett sätt som också stöder behovet av information i kommunerna .
det är lätt att på ett pålitligt sätt hitta väsentlig information om integration av invandrare och om att bo i Finland på ett ställe , www.infofinland.fi .
Avtalsparterna driver och utvecklar tjänsten tillsammans .
de vill dessutom stärka InfoFinlands riksomfattande ställning , så att det är möjligt för nya kommuner och andra organisationer att ansluta sig till tjänsten också i fortsättningen .
Kommunernas finansieringsandelar fastställs utgående från antalet invånare .
genomförandet av avtalet följs upp av en styrgrupp .
nya aktörer är välkomna att utveckla den flerspråkiga informationen till invandrare och ansluta sig till InfoFinlands samarbetsavtal .
närmare information om hur man ansluter sig till avtalet ger InfoFinlands chefredaktör Eija Kyllönen @-@ Saarnio , eija.kyllonen @-@ saarnio ( snabel @-@ a ) hel.fi , tfn 050.363.3285 .
InfoFinland finansieras av Samarbetskommunerna och staten .
åren 2017 @-@ 2020 var statens finansiärer arbets- och näringsministeriet , undervisnings- och kulturministeriet , miljöministeriet , FPA och Skatteförvaltningen .
InfoFinland utvecklas i samarbete med finansiärerna .
den som planerar att flytta till Finland med hjälp av Infobanken hittar lätt information om att leva , bo , arbeta och studera i Finland på många olika språk .
staten
arbets- och näringsministeriet
arbets- och näringsministeriet svarar för beredningen av ärenden i anslutning till integrationen av invandrare i Finland .
Kompetenscentret för integration av invandrare stöder arbete som främjar integrationen av invandrare lokalt , regionalt och riksomfattande .
linkkiArbets- och näringsministeriet :
integration av invandrarefinska _ svenska _ engelska
undervisnings- och kulturministeriet
undervisnings- och kulturministeriet svarar för utvecklingen av och det internationella samarbetet inom utbildnings- , vetenskaps- , kultur- , motions- och ungdomspolitiken .
linkkiUndervisnings- och kulturministeriet :
Webbsidorfinska _ svenska _ engelska
miljöministeriet
linkkiMiljöministeriet :
Webbsidorfinska _ svenska _ engelska
FPA
FPA sköter grundtryggheten i olika skeden av livet för dem som bor i Finland .
FPA:s kunder är alla personer som bor i Finland och utomlands och som omfattas av socialskyddet i Finland .
FPA och Skatteförvaltningen erbjuder information till utländska anställda på servicestället In To Finland i Helsingfors .
Flyttning till eller från Finlandfinska _ svenska _ engelska
Skatteförvaltningen
linkkiSkatteförvaltningen :
Webbsidorfinska _ svenska _ engelska
kommunerna
Helsingfors stad
Publicerar och administrerar InfoFinland .
kommuner som är med i samarbetsavtalet
InfoFinlands samarbetsavtal
InfoFinlands finansiärer har ingått ett samarbetsavtal med vilket man överenskommit om principerna för genomförandet och finansieringen av nättjänsten InfoFinland ( tidigare Infobanken ) för åren 2017 @-@ 2020 .
samarbetet möjliggör riksomfattande webbinformation för invandrare och personer som planerar att flytta till Finland och för myndigheter inom invandrarsektorn på ett sätt som också stöder behovet av information i kommunerna .
det är lätt att på ett pålitligt sätt hitta väsentlig information om integration av invandrare och om att bo i Finland på ett ställe , www.infofinland.fi .
Avtalsparterna driver och utvecklar tjänsten tillsammans .
de vill dessutom stärka InfoFinlands riksomfattande ställning , så att det är möjligt för nya kommuner och andra organisationer att ansluta sig till tjänsten också i fortsättningen .
Kommunernas finansieringsandelar fastställs utgående från antalet invånare .
genomförandet av avtalet följs upp av en styrgrupp .
nya aktörer är välkomna att utveckla den flerspråkiga informationen till invandrare och ansluta sig till InfoFinlands samarbetsavtal .
närmare information om hur man ansluter sig till avtalet ger InfoFinlands chefredaktör Eija Kyllönen @-@ Saarnio , eija.kyllonen @-@ saarnio ( snabel @-@ a ) hel.fi , tfn 050.363.3285 .
alla texter som publicerats på InfoFinlands webbplats på alla språk är fritt tillgängliga i enlighet med licensen Creative Commons Erkännande 4.0 .
du har tillstånd att :
Dela - kopiera och vidaredistribuera materialet oavsett medium eller format
Bearbeta - remixa , transformera , och bygga vidare på materialet för alla ändamål , även kommersiellt .
på följande villkor :
Erkännande ( BY ) - Du måste nämna källan InfoFinland.fi .
Ange en länk till webbplatsen InfoFinland.fi och nämn licensen CC BY 4.0 .
Ange om bearbetningar är gjorda .
du behöver göra så i enlighet med god sed , och inte på ett sätt som ger en bild av att InfoFinland stödjer dig eller ditt användande .
Inga ytterligare begränsningar - Du får inte tillämpa lagliga begränsningar eller teknologiska metoder som juridiskt begränsar andra från att gör något som licensen tillåter .
Erkännande 4.0 Internationellfinska _ svenska _ engelska _ ryska _ franska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ japanska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ grekiska
_ tjeckiska
öppet programmeringsgränssnitt ( API )
Vi erbjuder allt textinnehåll i InfoFinland via ett öppet programmeringsgränssnitt ( API ) .
med hjälp av gränssnittet kan du visa InfoFinlands innehåll på andra webbplatser eller skapa olika applikationer .
information om gränssnittetfinska _ engelska
öppet programmeringsgränssnittfinska
alla texter som publicerats på InfoFinlands webbplats på alla språk är fritt tillgängliga i enlighet med licensen Creative Commons Erkännande 4.0 .
du har tillstånd att :
Dela - kopiera och vidaredistribuera materialet oavsett medium eller format
Bearbeta - remixa , transformera , och bygga vidare på materialet för alla ändamål , även kommersiellt .
på följande villkor :
Erkännande ( BY ) - Du måste nämna källan InfoFinland.fi .
Ange en länk till webbplatsen InfoFinland.fi och nämn licensen CC BY 4.0 .
Ange om bearbetningar är gjorda .
du behöver göra så i enlighet med god sed , och inte på ett sätt som ger en bild av att InfoFinland stödjer dig eller ditt användande .
Inga ytterligare begränsningar - Du får inte tillämpa lagliga begränsningar eller teknologiska metoder som juridiskt begränsar andra från att gör något som licensen tillåter .
Erkännande 4.0 Internationellfinska _ svenska _ engelska _ ryska _ franska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ japanska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ grekiska
_ tjeckiska
öppet programmeringsgränssnitt ( API )
Vi erbjuder allt textinnehåll i InfoFinland via ett öppet programmeringsgränssnitt ( API ) .
med hjälp av gränssnittet kan du visa InfoFinlands innehåll på andra webbplatser eller skapa olika applikationer .
information om gränssnittetfinska _ engelska
öppet programmeringsgränssnittfinska
Användning av InfoFinland @-@ texterna på andra ställen
texterna ur webbtjänsten InfoFinland.fi används i följande tjänster :
linkkiArbets- och näringsministeriet :
guiden Välkommen till Finland ( pdf , 3,40 MB ) finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
alla texter som publicerats på InfoFinlands webbplats på alla språk är fritt tillgängliga i enlighet med licensen Creative Commons Erkännande 4.0 .
du har tillstånd att :
Dela - kopiera och vidaredistribuera materialet oavsett medium eller format
Bearbeta - remixa , transformera , och bygga vidare på materialet för alla ändamål , även kommersiellt .
på följande villkor :
Erkännande ( BY ) - Du måste nämna källan InfoFinland.fi .
Ange en länk till webbplatsen InfoFinland.fi och nämn licensen CC BY 4.0 .
Ange om bearbetningar är gjorda .
du behöver göra så i enlighet med god sed , och inte på ett sätt som ger en bild av att InfoFinland stödjer dig eller ditt användande .
Inga ytterligare begränsningar - Du får inte tillämpa lagliga begränsningar eller teknologiska metoder som juridiskt begränsar andra från att gör något som licensen tillåter .
Erkännande 4.0 Internationellfinska _ svenska _ engelska _ ryska _ franska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ japanska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ grekiska
_ tjeckiska
öppet programmeringsgränssnitt ( API )
Vi erbjuder allt textinnehåll i InfoFinland via ett öppet programmeringsgränssnitt ( API ) .
med hjälp av gränssnittet kan du visa InfoFinlands innehåll på andra webbplatser eller skapa olika applikationer .
information om gränssnittetfinska _ engelska
öppet programmeringsgränssnittfinska
Användning av InfoFinland @-@ texterna på andra ställen
texterna ur webbtjänsten InfoFinland.fi används i följande tjänster :
linkkiArbets- och näringsministeriet :
guiden Välkommen till Finland ( pdf , 3,40 MB ) finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
Medlemskommunerna har själv hand om översättningen av de övriga kommunsidorna .
Översättningsanvisning :
Översättningsanvisningen är på finska .
Översättningsanvisning :
Översättningsanvisningen är på finska .
Översättningsanvisning :
Översättningsanvisningen är på finska .
trafik
beslutsfattande och påverkan
religion
grundläggande information
historia
trafik
huvudstadsregionen har goda kollektivtrafikförbindelser .
i Grankulla finns en järnvägsstation och i staden finns många busslinjer .
du kan söka information om rutterna i tjänsten Reseplaneraren .
tjänsten ger dig förslag på olika kollektivtrafikförbindelser från ett ställe till ett annat .
Reseplanerarefinska _ svenska _ engelska _ ryska
inom kollektivtrafiken kan du betala med kontanter eller resekort .
i närtågen måste du köpa biljetten i förväg .
du kan köpa resekortet på Grankulla stadshus .
du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat .
stadshuset
Grankullavägen 10
mån @-@ fre kl . 8.00 @-@ 15.00 ; tis , ons , tors även kl . 17.00 @-@ 19.30
den närmaste flygstationen är Helsingfors @-@ Vanda flygplats .
Flygplatsenfinska _ svenska _ engelska _ ryska _ kinesiska
Läs mer :
trafiken i Finland .
beslutsfattande och påverkan
i Grankulla beslutas ärenden av stadsfullmäktige .
i stadsfullmäktige sitter 35 ledamöter som representerar olika politiska grupper .
Fullmäktige väljs var fjärde år genom kommunalval .
på Grankulla stads webbplats kan du skicka respons till förvaltningen .
du kan också lämna initiativ och ställa frågor samt kommentera ärenden på finska och på svenska .
även engelskspråkiga frågor besvaras .
delta och påverkafinska _ svenska
religion
många religiösa samfund är verksamma i Esbo och Helsingfors .
i tjänsten Uskonnot Suomessa kan du söka information enligt det religiösa samfundet och orten .
religiösa samfundfinska _ engelska
linkkiHelsingfors ortodoxa församling :
ortodoxa församlingenfinska _ ryska
i Grankulla finns en evangelisk @-@ luthersk kyrka med två församlingar , en finskspråkig och en svenskspråkig .
församlingarfinska _ svenska
Läs mer : kulturer och religioner i Finland .
grundläggande information
Grankulla är en av de fyra kommunerna i huvudstadsregionen .
den ligger mitt i Esbo , 15 kilometer västerut från Helsingfors .
Grankulla har cirka 9.600 invånare , varav 60 procent har finska , 36 procent svenska och 4 procent ett annat språk som modersmål .
Grankullas areal är 6,0 km2 .
information om stadenfinska _ svenska _ engelska
historia
år 1906 grundades ett aktiebolag i Grankulla som sålde villatomter till invånarna i huvudstadsregionen .
området hade en direkt förbindelse till Helsingfors .
år 1920 blev villasamhället en köping .
till en början var största delen av invånarna svenskspråkiga .
år 1972 fick köpingen stadsrättigheter .
Nätmuseetfinska _ svenska
trafik
beslutsfattande och påverkan
religion
grundläggande information
historia
trafik
huvudstadsregionen har goda kollektivtrafikförbindelser .
i Grankulla finns en järnvägsstation och i staden finns många busslinjer .
du kan söka information om rutterna i tjänsten Reseplaneraren .
tjänsten ger dig förslag på olika kollektivtrafikförbindelser från ett ställe till ett annat .
Reseplanerarefinska _ svenska _ engelska _ ryska
inom kollektivtrafiken kan du betala med kontanter eller resekort .
i närtågen måste du köpa biljetten i förväg .
du kan köpa resekortet på Grankulla stadshus .
du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat .
stadshuset
Grankullavägen 10
mån @-@ fre kl . 8.00 @-@ 15.00 ; tis , ons , tors även kl . 17.00 @-@ 19.30
den närmaste flygstationen är Helsingfors @-@ Vanda flygplats .
Flygplatsenfinska _ svenska _ engelska _ ryska _ kinesiska
Läs mer :
trafiken i Finland .
beslutsfattande och påverkan
i Grankulla beslutas ärenden av stadsfullmäktige .
i stadsfullmäktige sitter 35 ledamöter som representerar olika politiska grupper .
Fullmäktige väljs var fjärde år genom kommunalval .
på Grankulla stads webbplats kan du skicka respons till förvaltningen .
du kan också lämna initiativ och ställa frågor samt kommentera ärenden på finska och på svenska .
även engelskspråkiga frågor besvaras .
delta och påverkafinska _ svenska
religion
många religiösa samfund är verksamma i Esbo och Helsingfors .
i tjänsten Uskonnot Suomessa kan du söka information enligt det religiösa samfundet och orten .
religiösa samfundfinska _ engelska
linkkiHelsingfors ortodoxa församling :
ortodoxa församlingenfinska _ ryska
i Grankulla finns en evangelisk @-@ luthersk kyrka med två församlingar , en finskspråkig och en svenskspråkig .
församlingarfinska _ svenska
Läs mer : kulturer och religioner i Finland .
grundläggande information
Grankulla är en av de fyra kommunerna i huvudstadsregionen .
den ligger mitt i Esbo , 15 kilometer västerut från Helsingfors .
Grankulla har cirka 9.600 invånare , varav 60 procent har finska , 36 procent svenska och 4 procent ett annat språk som modersmål .
Grankullas areal är 6,0 km2 .
information om stadenfinska _ svenska _ engelska
historia
år 1906 grundades ett aktiebolag i Grankulla som sålde villatomter till invånarna i huvudstadsregionen .
området hade en direkt förbindelse till Helsingfors .
år 1920 blev villasamhället en köping .
till en början var största delen av invånarna svenskspråkiga .
år 1972 fick köpingen stadsrättigheter .
Nätmuseetfinska _ svenska
trafik
beslutsfattande och påverkan
religion
grundläggande information
historia
trafik
huvudstadsregionen har goda kollektivtrafikförbindelser .
i Grankulla finns en järnvägsstation och i staden finns många busslinjer .
du kan söka information om rutterna i tjänsten Reseplaneraren .
tjänsten ger dig förslag på olika kollektivtrafikförbindelser från ett ställe till ett annat .
Reseplanerarefinska _ svenska _ engelska
inom kollektivtrafiken kan du betala med kontanter eller resekort .
i närtågen måste du köpa biljetten i förväg .
du kan köpa resekortet på Grankulla stadshus .
du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat .
stadshuset
Grankullavägen 10
mån @-@ fre kl . 8.00 @-@ 15.00 ; tis , ons , tors även kl . 17.00 @-@ 19.30
den närmaste flygstationen är Helsingfors @-@ Vanda flygplats .
Flygplatsenfinska _ svenska _ engelska _ ryska _ kinesiska
Läs mer :
trafiken i Finland .
beslutsfattande och påverkan
i Grankulla beslutas ärenden av stadsfullmäktige .
i stadsfullmäktige sitter 35 ledamöter som representerar olika politiska grupper .
Fullmäktige väljs var fjärde år genom kommunalval .
på Grankulla stads webbplats kan du skicka respons till förvaltningen .
du kan också lämna initiativ och ställa frågor samt kommentera ärenden på finska och på svenska .
även engelskspråkiga frågor besvaras .
delta och påverkafinska _ svenska
religion
många religiösa samfund är verksamma i Esbo och Helsingfors .
i tjänsten Uskonnot Suomessa kan du söka information enligt det religiösa samfundet och orten .
religiösa samfundfinska _ engelska
linkkiHelsingfors ortodoxa församling :
ortodoxa församlingenfinska _ ryska
i Grankulla finns en evangelisk @-@ luthersk kyrka med två församlingar , en finskspråkig och en svenskspråkig .
församlingarfinska _ svenska
Läs mer : kulturer och religioner i Finland .
grundläggande information
Grankulla är en av de fyra kommunerna i huvudstadsregionen .
den ligger mitt i Esbo , 15 kilometer västerut från Helsingfors .
Grankulla har cirka 9.600 invånare , varav 60 procent har finska , 36 procent svenska och 4 procent ett annat språk som modersmål .
Grankullas areal är 6,0 km2 .
information om stadenfinska _ svenska _ engelska
historia
år 1906 grundades ett aktiebolag i Grankulla som sålde villatomter till invånarna i huvudstadsregionen .
området hade en direkt förbindelse till Helsingfors .
år 1920 blev villasamhället en köping .
till en början var största delen av invånarna svenskspråkiga .
år 1972 fick köpingen stadsrättigheter .
Nätmuseetfinska _ svenska
evenemang
bibliotek
Fritidsverksamhet för barn och unga
föreningar
evenemang
evenemang i Grankullafinska _ svenska _ engelska
vid medborgarinstitutet kan man till exempel skapa konst , göra handarbeten , laga mat , dansa eller motionera .
man kan även studera språk .
Medborgarinstitutetfinska _ svenska _ engelska
vid musikinstitutet kan man musicera .
information om Musikinstitutetfinska _ svenska
Grankulla stad ordnar mångsidig kulturverksamhet .
Kulturtjänsterfinska _ svenska _ engelska
i staden finns också många idrottsmöjligheter .
Idrottstjänsterfinska _ svenska _ engelska
det finns en biograf i Grankulla .
linkkiBio Grani :
Biograffinska
Läs mer : Fritid .
bibliotek
på Grankulla stadsbibliotek kan du låna böcker , tidningar , musik , filmer , spel och mycket annat .
i biblioteket kan du också använda dator .
Stadsbiblioteketfinska _ svenska _ engelska
huvudstadsregionens gemensamma bibliotekstjänstfinska _ svenska _ engelska _ somaliska _ persiska _ arabiska
Läs mer : bibliotek
Flerspråkiga biblioteket
Flerspråkiga biblioteket ligger i Böle i Helsingfors
här finns böcker , musik , tidningar och tidskrifter samt ljudböcker på flera olika språk .
du kan åka till Böle eller beställa material till ditt eget närbibliotek .
linkkiHelsingfors stadsbibliotek :
Flerspråkiga biblioteketfinska _ svenska _ engelska
hobbyer för barn och unga
barn och ungdomar kan studera musik vid Grankulla musikinstitut och bildkonst vid Grankulla konstskola .
i Grankulla kan man också motionera på många olika sätt .
på Grankulla ungdomsgård ordnas många olika slags verksamheter .
Ungdomsgårdenfinska _ svenska _ engelska
Läs mer : hobbyer för barn och unga
föreningar
i Grankulla finns många olika föreningar , till exempel kulturföreningar och idrottsklubbar .
Föreningarfinska _ svenska
Läs mer : föreningar .
Läs mer : Fritid i Esbo
evenemang
bibliotek
Fritidsverksamhet för barn och unga
föreningar
evenemang
evenemang i Grankullafinska _ svenska _ engelska
vid medborgarinstitutet kan man till exempel skapa konst , göra handarbeten , laga mat , dansa eller motionera .
man kan även studera språk .
Medborgarinstitutetfinska _ svenska _ engelska
vid musikinstitutet kan man musicera .
information om Musikinstitutetfinska _ svenska
Grankulla stad ordnar mångsidig kulturverksamhet .
Kulturtjänsterfinska _ svenska _ engelska
i staden finns också många idrottsmöjligheter .
Idrottstjänsterfinska _ svenska _ engelska
det finns en biograf i Grankulla .
linkkiBio Grani :
Biograffinska
Läs mer : Fritid .
bibliotek
på Grankulla stadsbibliotek kan du låna böcker , tidningar , musik , filmer , spel och mycket annat .
i biblioteket kan du också använda dator .
Stadsbiblioteketfinska _ svenska _ engelska
huvudstadsregionens gemensamma bibliotekstjänstfinska _ svenska _ engelska _ somaliska _ persiska _ arabiska
Läs mer : bibliotek
Flerspråkiga biblioteket
Flerspråkiga biblioteket ligger i Böle i Helsingfors
här finns böcker , musik , tidningar och tidskrifter samt ljudböcker på flera olika språk .
du kan åka till Böle eller beställa material till ditt eget närbibliotek .
linkkiHelsingfors stadsbibliotek :
Flerspråkiga biblioteketfinska _ svenska _ engelska
hobbyer för barn och unga
barn och ungdomar kan studera musik vid Grankulla musikinstitut och bildkonst vid Grankulla konstskola .
i Grankulla kan man också motionera på många olika sätt .
på Grankulla ungdomsgård ordnas många olika slags verksamheter .
Ungdomsgårdenfinska _ svenska _ engelska
Läs mer : hobbyer för barn och unga
föreningar
i Grankulla finns många olika föreningar , till exempel kulturföreningar och idrottsklubbar .
Föreningarfinska _ svenska
Läs mer : föreningar .
Läs mer : Fritid i Esbo
evenemang
bibliotek
Fritidsverksamhet för barn och unga
föreningar
evenemang
evenemang i Grankullafinska _ svenska _ engelska
vid medborgarinstitutet kan man till exempel skapa konst , göra handarbeten , laga mat , dansa eller motionera .
man kan även studera språk .
Medborgarinstitutetfinska _ svenska _ engelska
vid musikinstitutet kan man musicera .
information om Musikinstitutetfinska _ svenska
Grankulla stad ordnar mångsidig kulturverksamhet .
Kulturtjänsterfinska _ svenska _ engelska
i staden finns också många idrottsmöjligheter .
Idrottstjänsterfinska _ svenska _ engelska
det finns en biograf i Grankulla .
linkkiBio Grani :
Biograffinska
Läs mer : Fritid .
bibliotek
på Grankulla stadsbibliotek kan du låna böcker , tidningar , musik , filmer , spel och mycket annat .
i biblioteket kan du också använda dator .
Stadsbiblioteketfinska _ svenska _ engelska
huvudstadsregionens gemensamma bibliotekstjänstfinska _ svenska _ engelska _ somaliska _ persiska _ arabiska
Läs mer : bibliotek
Flerspråkiga biblioteket
Flerspråkiga biblioteket ligger i Böle i Helsingfors
här finns böcker , musik , tidningar och tidskrifter samt ljudböcker på flera olika språk .
du kan åka till Böle eller beställa material till ditt eget närbibliotek .
linkkiHelsingfors stadsbibliotek :
Flerspråkiga biblioteketfinska _ svenska _ engelska
hobbyer för barn och unga
barn och ungdomar kan studera musik vid Grankulla musikinstitut och bildkonst vid Grankulla konstskola .
i Grankulla kan man också motionera på många olika sätt .
på Grankulla ungdomsgård ordnas många olika slags verksamheter .
Ungdomsgårdenfinska _ svenska _ engelska
Läs mer : hobbyer för barn och unga
föreningar
i Grankulla finns många olika föreningar , till exempel kulturföreningar och idrottsklubbar .
Föreningarfinska _ svenska
Läs mer : föreningar .
Läs mer : Fritid i Esbo
social- och krisjouren
problem med uppehållstillstånd
brott
våld
problem i äktenskap och parförhållande
behöver du juristhjälp ? barns och ungas problem
Död
ring nödnumret 112 om det är fråga om en nödsituation .
via nödnumret kan du tillkalla polis , ambulans eller brandkår .
ring inte nödnumret om det inte är en nödsituation .
social- och krisjouren
social- och krisjouren vid Jorv sjukhus i Esbo hjälper dygnet runt om du eller din familj behöver hjälp i en akut krissituation , till exempel vid våld , problem med barnen eller psykiska problem .
i krissituationer kan du ringa eller åka till jouren .
Esbo social- och krisjour
Jorv sjukhus , Åbovägen 150 , Esbo
tfn ( 09 ) 816.42439
vardagar kl . 15 @-@ 08 , fre @-@ sön och helgdagar dygnet runt
linkkiEsbo stad :
social- och krisjourenfinska _ svenska _ engelska
linkkiFöreningen för mental hälsa i Finland :
krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
problem med uppehållstillstånd
om du har problem med eller det råder oklarheter kring uppehållstillståndet kan du ta kontakt med Migrationsverket , Flyktingrådgivningen eller Helsingfors stads Helsinki @-@ info .
Läs mer : problem med uppehållstillstånd
information om uppehållstillståndfinska _ svenska _ engelska
linkkiFlyktingrådgivningen r.f. :
rättshjälp till flyktingarfinska _ svenska _ engelska
Helsingfors @-@ infofinska _ svenska _ engelska
brott
om du blir utsatt för ett brott , gör en brottsanmälan hos polisen .
du kan göra brottsanmälan på internet .
du kan även fylla i en blankett och lämna den till Esbo huvudpolisstation .
Esbo huvudpolisstation
Knektbrovägen 4
Läs mer : brott
kontaktuppgifterfinska _ svenska _ engelska
elektronisk polisanmälanfinska _ svenska _ engelska
behöver du en jurist ?
Västra Nylands rättshjälpsbyrå betjänar invånarna i Grankulla .
Västra Nylands rättshjälpsbyrå
Östanvindsvägen 1 A
tfn 029.56.61820 .
linkkiVästra Nylands rättshjälpsbyrå :
Läs mer :
behöver du en jurist ?
våld
om du behöver brådskande hjälp av polisen i nödsituationer , ring nödnumret 112 .
om någon i din familj utövar våld mot dig eller hotar dig med våld , kontakta ett skyddshem .
tfn ( 09 ) 4777.180 ( 24h )
hjälp till offer för familjevåldfinska
föreningen Monika @-@ Naiset Liitto har en jourtelefon för invandrarkvinnor som blivit utsatta för våld .
tfn 0800.05058
hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
invandrarmän som har problem med våld kan få hjälp via tjänsten Miehen linja .
tfn ( 09 ) 276.62899
hjälp för invandrarmänfinska _ engelska
Läs mer : våld
problem i äktenskap och parförhållande
vid problem i äktenskap och parförhållande kan du få hjälp vid familjerådgivningen .
familjerådgivningen betjänar invånarna i Grankulla .
familjerådgivningen
tfn ( 09 ) 5056.297
familjerådgivningfinska _ svenska
problem i äktenskap och parförhållande
barns och ungas problem
vid problem som gäller barn under skolåldern , kontakta barnrådgivningen .
barnrådgivningen
tfn ( 09 ) 5056.357 eller ( 09 ) 5056.358
Rådgivningsbyråerfinska _ svenska _ engelska
vid problem som gäller barn i skolåldern hjälper till exempel skolans hälsovårdare .
skolhälsovårdenfinska _ svenska
om du behöver råd i frågor kring barns psykiska tillväxt och utveckling , kan du boka en tid hos familjerådgivningen .
familjerådgivningfinska _ svenska
du kan prata om dina problem med skolans eller läroanstaltens hälsovårdare eller de vuxna vid ungdomsgården .
den unga själv eller föräldrarna kan också kontakta familjerådgivningen .
en ung som inte är trygg i sitt eget hem kan kontakta Finlands Röda Kors De ungas skyddshus .
skyddshuset finns i Stensvik .
de ungas skyddshus
tfn ( 09 ) 8195.5360
linkkiFinlands Röda Kors :
de ungas skyddshusfinska
Läs mer : barns och ungas problem
Död
om en nära anhörig till dig avlider oväntat , kan du få stöd av Grankullas grupp för krisbearbetning , tfn 050.344.6652 .
Grankulla stad har en egen begravningsplats i Kasabergsområdet .
den är avsedd för stadens invånare .
Läs mer : Död
social- och krisjouren
problem med uppehållstillstånd
brott
våld
problem i äktenskap och parförhållande
behöver du juristhjälp ? barns och ungas problem
Död
ring nödnumret 112 om det är fråga om en nödsituation .
via nödnumret kan du tillkalla polis , ambulans eller brandkår .
ring inte nödnumret om det inte är en nödsituation .
social- och krisjouren
social- och krisjouren vid Jorv sjukhus i Esbo hjälper dygnet runt om du eller din familj behöver hjälp i en akut krissituation , till exempel vid våld , problem med barnen eller psykiska problem .
i krissituationer kan du ringa eller åka till jouren .
Esbo social- och krisjour
Jorv sjukhus , Åbovägen 150 , Esbo
tfn ( 09 ) 816.42439
vardagar kl . 15 @-@ 08 , fre @-@ sön och helgdagar dygnet runt
linkkiEsbo stad :
social- och krisjourenfinska _ svenska _ engelska
linkkiFöreningen för mental hälsa i Finland :
krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
problem med uppehållstillstånd
om du har problem med eller det råder oklarheter kring uppehållstillståndet kan du ta kontakt med Migrationsverket , Flyktingrådgivningen eller Helsingfors stads Helsinki @-@ info .
Läs mer : problem med uppehållstillstånd
information om uppehållstillståndfinska _ svenska _ engelska
linkkiFlyktingrådgivningen r.f. :
rättshjälp till flyktingarfinska _ svenska _ engelska
Helsingfors @-@ infofinska _ svenska _ engelska
brott
om du blir utsatt för ett brott , gör en brottsanmälan hos polisen .
du kan göra brottsanmälan på internet .
du kan även fylla i en blankett och lämna den till Esbo huvudpolisstation .
Esbo huvudpolisstation
Knektbrovägen 4
Läs mer : brott
kontaktuppgifterfinska _ svenska _ engelska
elektronisk polisanmälanfinska _ svenska _ engelska
behöver du en jurist ?
Västra Nylands rättshjälpsbyrå betjänar invånarna i Grankulla .
Västra Nylands rättshjälpsbyrå
Östanvindsvägen 1 A
tfn 029.56.61820 .
linkkiVästra Nylands rättshjälpsbyrå :
Läs mer :
behöver du en jurist ?
våld
om du behöver brådskande hjälp av polisen i nödsituationer , ring nödnumret 112 .
om någon i din familj utövar våld mot dig eller hotar dig med våld , kontakta ett skyddshem .
tfn ( 09 ) 4777.180 ( 24h )
hjälp till offer för familjevåldfinska
föreningen Monika @-@ Naiset Liitto har en jourtelefon för invandrarkvinnor som blivit utsatta för våld .
tfn 0800.05058
hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
invandrarmän som har problem med våld kan få hjälp via tjänsten Miehen linja .
tfn ( 09 ) 276.62899
hjälp för invandrarmänfinska _ engelska
Läs mer : våld
problem i äktenskap och parförhållande
vid problem i äktenskap och parförhållande kan du få hjälp vid familjerådgivningen .
familjerådgivningen betjänar invånarna i Grankulla .
familjerådgivningen
tfn ( 09 ) 5056.297
familjerådgivningfinska _ svenska
problem i äktenskap och parförhållande
barns och ungas problem
vid problem som gäller barn under skolåldern , kontakta barnrådgivningen .
barnrådgivningen
tfn ( 09 ) 5056.357 eller ( 09 ) 5056.358
Rådgivningsbyråerfinska _ svenska _ engelska
vid problem som gäller barn i skolåldern hjälper till exempel skolans hälsovårdare .
skolhälsovårdenfinska _ svenska
om du behöver råd i frågor kring barns psykiska tillväxt och utveckling , kan du boka en tid hos familjerådgivningen .
familjerådgivningfinska _ svenska
du kan prata om dina problem med skolans eller läroanstaltens hälsovårdare eller de vuxna vid ungdomsgården .
den unga själv eller föräldrarna kan också kontakta familjerådgivningen .
en ung som inte är trygg i sitt eget hem kan kontakta Finlands Röda Kors De ungas skyddshus .
skyddshuset finns i Stensvik .
de ungas skyddshus
tfn ( 09 ) 8195.5360
linkkiFinlands Röda Kors :
de ungas skyddshusfinska
Läs mer : barns och ungas problem
Död
om en nära anhörig till dig avlider oväntat , kan du få stöd av Grankullas grupp för krisbearbetning , tfn 050.344.6652 .
Grankulla stad har en egen begravningsplats i Kasabergsområdet .
den är avsedd för stadens invånare .
Läs mer : Död
social- och krisjouren
problem med uppehållstillstånd
brott
våld
problem i äktenskap och parförhållande
behöver du juristhjälp ? barns och ungas problem
Död
ring nödnumret 112 om det är fråga om en nödsituation .
via nödnumret kan du tillkalla polis , ambulans eller brandkår .
ring inte nödnumret om det inte är en nödsituation .
social- och krisjouren
social- och krisjouren vid Jorv sjukhus i Esbo hjälper dygnet runt om du eller din familj behöver hjälp i en akut krissituation , till exempel vid våld , problem med barnen eller psykiska problem .
i krissituationer kan du ringa eller åka till jouren .
Esbo social- och krisjour
Jorv sjukhus , Åbovägen 150 , Esbo
tfn ( 09 ) 816.42439
vardagar kl . 15 @-@ 08 , fre @-@ sön och helgdagar dygnet runt
linkkiEsbo stad :
social- och krisjourenfinska _ svenska _ engelska
linkkiFöreningen för mental hälsa i Finland :
krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
problem med uppehållstillstånd
om du har problem med eller det råder oklarheter kring uppehållstillståndet kan du ta kontakt med Migrationsverket , Flyktingrådgivningen eller Helsingfors stads Helsinki @-@ info .
Läs mer : problem med uppehållstillstånd
information om uppehållstillståndfinska _ svenska _ engelska
linkkiFlyktingrådgivningen r.f. :
rättshjälp till flyktingarfinska _ svenska _ engelska
Helsingfors @-@ infofinska _ svenska _ engelska
brott
om du blir utsatt för ett brott , gör en brottsanmälan hos polisen .
du kan göra brottsanmälan på internet .
du kan även fylla i en blankett och lämna den till Esbo huvudpolisstation .
Esbo huvudpolisstation
Knektbrovägen 4
Läs mer : brott
kontaktuppgifterfinska _ svenska _ engelska
elektronisk polisanmälanfinska _ svenska _ engelska
behöver du en jurist ?
Västra Nylands rättshjälpsbyrå betjänar invånarna i Grankulla .
Västra Nylands rättshjälpsbyrå
Östanvindsvägen 1 A
tfn 029.56.61820 .
linkkiVästra Nylands rättshjälpsbyrå :
Läs mer :
behöver du en jurist ?
våld
om du behöver brådskande hjälp av polisen i nödsituationer , ring nödnumret 112 .
om någon i din familj utövar våld mot dig eller hotar dig med våld , kontakta ett skyddshem .
tfn ( 09 ) 4777.180 ( 24h )
hjälp till offer för familjevåldfinska
föreningen Monika @-@ Naiset Liitto har en jourtelefon för invandrarkvinnor som blivit utsatta för våld .
tfn 0800.05058
hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
invandrarmän som har problem med våld kan få hjälp via tjänsten Miehen linja .
tfn ( 09 ) 276.62899
hjälp för invandrarmänfinska _ engelska
Läs mer : våld
problem i äktenskap och parförhållande
vid problem i äktenskap och parförhållande kan du få hjälp vid familjerådgivningen .
familjerådgivningen betjänar invånarna i Grankulla .
familjerådgivningen
tfn ( 09 ) 5056.297
familjerådgivningfinska _ svenska
problem i äktenskap och parförhållande
barns och ungas problem
vid problem som gäller barn under skolåldern , kontakta barnrådgivningen .
barnrådgivningen
tfn ( 09 ) 5056.357 eller ( 09 ) 5056.358
Rådgivningsbyråerfinska _ svenska _ engelska
vid problem som gäller barn i skolåldern hjälper till exempel skolans hälsovårdare .
skolhälsovårdenfinska _ svenska
om du behöver råd i frågor kring barns psykiska tillväxt och utveckling , kan du boka en tid hos familjerådgivningen .
familjerådgivningfinska _ svenska
du kan prata om dina problem med skolans eller läroanstaltens hälsovårdare eller de vuxna vid ungdomsgården .
den unga själv eller föräldrarna kan också kontakta familjerådgivningen .
en ung som inte är trygg i sitt eget hem kan kontakta Finlands Röda Kors De ungas skyddshus .
skyddshuset finns i Stensvik .
de ungas skyddshus
tfn ( 09 ) 8195.5360
linkkiFinlands Röda Kors :
de ungas skyddshusfinska
Läs mer : barns och ungas problem
Död
om en nära anhörig till dig avlider oväntat , kan du få stöd av Grankullas grupp för krisbearbetning , tfn 050.344.6652 .
Grankulla stad har en egen begravningsplats i Kasabergsområdet .
den är avsedd för stadens invånare .
Läs mer : Död
äktenskap
skilsmässa
barn vid skilsmässa
vård av barnet
äktenskap
före äktenskapet ska du skriftligt begära prövning av hinder mot äktenskap .
Hindersprövningen görs i magistraten .
Läs mer : prövning av hinder mot äktenskap , Äktenskap
kontaktuppgifter till magistratfinska _ svenska _ engelska
skilsmässa
kvinnan eller mannen kan lämna in skilsmässoansökan i Västra Nylands tingsrätts kansli .
du kan också söka skilsmässa ensam , utan din makes eller makas samtycke .
du kan skicka in ansökan till tingsrättens kansli per post , fax eller via e @-@ post .
Västra Nylands tingsrätt
tfn 029.5645.000
Läs mer : skilsmässa
linkkiVästra Nylands tingsrätt :
kontaktuppgifterfinska _ svenska
barn vid skilsmässa
om du har barn och ska skilja dig , ta kontakt med barnatillsyningsmannen .
Socialväsendet bekräftar ett avtal om barnens boende , vårdnad , umgängesrätt och underhållsbidrag .
Läs mer : barn vid skilsmässa
vårdnad om barn och umgängesrättfinska _ svenska
vård av barnet
på InfoFinlands sida Utbildning i Grankulla finns information om dagvård för barn .
vård av barnet i hemmet
om du sköter ditt barn hemma kan du delta i Grankulla stads öppna familjeverksamhet . där kan du träffa andra barnfamiljer .
Läs mer : stöd för vård av barn i hemmet
öppen familjeverksamhetfinska _ svenska
stöd för hemvård av barnfinska _ svenska
äktenskap
skilsmässa
barn vid skilsmässa
vård av barnet
äktenskap
före äktenskapet ska du skriftligt begära prövning av hinder mot äktenskap .
Hindersprövningen görs i magistraten .
Läs mer : prövning av hinder mot äktenskap , Äktenskap
kontaktuppgifter till magistratfinska _ svenska _ engelska
skilsmässa
kvinnan eller mannen kan lämna in skilsmässoansökan i Västra Nylands tingsrätts kansli .
du kan också söka skilsmässa ensam , utan din makes eller makas samtycke .
du kan skicka in ansökan till tingsrättens kansli per post , fax eller via e @-@ post .
Västra Nylands tingsrätt
tfn 029.5645.000
Läs mer : skilsmässa
linkkiVästra Nylands tingsrätt :
kontaktuppgifterfinska _ svenska
barn vid skilsmässa
om du har barn och ska skilja dig , ta kontakt med barnatillsyningsmannen .
Socialväsendet bekräftar ett avtal om barnens boende , vårdnad , umgängesrätt och underhållsbidrag .
Läs mer : barn vid skilsmässa
vårdnad om barn och umgängesrättfinska _ svenska
vård av barnet
på InfoFinlands sida Utbildning i Grankulla finns information om dagvård för barn .
vård av barnet i hemmet
om du sköter ditt barn hemma kan du delta i Grankulla stads öppna familjeverksamhet . där kan du träffa andra barnfamiljer .
Läs mer : stöd för vård av barn i hemmet
öppen familjeverksamhetfinska _ svenska
stöd för hemvård av barnfinska _ svenska
äktenskap
skilsmässa
barn vid skilsmässa
vård av barnet
äktenskap
före äktenskapet ska du skriftligt begära prövning av hinder mot äktenskap .
Hindersprövningen görs i magistraten .
Läs mer : prövning av hinder mot äktenskap , Äktenskap
kontaktuppgifter till magistratfinska _ svenska _ engelska
skilsmässa
kvinnan eller mannen kan lämna in skilsmässoansökan i Västra Nylands tingsrätts kansli .
du kan också söka skilsmässa ensam , utan din makes eller makas samtycke .
du kan skicka in ansökan till tingsrättens kansli per post , fax eller via e @-@ post .
Västra Nylands tingsrätt
tfn 029.5645.000
Läs mer : skilsmässa
linkkiVästra Nylands tingsrätt :
kontaktuppgifterfinska _ svenska
barn vid skilsmässa
om du har barn och ska skilja dig , ta kontakt med barnatillsyningsmannen .
Socialväsendet bekräftar ett avtal om barnens boende , vårdnad , umgängesrätt och underhållsbidrag .
Läs mer : barn vid skilsmässa
vårdnad om barn och umgängesrättfinska _ svenska
vård av barnet
på InfoFinlands sida Utbildning i Grankulla finns information om dagvård för barn .
vård av barnet i hemmet
om du sköter ditt barn hemma kan du delta i Grankulla stads öppna familjeverksamhet . där kan du träffa andra barnfamiljer .
Läs mer : stöd för vård av barn i hemmet
öppen familjeverksamhetfinska _ svenska
stöd för hemvård av barnfinska _ svenska
hälsovårdstjänsterna i Grankulla
barns hälsa
äldre människors hälsa
tandvård
mental hälsa
Sexualhälsa
när du väntar barn
handikappade personer
ring nödnumret 112 om det är fråga om en brådskande nödsituation .
ring nödnumret till exempel vid en allvarlig olycka eller när någon drabbas av en sjukdomsattack .
ring inte nödnumret om det inte är en nödsituation .
om du har din hemkommun i Grankulla , kan du utnyttja de offentliga hälso- och sjukvårdstjänsterna .
offentliga hälso- och sjukvårdstjänster tillhandahålls till exempel vid hälsostationer , tandkliniker , rådgivningsbyråer och sjukhus .
om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna , kan du söka dig till en privat läkarstation .
på en privat läkarstation måste du betala samtliga kostnader själv .
Läs mer : hälsa
hälsovårdstjänsterna i Grankulla
i Grankulla tillhandahålls offentliga hälso- och sjukvårdstjänster på hälsostationen .
på hälsostationen finns läkarens , sjukskötarens och hälsovårdarens mottagningar .
hälsostationen har öppet vardagar kl . 8.00 @-@ 16.00 .
om du behöver vård under samma dag ska du kontakta hälsostationen direkt på morgonen när hälsostationen öppnar .
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
tfn ( 09 ) 8789.1300
Hälsostationenfinska _ svenska _ engelska
privata hälsotjänster
information om privata hälsotjänster hittar du på sidorna Hälsa i Esbo och Hälsa i Helsingfors .
läkemedel
du kan köpa läkemedel på apoteket .
adressen till apoteket i Grankulla är Kyrkovägen 15 , Grankulla .
Läs mer : läkemedel .
Apotekfinska _ svenska
linkkiApotekareförbundet :
hälsovård för papperslösa
i Helsingfors finns Global Clinic , där personer som vistas i Finland utan tillstånd kan få primärvård .
tfn 044.977.4547
kontaktuppgifterfinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Läs mer : hälsovårdstjänster i Finland
kvällstid och under veckoslut har hälsostationen stängt .
då vårdas akuta sjukdomar och olycksfall på jourmottagningen .
den närmaste jourmottagningen finns vid Jorv sjukhus i Esbo .
ring den kostnadsfria Jourhjälpen på tfn 116.117 innan du kommer till jourmottagningen .
jouren vid Jorv sjukhus
Åbovägen 150
tfn ( 09 ) 4711
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS :
Jourfinska _ svenska _ engelska
Läs mer : hälsovårdstjänster i Finland
barns hälsa
i hälso- och sjukvården av barn under skolåldern får man hjälp av rådgivningens hälsovårdare och läkare .
dem kan du fråga om råd och få stöd i föräldraskapet och fostran av barn .
på rådgivningsbyrån följs barnets hälsa och tillväxt .
Rådgivningsbyråerfinska _ svenska _ engelska
när barnet blir sjukt ska du vid behov kontakta Grankulla hälsostation .
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
tfn ( 09 ) 8789.1300
Hälsostationenfinska _ svenska _ engelska
Skolhälsovårdaren tar hand om skolbarns hälsa .
skolhälsovårdenfinska _ svenska
under kvällar och veckoslut finns jourmottagningen för barn under 16 år vid Jorv sjukhus i Esbo och på Barnkliniken i Helsingfors .
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS :
jourmottagning för barnfinska _ svenska _ engelska
Läs mer : barns hälsa
äldre människors hälsa
om du är över 65 år kan du kontakta seniorrådgivningen vid Grankulla hälsostation .
Seniorrådgivningenfinska _ svenska
Serviceguide för seniorer ( pdf , 1,8 MB ) finska _ svenska
tandvård
Tidsbeställningen till tandkliniken vid Grankulla hälsostation mån @-@ fre :
tfn ( 09 ) 505.6379
jourmottagningen vid Haartmanska sjukhuset har öppet vardagar kl . 14 @-@ 21 och lör @-@ sön kl . 8 @-@ 21 .
tfn ( 09 ) 310.49999
Mun- och tandhälsovårdenfinska _ svenska
privat tandvård
i Grankulla finns också privata tandläkare .
om om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna , kan du gå till en privat tandläkare .
privat tandvård är dyrare än offentlig tandvård .
privat tandläkarefinska _ svenska
Läs mer : tandvård
mental hälsa
om du behöver psykisk hjälp och psykiskt stöd kan du kontakta hälsostationen .
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
tfn ( 09 ) 5056.600
mental hälsafinska _ svenska
Esbo social- och krisjour vid Jorv sjukhus betjänar personer som bor i Grankulla .
i krissituationer kan du ringa eller åka till jouren .
Esbo social- och krisjour
Jorv sjukhus , Åbovägen 150 , Esbo
tfn ( 09 ) 816.42439
vardagar kl . 15 @-@ 08 , fre @-@ sön och helgdagar dygnet runt
Kristjänsterfinska _ svenska
Läs mer : mental hälsa
Sexualhälsa
vid mödra- och preventivrådgivningen får du hjälp med graviditetsprevention och familjeplanering .
könssjukdomar behandlas på hälsostationen och på polikliniken för könssjukdomar i Helsingfors . .
Hälsostationenfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS :
polikliniken för könssjukdomarfinska _ svenska _ engelska
när du väntar barn
vid mödrarådgivningen följs moderns , fostrets och hela familjens hälsotillstånd under graviditeten .
kontakta rådgivningsbyrån när du upptäcker att du är gravid .
tidsbokning vardagar kl . 12 @-@ 13
tfn ( 09 ) 8789.1344
Rådgivningsbyråerfinska _ svenska _ engelska
det närmaste förlossningssjukhuset är Jorv sjukhus i Esbo .
om du vill kan du även föda barnet på något annat sjukhus inom Helsingfors och Nylands sjukvårdsdistrikt ( HNS ) .
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS :
Val av förlossningssjukhusfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt :
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Läs mer : förlossning
handikappade personer
Grankulla stad erbjuder olika tjänster för handikappade , till exempel hjälpmedel och dagverksamhet .
du kan fråga om tjänsterna för handikappade hos socialarbetaren för ditt område .
tjänster inom handikappvårdenfinska _ svenska
Läs mer : handikappade personer
hälsovårdstjänsterna i Grankulla
barns hälsa
äldre människors hälsa
tandvård
mental hälsa
Sexualhälsa
när du väntar barn
handikappade personer
ring nödnumret 112 om det är fråga om en brådskande nödsituation .
ring nödnumret till exempel vid en allvarlig olycka eller när någon drabbas av en sjukdomsattack .
ring inte nödnumret om det inte är en nödsituation .
om du har din hemkommun i Grankulla , kan du utnyttja de offentliga hälso- och sjukvårdstjänsterna .
offentliga hälso- och sjukvårdstjänster tillhandahålls till exempel vid hälsostationer , tandkliniker , rådgivningsbyråer och sjukhus .
om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna , kan du söka dig till en privat läkarstation .
på en privat läkarstation måste du betala samtliga kostnader själv .
Läs mer : hälsa
hälsovårdstjänsterna i Grankulla
i Grankulla tillhandahålls offentliga hälso- och sjukvårdstjänster på hälsostationen .
på hälsostationen finns läkarens , sjukskötarens och hälsovårdarens mottagningar .
hälsostationen har öppet vardagar kl . 8.00 @-@ 16.00 .
om du behöver vård under samma dag ska du kontakta hälsostationen direkt på morgonen när hälsostationen öppnar .
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
tfn ( 09 ) 8789.1300
Hälsostationenfinska _ svenska _ engelska
privata hälsotjänster
information om privata hälsotjänster hittar du på sidorna Hälsa i Esbo och Hälsa i Helsingfors .
läkemedel
du kan köpa läkemedel på apoteket .
adressen till apoteket i Grankulla är Kyrkovägen 15 , Grankulla .
Läs mer : läkemedel .
Apotekfinska _ svenska
linkkiApotekareförbundet :
hälsovård för papperslösa
i Helsingfors finns Global Clinic , där personer som vistas i Finland utan tillstånd kan få primärvård .
tfn 044.977.4547
kontaktuppgifterfinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Läs mer : hälsovårdstjänster i Finland
kvällstid och under veckoslut har hälsostationen stängt .
då vårdas akuta sjukdomar och olycksfall på jourmottagningen .
den närmaste jourmottagningen finns vid Jorv sjukhus i Esbo .
ring den kostnadsfria Jourhjälpen på tfn 116.117 innan du kommer till jourmottagningen .
jouren vid Jorv sjukhus
Åbovägen 150
tfn ( 09 ) 4711
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS :
Jourfinska _ svenska _ engelska
Läs mer : hälsovårdstjänster i Finland
barns hälsa
i hälso- och sjukvården av barn under skolåldern får man hjälp av rådgivningens hälsovårdare och läkare .
dem kan du fråga om råd och få stöd i föräldraskapet och fostran av barn .
på rådgivningsbyrån följs barnets hälsa och tillväxt .
Rådgivningsbyråerfinska _ svenska _ engelska
när barnet blir sjukt ska du vid behov kontakta Grankulla hälsostation .
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
tfn ( 09 ) 8789.1300
Hälsostationenfinska _ svenska _ engelska
Skolhälsovårdaren tar hand om skolbarns hälsa .
skolhälsovårdenfinska _ svenska
under kvällar och veckoslut finns jourmottagningen för barn under 16 år vid Jorv sjukhus i Esbo och på Barnkliniken i Helsingfors .
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS :
jourmottagning för barnfinska _ svenska _ engelska
Läs mer : barns hälsa
äldre människors hälsa
om du är över 65 år kan du kontakta seniorrådgivningen vid Grankulla hälsostation .
information om tjänster för äldrefinska _ svenska
Serviceguide för seniorer ( pdf , 1,8 MB ) finska _ svenska
äldre människor
tandvård
Tidsbeställningen till tandkliniken vid Grankulla hälsostation mån @-@ fre :
tfn ( 09 ) 505.6379
jourmottagningen vid Haartmanska sjukhuset har öppet vardagar kl . 14 @-@ 21 och lör @-@ sön kl . 8 @-@ 21 .
tfn ( 09 ) 310.49999
Mun- och tandhälsovårdenfinska _ svenska
privat tandvård
i Grankulla finns också privata tandläkare .
om om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna , kan du gå till en privat tandläkare .
privat tandvård är dyrare än offentlig tandvård .
privat tandläkarefinska _ svenska
Läs mer : tandvård
mental hälsa
om du behöver psykisk hjälp och psykiskt stöd kan du kontakta hälsostationen .
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
tfn ( 09 ) 5056.600
mental hälsafinska _ svenska
Esbo social- och krisjour vid Jorv sjukhus betjänar personer som bor i Grankulla .
i krissituationer kan du ringa eller åka till jouren .
Esbo social- och krisjour
Jorv sjukhus , Åbovägen 150 , Esbo
tfn ( 09 ) 816.42439
vardagar kl . 15 @-@ 08 , fre @-@ sön och helgdagar dygnet runt
Kristjänsterfinska _ svenska
Läs mer : mental hälsa
Sexualhälsa
vid mödra- och preventivrådgivningen får du hjälp med graviditetsprevention och familjeplanering .
könssjukdomar behandlas på hälsostationen och på polikliniken för könssjukdomar i Helsingfors . .
Hälsostationenfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS :
polikliniken för könssjukdomarfinska _ svenska _ engelska
när du väntar barn
vid mödrarådgivningen följs moderns , fostrets och hela familjens hälsotillstånd under graviditeten .
kontakta rådgivningsbyrån när du upptäcker att du är gravid .
tidsbokning vardagar kl . 12 @-@ 13
tfn ( 09 ) 8789.1344
Rådgivningsbyråerfinska _ svenska _ engelska
det närmaste förlossningssjukhuset är Jorv sjukhus i Esbo .
om du vill kan du även föda barnet på något annat sjukhus inom Helsingfors och Nylands sjukvårdsdistrikt ( HNS ) .
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS :
Val av förlossningssjukhusfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt :
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Läs mer : förlossning
handikappade personer
Grankulla stad erbjuder olika tjänster för handikappade , till exempel hjälpmedel och dagverksamhet .
du kan fråga om tjänsterna för handikappade hos socialarbetaren för ditt område .
tjänster inom handikappvårdenfinska _ svenska
Läs mer : handikappade personer
hälsovårdstjänsterna i Grankulla
barns hälsa
äldre människors hälsa
tandvård
mental hälsa
Sexualhälsa
när du väntar barn
handikappade personer
ring nödnumret 112 om det är fråga om en brådskande nödsituation .
ring nödnumret till exempel vid en allvarlig olycka eller när någon drabbas av en sjukdomsattack .
ring inte nödnumret om det inte är en nödsituation .
om du har din hemkommun i Grankulla , kan du utnyttja de offentliga hälso- och sjukvårdstjänsterna .
offentliga hälso- och sjukvårdstjänster tillhandahålls till exempel vid hälsostationer , tandkliniker , rådgivningsbyråer och sjukhus .
om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna , kan du söka dig till en privat läkarstation .
på en privat läkarstation måste du betala samtliga kostnader själv .
Läs mer : hälsa
hälsovårdstjänsterna i Grankulla
i Grankulla tillhandahålls offentliga hälso- och sjukvårdstjänster på hälsostationen .
på hälsostationen finns läkarens , sjukskötarens och hälsovårdarens mottagningar .
hälsostationen har öppet vardagar kl . 8.00 @-@ 16.00 .
om du behöver vård under samma dag ska du kontakta hälsostationen direkt på morgonen när hälsostationen öppnar .
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
tfn ( 09 ) 8789.1300
Hälsostationenfinska _ svenska
privata hälsotjänster
information om privata hälsotjänster hittar du på sidorna Hälsa i Esbo och Hälsa i Helsingfors .
läkemedel
du kan köpa läkemedel på apoteket .
adressen till apoteket i Grankulla är Kyrkovägen 15 , Grankulla .
Läs mer : läkemedel .
Apotekfinska _ svenska
linkkiApotekareförbundet :
hälsovård för papperslösa
i Helsingfors finns Global Clinic , där personer som vistas i Finland utan tillstånd kan få primärvård .
tfn 044.977.4547
kontaktuppgifterfinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Läs mer : hälsovårdstjänster i Finland
kvällstid och under veckoslut har hälsostationen stängt .
då vårdas akuta sjukdomar och olycksfall på jourmottagningen .
den närmaste jourmottagningen finns vid Jorv sjukhus i Esbo .
ring den kostnadsfria Jourhjälpen på tfn 116.117 innan du kommer till jourmottagningen .
jouren vid Jorv sjukhus
Åbovägen 150
tfn ( 09 ) 4711
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS :
Jourfinska _ svenska _ engelska
Läs mer : hälsovårdstjänster i Finland
barns hälsa
i hälso- och sjukvården av barn under skolåldern får man hjälp av rådgivningens hälsovårdare och läkare .
dem kan du fråga om råd och få stöd i föräldraskapet och fostran av barn .
på rådgivningsbyrån följs barnets hälsa och tillväxt .
Rådgivningsbyråerfinska _ svenska _ engelska
när barnet blir sjukt ska du vid behov kontakta Grankulla hälsostation .
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
tfn ( 09 ) 8789.1300
Hälsostationenfinska _ svenska
Skolhälsovårdaren tar hand om skolbarns hälsa .
skolhälsovårdenfinska _ svenska
under kvällar och veckoslut finns jourmottagningen för barn under 16 år vid Jorv sjukhus i Esbo och på Barnkliniken i Helsingfors .
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS :
jourmottagning för barnfinska _ svenska _ engelska
Läs mer : barns hälsa
äldre människors hälsa
om du är över 65 år kan du kontakta seniorrådgivningen vid Grankulla hälsostation .
information om tjänster för äldrefinska _ svenska
äldre människor
tandvård
Tidsbeställningen till tandkliniken vid Grankulla hälsostation mån @-@ fre :
tfn ( 09 ) 505.6379
jourmottagningen vid Haartmanska sjukhuset har öppet vardagar kl . 14 @-@ 21 och lör @-@ sön kl . 8 @-@ 21 .
tfn ( 09 ) 310.49999
Mun- och tandhälsovårdenfinska _ svenska
privat tandvård
i Grankulla finns också privata tandläkare .
om om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna , kan du gå till en privat tandläkare .
privat tandvård är dyrare än offentlig tandvård .
privat tandläkarefinska _ svenska
Läs mer : tandvård
mental hälsa
om du behöver psykisk hjälp och psykiskt stöd kan du kontakta hälsostationen .
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
tfn ( 09 ) 5056.600
mental hälsafinska _ svenska
Esbo social- och krisjour vid Jorv sjukhus betjänar personer som bor i Grankulla .
i krissituationer kan du ringa eller åka till jouren .
Esbo social- och krisjour
Jorv sjukhus , Åbovägen 150 , Esbo
tfn ( 09 ) 816.42439
vardagar kl . 15 @-@ 08 , fre @-@ sön och helgdagar dygnet runt
Kristjänsterfinska _ svenska
Läs mer : mental hälsa
Sexualhälsa
vid mödra- och preventivrådgivningen får du hjälp med graviditetsprevention och familjeplanering .
könssjukdomar behandlas på hälsostationen och på polikliniken för könssjukdomar i Helsingfors . .
Hälsostationenfinska _ svenska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS :
polikliniken för könssjukdomarfinska _ svenska _ engelska
när du väntar barn
vid mödrarådgivningen följs moderns , fostrets och hela familjens hälsotillstånd under graviditeten .
kontakta rådgivningsbyrån när du upptäcker att du är gravid .
tidsbokning vardagar kl . 12 @-@ 13
tfn ( 09 ) 8789.1344
Rådgivningsbyråerfinska _ svenska _ engelska
det närmaste förlossningssjukhuset är Jorv sjukhus i Esbo .
om du vill kan du även föda barnet på något annat sjukhus inom Helsingfors och Nylands sjukvårdsdistrikt ( HNS ) .
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS :
Val av förlossningssjukhusfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt :
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Läs mer : förlossning
handikappade personer
Grankulla stad erbjuder olika tjänster för handikappade , till exempel hjälpmedel och dagverksamhet .
du kan fråga om tjänsterna för handikappade hos socialarbetaren för ditt område .
tjänster inom handikappvårdenfinska _ svenska
Läs mer : handikappade personer
dagvård
förskoleundervisning
grundläggande utbildning
yrkesutbildning
gymnasium
Högskoleutbildning
andra studiemöjligheter
dagvård
i Grankulla finns stadens egna daghem , privata daghem och privata familjedagvårdare .
dagvård fås på finska och på svenska .
i Grankulla finns också ett engelskspråkigt daghem .
Ansök om dagvårdsplats för ditt barn minst fyra månader innan barnet ska börja i dagvården .
om du ansöker om dagvårdplats för första gången ska du använda den elektroniska ansökan .
du kan också hämta ansökningsblanketten på daghemmet eller vid informationen i stadshuset .
lämna in ansökan till daghemmet eller stadshuset .
familjer som bor i Grankulla kan också söka dagvårdsplats till sitt barn i Esbo , Helsingfors eller Vanda .
du ska ändå lämna in din ansökan i Grankulla .
mer information finns på tjänsten HelsingforsRegionen.fi .
Läs mer : dagvård
dagvård och förskoleundervisningfinska _ svenska _ engelska
ansökan om dagvårdsplatsfinska _ svenska
Engelsk @-@ finskspråkigt daghemfinska _ engelska
Dagvårdens samanvändningsområdefinska _ svenska _ engelska
förskoleundervisning
i Grankulla anordnas förskoleundervisningen i daghemmen .
förskoleundervisningen börjar i augusti och ansökningstiden är i januari .
Läs mer : förskoleundervisning
information om förskoleundervisningenfinska _ svenska _ engelska
grundläggande utbildning
i Grankulla finns både en finsk- och en svenskspråkig grundskola . anmälan till grundskolan ska ske i början av året .
om du har frågor om den grundläggande utbildningen kan du kontakta skolbyrån .
skolbyrån
Grankulla stadshus
Grankullavägen 10
02700 Grankulla
tfn ( 09 ) 50.561 ( växel )
grundläggande utbildning
grundläggande utbildning och gymnasiumfinska _ svenska _ engelska
internationella skolor i huvudstadsregionenfinska
linkkiExpatFinland.fi :
internationella skolor i huvudstadsregionenengelska
yrkesutbildning
de närmaste yrkesläroanstalterna finns i Esbo och Helsingfors .
Läs mer : yrkesutbildning
yrkesutbildningfinska _ engelska
Yrkesinriktad utbildningfinska
gymnasium
i Grankulla finns två gymnasier , ett finskspråkigt och ett svenskspråkigt .
i Esbo finns ett vuxengymnasium där vuxna kan avlägga gymnasiet och studentexamen .
Läs mer : gymnasium
grundläggande utbildning och gymnasiumfinska _ svenska _ engelska
linkkiEsbo stad :
Vuxengymnasietfinska
Högskoleutbildning
i anslutning till folkhögskolan Työväen Akatemia i Grankulla finns en enhet för Humanistiska Yrkeshögskolan , där du kan avlägga yrkeshögskoleexamen för kulturproducenter .
vid yrkeshögskolorna och universiteten i Esbo och Helsingfors kan du studera inom många områden .
mer information om högskolorna i Esbo och Helsingfors hittar du på städernas webbplatser .
Läs mer : Högskoleutbildning
linkkiHumanistiska yrkeshögskolan :
information om Humanistiska yrkeshögskolanfinska _ engelska
linkkiEsbo stad :
Högskolorfinska _ engelska
Högskolorfinska
andra studiemöjligheter
vid Grankulla medborgarinstitut kan du studera till exempel språk , handarbete och matlagning eller delta i ledd motion .
Medborgarinstitutetfinska _ svenska _ engelska
vid Grankulla konstskola kan barn och unga studera bildkonst och vid Grankulla musikinstitut kan barn och vuxna studera musik .
information om Konstskolanfinska _ svenska
information om Musikinstitutetfinska _ svenska
i Grankulla ligger Finska Bibelinstitutet .
vid institutet kan du avlägga enskilda kurser eller studera på någon av institutets studielinjer .
studierna på studielinjerna pågår i 1 @-@ 2 år .
vid bibelinstitutet finns även en studielinje som är särskilt avsedd för invandrare .
Kristliga folkhögskolanfinska _ engelska
folkhögskolan Työväen Akatemia tillhandahåller undervisning inom många akademiska discipliner samt träning för dem som vill läsa på universitet .
information om Työväen Akatemiafinska _ engelska
Läs mer : andra studiemöjligheter
dagvård
förskoleundervisning
grundläggande utbildning
yrkesutbildning
gymnasium
Högskoleutbildning
andra studiemöjligheter
dagvård
i Grankulla finns stadens egna daghem , privata daghem och privata familjedagvårdare .
dagvård fås på finska och på svenska .
i Grankulla finns också ett engelskspråkigt daghem .
Ansök om dagvårdsplats för ditt barn minst fyra månader innan barnet ska börja i dagvården .
om du ansöker om dagvårdplats för första gången ska du använda den elektroniska ansökan .
du kan också hämta ansökningsblanketten på daghemmet eller vid informationen i stadshuset .
lämna in ansökan till daghemmet eller stadshuset .
familjer som bor i Grankulla kan också söka dagvårdsplats till sitt barn i Esbo , Helsingfors eller Vanda .
du ska ändå lämna in din ansökan i Grankulla .
mer information finns på tjänsten HelsingforsRegionen.fi .
Läs mer : dagvård
dagvård och förskoleundervisningfinska _ svenska _ engelska
ansökan om dagvårdsplatsfinska _ svenska
Engelsk @-@ finskspråkigt daghemfinska _ engelska
Dagvårdens samanvändningsområdefinska _ svenska _ engelska
förskoleundervisning
i Grankulla anordnas förskoleundervisningen i daghemmen .
förskoleundervisningen börjar i augusti och ansökningstiden är i januari .
Läs mer : förskoleundervisning
information om förskoleundervisningenfinska _ svenska _ engelska
grundläggande utbildning
i Grankulla finns både en finsk- och en svenskspråkig grundskola . anmälan till grundskolan ska ske i början av året .
om du har frågor om den grundläggande utbildningen kan du kontakta skolbyrån .
skolbyrån
Grankulla stadshus
Grankullavägen 10
02700 Grankulla
tfn ( 09 ) 50.561 ( växel )
grundläggande utbildning
grundläggande utbildning och gymnasiumfinska _ svenska _ engelska
internationella skolor i huvudstadsregionenfinska
linkkiExpatFinland.fi :
internationella skolor i huvudstadsregionenengelska
yrkesutbildning
de närmaste yrkesläroanstalterna finns i Esbo och Helsingfors .
Läs mer : yrkesutbildning
yrkesutbildningfinska _ engelska
Yrkesinriktad utbildningfinska
gymnasium
i Grankulla finns två gymnasier , ett finskspråkigt och ett svenskspråkigt .
i Esbo finns ett vuxengymnasium där vuxna kan avlägga gymnasiet och studentexamen .
Läs mer : gymnasium
grundläggande utbildning och gymnasiumfinska _ svenska _ engelska
linkkiEsbo stad :
Vuxengymnasietfinska
Högskoleutbildning
i anslutning till folkhögskolan Työväen Akatemia i Grankulla finns en enhet för Humanistiska Yrkeshögskolan , där du kan avlägga yrkeshögskoleexamen för kulturproducenter .
vid yrkeshögskolorna och universiteten i Esbo och Helsingfors kan du studera inom många områden .
mer information om högskolorna i Esbo och Helsingfors hittar du på städernas webbplatser .
Läs mer : Högskoleutbildning
linkkiHumanistiska yrkeshögskolan :
information om Humanistiska yrkeshögskolanfinska _ engelska
linkkiEsbo stad :
Högskolorfinska _ engelska
Högskolorfinska
andra studiemöjligheter
vid Grankulla medborgarinstitut kan du studera till exempel språk , handarbete och matlagning eller delta i ledd motion .
Medborgarinstitutetfinska _ svenska _ engelska
vid Grankulla konstskola kan barn och unga studera bildkonst och vid Grankulla musikinstitut kan barn och vuxna studera musik .
information om Konstskolanfinska _ svenska
information om Musikinstitutetfinska _ svenska
i Grankulla ligger Finska Bibelinstitutet .
vid institutet kan du avlägga enskilda kurser eller studera på någon av institutets studielinjer .
studierna på studielinjerna pågår i 1 @-@ 2 år .
vid bibelinstitutet finns även en studielinje som är särskilt avsedd för invandrare .
Kristliga folkhögskolanfinska _ engelska
folkhögskolan Työväen Akatemia tillhandahåller undervisning inom många akademiska discipliner samt träning för dem som vill läsa på universitet .
information om Työväen Akatemiafinska _ engelska
Läs mer : andra studiemöjligheter
dagvård
förskoleundervisning
grundläggande utbildning
yrkesutbildning
gymnasium
Högskoleutbildning
andra studiemöjligheter
dagvård
i Grankulla finns stadens egna daghem , privata daghem och privata familjedagvårdare .
dagvård fås på finska och på svenska .
i Grankulla finns också ett engelskspråkigt daghem .
Ansök om dagvårdsplats för ditt barn minst fyra månader innan barnet ska börja i dagvården .
om du ansöker om dagvårdplats för första gången ska du använda den elektroniska ansökan .
du kan också hämta ansökningsblanketten på daghemmet eller vid informationen i stadshuset .
lämna in ansökan till daghemmet eller stadshuset .
familjer som bor i Grankulla kan också söka dagvårdsplats till sitt barn i Esbo , Helsingfors eller Vanda .
du ska ändå lämna in din ansökan i Grankulla .
mer information finns på tjänsten HelsingforsRegionen.fi .
Läs mer : dagvård
dagvård och förskoleundervisningfinska _ svenska _ engelska
ansökan om dagvårdsplatsfinska _ svenska
Engelsk @-@ finskspråkigt daghemfinska _ engelska
Dagvårdens samanvändningsområdefinska _ svenska _ engelska
förskoleundervisning
i Grankulla anordnas förskoleundervisningen i daghemmen .
förskoleundervisningen börjar i augusti och ansökningstiden är i januari .
Läs mer : förskoleundervisning
information om förskoleundervisningenfinska _ svenska _ engelska
grundläggande utbildning
i Grankulla finns både en finsk- och en svenskspråkig grundskola . anmälan till grundskolan ska ske i början av året .
om du har frågor om den grundläggande utbildningen kan du kontakta skolbyrån .
skolbyrån
Grankulla stadshus
Grankullavägen 10
02700 Grankulla
tfn ( 09 ) 50.561 ( växel )
grundläggande utbildning
grundläggande utbildning och gymnasiumfinska _ svenska _ engelska
internationella skolor i huvudstadsregionenfinska
linkkiExpatFinland.fi :
internationella skolor i huvudstadsregionenengelska
yrkesutbildning
de närmaste yrkesläroanstalterna finns i Esbo och Helsingfors .
Läs mer : yrkesutbildning
yrkesutbildningfinska _ engelska
Yrkesinriktad utbildningfinska
gymnasium
i Grankulla finns två gymnasier , ett finskspråkigt och ett svenskspråkigt .
i Esbo finns ett vuxengymnasium där vuxna kan avlägga gymnasiet och studentexamen .
Läs mer : gymnasium
grundläggande utbildning och gymnasiumfinska _ svenska _ engelska
linkkiEsbo stad :
Vuxengymnasietfinska
Högskoleutbildning
i anslutning till folkhögskolan Työväen Akatemia i Grankulla finns en enhet för Humanistiska Yrkeshögskolan , där du kan avlägga yrkeshögskoleexamen för kulturproducenter .
vid yrkeshögskolorna och universiteten i Esbo och Helsingfors kan du studera inom många områden .
mer information om högskolorna i Esbo och Helsingfors hittar du på städernas webbplatser .
Läs mer : Högskoleutbildning
linkkiHumanistiska yrkeshögskolan :
information om Humanistiska yrkeshögskolanfinska _ engelska
linkkiEsbo stad :
Högskolorfinska _ engelska
Högskolorfinska
andra studiemöjligheter
vid Grankulla medborgarinstitut kan du studera till exempel språk , handarbete och matlagning eller delta i ledd motion .
Medborgarinstitutetfinska _ svenska _ engelska
vid Grankulla konstskola kan barn och unga studera bildkonst och vid Grankulla musikinstitut kan barn och vuxna studera musik .
information om Konstskolanfinska _ svenska
information om Musikinstitutetfinska _ svenska
i Grankulla ligger Finska Bibelinstitutet .
vid institutet kan du avlägga enskilda kurser eller studera på någon av institutets studielinjer .
studierna på studielinjerna pågår i 1 @-@ 2 år .
vid bibelinstitutet finns även en studielinje som är särskilt avsedd för invandrare .
Kristliga folkhögskolanfinska _ engelska
folkhögskolan Työväen Akatemia tillhandahåller undervisning inom många akademiska discipliner samt träning för dem som vill läsa på universitet .
information om Työväen Akatemiafinska _ engelska
Läs mer : andra studiemöjligheter
hyresbostad
Ägarbostad
Stöd- och serviceboende
avfallshantering i bostaden
hyresbostad
Hyresbostäderna är dyra i huvudstadsregionen .
stadens hyresbostäder är förmånligare än bostäder som hyrs ut av företag och privatpersoner .
privata hyresbostäder
du hittar bostäder som hyrs ut av företag och privatpersoner via bostadssidor på internet .
Sökning av hyresbostäderfinska
Sökning av hyresbostäderfinska _ engelska
stadens hyresbostäder
om du vill söka en av stadens hyresbostäder ska du fylla i en ansökningsblankett för hyresbostäder .
blanketten får du antingen vid informationen på Grankulla stadshus , på socialbyrån eller på Grankulla stads webbplats .
på stadens webbplats hittar du också anvisningar om hur du söker hyresbostad .
skicka din ansökan till adressen :
PB 52
02701 Grankulla
stadens hyresbostäderfinska _ svenska _ engelska
om du är studerande kan du få en hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS .
linkkiHOAS :
hyresbostäder för studerandefinska _ svenska _ engelska
Läs mer : hyresbostad
Ägarbostad
på internet finns många annonser om bostäder som är till salu .
bostäderna i Grankulla är tämligen dyra .
information om köp av bostad hittar du på InfoFinlands sida Ägarbostad .
om du blir bostadslös på grund av en kris eller en olycka , ska du kontakta socialbyrån .
om någon i din familj utövar våld mot dig eller hotar dig med våld , kan du kontakta ett skyddshem .
Steniusvägen 20
du kan ringa skyddshemmet dygnet runt , telefonnumret är 09.4777.180 .
du behöver inte uppge ditt namn när du ringer .
om du är ung och har problem hemma , kan du kontakta Finlands Röda Kors De ungas skyddshus .
det närmaste skyddshuset finns i Esbo .
de ungas skyddshus
tfn 09.819.55360
hjälp till offer för familjevåldfinska
linkkiFörbundet för mödra- och skyddshem :
information om skyddshem och mödrahemfinska
linkkiFinlands Röda Kors :
de ungas skyddshusfinska _ svenska _ engelska
Stöd- och serviceboende
personer som har svårt att klara av de dagliga sysslorna utan hjälp , till exempel äldre eller personer med funktionsnedsättning , kan få ta del av hemvårdens stödtjänster .
en person som inte kan bo på egen hand kan bo på en anstalt .
på Grankulla socialbyrå kan du fråga mer om hemvårdens stödtjänster och boende på anstalt .
Grankulla socialbyrå
Köpcentret Grani
Grankullavägen 7.02700 Grankulla
tfn 09.505.61
Läs mer : Stöd- och serviceboende
information om hemvårdens stödtjänsterfinska _ svenska
information om boende på anstaltfinska _ svenska
avfallshantering och återvinning
på InfoFinlands sida Avfallshantering och återvinning hittar du information om sopsortering .
linkkiHelsingforsregionens miljötjänster :
Sopsorteringsanvisningarfinska _ svenska _ engelska
Avfallsinsamlingsstationerfinska
hyresbostad
Ägarbostad
Stöd- och serviceboende
avfallshantering i bostaden
hyresbostad
Hyresbostäderna är dyra i huvudstadsregionen .
stadens hyresbostäder är förmånligare än bostäder som hyrs ut av företag och privatpersoner .
privata hyresbostäder
du hittar bostäder som hyrs ut av företag och privatpersoner via bostadssidor på internet .
Sökning av hyresbostäderfinska
Sökning av hyresbostäderfinska _ engelska
stadens hyresbostäder
om du vill söka en av stadens hyresbostäder ska du fylla i en ansökningsblankett för hyresbostäder .
blanketten får du antingen vid informationen på Grankulla stadshus , på socialbyrån eller på Grankulla stads webbplats .
på stadens webbplats hittar du också anvisningar om hur du söker hyresbostad .
skicka din ansökan till adressen :
PB 52
02701 Grankulla
stadens hyresbostäderfinska _ svenska _ engelska
om du är studerande kan du få en hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS .
linkkiHOAS :
hyresbostäder för studerandefinska _ svenska _ engelska
Läs mer : hyresbostad
Ägarbostad
på internet finns många annonser om bostäder som är till salu .
bostäderna i Grankulla är tämligen dyra .
information om köp av bostad hittar du på InfoFinlands sida Ägarbostad .
om du blir bostadslös på grund av en kris eller en olycka , ska du kontakta socialbyrån .
om någon i din familj utövar våld mot dig eller hotar dig med våld , kan du kontakta ett skyddshem .
Steniusvägen 20
du kan ringa skyddshemmet dygnet runt , telefonnumret är 09.4777.180 .
du behöver inte uppge ditt namn när du ringer .
om du är ung och har problem hemma , kan du kontakta Finlands Röda Kors De ungas skyddshus .
det närmaste skyddshuset finns i Esbo .
de ungas skyddshus
tfn 09.819.55360
hjälp till offer för familjevåldfinska
linkkiFörbundet för mödra- och skyddshem :
information om skyddshem och mödrahemfinska
linkkiFinlands Röda Kors :
de ungas skyddshusfinska _ svenska _ engelska
Stöd- och serviceboende
personer som har svårt att klara av de dagliga sysslorna utan hjälp , till exempel äldre eller personer med funktionsnedsättning , kan få ta del av hemvårdens stödtjänster .
en person som inte kan bo på egen hand kan bo på en anstalt .
på Grankulla socialbyrå kan du fråga mer om hemvårdens stödtjänster och boende på anstalt .
Grankulla socialbyrå
Köpcentret Grani
Grankullavägen 7.02700 Grankulla
tfn 09.505.61
Läs mer : Stöd- och serviceboende
information om hemvårdens stödtjänsterfinska _ svenska
information om boende på anstaltfinska _ svenska
avfallshantering och återvinning
på InfoFinlands sida Avfallshantering och återvinning hittar du information om sopsortering .
linkkiHelsingforsregionens miljötjänster :
Sopsorteringsanvisningarfinska _ svenska _ engelska
Avfallsinsamlingsstationerfinska
hyresbostad
Ägarbostad
Stöd- och serviceboende
avfallshantering i bostaden
hyresbostad
Hyresbostäderna är dyra i huvudstadsregionen .
stadens hyresbostäder är förmånligare än bostäder som hyrs ut av företag och privatpersoner .
privata hyresbostäder
du hittar bostäder som hyrs ut av företag och privatpersoner via bostadssidor på internet .
Sökning av hyresbostäderfinska
Sökning av hyresbostäderfinska _ engelska
stadens hyresbostäder
om du vill söka en av stadens hyresbostäder ska du fylla i en ansökningsblankett för hyresbostäder .
blanketten får du antingen vid informationen på Grankulla stadshus , på socialbyrån eller på Grankulla stads webbplats .
på stadens webbplats hittar du också anvisningar om hur du söker hyresbostad .
skicka din ansökan till adressen :
PB 52
02701 Grankulla
stadens hyresbostäderfinska _ svenska _ engelska
om du är studerande kan du få en hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS .
linkkiHOAS :
hyresbostäder för studerandefinska _ svenska _ engelska
Läs mer : hyresbostad
Ägarbostad
på internet finns många annonser om bostäder som är till salu .
bostäderna i Grankulla är tämligen dyra .
information om köp av bostad hittar du på InfoFinlands sida Ägarbostad .
om du blir bostadslös på grund av en kris eller en olycka , ska du kontakta socialbyrån .
om någon i din familj utövar våld mot dig eller hotar dig med våld , kan du kontakta ett skyddshem .
Steniusvägen 20
du kan ringa skyddshemmet dygnet runt , telefonnumret är 09.4777.180 .
du behöver inte uppge ditt namn när du ringer .
om du är ung och har problem hemma , kan du kontakta Finlands Röda Kors De ungas skyddshus .
det närmaste skyddshuset finns i Esbo .
de ungas skyddshus
tfn 09.819.55360
hjälp till offer för familjevåldfinska
linkkiFörbundet för mödra- och skyddshem :
information om skyddshem och mödrahemfinska
linkkiFinlands Röda Kors :
de ungas skyddshusfinska _ svenska _ engelska
Stöd- och serviceboende
personer som har svårt att klara av de dagliga sysslorna utan hjälp , till exempel äldre eller personer med funktionsnedsättning , kan få ta del av hemvårdens stödtjänster .
en person som inte kan bo på egen hand kan bo på en anstalt .
på Grankulla socialbyrå kan du fråga mer om hemvårdens stödtjänster och boende på anstalt .
Grankulla socialbyrå
Köpcentret Grani
Grankullavägen 7.02700 Grankulla
tfn 09.505.61
Läs mer : Stöd- och serviceboende
information om hemvårdens stödtjänsterfinska _ svenska
information om boende på anstaltfinska _ svenska
avfallshantering och återvinning
på InfoFinlands sida Avfallshantering och återvinning hittar du information om sopsortering .
linkkiHelsingforsregionens miljötjänster :
Sopsorteringsanvisningarfinska _ svenska _ engelska
Avfallsinsamlingsstationerfinska
språkkurser
med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors , Vanda , Esbo eller Grankulla .
i tjänsten finns också information om kurser i svenska .
kurser i finska och svenska språketfinska _ engelska _ ryska
i Grankulla ordnas kurser i finska och svenska av Grankulla medborgarinstitut .
du kan anmäla dig till medborgarinstitutets kurser per telefon eller via internet .
Medborgarinstitutetfinska _ svenska _ engelska
Läs mer : studier i finska och svenska
svenska språket i Finland .
diskutera på finska
information om bibliotekens språkkaféer och andra finska samtalsgrupper hittar du på InfoFinlands sidor Finska och svenska språket i Esbo och Finska och svenska språket i Helsingfors .
allmän språkexamen
du kan avlägga allmän språkexamen i finska eller svenska till exempel i Esbo och Helsingfors .
på Utbildningsstyrelsens webbplats finns en sökmotor med vilken du kan kontrollera var och när du kan avlägga examen .
Läs mer : Officiellt intyg på språkkunskaper .
linkkiUtbildningsstyrelsen :
allmänna språkexaminafinska _ svenska _ engelska
språkkurser
med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors , Vanda , Esbo eller Grankulla .
i tjänsten finns också information om kurser i svenska .
kurser i finska och svenska språketfinska _ engelska _ ryska
i Grankulla ordnas kurser i finska och svenska av Grankulla medborgarinstitut .
du kan anmäla dig till medborgarinstitutets kurser per telefon eller via internet .
Medborgarinstitutetfinska _ svenska _ engelska
Läs mer : studier i finska och svenska
svenska språket i Finland .
diskutera på finska
information om bibliotekens språkkaféer och andra finska samtalsgrupper hittar du på InfoFinlands sidor Finska och svenska språket i Esbo och Finska och svenska språket i Helsingfors .
allmän språkexamen
du kan avlägga allmän språkexamen i finska eller svenska till exempel i Esbo och Helsingfors .
på Utbildningsstyrelsens webbplats finns en sökmotor med vilken du kan kontrollera var och när du kan avlägga examen .
Läs mer : Officiellt intyg på språkkunskaper .
linkkiUtbildningsstyrelsen :
allmänna språkexaminafinska _ svenska _ engelska
språkkurser
med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors , Vanda , Esbo eller Grankulla .
i tjänsten finns också information om kurser i svenska .
kurser i finska och svenska språketfinska _ engelska _ ryska
i Grankulla ordnas kurser i finska och svenska av Grankulla medborgarinstitut .
du kan anmäla dig till medborgarinstitutets kurser per telefon eller via internet .
Medborgarinstitutetfinska _ svenska _ engelska
Läs mer : studier i finska och svenska
svenska språket i Finland .
diskutera på finska
information om bibliotekens språkkaféer och andra finska samtalsgrupper hittar du på InfoFinlands sidor Finska och svenska språket i Esbo och Finska och svenska språket i Helsingfors .
allmän språkexamen
du kan avlägga allmän språkexamen i finska eller svenska till exempel i Esbo och Helsingfors .
på Utbildningsstyrelsens webbplats finns en sökmotor med vilken du kan kontrollera var och när du kan avlägga examen .
Läs mer : Officiellt intyg på språkkunskaper .
linkkiUtbildningsstyrelsen :
allmänna språkexaminafinska _ svenska _ engelska
var hittar jag jobb ?
att grunda ett företag
beskattning
var hittar jag jobb ?
Nylands arbets- och näringsbyrå hjälper invånare i Grankulla att söka jobb .
den närmaste byrån finns i Esbo .
Nylands arbets- och näringsbyrå , Esbo
Läs mer : arbete och entreprenörskap i Esbo
information om arbets- och näringsbyråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös .
information om jobbsökning i Finland hittar du på InfoFinlands sida Var hittar jag jobb ?
Seure erbjuder kortvariga jobb vid Helsingfors , Vanda , Esbo och Grankulla städer .
Jobben finns till exempel på skolor , daghem och sjukhus .
arbetsplatser i kommunernafinska _ svenska
lediga jobbfinska _ svenska _ engelska
arbetslöshetsersättning
information om att ansöka om arbetslöshetsersättning hittar du på InfoFinlands sida Arbetslöshetsförsäkring .
att grunda ett företag
på InfoFinlands sida Att grunda ett företag hittar du information om hur man grundar ett företag i Finland .
Bekanta dig med de lokala tjänsterna på sidorna Arbete och entreprenörskap i Esbo och Arbete och entreprenörskap i Helsingfors .
om du är företagare kan du bli medlem i företagarnas intressebevakningsorganisation Grankulla företagare rf som erbjuder sina medlemmar utbildning , nätverk och rådgivning .
information för företagarefinska
beskattning
huvudstadsregionens skattebyrå ligger på Alexandersgatan 9 i Gloet i Helsingfors .
linkkiSkatteförvaltningen :
kontaktuppgifter till skattebyråerfinska _ svenska _ engelska
du kan även besöka servicestället In To Finland i Kampen i Helsingfors för att fråga om beskattningen .
servicestället betjänar invandrare som kommer till Finland för att arbeta i ärenden som berör beskattning och social trygghet .
Albertsgatan 25
lär mer Beskattning
var hittar jag jobb ?
att grunda ett företag
beskattning
var hittar jag jobb ?
Nylands arbets- och näringsbyrå hjälper invånare i Grankulla att söka jobb .
den närmaste byrån finns i Esbo .
Nylands arbets- och näringsbyrå , Esbo
Läs mer : arbete och entreprenörskap i Esbo
information om arbets- och näringsbyråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös .
information om jobbsökning i Finland hittar du på InfoFinlands sida Var hittar jag jobb ?
Seure erbjuder kortvariga jobb vid Helsingfors , Vanda , Esbo och Grankulla städer .
Jobben finns till exempel på skolor , daghem och sjukhus .
arbetsplatser i kommunernafinska _ svenska
lediga jobbfinska _ svenska _ engelska
arbetslöshetsersättning
information om att ansöka om arbetslöshetsersättning hittar du på InfoFinlands sida Arbetslöshetsförsäkring .
att grunda ett företag
på InfoFinlands sida Att grunda ett företag hittar du information om hur man grundar ett företag i Finland .
Bekanta dig med de lokala tjänsterna på sidorna Arbete och entreprenörskap i Esbo och Arbete och entreprenörskap i Helsingfors .
om du är företagare kan du bli medlem i företagarnas intressebevakningsorganisation Grankulla företagare rf som erbjuder sina medlemmar utbildning , nätverk och rådgivning .
information för företagarefinska
beskattning
huvudstadsregionens skattebyrå ligger på Alexandersgatan 9 i Gloet i Helsingfors .
linkkiSkatteförvaltningen :
kontaktuppgifter till skattebyråerfinska _ svenska _ engelska
invandrare kan även sköta ärenden vid servicestället International House Helsinki .
på servicestället hjälper FPA:s och Skatteförvaltningens experter invandrare som kommer till Finland för att arbeta i frågor som rör beskattning och social trygghet .
lär mer Beskattning
var hittar jag jobb ?
att grunda ett företag
beskattning
var hittar jag jobb ?
Nylands arbets- och näringsbyrå hjälper invånare i Grankulla att söka jobb .
den närmaste byrån finns i Esbo .
Nylands arbets- och näringsbyrå , Esbo
Läs mer : arbete och entreprenörskap i Esbo
information om arbets- och näringsbyråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös .
information om jobbsökning i Finland hittar du på InfoFinlands sida Var hittar jag jobb ?
Seure erbjuder kortvariga jobb vid Helsingfors , Vanda , Esbo och Grankulla städer .
Jobben finns till exempel på skolor , daghem och sjukhus .
arbetsplatser i kommunernafinska _ svenska _ engelska
lediga jobbfinska _ svenska _ engelska
arbetslöshetsersättning
information om att ansöka om arbetslöshetsersättning hittar du på InfoFinlands sida Arbetslöshetsförsäkring .
att grunda ett företag
på InfoFinlands sida Att grunda ett företag hittar du information om hur man grundar ett företag i Finland .
Bekanta dig med de lokala tjänsterna på sidorna Arbete och entreprenörskap i Esbo och Arbete och entreprenörskap i Helsingfors .
om du är företagare kan du bli medlem i företagarnas intressebevakningsorganisation Grankulla företagare rf som erbjuder sina medlemmar utbildning , nätverk och rådgivning .
information för företagarefinska
beskattning
huvudstadsregionens skattebyrå ligger på Alexandersgatan 9 i Gloet i Helsingfors .
linkkiSkatteförvaltningen :
kontaktuppgifter till skattebyråerfinska _ svenska _ engelska
invandrare kan även sköta ärenden vid servicestället International House Helsinki .
på servicestället hjälper FPA:s och Skatteförvaltningens experter invandrare som kommer till Finland för att arbeta i frågor som rör beskattning och social trygghet .
IHH - serviceställe för dig som flyttar till Finland engelska
lär mer Beskattning
rådgivning för och integration av invandrare
inledande kartläggning och integrationsplan
behöver du en tolk ?
rådgivning för och integration av invandrare
om du har frågor om tjänsterna vid Grankulla stad kan du kontakta stadens rådgivningstjänst via e @-@ post på adressen neuvontapalvelu ( at ) kauniainen.fi .
du kan skriva på finska , svenska eller engelska .
Helsingfors stads rådgivning för invandrare , Helsingfors @-@ info , betjänar alla invandrare i huvudstadsregionen .
Helsingfors @-@ infofinska _ svenska _ engelska
om du har flyttat till huvudstadsregionen nyligen , kan du vid International House Helsinki ( IHH ) få rådgivning och myndighetstjänster på ett och samma besök .
IHH - serviceställe för dig som flyttar till Finland engelska
inledande kartläggning och integrationsplan
tillsammans med en anställd vid arbets- och näringsbyrån ( TE @-@ byrån ) gör du en inledande kartläggning och en integrationsplan i samband med att du registrerar dig som arbetssökande .
linkkiArbets- och näringsministeriet :
arbets- och näringsbyråerna i Nylandfinska _ svenska
om du inte är kund hos arbets- och näringsbyrån görs den inledande kartläggningen och integrationsplanen på socialbyrån .
kontaktuppgifter till socialbyrån :
Köpcentret Grani
Grankullavägen 7
02700 Grankulla
tfn ( 09 ) 50.561
Socialbyrånfinska _ svenska
behöver du en tolk ?
om du inte kan finska eller svenska kan du anlita en tolk när du sköter ärenden med myndigheter .
du kan anlita en tolk när som helst om du bokar tolken och betalar kostnaderna själv .
i vissa fall får du en tolk via myndigheten .
då är tolkningen avgiftsfri för dig .
Läs mer : behöver du en tolk ?
linkkiFinlands översättar- och tolkförbund :
Sök tolk eller översättarefinska _ svenska _ engelska
rådgivning för och integration av invandrare
inledande kartläggning och integrationsplan
behöver du en tolk ?
rådgivning för och integration av invandrare
om du har frågor om tjänsterna vid Grankulla stad kan du kontakta stadens rådgivningstjänst via e @-@ post på adressen neuvontapalvelu ( at ) kauniainen.fi .
du kan skriva på finska , svenska eller engelska .
Helsingfors stads rådgivning för invandrare , Helsingfors @-@ info , betjänar alla invandrare i huvudstadsregionen .
Helsingfors @-@ infofinska _ svenska _ engelska
om du har flyttat till huvudstadsregionen nyligen , kan du vid International House Helsinki ( IHH ) få rådgivning och myndighetstjänster på ett och samma besök .
IHH - serviceställe för dig som flyttar till Finland engelska
inledande kartläggning och integrationsplan
tillsammans med en anställd vid arbets- och näringsbyrån ( TE @-@ byrån ) gör du en inledande kartläggning och en integrationsplan i samband med att du registrerar dig som arbetssökande .
linkkiArbets- och näringsministeriet :
arbets- och näringsbyråerna i Nylandfinska _ svenska
om du inte är kund hos arbets- och näringsbyrån görs den inledande kartläggningen och integrationsplanen på socialbyrån .
kontaktuppgifter till socialbyrån :
Köpcentret Grani
Grankullavägen 7
02700 Grankulla
tfn ( 09 ) 50.561
Socialbyrånfinska _ svenska
behöver du en tolk ?
om du inte kan finska eller svenska kan du anlita en tolk när du sköter ärenden med myndigheter .
du kan anlita en tolk när som helst om du bokar tolken och betalar kostnaderna själv .
i vissa fall får du en tolk via myndigheten .
då är tolkningen avgiftsfri för dig .
Läs mer : behöver du en tolk ?
linkkiFinlands översättar- och tolkförbund :
Sök tolk eller översättarefinska _ svenska _ engelska
rådgivning för och integration av invandrare
inledande kartläggning och integrationsplan
behöver du en tolk ?
rådgivning för och integration av invandrare
om du har frågor om tjänsterna vid Grankulla stad kan du kontakta stadens rådgivningstjänst via e @-@ post på adressen neuvontapalvelu ( at ) kauniainen.fi .
du kan skriva på finska , svenska eller engelska .
Helsingfors stads rådgivning för invandrare , Helsingfors @-@ info , betjänar alla invandrare i huvudstadsregionen .
Helsingfors @-@ infofinska _ svenska _ engelska
om du har flyttat till huvudstadsregionen nyligen , kan du vid International House Helsinki ( IHH ) få rådgivning och myndighetstjänster på ett och samma besök .
IHH - serviceställe för dig som flyttar till Finland engelska
inledande kartläggning och integrationsplan
tillsammans med en anställd vid arbets- och näringsbyrån ( TE @-@ byrån ) gör du en inledande kartläggning och en integrationsplan i samband med att du registrerar dig som arbetssökande .
linkkiArbets- och näringsministeriet :
arbets- och näringsbyråerna i Nylandfinska _ svenska
om du inte är kund hos arbets- och näringsbyrån görs den inledande kartläggningen och integrationsplanen på socialbyrån .
kontaktuppgifter till socialbyrån :
Köpcentret Grani
Grankullavägen 7
02700 Grankulla
tfn ( 09 ) 50.561
Socialbyrånfinska _ svenska
behöver du en tolk ?
om du inte kan finska eller svenska kan du anlita en tolk när du sköter ärenden med myndigheter .
du kan anlita en tolk när som helst om du bokar tolken och betalar kostnaderna själv .
i vissa fall får du en tolk via myndigheten .
då är tolkningen avgiftsfri för dig .
Läs mer : behöver du en tolk ?
linkkiFinlands översättar- och tolkförbund :
Sök tolk eller översättarefinska _ svenska _ engelska
tillståndsärenden
på Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU @-@ medborgarens uppehållsrätt .
boka en tid i förväg .
adress :
Göksgränd 3A
elektronisk tidsbokningfinska _ svenska _ engelska
du kan också ansöka om många slags uppehållstillstånd och EU @-@ registrering på internet i tjänsten Enter Finland .
linkkiEnterfinland.fi :
elektronisk ansökanfinska _ svenska _ engelska
Läs mer : flytta till Finland .
registrering som invånare
om du flyttar ditt stadigvarande boende till Grankulla , ska du registrera dig som invånare i kommunen .
du kan registrera dig vid Helsingfors enhet vid magistraten i Nyland .
Helsingfors enhet
Albertsgatan 25
tfn 029.55.39391
när du går till magistraten ska du ta med dig
legitimation ( till exempel pass )
uppehållstillstånd och uppehållskort ( om du behöver uppehållstillstånd i Finland )
registreringsintyget över uppehållsrätten ( om du är EU @-@ medborgare )
äktenskapsintyg
dina barns födelseattester .
Observera att utländska handlingar ska vara legaliserade samt översatta till finska eller svenska .
Läs mer : registrering som invånare
hemkommun i Finland
registrering av utlänningarfinska _ svenska _ engelska
IHH - serviceställe för dig som flyttar till Finland engelska
tillståndsärenden
på Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU @-@ medborgarens uppehållsrätt .
boka en tid i förväg .
adress :
Göksgränd 3A
elektronisk tidsbokningfinska _ svenska _ engelska
du kan också ansöka om många slags uppehållstillstånd och EU @-@ registrering på internet i tjänsten Enter Finland .
linkkiEnterfinland.fi :
elektronisk ansökanfinska _ svenska _ engelska
Läs mer : flytta till Finland .
registrering som invånare
om du flyttar ditt stadigvarande boende till Grankulla , ska du registrera dig som invånare i kommunen .
du kan registrera dig vid Helsingfors enhet vid magistraten i Nyland .
Helsingfors enhet
tfn 029.55.39391
när du går till magistraten ska du ta med dig
legitimation ( till exempel pass )
uppehållstillstånd och uppehållskort ( om du behöver uppehållstillstånd i Finland )
registreringsintyget över uppehållsrätten ( om du är EU @-@ medborgare )
äktenskapsintyg
dina barns födelseattester .
Observera att utländska handlingar ska vara legaliserade samt översatta till finska eller svenska .
Läs mer : registrering som invånare
hemkommun i Finland
registrering av utlänningarfinska _ svenska _ engelska
IHH - serviceställe för dig som flyttar till Finland engelska
tillståndsärenden
på Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU @-@ medborgarens uppehållsrätt .
boka en tid i förväg .
adress :
Göksgränd 3A
elektronisk tidsbokningfinska _ svenska _ engelska
du kan också ansöka om många slags uppehållstillstånd och EU @-@ registrering på internet i tjänsten Enter Finland .
linkkiEnterfinland.fi :
elektronisk ansökanfinska _ svenska _ engelska
Läs mer : flytta till Finland .
registrering som invånare
om du flyttar ditt stadigvarande boende till Grankulla , ska du registrera dig som invånare i kommunen .
du kan registrera dig vid Helsingfors enhet vid magistraten i Nyland .
Helsingfors enhet
tfn 029.55.39391
när du går till magistraten ska du ta med dig
legitimation ( till exempel pass )
uppehållstillstånd och uppehållskort ( om du behöver uppehållstillstånd i Finland )
registreringsintyget över uppehållsrätten ( om du är EU @-@ medborgare )
äktenskapsintyg
dina barns födelseattester .
Observera att utländska handlingar ska vara legaliserade samt översatta till finska eller svenska .
Läs mer : registrering som invånare
hemkommun i Finland
registrering av utlänningarfinska _ svenska _ engelska
IHH - serviceställe för dig som flyttar till Finland engelska
trafik
beslutsfattande och påverkan
religion
grundläggande information
historia
trafik
kollektivtrafiken
Vanda och hela huvudstadsregionen har goda kollektivtrafikförbindelser .
längs stambanan och Mårtensdals bana finns flera tågstationer .
i staden finns flera busslinjer .
Vanda tillhör samkommunen Helsingforsregionens trafik ( HRT ) ( Helsingin seudun liikenne -kuntayhtymä ( HSL ) ) , som ordnar kollektivtrafiken i huvudstadsregionen .
mer information hittar du på HRT:s webbplats .
du kan söka information om rutterna i Reseplaneraren ( Reittiopas ) .
tjänsten ger dig förslag på olika kollektivtrafikförbindelser från ett ställe till ett annat .
i kollektivtrafiken kan du betala med kontanter eller resekort .
i närtågen måste du köpa biljetten i förväg .
du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat .
Reseplanerarefinska _ svenska _ engelska _ ryska
resekort
med ett resekort ( matkakortti ) reser du förmånligare än med kontanter .
resekortet gäller i lokaltrafikens bussar , närtågen , metron , spårvagnarna och Sveaborgsfärjorna .
det finns två slags resekort .
det är det billigaste sättet att resa .
ett innehavarkort ( haltijakohtainen kortti ) kan användas av flera personer .
innan du skaffar dig ett personligt kort ska du registrera dig som invånare i någon av kommunerna inom HRT @-@ området .
du kan köpa resekort vid HRT:s försäljningsställen ( myyntipiste ) eller serviceställen ( palvelupiste ) .
de finns runtom i huvudstadsregionen .
personligt resekort kan du köpa vid serviceställena .
ta med dig identitetsbevis om du ska köpa personligt resekort .
om du har finska nätbankskoder kan du även köpa personligt resekort på HRT:s webbplats .
du kan resa med resekortet när du laddar kortet med period ( kausi ) eller värde ( arvo ) .
en period betyder tid : till exempel en månad .
värde betyder pengar .
om du använder kollektivtrafiken ofta tjänar du på att ladda kortet med period .
du kan ladda resekortet på vilket serviceställe för resekort ( matkakortin latauspiste ) som helst .
du hittar mer information på HRT:s webbplats .
ansökan om försäljningsplatserfinska _ svenska _ engelska
information och råd till resenärerfinska _ svenska _ engelska
Biljetter och priserfinska _ svenska _ engelska
att gå och cykla
om du vill gå eller cykla i Vanda kan du söka en lämplig rutt i reseplaneraren för cykling och gång .
en cykelkarta i pappersformat för Vanda kan du hämta i Vandainfo .
Cykelkartorna är kostnadsfria .
linkkiVanda stad :
Vandainfofinska _ svenska _ engelska
bil och flyg
Helsingfors @-@ Vanda internationella flygplats ligger i Vanda .
Flygplatsen har goda trafikförbindelser till exempel med bil , buss och tåg .
du kan parkera bilen på många järnvägsstationer och fortsätta färden med kollektivtrafiken .
Tidtabellerna för bussar och tåg hittar du enkelt i reseplaneraren .
Läs mer : trafik .
Flygplatsenfinska _ svenska _ engelska _ ryska _ kinesiska
beslutsfattande och påverkan
i Vanda beslutas ärenden av stadsfullmäktige ( kaupunginvaltuusto ) .
i stadsfullmäktige sitter 67 ledamöter som representerar olika politiska grupper .
Fullmäktige väljs var fjärde år genom kommunalval ( kunnallisvaalit ) .
invånarna i Vanda kan påverka beslutsfattandet och beredning av ärenden på många olika sätt .
på Vandakanalen kan du följa fullmäktiges sammanträden och få mer information om beslutsfattandet .
i Vanda finns en delegation för mångkulturella frågor ( monikulttuurisuusasiain neuvottelukunta ) som lägger fram propositioner i ärenden som rör invandrare .
Läs mer på Vanda stads webbplats .
i Vanda finns många politiska föreningar , invandrarföreningar och andra föreningar via vilka du också kan påverka beslutsfattandet .
mer information om föreningarna hittar du på sidan Vantaalla.info .
linkkiVanda stad :
beslutsfattandefinska _ svenska _ engelska
linkkiVanda stad :
delta och påverkafinska
Stadsfullmäktiges sammanträden på Internetfinska
linkkiVanda stad :
Delegationen för mångkulturella frågorfinska
religion
många religiösa samfund är verksamma i Vanda och Helsingfors .
via tjänsten Uskonnot Suomessa kan du söka information efter det religiösa samfundet och orten .
den evangelisk @-@ lutherska kyrkan har sex finskspråkiga församlingar och en svenskspråkig församling i Vanda .
Läs mer på Vanda kyrkliga samfällighets webbplats .
i Dickursby finns en ortodox kyrka .
mer information om verksamheten vid den ortodoxa kyrkan i Vanda hittar du på Helsingfors ortodoxa församlings webbplats .
Läs mer : kulturer och religioner i Finland .
linkkiVanda kyrkliga samfällighet :
evangelisk @-@ lutherska församlingarfinska
linkkiHelsingfors ortodoxa församling :
ortodoxa församlingenfinska _ ryska
religiösa samfundfinska _ engelska
grundläggande information
Vanda är en av de fyra kommunerna i huvudstadsregionen .
den ligger intill Esbo och Helsingfors .
Vanda centrum ligger i Dickursby .
Därtill finns det andra stora tätorter i Vanda , till exempel Korso , Björkby @-@ Havukoski , Myrbacka , Mårtensdal , Håkansböle , Västerkulla och Backas .
Vanda har drygt 205.000 invånare .
av dem är cirka 2,8 procent svenskspråkiga och 11 procent har något annat modersmål än finska eller svenska .
Arealen är cirka 240 km2 , varav cirka 2 km2 består av vatten .
linkkiVanda stad :
grundläggande informationfinska _ svenska _ engelska
historia
Vanda område har varit bebott länge .
man har hittat upp till 7.000 år gamla lämningar efter bosättning .
Nuvarande Vanda har uppstått på ett område som förr var Helsingfors socken .
Helsingfors sockens historia sträcker sig ända till 1300 @-@ talet .
Helsingfors socken blev först Helsingfors landskommun , sedan Vanda köping år 1972 och till slut Vanda stad år 1974 .
Läget som granne till huvudstaden Helsingfors har varit viktigt för Vanda .
viktiga vägar , såsom vägen från Åbo via Helsingfors till Viborg och senare järnvägen norrut från Helsingfors , har gått genom Vanda .
längs med vägarna och järnvägen har det utvecklats industrier och bostadsområden .
Vanda är än idag en viktig trafikknutpunkt .
till exempel ligger Helsingfors @-@ Vanda flygplats i Vanda .
linkkiVanda stad :
information om Vandafinska
linkkiVanda stad :
Stadsmuseetfinska _ svenska _ engelska
trafik
beslutsfattande och påverkan
religion
grundläggande information
historia
trafik
kollektivtrafiken
Vanda och hela huvudstadsregionen har goda kollektivtrafikförbindelser .
längs stambanan och Mårtensdals bana finns flera tågstationer .
i staden finns flera busslinjer .
Vanda tillhör samkommunen Helsingforsregionens trafik ( HRT ) ( Helsingin seudun liikenne -kuntayhtymä ( HSL ) ) , som ordnar kollektivtrafiken i huvudstadsregionen .
mer information hittar du på HRT:s webbplats .
du kan söka information om rutterna i Reseplaneraren ( Reittiopas ) .
tjänsten ger dig förslag på olika kollektivtrafikförbindelser från ett ställe till ett annat .
i kollektivtrafiken kan du betala med kontanter eller resekort .
i närtågen måste du köpa biljetten i förväg .
du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat .
Reseplanerarefinska _ svenska _ engelska _ ryska
resekort
med ett resekort ( matkakortti ) reser du förmånligare än med kontanter .
resekortet gäller i lokaltrafikens bussar , närtågen , metron , spårvagnarna och Sveaborgsfärjorna .
det finns två slags resekort .
det är det billigaste sättet att resa .
ett innehavarkort ( haltijakohtainen kortti ) kan användas av flera personer .
innan du skaffar dig ett personligt kort ska du registrera dig som invånare i någon av kommunerna inom HRT @-@ området .
du kan köpa resekort vid HRT:s försäljningsställen ( myyntipiste ) eller serviceställen ( palvelupiste ) .
de finns runtom i huvudstadsregionen .
personligt resekort kan du köpa vid serviceställena .
ta med dig identitetsbevis om du ska köpa personligt resekort .
om du har finska nätbankskoder kan du även köpa personligt resekort på HRT:s webbplats .
du kan resa med resekortet när du laddar kortet med period ( kausi ) eller värde ( arvo ) .
en period betyder tid : till exempel en månad .
värde betyder pengar .
om du använder kollektivtrafiken ofta tjänar du på att ladda kortet med period .
du kan ladda resekortet på vilket serviceställe för resekort ( matkakortin latauspiste ) som helst .
du hittar mer information på HRT:s webbplats .
ansökan om försäljningsplatserfinska _ svenska _ engelska
information och råd till resenärerfinska _ svenska _ engelska
Biljetter och priserfinska _ svenska _ engelska
att gå och cykla
om du vill gå eller cykla i Vanda kan du söka en lämplig rutt i reseplaneraren för cykling och gång .
en cykelkarta i pappersformat för Vanda kan du hämta i Vandainfo .
Cykelkartorna är kostnadsfria .
linkkiVanda stad :
Vandainfofinska _ svenska _ engelska
bil och flyg
Helsingfors @-@ Vanda internationella flygplats ligger i Vanda .
Flygplatsen har goda trafikförbindelser till exempel med bil , buss och tåg .
du kan parkera bilen på många järnvägsstationer och fortsätta färden med kollektivtrafiken .
Tidtabellerna för bussar och tåg hittar du enkelt i reseplaneraren .
Läs mer : trafik .
Flygplatsenfinska _ svenska _ engelska _ ryska _ kinesiska
beslutsfattande och påverkan
i Vanda beslutas ärenden av stadsfullmäktige ( kaupunginvaltuusto ) .
i stadsfullmäktige sitter 67 ledamöter som representerar olika politiska grupper .
Fullmäktige väljs var fjärde år genom kommunalval ( kunnallisvaalit ) .
invånarna i Vanda kan påverka beslutsfattandet och beredning av ärenden på många olika sätt .
på Vandakanalen kan du följa fullmäktiges sammanträden och få mer information om beslutsfattandet .
i Vanda finns en delegation för mångkulturella frågor ( monikulttuurisuusasiain neuvottelukunta ) som lägger fram propositioner i ärenden som rör invandrare .
Läs mer på Vanda stads webbplats .
i Vanda finns många politiska föreningar , invandrarföreningar och andra föreningar via vilka du också kan påverka beslutsfattandet .
mer information om föreningarna hittar du på sidan Vantaalla.info .
linkkiVanda stad :
beslutsfattandefinska _ svenska _ engelska
linkkiVanda stad :
delta och påverkafinska
Stadsfullmäktiges sammanträden på Internetfinska
linkkiVanda stad :
Delegationen för mångkulturella frågorfinska
religion
många religiösa samfund är verksamma i Vanda och Helsingfors .
via tjänsten Uskonnot Suomessa kan du söka information efter det religiösa samfundet och orten .
den evangelisk @-@ lutherska kyrkan har sex finskspråkiga församlingar och en svenskspråkig församling i Vanda .
Läs mer på Vanda kyrkliga samfällighets webbplats .
i Dickursby finns en ortodox kyrka .
mer information om verksamheten vid den ortodoxa kyrkan i Vanda hittar du på Helsingfors ortodoxa församlings webbplats .
Läs mer : kulturer och religioner i Finland .
linkkiVanda kyrkliga samfällighet :
evangelisk @-@ lutherska församlingarfinska
linkkiHelsingfors ortodoxa församling :
ortodoxa församlingenfinska _ ryska
religiösa samfundfinska _ engelska
grundläggande information
Vanda är en av de fyra kommunerna i huvudstadsregionen .
den ligger intill Esbo och Helsingfors .
Vanda centrum ligger i Dickursby .
Därtill finns det andra stora tätorter i Vanda , till exempel Korso , Björkby @-@ Havukoski , Myrbacka , Mårtensdal , Håkansböle , Västerkulla och Backas .
Vanda har drygt 205.000 invånare .
av dem är cirka 2,8 procent svenskspråkiga och 11 procent har något annat modersmål än finska eller svenska .
Arealen är cirka 240 km2 , varav cirka 2 km2 består av vatten .
linkkiVanda stad :
grundläggande informationfinska _ svenska _ engelska
historia
Vanda område har varit bebott länge .
man har hittat upp till 7.000 år gamla lämningar efter bosättning .
Nuvarande Vanda har uppstått på ett område som förr var Helsingfors socken .
Helsingfors sockens historia sträcker sig ända till 1300 @-@ talet .
Helsingfors socken blev först Helsingfors landskommun , sedan Vanda köping år 1972 och till slut Vanda stad år 1974 .
Läget som granne till huvudstaden Helsingfors har varit viktigt för Vanda .
viktiga vägar , såsom vägen från Åbo via Helsingfors till Viborg och senare järnvägen norrut från Helsingfors , har gått genom Vanda .
längs med vägarna och järnvägen har det utvecklats industrier och bostadsområden .
Vanda är än idag en viktig trafikknutpunkt .
till exempel ligger Helsingfors @-@ Vanda flygplats i Vanda .
linkkiVanda stad :
information om Vandafinska
linkkiVanda stad :
Stadsmuseetfinska _ svenska _ engelska
trafik
beslutsfattande och påverkan
religion
grundläggande information
historia
trafik
kollektivtrafiken
Vanda och hela huvudstadsregionen har goda kollektivtrafikförbindelser .
längs stambanan och Mårtensdals bana finns flera tågstationer .
i staden finns flera busslinjer .
Vanda tillhör samkommunen Helsingforsregionens trafik ( HRT ) ( Helsingin seudun liikenne -kuntayhtymä ( HSL ) ) , som ordnar kollektivtrafiken i huvudstadsregionen .
mer information hittar du på HRT:s webbplats .
du kan söka information om rutterna i Reseplaneraren ( Reittiopas ) .
tjänsten ger dig förslag på olika kollektivtrafikförbindelser från ett ställe till ett annat .
i kollektivtrafiken kan du betala med kontanter eller resekort .
i närtågen måste du köpa biljetten i förväg .
du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat .
Reseplanerarefinska _ svenska _ engelska
resekort
med ett resekort ( matkakortti ) reser du förmånligare än med kontanter .
resekortet gäller i lokaltrafikens bussar , närtågen , metron , spårvagnarna och Sveaborgsfärjorna .
det finns två slags resekort .
det är det billigaste sättet att resa .
ett innehavarkort ( haltijakohtainen kortti ) kan användas av flera personer .
innan du skaffar dig ett personligt kort ska du registrera dig som invånare i någon av kommunerna inom HRT @-@ området .
du kan köpa resekort vid HRT:s försäljningsställen ( myyntipiste ) eller serviceställen ( palvelupiste ) .
de finns runtom i huvudstadsregionen .
personligt resekort kan du köpa vid serviceställena .
ta med dig identitetsbevis om du ska köpa personligt resekort .
om du har finska nätbankskoder kan du även köpa personligt resekort på HRT:s webbplats .
du kan resa med resekortet när du laddar kortet med period ( kausi ) eller värde ( arvo ) .
en period betyder tid : till exempel en månad .
värde betyder pengar .
om du använder kollektivtrafiken ofta tjänar du på att ladda kortet med period .
du kan ladda resekortet på vilket serviceställe för resekort ( matkakortin latauspiste ) som helst .
du hittar mer information på HRT:s webbplats .
ansökan om försäljningsplatserfinska _ svenska _ engelska
information och råd till resenärerfinska _ svenska _ engelska
Biljetter och priserfinska _ svenska _ engelska
att gå och cykla
om du vill gå eller cykla i Vanda kan du söka en lämplig rutt i reseplaneraren för cykling och gång .
en cykelkarta i pappersformat för Vanda kan du hämta i Vandainfo .
Cykelkartorna är kostnadsfria .
linkkiVanda stad :
Vandainfofinska _ svenska _ engelska
bil och flyg
Helsingfors @-@ Vanda internationella flygplats ligger i Vanda .
Flygplatsen har goda trafikförbindelser till exempel med bil , buss och tåg .
du kan parkera bilen på många järnvägsstationer och fortsätta färden med kollektivtrafiken .
Tidtabellerna för bussar och tåg hittar du enkelt i reseplaneraren .
Läs mer : trafik .
Flygplatsenfinska _ svenska _ engelska _ ryska _ kinesiska
beslutsfattande och påverkan
i Vanda beslutas ärenden av stadsfullmäktige ( kaupunginvaltuusto ) .
i stadsfullmäktige sitter 67 ledamöter som representerar olika politiska grupper .
Fullmäktige väljs var fjärde år genom kommunalval ( kunnallisvaalit ) .
invånarna i Vanda kan påverka beslutsfattandet och beredning av ärenden på många olika sätt .
på Vandakanalen kan du följa fullmäktiges sammanträden och få mer information om beslutsfattandet .
i Vanda finns en delegation för mångkulturella frågor ( monikulttuurisuusasiain neuvottelukunta ) som lägger fram propositioner i ärenden som rör invandrare .
Läs mer på Vanda stads webbplats .
i Vanda finns många politiska föreningar , invandrarföreningar och andra föreningar via vilka du också kan påverka beslutsfattandet .
mer information om föreningarna hittar du på sidan Vantaalla.info .
linkkiVanda stad :
beslutsfattandefinska _ svenska _ engelska
linkkiVanda stad :
delta och påverkafinska
Stadsfullmäktiges sammanträden på Internetfinska
linkkiVanda stad :
Delegationen för mångkulturella frågorfinska
religion
många religiösa samfund är verksamma i Vanda och Helsingfors .
via tjänsten Uskonnot Suomessa kan du söka information efter det religiösa samfundet och orten .
den evangelisk @-@ lutherska kyrkan har sex finskspråkiga församlingar och en svenskspråkig församling i Vanda .
Läs mer på Vanda kyrkliga samfällighets webbplats .
i Dickursby finns en ortodox kyrka .
mer information om verksamheten vid den ortodoxa kyrkan i Vanda hittar du på Helsingfors ortodoxa församlings webbplats .
Läs mer : kulturer och religioner i Finland .
linkkiVanda kyrkliga samfällighet :
evangelisk @-@ lutherska församlingarfinska
linkkiHelsingfors ortodoxa församling :
ortodoxa församlingenfinska _ ryska
religiösa samfundfinska _ engelska
grundläggande information
Vanda är en av de fyra kommunerna i huvudstadsregionen .
den ligger intill Esbo och Helsingfors .
Vanda centrum ligger i Dickursby .
Därtill finns det andra stora tätorter i Vanda , till exempel Korso , Björkby @-@ Havukoski , Myrbacka , Mårtensdal , Håkansböle , Västerkulla och Backas .
Vanda har drygt 205.000 invånare .
av dem är cirka 2,8 procent svenskspråkiga och 11 procent har något annat modersmål än finska eller svenska .
Arealen är cirka 240 km2 , varav cirka 2 km2 består av vatten .
linkkiVanda stad :
grundläggande informationfinska _ svenska _ engelska
historia
Vanda område har varit bebott länge .
man har hittat upp till 7.000 år gamla lämningar efter bosättning .
Nuvarande Vanda har uppstått på ett område som förr var Helsingfors socken .
Helsingfors sockens historia sträcker sig ända till 1300 @-@ talet .
Helsingfors socken blev först Helsingfors landskommun , sedan Vanda köping år 1972 och till slut Vanda stad år 1974 .
Läget som granne till huvudstaden Helsingfors har varit viktigt för Vanda .
viktiga vägar , såsom vägen från Åbo via Helsingfors till Viborg och senare järnvägen norrut från Helsingfors , har gått genom Vanda .
längs med vägarna och järnvägen har det utvecklats industrier och bostadsområden .
Vanda är än idag en viktig trafikknutpunkt .
till exempel ligger Helsingfors @-@ Vanda flygplats i Vanda .
linkkiVanda stad :
information om Vandafinska
linkkiVanda stad :
Stadsmuseetfinska _ svenska _ engelska
bibliotek
motion
att röra sig i naturen
teater och film
museer
Fritidsverksamhet för barn och unga
Fritidsverksamhet för seniorer
föreningar
vid Vanda vuxenutbildningsinstitut ( Vantaan Aikuisopisto ) kan man till exempel skapa konst , handarbeten , laga mat eller dansa .
man kan även studera språk .
i Vanda finns två kulturhus : konserthuset Martinus och allaktivitetscentret Myrbackahuset .
dessutom ordnar allaktivitetscentret LUMO många evenemang .
Kulturhuset för barn och unga Fernissan , Konsthuset Pessi och Konsthuset Totem ordnar kulturevenemang för barn .
Läs mer : Fritid .
linkkiVanda vuxenutbildningsinstitut :
Studiehandbokfinska
linkkiVanda stad :
Kulturevenemangfinska _ svenska _ engelska
Konserterfinska _ svenska _ engelska
Evenemangfinska _ engelska
linkkiKulturhuset för barn och unga Fernissan :
kulturevenemang för barnfinska
kulturevenemang för barnfinska
kulturevenemang för barnfinska _ svenska
linkkiVanda stad :
evenemang och festivalerfinska _ engelska
bibliotek
i Vanda finns 10 bibliotek ( kirjasto ) och två bokbussar ( kirjastoauto ) .
på biblioteket kan du låna böcker , tidningar , musik , filmer , spel och mycket annat .
böcker och annat material finns på flera olika språk .
på biblioteket kan du också använda dator .
på vissa bibliotek ordnas även språkcaféer i det finska språket för invandrare .
biblioteken i Vanda är med i huvudstadsregionens bibliotekstjänst HelMet .
du kan alltså använda samma bibliotekskort på stadsbiblioteken i Vanda , Esbo , Grankulla och Helsingfors .
i Helsingfors huvudbibliotek i Böle finns Flerspråkigt bibliotek .
där hittar man böcker på över 60 olika språk .
om du har ett Helmet @-@ lånekort , kan du också låna böcker i Flerspråkiga biblioteket .
Läs mer : bibliotek
linkkiVanda stad :
information om bibliotekenfinska _ svenska _ engelska
linkkiHelsingfors stadsbibliotek :
Flerspråkiga biblioteketfinska _ svenska _ engelska
motion
i Vanda finns fem kommunala simhallar .
Simhallen i Korso har ett eget simpass för invandrarkvinnor och -flickor .
i Vanda finns flera idrottshallar , idrottsplaner och andra idrottsplatser för olika idrottsgrenar .
på motionsslingorna kan man springa på somrarna och åka skidor på vintrarna .
Läs mer : motion .
linkkiVanda stad :
Simhallarnas kontaktuppgifterfinska _ svenska _ engelska
linkkiVanda stad :
simpass för invandrarkvinnorfinska _ engelska
linkkiVanda stad :
Idrottsklubbarfinska
att röra sig i naturen
i Vanda finns många motionsslingor och naturstigar .
du kan även röra dig i naturen i Petikkos rekreationsområde .
du kan fiska på Vanda stads fiskeområden i Vanda å , Kervo å och på Finska viken .
Läs mer : att röra sig i naturen .
linkkiVanda stad :
Rekreations- och campingområdenfinska _ svenska
linkkiVanda stad :
idrottsplatser och friluftsområdenfinska _ svenska
friluftsområdenfinska
linkkiVanda stad :
fiske och båtlivfinska
teater och film
i Vanda finns flera yrkes- och amatörteatrar .
i Vanda finns fyra biografer .
mer information om filmerna hittar du på biografernas webbplatser .
Därtill ordnar Vanda stad filmvisningar .
Läs mer : teater och film .
linkkiVanda stad :
film , dans och teaterfinska _ engelska
museer
i Vanda finns flera museer .
på Vanda konstmuseum ordnas växlande utställningar med inhemsk och utländsk modern konst .
om de övriga museerna hittar du information på Vanda stads webbplats .
Läs mer : museer .
linkkiVanda stad :
Museerfinska _ engelska
linkkiVanda stad :
Stadsmuseetfinska _ svenska _ engelska
linkkiVanda stad :
Konstmuseetfinska _ svenska _ engelska
Fritidsverksamhet för barn och unga
i Vanda finns flera läroanstalter som ger grundundervisning i konst speciellt för barn och unga .
olika konstarter är musik , bildkonst , dans , teater , cirkuskonst , ordkonst , handarbete och arkitektur .
stadens ungdomsgårdar är öppna för alla ungdomar i åldrarna 10 @-@ 17 år .
Projektet Sport för alla ( Sporttia kaikille @-@ hanke ) ordnar idrottsklubbar , turneringar och läger för barn och ungdomar med invandrarbakgrund .
också föreningar och idrottsklubbar ordnar mycket verksamhet för ungdomar .
mer information hittar du på Vanda stads webbplats .
Läs mer : Fritidsverksamhet för barn och unga .
linkkiVanda stad :
information om hobbymöjligheter för ungdomarfinska
linkkiVanda stad :
kultur för barn och ungafinska _ svenska _ engelska
linkkiVanda stad :
information om konstundervisningfinska _ engelska
Ungdomsgårdarfinska
Motionsmöjligheterfinska
Hobbysökningfinska
linkkiVanda stad :
delta och påverkafinska _ svenska
Fritidsverksamhet för seniorer
om du har fyllt 70 år och Vanda är din hemkommun kan du kostnadsfritt använda Vanda stads simhallar och gym . du kommer gratis in till idrottsanläggningarna om du har ett Sportkort ( Sporttikortti ) .
du kan avhämta Sportkortet kostnadsfritt vid Vanda @-@ informationspunkterna .
ta med dig identitetsbevis och ett foto när du ansöker om kortet .
på Seniorrådgivningen ( seniorineuvonta ) får du information om hobbyer och tjänster för seniorer som olika organisationer , företag och staden erbjuder .
seniorrådgivningen
tfn : ( 09 ) 8392.4202
Motionsmöjligheterfinska _ svenska
föreningar
i Vanda finns många olika föreningar , till exempel kulturföreningar och idrottsklubbar .
mer information hittar du på Vanda stads webbplats .
Läs mer : föreningar .
linkkiVanda stad :
Kulturföreningarfinska
linkkiVanda stad :
Idrottsklubbarfinska
bibliotek
motion
att röra sig i naturen
teater och film
museer
Fritidsverksamhet för barn och unga
Fritidsverksamhet för seniorer
föreningar
vid Vanda vuxenutbildningsinstitut ( Vantaan Aikuisopisto ) kan man till exempel skapa konst , handarbeten , laga mat eller dansa .
man kan även studera språk .
i Vanda finns två kulturhus : konserthuset Martinus och allaktivitetscentret Myrbackahuset .
dessutom ordnar allaktivitetscentret LUMO många evenemang .
Kulturhuset för barn och unga Fernissan , Konsthuset Pessi och Konsthuset Totem ordnar kulturevenemang för barn .
Läs mer : Fritid .
linkkiVanda vuxenutbildningsinstitut :
Studiehandbokfinska
linkkiVanda stad :
Kulturevenemangfinska _ svenska _ engelska
Konserterfinska _ svenska _ engelska
Evenemangfinska _ engelska
linkkiKulturhuset för barn och unga Fernissan :
kulturevenemang för barnfinska
kulturevenemang för barnfinska
kulturevenemang för barnfinska _ svenska
linkkiVanda stad :
evenemang och festivalerfinska _ engelska
bibliotek
i Vanda finns 10 bibliotek ( kirjasto ) och två bokbussar ( kirjastoauto ) .
på biblioteket kan du låna böcker , tidningar , musik , filmer , spel och mycket annat .
böcker och annat material finns på flera olika språk .
på biblioteket kan du också använda dator .
på vissa bibliotek ordnas även språkcaféer i det finska språket för invandrare .
biblioteken i Vanda är med i huvudstadsregionens bibliotekstjänst HelMet .
du kan alltså använda samma bibliotekskort på stadsbiblioteken i Vanda , Esbo , Grankulla och Helsingfors .
i Helsingfors huvudbibliotek i Böle finns Flerspråkigt bibliotek .
där hittar man böcker på över 60 olika språk .
om du har ett Helmet @-@ lånekort , kan du också låna böcker i Flerspråkiga biblioteket .
Läs mer : bibliotek
linkkiVanda stad :
information om bibliotekenfinska _ svenska _ engelska
linkkiHelsingfors stadsbibliotek :
Flerspråkiga biblioteketfinska _ svenska _ engelska
motion
i Vanda finns fem kommunala simhallar .
Simhallen i Korso har ett eget simpass för invandrarkvinnor och -flickor .
i Vanda finns flera idrottshallar , idrottsplaner och andra idrottsplatser för olika idrottsgrenar .
på motionsslingorna kan man springa på somrarna och åka skidor på vintrarna .
Läs mer : motion .
linkkiVanda stad :
Simhallarnas kontaktuppgifterfinska _ svenska _ engelska
linkkiVanda stad :
simpass för invandrarkvinnorfinska _ engelska
linkkiVanda stad :
Idrottsklubbarfinska
att röra sig i naturen
i Vanda finns många motionsslingor och naturstigar .
du kan även röra dig i naturen i Petikkos rekreationsområde .
du kan fiska på Vanda stads fiskeområden i Vanda å , Kervo å och på Finska viken .
Läs mer : att röra sig i naturen .
linkkiVanda stad :
Rekreations- och campingområdenfinska _ svenska
linkkiVanda stad :
idrottsplatser och friluftsområdenfinska _ svenska
friluftsområdenfinska
linkkiVanda stad :
fiske och båtlivfinska
teater och film
i Vanda finns flera yrkes- och amatörteatrar .
i Vanda finns fyra biografer .
mer information om filmerna hittar du på biografernas webbplatser .
Därtill ordnar Vanda stad filmvisningar .
Läs mer : teater och film .
linkkiVanda stad :
film , dans och teaterfinska _ engelska
museer
i Vanda finns flera museer .
på Vanda konstmuseum ordnas växlande utställningar med inhemsk och utländsk modern konst .
om de övriga museerna hittar du information på Vanda stads webbplats .
Läs mer : museer .
linkkiVanda stad :
Museerfinska _ engelska
linkkiVanda stad :
Stadsmuseetfinska _ svenska _ engelska
linkkiVanda stad :
Konstmuseetfinska _ svenska _ engelska
Fritidsverksamhet för barn och unga
i Vanda finns flera läroanstalter som ger grundundervisning i konst speciellt för barn och unga .
olika konstarter är musik , bildkonst , dans , teater , cirkuskonst , ordkonst , handarbete och arkitektur .
stadens ungdomsgårdar är öppna för alla ungdomar i åldrarna 10 @-@ 17 år .
Projektet Sport för alla ( Sporttia kaikille @-@ hanke ) ordnar idrottsklubbar , turneringar och läger för barn och ungdomar med invandrarbakgrund .
också föreningar och idrottsklubbar ordnar mycket verksamhet för ungdomar .
mer information hittar du på Vanda stads webbplats .
Läs mer : Fritidsverksamhet för barn och unga .
linkkiVanda stad :
information om hobbymöjligheter för ungdomarfinska
linkkiVanda stad :
kultur för barn och ungafinska _ svenska _ engelska
linkkiVanda stad :
information om konstundervisningfinska _ engelska
Ungdomsgårdarfinska
Motionsmöjligheterfinska
Hobbysökningfinska
linkkiVanda stad :
delta och påverkafinska _ svenska
Fritidsverksamhet för seniorer
om du har fyllt 70 år och Vanda är din hemkommun kan du kostnadsfritt använda Vanda stads simhallar och gym . du kommer gratis in till idrottsanläggningarna om du har ett Sportkort ( Sporttikortti ) .
du kan avhämta Sportkortet kostnadsfritt vid Vanda @-@ informationspunkterna .
ta med dig identitetsbevis och ett foto när du ansöker om kortet .
på Seniorrådgivningen ( seniorineuvonta ) får du information om hobbyer och tjänster för seniorer som olika organisationer , företag och staden erbjuder .
seniorrådgivningen
tfn : ( 09 ) 8392.4202
Motionsmöjligheterfinska _ svenska
föreningar
i Vanda finns många olika föreningar , till exempel kulturföreningar och idrottsklubbar .
mer information hittar du på Vanda stads webbplats .
Läs mer : föreningar .
linkkiVanda stad :
Kulturföreningarfinska
linkkiVanda stad :
Idrottsklubbarfinska
bibliotek
motion
att röra sig i naturen
teater och film
museer
Fritidsverksamhet för barn och unga
Fritidsverksamhet för seniorer
föreningar
vid Vanda vuxenutbildningsinstitut ( Vantaan Aikuisopisto ) kan man till exempel skapa konst , handarbeten , laga mat eller dansa .
man kan även studera språk .
i Vanda finns två kulturhus : konserthuset Martinus och allaktivitetscentret Myrbackahuset .
dessutom ordnar allaktivitetscentret LUMO många evenemang .
Kulturhuset för barn och unga Fernissan , Konsthuset Pessi och Konsthuset Totem ordnar kulturevenemang för barn .
Läs mer : Fritid .
linkkiVanda vuxenutbildningsinstitut :
Studiehandbokfinska
linkkiVanda stad :
Kulturevenemangfinska _ svenska _ engelska
Konserterfinska _ svenska _ engelska
Evenemangfinska _ engelska
linkkiKulturhuset för barn och unga Fernissan :
kulturevenemang för barnfinska
kulturevenemang för barnfinska
kulturevenemang för barnfinska _ svenska
linkkiVanda stad :
evenemang och festivalerfinska _ engelska
bibliotek
i Vanda finns 10 bibliotek ( kirjasto ) och två bokbussar ( kirjastoauto ) .
på biblioteket kan du låna böcker , tidningar , musik , filmer , spel och mycket annat .
böcker och annat material finns på flera olika språk .
på biblioteket kan du också använda dator .
på vissa bibliotek ordnas även språkcaféer i det finska språket för invandrare .
biblioteken i Vanda är med i huvudstadsregionens bibliotekstjänst HelMet .
du kan alltså använda samma bibliotekskort på stadsbiblioteken i Vanda , Esbo , Grankulla och Helsingfors .
i Helsingfors huvudbibliotek i Böle finns Flerspråkigt bibliotek .
där hittar man böcker på över 60 olika språk .
om du har ett Helmet @-@ lånekort , kan du också låna böcker i Flerspråkiga biblioteket .
Läs mer : bibliotek
linkkiVanda stad :
information om bibliotekenfinska _ svenska _ engelska
linkkiHelsingfors stadsbibliotek :
Flerspråkiga biblioteketfinska _ svenska _ engelska
motion
i Vanda finns fem kommunala simhallar .
Simhallen i Korso har ett eget simpass för invandrarkvinnor och -flickor .
i Vanda finns flera idrottshallar , idrottsplaner och andra idrottsplatser för olika idrottsgrenar .
på motionsslingorna kan man springa på somrarna och åka skidor på vintrarna .
Läs mer : motion .
linkkiVanda stad :
Simhallarnas kontaktuppgifterfinska _ svenska _ engelska
linkkiVanda stad :
simpass för invandrarkvinnorfinska _ engelska
linkkiVanda stad :
Idrottsklubbarfinska
att röra sig i naturen
i Vanda finns många motionsslingor och naturstigar .
du kan även röra dig i naturen i Petikkos rekreationsområde .
du kan fiska på Vanda stads fiskeområden i Vanda å , Kervo å och på Finska viken .
Läs mer : att röra sig i naturen .
linkkiVanda stad :
Rekreations- och campingområdenfinska _ svenska
linkkiVanda stad :
idrottsplatser och friluftsområdenfinska _ svenska
friluftsområdenfinska
linkkiVanda stad :
fiske och båtlivfinska
teater och film
i Vanda finns flera yrkes- och amatörteatrar .
i Vanda finns fyra biografer .
mer information om filmerna hittar du på biografernas webbplatser .
Därtill ordnar Vanda stad filmvisningar .
Läs mer : teater och film .
linkkiVanda stad :
film , dans och teaterfinska _ engelska
museer
i Vanda finns flera museer .
på Vanda konstmuseum ordnas växlande utställningar med inhemsk och utländsk modern konst .
om de övriga museerna hittar du information på Vanda stads webbplats .
Läs mer : museer .
linkkiVanda stad :
Museerfinska _ engelska
linkkiVanda stad :
Stadsmuseetfinska _ svenska _ engelska
linkkiVanda stad :
Konstmuseetfinska _ svenska _ engelska
Fritidsverksamhet för barn och unga
i Vanda finns flera läroanstalter som ger grundundervisning i konst speciellt för barn och unga .
olika konstarter är musik , bildkonst , dans , teater , cirkuskonst , ordkonst , handarbete och arkitektur .
stadens ungdomsgårdar är öppna för alla ungdomar i åldrarna 10 @-@ 17 år .
Projektet Sport för alla ( Sporttia kaikille @-@ hanke ) ordnar idrottsklubbar , turneringar och läger för barn och ungdomar med invandrarbakgrund .
också föreningar och idrottsklubbar ordnar mycket verksamhet för ungdomar .
mer information hittar du på Vanda stads webbplats .
Läs mer : Fritidsverksamhet för barn och unga .
linkkiVanda stad :
information om hobbymöjligheter för ungdomarfinska
linkkiVanda stad :
kultur för barn och ungafinska _ svenska _ engelska
linkkiVanda stad :
information om konstundervisningfinska _ engelska
Ungdomsgårdarfinska
Motionsmöjligheterfinska
Hobbysökningfinska
linkkiVanda stad :
delta och påverkafinska _ svenska
Fritidsverksamhet för seniorer
om du har fyllt 70 år och Vanda är din hemkommun kan du kostnadsfritt använda Vanda stads simhallar och gym . du kommer gratis in till idrottsanläggningarna om du har ett Sportkort ( Sporttikortti ) .
du kan avhämta Sportkortet kostnadsfritt vid Vanda @-@ informationspunkterna .
ta med dig identitetsbevis och ett foto när du ansöker om kortet .
på Seniorrådgivningen ( seniorineuvonta ) får du information om hobbyer och tjänster för seniorer som olika organisationer , företag och staden erbjuder .
seniorrådgivningen
tfn : ( 09 ) 8392.4202
Motionsmöjligheterfinska _ svenska
föreningar
i Vanda finns många olika föreningar , till exempel kulturföreningar och idrottsklubbar .
mer information hittar du på Vanda stads webbplats .
Läs mer : föreningar .
linkkiVanda stad :
Kulturföreningarfinska
linkkiVanda stad :
Idrottsklubbarfinska
problem med uppehållstillståndet
brott
behöver du en jurist ?
våld
missbruksproblem och spelberoende
Dödsfall
om du behöver brådskande hjälp av polisen , brandkåren eller ambulansen , ring nödnumret 112 .
du får ringa nödnumret endast i brådskande nödfall där liv , hälsa , egendom eller miljö är i fara .
om du drabbas av en akut krissituation , såsom att en närstående avlider eller på grund av familjevåld , kan du kontakta social- och krisjouren ( sosiaali- ja kriisipäivystys ) .
du kan också söka hjälp för en familjemedlem eller en vän .
social- och krisjouren har öppet dygnet runt varje dag .
social- och krisjouren
tfn ( 09 ) 8392.4005
linkkiNödcentralsverket :
hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
linkkiVanda stad :
social- och krisjourenfinska _ svenska _ engelska
problem med uppehållstillståndet
om du har problem eller oklarheter med uppehållstillståndet , kontakta Migrationsverket .
du kan även fråga om råd på rådgivningstjänsterna för invandrare .
information om tjänsterna finns på sidan Som invandrare i Vanda .
Migrationsverkets närmaste tjänsteställe finns i Helsingfors :
Göksgränd 3A
Läs mer : problem med uppehållstillståndet
olika tillståndfinska _ svenska _ engelska
hälsovård för papperslösa
i Helsingfors finns Global Clinic , där personer som vistas i Finland utan tillstånd kan få primärhälsovård .
tjänsterna vid Global Clinic är avgiftsfria för kunderna .
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter .
för att skydda kunderna uppges inte klinikens adress eller öppettider offentligt .
telefonnumret till Global Clinic i Helsingfors är 044.977.4547 .
Samtalet besvaras av en sjukskötare eller en läkare .
e @-@ postadressen är globalclinic.finland ( at ) gmail.com .
Läs mer : problem med uppehållstillstånd
hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
brott
brottsanmälan ( rikosilmoitus ) kan göras per telefon eller personligen på polisstationen .
du kan också göra brottsanmälan på internet om brottet i fråga är ringa och du inte behöver omedelbar hjälp av polisen .
Konvaljvägen 21
tfn 0295.430291
Läs mer : brott .
kontaktuppgifterfinska _ svenska
elektronisk polisanmälanfinska _ svenska _ engelska
behöver du en jurist ?
östra Nylands rättshjälpsbyrå ( Itä @-@ Uudenmaan oikeusaputoimisto ) betjänar invånarna i Vanda .
Pyrolavägen 37
tfn 029.5660.160
du kan också söka information om privata jurister på till exempel Finlands Juristförbunds ( Suomen Asianajajaliitto ) webbplats .
Läs mer : behöver du en jurist ?
linkkiÖstra Nylands rättshjälpsbyrå :
information om rättshjälpfinska _ svenska _ engelska
linkkiFinlands Advokatförbund :
Advokaterfinska _ svenska _ engelska
våld
i nödsituationer ringer du nödnumret 112 .
i krissituationer får man även hjälp vid Vanda stads social- och krisjour ( sosiaali- ja kriisipäivystys ) , som har öppet dygnet runt .
social- och krisjouren
tfn ( 09 ) 8392.4005
linkkiNödcentralsverket :
hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
skyddshem
om någon i din familj utövar våld mot dig eller hotar dig med våld , kan du kontakta ett skyddshem ( turvakoti ) .
Skyddshemmen har jourmottagning dygnet runt .
skyddshemmet Mona ( turvakoti Mona ) är ett skyddshem avsett för invandrarkvinnor och deras barn .
tfn 045.639.6274
linkkiTurvakoti Mona :
skyddshemfinska
du kan även gå till Vanda skyddshem ( Vantaan turvakoti ) eller huvudstadsregionens skyddshem ( pääkaupunkiseudun turvakoti ) .
Puh . ( 09 ) 8392.0071
skyddshemfinska _ engelska
Steniusvägen 20
tfn ( 09 ) 4777.180
hjälp till offer för familjevåldfinska
hjälp för invandrarkvinnor
föreningen Monika @-@ Naiset liitto ( Monika @-@ Naiset Liitto ) ger råd och stöd till invandrarkvinnor .
föreningen har ett resurscenter ( voimavarakeskus ) i Vanda där man får stöd och råd .
tfn ( 09 ) 839.35013
hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
hjälp för män
män som har utövat våld mot sina familjemedlemmar eller har själva blivit offer för våld i hemmet , kan få hjälp från Jussi @-@ arbetet i Vanda ( Vantaan Jussi @-@ työ ) .
hjälp för män att sluta med våldsamt beteendefinska
Miehen linja ( Miehen linja ) hjälper invandrarmän som har problem med våld .
tfn ( 09 ) 276.62899
hjälp för män för att sluta med våldsamt beteendefinska _ engelska
hjälp för unga
Finlands Röda Kors De ungas skyddshus ( Suomen Punaisen Ristin Nuorten turvatalo ) ger stöd och hjälp i krissituationer för 12 @-@ 19 @-@ åringar .
skyddshuset har öppet kl . 17 @-@ 10 , telefonjouren betjänar dygnet runt .
Sjukhusgatan 3 ( Räckhals gård )
tfn ( 09 ) 871.4043
linkkiFinlands Röda Kors :
de ungas skyddshusfinska _ svenska _ engelska
Läs mer : våld
problem i äktenskap eller parförhållande
par med barn under 13 år kan vid problem i äktenskap och parförhållande få hjälp vid familjerådgivningen ( perheneuvola ) .
kontaktuppgifterna hittar du på Vanda stads webbplats .
Familjerådgivningens tjänster är konfidentiella och avgiftsfria .
vid akuta krissituationer inom familjen kan du kontakta social- och krisjouren ( sosiaali- ja kriisipäivystys ) , som har öppet dygnet runt varje dag .
social- och krisjouren
tfn ( 09 ) 8392.4005
vid problem i parförhållandet och familjen får man även hjälp av familjerådgivningen vid Vanda församlingar ( Vantaan seurakunnan perheneuvonta ) .
Läs mer : problem i äktenskap och parförhållande
linkkiVanda stad :
Familjerådgivningarfinska _ svenska
linkkiVanda kyrkliga samfällighet :
familjerådgivningfinska _ engelska
Barnrådgivningsbyråerna ( lastenneuvola ) och familjerådgivningsbyråerna ( perheneuvola ) ger råd i frågor som rör barns hälsa , uppväxt och utveckling .
vid problem hos barn i skolåldern får man hjälp hos skolhälsovårdarna ( kouluterveydenhoitaja ) , skolkuratorerna ( koulukuraattori ) och socialhandledarna ( sosiaaliohjaaja ) .
mer information hittar du på Vanda stads webbplats .
Läs mer : barns och ungas problem
linkkiVanda stad :
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad :
Familjerådgivningarfinska _ svenska
linkkiVanda stad :
information om tjänster för barn , ungdomar och familjerfinska _ svenska _ engelska
i skolan får de unga hjälp av skol- och studenthälsovårdarna ( koulu- ja opiskeluterveydenhoitajat ) , skolkuratorerna ( koulukuraattorit ) och skolpsykologerna ( koulupsykologit ) .
linkkiVanda stad :
information om skolhälsovårdenfinska _ svenska _ engelska
linkkiVanda stad :
Skolkuratorerfinska _ svenska
linkkiVanda stad :
Skolpsykologerfinska _ svenska
Nuppi
13 @-@ 21 @-@ åriga barn och ungdomar samt deras familjer kan få hjälp hos ungdomscentralen ( nuortenkeskus ) .
på Nuppi kan du till exempel få hjälp med mentala problem och missbruksproblem .
hjälp för ungafinska _ svenska _ engelska
om du är under 30 år , kan du få råd och handledning via tjänsten Navigatorn .
Personalen vid Navigatorn hjälper dig om du inte har något arbete eller en studieplats .
du kan även be om råd gällande andra saker , till exempel boende och ekonomi .
de ungas skyddshus
Finlands Röda Kors De ungas skyddshus ( Suomen Punaisen Ristin Nuorten turvatalo ) ger stöd och hjälp i krissituationer för 12 @-@ 19 @-@ åringar .
skyddshuset har öppet kl . 17 @-@ 10 , telefonjouren betjänar dygnet runt .
Sjukhusgatan 3
tfn ( 09 ) 871.4043
Läs mer : barns och ungas problem
linkkiFinlands Röda Kors :
de ungas skyddshusfinska _ svenska _ engelska
vägledning och stöd för ungafinska _ svenska
Socialrådgivningen ( sosiaalineuvonta ) ger information om utkomststöd ( toimeentulotuki ) och andra bidrag om du har ekonomiska problem .
tfn ( 09 ) 83.911 .
linkkiVanda stad :
Socialrådgivningenfinska _ svenska _ engelska
utkomststöd
Utkomststödet ( toimeentulotuki ) är avsett som en sista utväg då du inte har några andra inkomster eller medel , eller om dina inkomster är mycket låga .
utkomststöd kan du få om du inte lyckas få tillräckliga inkomster genom eget arbete , andras omsorg eller på något annat sätt .
du kan be om råd gällande ansökan om utkomststöd via den centraliserade telefontjänsten tfn ( 09 ) 8392.1119 .
linkkiVanda stad :
information om utkomststödfinska _ svenska _ engelska
ekonomi- och skuldrådgivning
om du inte kan betala dina räkningar eller skulder då de förfaller , ska du kontakta skuldrådgivningen ( velkaneuvonta ) .
tfn ( 09 ) 8392.2120 .
linkkiVanda ekonomi- och skuldrådgivning :
ekonomi- och skuldrådgivningfinska _ svenska _ engelska
social kreditgivning
om du har låga inkomster och är medellös samt har svårt att få lån , kan du ansöka om lån via den sociala kreditgivningen ( sosiaalinen luototus ) .
telefonnumret till kundrådgivningen och tidsbokningen är ( 09 ) 8392.0173 .
linkkiVanda stad :
information om social kreditgivningfinska _ svenska _ engelska
missbruksproblem och spelberoende
Itä @-@ Vantaan A @-@ klinikka
Konvaljvägen 20 C vån .
tfn ( 09 ) 8392.3415
Länsi @-@ Vantaan A @-@ klinikka
tfn ( 09 ) 8393.5534
H @-@ klinikka
Eldstadsvägen 7 B , vån .
tfn ( 09 ) 839.21064
H @-@ kliniken har också verksamhetsställen på Dickursby och Myrbacka hälsostationer .
om du har spelproblem kan du söka hjälp vid Spelkliniken ( Peliklinikka ) , som finns i centrala Helsingfors .
Peliklinikka
tfn 040.152.3918 .
ungdomscentralen Nuppi ( nuortenkeskus Nuppi ) hjälper ungdomar med missbruksproblem , Internetberoende eller spelberoende .
Nuppi ger också stöd till ungdomar som oroar sig för rusmedelsbruket hos någon närstående person .
Läs mer : missbruksproblem .
linkkiVanda stad :
hjälp med missbruksproblemfinska _ svenska _ engelska
linkkiVanda stad :
information om vård av drogproblemfinska _ svenska _ engelska
hjälp med penningspelproblemfinska
hjälp för ungafinska _ svenska _ engelska
Dödsfall
i Vanda finns fyra begravningsplatser som tillhör de evangelisk @-@ lutherska församlingarna .
i Furumo i Vanda finns dessutom Vandas och Helsingfors gemensamma begravningsplats för avlidna personer som inte har varit medlemmar i något religionssamfund .
information om begravning får du på Vanda församlingars gravkontor ( Vantaan seurakuntien hautaustoimisto ) och vid privata begravningsbyråer ( hautaustoimisto ) .
Vanda församlingars gravkontor
Prästgårdsgränden 5
tfn ( 09 ) 8306.220
om din närstående avlider plötsligt , kan du få hjälp med att återhämta dig från den chockartade upplevelsen och stöd i att klara dig efter förlusten av Vandas social- och krisjour ( sosiaali- ja kriisipäivystys ) .
jouren har öppet varje dag dygnet runt .
social- och krisjouren
tfn ( 09 ) 8392.4005
Läs mer : Död
linkkiVanda kyrkliga samfällighet :
Begravningsplatserfinska
linkkiHelsingfors kyrkliga samfällighet :
Konfessionslös begravningsplatsfinska
linkkiFinlands Begravningbyråers Förbund :
Begravningsbyråerfinska _ svenska _ engelska
när en närstående har avliditfinska _ svenska _ engelska
linkkiVanda stad :
social- och krisjourenfinska _ svenska _ engelska
problem med uppehållstillståndet
brott
behöver du en jurist ?
våld
missbruksproblem och spelberoende
Dödsfall
om du behöver brådskande hjälp av polisen , brandkåren eller ambulansen , ring nödnumret 112 .
du får ringa nödnumret endast i brådskande nödfall där liv , hälsa , egendom eller miljö är i fara .
om du drabbas av en akut krissituation , såsom att en närstående avlider eller på grund av familjevåld , kan du kontakta social- och krisjouren ( sosiaali- ja kriisipäivystys ) .
du kan också söka hjälp för en familjemedlem eller en vän .
social- och krisjouren har öppet dygnet runt varje dag .
social- och krisjouren
tfn ( 09 ) 8392.4005
linkkiNödcentralsverket :
hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
linkkiVanda stad :
social- och krisjourenfinska _ svenska _ engelska
problem med uppehållstillståndet
om du har problem eller oklarheter med uppehållstillståndet , kontakta Migrationsverket .
du kan även fråga om råd på rådgivningstjänsterna för invandrare .
information om tjänsterna finns på sidan Som invandrare i Vanda .
Migrationsverkets närmaste tjänsteställe finns i Helsingfors :
Göksgränd 3A
Läs mer : problem med uppehållstillståndet
olika tillståndfinska _ svenska _ engelska
hälsovård för papperslösa
i Helsingfors finns Global Clinic , där personer som vistas i Finland utan tillstånd kan få primärhälsovård .
tjänsterna vid Global Clinic är avgiftsfria för kunderna .
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter .
för att skydda kunderna uppges inte klinikens adress eller öppettider offentligt .
telefonnumret till Global Clinic i Helsingfors är 044.977.4547 .
Samtalet besvaras av en sjukskötare eller en läkare .
e @-@ postadressen är globalclinic.finland ( at ) gmail.com .
Läs mer : problem med uppehållstillstånd
hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
brott
brottsanmälan ( rikosilmoitus ) kan göras per telefon eller personligen på polisstationen .
du kan också göra brottsanmälan på internet om brottet i fråga är ringa och du inte behöver omedelbar hjälp av polisen .
Konvaljvägen 21
tfn 0295.430291
Läs mer : brott .
kontaktuppgifterfinska _ svenska
elektronisk polisanmälanfinska _ svenska _ engelska
behöver du en jurist ?
östra Nylands rättshjälpsbyrå ( Itä @-@ Uudenmaan oikeusaputoimisto ) betjänar invånarna i Vanda .
Pyrolavägen 37
tfn 029.5660.160
du kan också söka information om privata jurister på till exempel Finlands Juristförbunds ( Suomen Asianajajaliitto ) webbplats .
Läs mer : behöver du en jurist ?
linkkiÖstra Nylands rättshjälpsbyrå :
information om rättshjälpfinska _ svenska _ engelska
linkkiFinlands Advokatförbund :
Advokaterfinska _ svenska _ engelska
våld
i nödsituationer ringer du nödnumret 112 .
i krissituationer får man även hjälp vid Vanda stads social- och krisjour ( sosiaali- ja kriisipäivystys ) , som har öppet dygnet runt .
social- och krisjouren
tfn ( 09 ) 8392.4005
linkkiNödcentralsverket :
hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
skyddshem
om någon i din familj utövar våld mot dig eller hotar dig med våld , kan du kontakta ett skyddshem ( turvakoti ) .
Skyddshemmen har jourmottagning dygnet runt .
skyddshemmet Mona ( turvakoti Mona ) är ett skyddshem avsett för invandrarkvinnor och deras barn .
tfn 045.639.6274
linkkiTurvakoti Mona :
skyddshemfinska
du kan även gå till Vanda skyddshem ( Vantaan turvakoti ) eller huvudstadsregionens skyddshem ( pääkaupunkiseudun turvakoti ) .
Puh . ( 09 ) 8392.0071
skyddshemfinska _ engelska
Steniusvägen 20
tfn ( 09 ) 4777.180
hjälp till offer för familjevåldfinska
hjälp för invandrarkvinnor
föreningen Monika @-@ Naiset liitto ( Monika @-@ Naiset Liitto ) ger råd och stöd till invandrarkvinnor .
föreningen har ett resurscenter ( voimavarakeskus ) i Vanda där man får stöd och råd .
tfn ( 09 ) 839.35013
hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
hjälp för män
män som har utövat våld mot sina familjemedlemmar eller har själva blivit offer för våld i hemmet , kan få hjälp från Jussi @-@ arbetet i Vanda ( Vantaan Jussi @-@ työ ) .
hjälp för män att sluta med våldsamt beteendefinska
Miehen linja ( Miehen linja ) hjälper invandrarmän som har problem med våld .
tfn ( 09 ) 276.62899
hjälp för män för att sluta med våldsamt beteendefinska _ engelska
hjälp för unga
Finlands Röda Kors De ungas skyddshus ( Suomen Punaisen Ristin Nuorten turvatalo ) ger stöd och hjälp i krissituationer för 12 @-@ 19 @-@ åringar .
skyddshuset har öppet kl . 17 @-@ 10 , telefonjouren betjänar dygnet runt .
Sjukhusgatan 3 ( Räckhals gård )
tfn ( 09 ) 871.4043
linkkiFinlands Röda Kors :
de ungas skyddshusfinska _ svenska _ engelska
Läs mer : våld
problem i äktenskap eller parförhållande
par med barn under 13 år kan vid problem i äktenskap och parförhållande få hjälp vid familjerådgivningen ( perheneuvola ) .
kontaktuppgifterna hittar du på Vanda stads webbplats .
Familjerådgivningens tjänster är konfidentiella och avgiftsfria .
vid akuta krissituationer inom familjen kan du kontakta social- och krisjouren ( sosiaali- ja kriisipäivystys ) , som har öppet dygnet runt varje dag .
social- och krisjouren
tfn ( 09 ) 8392.4005
vid problem i parförhållandet och familjen får man även hjälp av familjerådgivningen vid Vanda församlingar ( Vantaan seurakunnan perheneuvonta ) .
Läs mer : problem i äktenskap och parförhållande
linkkiVanda stad :
Familjerådgivningarfinska _ svenska
linkkiVanda kyrkliga samfällighet :
familjerådgivningfinska _ engelska
Barnrådgivningsbyråerna ( lastenneuvola ) och familjerådgivningsbyråerna ( perheneuvola ) ger råd i frågor som rör barns hälsa , uppväxt och utveckling .
vid problem hos barn i skolåldern får man hjälp hos skolhälsovårdarna ( kouluterveydenhoitaja ) , skolkuratorerna ( koulukuraattori ) och socialhandledarna ( sosiaaliohjaaja ) .
mer information hittar du på Vanda stads webbplats .
Läs mer : barns och ungas problem
linkkiVanda stad :
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad :
Familjerådgivningarfinska _ svenska
linkkiVanda stad :
information om tjänster för barn , ungdomar och familjerfinska _ svenska _ engelska
i skolan får de unga hjälp av skol- och studenthälsovårdarna ( koulu- ja opiskeluterveydenhoitajat ) , skolkuratorerna ( koulukuraattorit ) och skolpsykologerna ( koulupsykologit ) .
linkkiVanda stad :
information om skolhälsovårdenfinska _ svenska _ engelska
linkkiVanda stad :
Skolkuratorerfinska _ svenska
linkkiVanda stad :
Skolpsykologerfinska _ svenska
Nuppi
13 @-@ 21 @-@ åriga barn och ungdomar samt deras familjer kan få hjälp hos ungdomscentralen ( nuortenkeskus ) .
på Nuppi kan du till exempel få hjälp med mentala problem och missbruksproblem .
hjälp för ungafinska _ svenska _ engelska
om du är under 30 år , kan du få råd och handledning via tjänsten Navigatorn .
Personalen vid Navigatorn hjälper dig om du inte har något arbete eller en studieplats .
du kan även be om råd gällande andra saker , till exempel boende och ekonomi .
de ungas skyddshus
Finlands Röda Kors De ungas skyddshus ( Suomen Punaisen Ristin Nuorten turvatalo ) ger stöd och hjälp i krissituationer för 12 @-@ 19 @-@ åringar .
skyddshuset har öppet kl . 17 @-@ 10 , telefonjouren betjänar dygnet runt .
Sjukhusgatan 3
tfn ( 09 ) 871.4043
Läs mer : barns och ungas problem
linkkiFinlands Röda Kors :
de ungas skyddshusfinska _ svenska _ engelska
vägledning och stöd för ungafinska _ svenska
Socialrådgivningen ( sosiaalineuvonta ) ger information om utkomststöd ( toimeentulotuki ) och andra bidrag om du har ekonomiska problem .
tfn ( 09 ) 83.911 .
linkkiVanda stad :
Socialrådgivningenfinska _ svenska _ engelska
utkomststöd
Utkomststödet ( toimeentulotuki ) är avsett som en sista utväg då du inte har några andra inkomster eller medel , eller om dina inkomster är mycket låga .
utkomststöd kan du få om du inte lyckas få tillräckliga inkomster genom eget arbete , andras omsorg eller på något annat sätt .
du kan be om råd gällande ansökan om utkomststöd via den centraliserade telefontjänsten tfn ( 09 ) 8392.1119 .
linkkiVanda stad :
information om utkomststödfinska _ svenska _ engelska
ekonomi- och skuldrådgivning
om du inte kan betala dina räkningar eller skulder då de förfaller , ska du kontakta skuldrådgivningen ( velkaneuvonta ) .
tfn ( 09 ) 8392.2120 .
linkkiVanda ekonomi- och skuldrådgivning :
ekonomi- och skuldrådgivningfinska _ svenska _ engelska
social kreditgivning
om du har låga inkomster och är medellös samt har svårt att få lån , kan du ansöka om lån via den sociala kreditgivningen ( sosiaalinen luototus ) .
telefonnumret till kundrådgivningen och tidsbokningen är ( 09 ) 8392.0173 .
linkkiVanda stad :
information om social kreditgivningfinska _ svenska _ engelska
missbruksproblem och spelberoende
Itä @-@ Vantaan A @-@ klinikka
Konvaljvägen 20 C vån .
tfn ( 09 ) 8392.3415
Länsi @-@ Vantaan A @-@ klinikka
tfn ( 09 ) 8393.5534
H @-@ klinikka
Eldstadsvägen 7 B , vån .
tfn ( 09 ) 839.21064
H @-@ kliniken har också verksamhetsställen på Dickursby och Myrbacka hälsostationer .
om du har spelproblem kan du söka hjälp vid Spelkliniken ( Peliklinikka ) , som finns i centrala Helsingfors .
Peliklinikka
tfn 040.152.3918 .
ungdomscentralen Nuppi ( nuortenkeskus Nuppi ) hjälper ungdomar med missbruksproblem , Internetberoende eller spelberoende .
Nuppi ger också stöd till ungdomar som oroar sig för rusmedelsbruket hos någon närstående person .
Läs mer : missbruksproblem .
linkkiVanda stad :
hjälp med missbruksproblemfinska _ svenska _ engelska
linkkiVanda stad :
information om vård av drogproblemfinska _ svenska _ engelska
hjälp med penningspelproblemfinska
hjälp för ungafinska _ svenska _ engelska
Dödsfall
i Vanda finns fyra begravningsplatser som tillhör de evangelisk @-@ lutherska församlingarna .
i Furumo i Vanda finns dessutom Vandas och Helsingfors gemensamma begravningsplats för avlidna personer som inte har varit medlemmar i något religionssamfund .
information om begravning får du på Vanda församlingars gravkontor ( Vantaan seurakuntien hautaustoimisto ) och vid privata begravningsbyråer ( hautaustoimisto ) .
Vanda församlingars gravkontor
Prästgårdsgränden 5
tfn ( 09 ) 8306.220
om din närstående avlider plötsligt , kan du få hjälp med att återhämta dig från den chockartade upplevelsen och stöd i att klara dig efter förlusten av Vandas social- och krisjour ( sosiaali- ja kriisipäivystys ) .
jouren har öppet varje dag dygnet runt .
social- och krisjouren
tfn ( 09 ) 8392.4005
Läs mer : Död
linkkiVanda kyrkliga samfällighet :
Begravningsplatserfinska
linkkiHelsingfors kyrkliga samfällighet :
Konfessionslös begravningsplatsfinska
linkkiFinlands Begravningbyråers Förbund :
Begravningsbyråerfinska
när en närstående har avliditfinska _ svenska _ engelska
linkkiVanda stad :
social- och krisjourenfinska _ svenska _ engelska
problem med uppehållstillståndet
brott
behöver du en jurist ?
våld
missbruksproblem och spelberoende
Dödsfall
om du behöver brådskande hjälp av polisen , brandkåren eller ambulansen , ring nödnumret 112 .
du får ringa nödnumret endast i brådskande nödfall där liv , hälsa , egendom eller miljö är i fara .
om du drabbas av en akut krissituation , såsom att en närstående avlider eller på grund av familjevåld , kan du kontakta social- och krisjouren ( sosiaali- ja kriisipäivystys ) .
du kan också söka hjälp för en familjemedlem eller en vän .
social- och krisjouren har öppet dygnet runt varje dag .
social- och krisjouren
tfn ( 09 ) 8392.4005
linkkiNödcentralsverket :
hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
linkkiVanda stad :
social- och krisjourenfinska _ svenska _ engelska
problem med uppehållstillståndet
om du har problem eller oklarheter med uppehållstillståndet , kontakta Migrationsverket .
du kan även fråga om råd på rådgivningstjänsterna för invandrare .
information om tjänsterna finns på sidan Som invandrare i Vanda .
Migrationsverkets närmaste tjänsteställe finns i Helsingfors :
Göksgränd 3A
Läs mer : problem med uppehållstillståndet
olika tillståndfinska _ svenska _ engelska
hälsovård för papperslösa
i Helsingfors finns Global Clinic , där personer som vistas i Finland utan tillstånd kan få primärhälsovård .
tjänsterna vid Global Clinic är avgiftsfria för kunderna .
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter .
för att skydda kunderna uppges inte klinikens adress eller öppettider offentligt .
telefonnumret till Global Clinic i Helsingfors är 044.977.4547 .
Samtalet besvaras av en sjukskötare eller en läkare .
e @-@ postadressen är globalclinic.finland ( at ) gmail.com .
Läs mer : problem med uppehållstillstånd
hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
brott
brottsanmälan ( rikosilmoitus ) kan göras per telefon eller personligen på polisstationen .
du kan också göra brottsanmälan på internet om brottet i fråga är ringa och du inte behöver omedelbar hjälp av polisen .
Konvaljvägen 21
tfn 0295.430291
Läs mer : brott .
kontaktuppgifterfinska _ svenska
elektronisk polisanmälanfinska _ svenska _ engelska
behöver du en jurist ?
östra Nylands rättshjälpsbyrå ( Itä @-@ Uudenmaan oikeusaputoimisto ) betjänar invånarna i Vanda .
Pyrolavägen 37
tfn 029.5660.160
du kan också söka information om privata jurister på till exempel Finlands Juristförbunds ( Suomen Asianajajaliitto ) webbplats .
Läs mer : behöver du en jurist ?
linkkiÖstra Nylands rättshjälpsbyrå :
information om rättshjälpfinska _ svenska _ engelska
linkkiFinlands Advokatförbund :
Advokaterfinska _ svenska _ engelska
våld
i nödsituationer ringer du nödnumret 112 .
i krissituationer får man även hjälp vid Vanda stads social- och krisjour ( sosiaali- ja kriisipäivystys ) , som har öppet dygnet runt .
social- och krisjouren
tfn ( 09 ) 8392.4005
linkkiNödcentralsverket :
hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
skyddshem
om någon i din familj utövar våld mot dig eller hotar dig med våld , kan du kontakta ett skyddshem ( turvakoti ) .
Skyddshemmen har jourmottagning dygnet runt .
skyddshemmet Mona ( turvakoti Mona ) är ett skyddshem avsett för invandrarkvinnor och deras barn .
tfn 045.639.6274
linkkiTurvakoti Mona :
skyddshemfinska
du kan även gå till Vanda skyddshem ( Vantaan turvakoti ) eller huvudstadsregionens skyddshem ( pääkaupunkiseudun turvakoti ) .
Puh . ( 09 ) 8392.0071
skyddshemfinska _ engelska
Steniusvägen 20
tfn ( 09 ) 4777.180
hjälp till offer för familjevåldfinska
hjälp för invandrarkvinnor
föreningen Monika @-@ Naiset liitto ( Monika @-@ Naiset Liitto ) ger råd och stöd till invandrarkvinnor .
föreningen har ett resurscenter ( voimavarakeskus ) i Vanda där man får stöd och råd .
tfn ( 09 ) 839.35013
hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
hjälp för män
män som har utövat våld mot sina familjemedlemmar eller har själva blivit offer för våld i hemmet , kan få hjälp från Jussi @-@ arbetet i Vanda ( Vantaan Jussi @-@ työ ) .
hjälp för män att sluta med våldsamt beteendefinska
Miehen linja ( Miehen linja ) hjälper invandrarmän som har problem med våld .
tfn ( 09 ) 276.62899
hjälp för män för att sluta med våldsamt beteendefinska _ engelska
hjälp för unga
Finlands Röda Kors De ungas skyddshus ( Suomen Punaisen Ristin Nuorten turvatalo ) ger stöd och hjälp i krissituationer för 12 @-@ 19 @-@ åringar .
skyddshuset har öppet kl . 17 @-@ 10 , telefonjouren betjänar dygnet runt .
Sjukhusgatan 3 ( Räckhals gård )
tfn ( 09 ) 871.4043
linkkiFinlands Röda Kors :
de ungas skyddshusfinska _ svenska _ engelska
Läs mer : våld
problem i äktenskap eller parförhållande
par med barn under 13 år kan vid problem i äktenskap och parförhållande få hjälp vid familjerådgivningen ( perheneuvola ) .
kontaktuppgifterna hittar du på Vanda stads webbplats .
Familjerådgivningens tjänster är konfidentiella och avgiftsfria .
vid akuta krissituationer inom familjen kan du kontakta social- och krisjouren ( sosiaali- ja kriisipäivystys ) , som har öppet dygnet runt varje dag .
social- och krisjouren
tfn ( 09 ) 8392.4005
vid problem i parförhållandet och familjen får man även hjälp av familjerådgivningen vid Vanda församlingar ( Vantaan seurakunnan perheneuvonta ) .
Läs mer : problem i äktenskap och parförhållande
linkkiVanda stad :
Familjerådgivningarfinska _ svenska
linkkiVanda kyrkliga samfällighet :
familjerådgivningfinska _ engelska
Barnrådgivningsbyråerna ( lastenneuvola ) och familjerådgivningsbyråerna ( perheneuvola ) ger råd i frågor som rör barns hälsa , uppväxt och utveckling .
vid problem hos barn i skolåldern får man hjälp hos skolhälsovårdarna ( kouluterveydenhoitaja ) , skolkuratorerna ( koulukuraattori ) och socialhandledarna ( sosiaaliohjaaja ) .
mer information hittar du på Vanda stads webbplats .
Läs mer : barns och ungas problem
linkkiVanda stad :
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad :
Familjerådgivningarfinska _ svenska
linkkiVanda stad :
information om tjänster för barn , ungdomar och familjerfinska _ svenska _ engelska
i skolan får de unga hjälp av skol- och studenthälsovårdarna ( koulu- ja opiskeluterveydenhoitajat ) , skolkuratorerna ( koulukuraattorit ) och skolpsykologerna ( koulupsykologit ) .
linkkiVanda stad :
information om skolhälsovårdenfinska _ svenska _ engelska
linkkiVanda stad :
Skolkuratorerfinska _ svenska
linkkiVanda stad :
Skolpsykologerfinska _ svenska
Nuppi
13 @-@ 21 @-@ åriga barn och ungdomar samt deras familjer kan få hjälp hos ungdomscentralen ( nuortenkeskus ) .
på Nuppi kan du till exempel få hjälp med mentala problem och missbruksproblem .
hjälp för ungafinska _ svenska _ engelska
om du är under 30 år , kan du få råd och handledning via tjänsten Navigatorn .
Personalen vid Navigatorn hjälper dig om du inte har något arbete eller en studieplats .
du kan även be om råd gällande andra saker , till exempel boende och ekonomi .
de ungas skyddshus
Finlands Röda Kors De ungas skyddshus ( Suomen Punaisen Ristin Nuorten turvatalo ) ger stöd och hjälp i krissituationer för 12 @-@ 19 @-@ åringar .
skyddshuset har öppet kl . 17 @-@ 10 , telefonjouren betjänar dygnet runt .
Sjukhusgatan 3
tfn ( 09 ) 871.4043
Läs mer : barns och ungas problem
linkkiFinlands Röda Kors :
de ungas skyddshusfinska _ svenska _ engelska
vägledning och stöd för ungafinska _ svenska
Socialrådgivningen ( sosiaalineuvonta ) ger information om utkomststöd ( toimeentulotuki ) och andra bidrag om du har ekonomiska problem .
tfn ( 09 ) 83.911 .
linkkiVanda stad :
Socialrådgivningenfinska _ svenska _ engelska
utkomststöd
Utkomststödet ( toimeentulotuki ) är avsett som en sista utväg då du inte har några andra inkomster eller medel , eller om dina inkomster är mycket låga .
utkomststöd kan du få om du inte lyckas få tillräckliga inkomster genom eget arbete , andras omsorg eller på något annat sätt .
du kan be om råd gällande ansökan om utkomststöd via den centraliserade telefontjänsten tfn ( 09 ) 8392.1119 .
linkkiVanda stad :
information om utkomststödfinska _ svenska _ engelska
ekonomi- och skuldrådgivning
om du inte kan betala dina räkningar eller skulder då de förfaller , ska du kontakta skuldrådgivningen ( velkaneuvonta ) .
tfn 029.566.0175 .
linkkiVanda ekonomi- och skuldrådgivning :
ekonomi- och skuldrådgivningfinska _ svenska _ engelska
social kreditgivning
om du har låga inkomster och är medellös samt har svårt att få lån , kan du ansöka om lån via den sociala kreditgivningen ( sosiaalinen luototus ) .
telefonnumret till kundrådgivningen och tidsbokningen är ( 09 ) 8392.0173 .
linkkiVanda stad :
information om social kreditgivningfinska _ svenska _ engelska
missbruksproblem och spelberoende
Itä @-@ Vantaan A @-@ klinikka
Konvaljvägen 20 C vån .
tfn ( 09 ) 8392.3415
Länsi @-@ Vantaan A @-@ klinikka
tfn ( 09 ) 8393.5534
H @-@ klinikka
Eldstadsvägen 7 B , vån .
tfn ( 09 ) 839.21064
H @-@ kliniken har också verksamhetsställen på Dickursby och Myrbacka hälsostationer .
om du har spelproblem kan du söka hjälp vid Spelkliniken ( Peliklinikka ) , som finns i centrala Helsingfors .
Peliklinikka
tfn 040.152.3918 .
ungdomscentralen Nuppi ( nuortenkeskus Nuppi ) hjälper ungdomar med missbruksproblem , Internetberoende eller spelberoende .
Nuppi ger också stöd till ungdomar som oroar sig för rusmedelsbruket hos någon närstående person .
Läs mer : missbruksproblem .
linkkiVanda stad :
hjälp med missbruksproblemfinska _ svenska _ engelska
linkkiVanda stad :
information om vård av drogproblemfinska _ svenska _ engelska
hjälp med penningspelproblemfinska
hjälp för ungafinska _ svenska _ engelska
Dödsfall
i Vanda finns fyra begravningsplatser som tillhör de evangelisk @-@ lutherska församlingarna .
i Furumo i Vanda finns dessutom Vandas och Helsingfors gemensamma begravningsplats för avlidna personer som inte har varit medlemmar i något religionssamfund .
information om begravning får du på Vanda församlingars gravkontor ( Vantaan seurakuntien hautaustoimisto ) och vid privata begravningsbyråer ( hautaustoimisto ) .
Vanda församlingars gravkontor
Prästgårdsgränden 5
tfn ( 09 ) 8306.220
om din närstående avlider plötsligt , kan du få hjälp med att återhämta dig från den chockartade upplevelsen och stöd i att klara dig efter förlusten av Vandas social- och krisjour ( sosiaali- ja kriisipäivystys ) .
jouren har öppet varje dag dygnet runt .
social- och krisjouren
tfn ( 09 ) 8392.4005
Läs mer : Död
linkkiVanda kyrkliga samfällighet :
Begravningsplatserfinska
linkkiHelsingfors kyrkliga samfällighet :
Konfessionslös begravningsplatsfinska
linkkiFinlands Begravningbyråers Förbund :
Begravningsbyråerfinska
när en närstående har avliditfinska _ svenska _ engelska
linkkiVanda stad :
social- och krisjourenfinska _ svenska _ engelska
äktenskap
skilsmässa
barnets födelse
vård av barn
problem i familjen
äktenskap
före äktenskapet ska du skriftligt begära hindersprövning ( avioliiton esteiden tutkiminen ) .
Hindersprövningen görs på magistraten ( maistraatti ) .
du kan begära hindersprövning på vilken magistrat som helst .
mer information hittar du på magistratens webbplats .
också borgerliga vigslar förrättas på magistraten .
Konvaljvägen 15 , PB 112
01301 Vanda
Läs mer : äktenskap .
Anhållan om prövning av hinder mot äktenskapfinska _ svenska
Ingående av äktenskapfinska _ svenska _ engelska
linkkiVanda församlingar :
information om kyrklig vigselfinska _ svenska _ engelska
linkkiHelsingfors ortodoxa församling :
information om ortodox vigselfinska _ ryska
skilsmässa
kvinnan eller mannen kan lämna in skilsmässoansökan i Vanda tingsrätts kansli .
makarna kan ansöka om skilsmässa tillsammans eller också kan den ena maken göra det ensam .
ansökan kan lämnas till tingsrättens kansli eller skickas dit per post , fax eller via e @-@ post .
tfn 029.56.45200
Läs mer : skilsmässa .
linkkiVanda stad :
information om skilsmässafinska _ engelska
att ansöka om skilsmässafinska _ svenska _ engelska
om du har barn och ska skilja dig tar du kontakt med barnatillsyningsmannen ( lastenvalvoja ) vid Vanda stad .
Socialväsendet bekräftar ett avtal om barnens boende , vårdnad , umgängesrätt och underhållsbidrag .
barnatillsyningsmännen ger även råd till föräldrar som ska skiljas .
kontaktuppgifterna till barnatillsyningsmannen hittar du på Vanda stads webbplats .
Läs mer :
barn vid skilsmässa .
linkkiVanda stad :
kontaktuppgifter till barnatillsyningsmännenfinska _ svenska _ engelska
barnets födelse
Uppgifterna om barnets födelse skickas från sjukhuset till befolkningsdataregistret i Finland .
du ska meddela barnets namn , modersmål och andra erforderliga uppgifter till magistraten ( Maistraatti ) med en separat blankett som skickas hem till dig .
du kan läsa mer om registrering av barnets födelse , faderskapserkännande och vårdnaden om barnet på InfoFinlands sida : när ett barn föds i Finland .
vård av barn
dagvård
på InfoFinlands sida Utbildning i Vanda hittar du information om dagvård för barn i Vanda .
hemvårdsstöd
om du tar hand om ett under treårigt barn , kan du få hemvårdsstöd ( kotihoidon tuki ) .
du ansöker om hemvårdsstödet hos FPA .
Vanda stad betalar dessutom ett kommuntillägg till hemvårdsstödet för barn till de familjer som vårdar ett under 1 ½ -årigt barn i hemmet .
du behöver inte ansöka separat om stödet , utan FPA betalar ut Vandatillägget ( Vantaa @-@ lisä ) med hemvårdsstödet .
information om hemvårdsstödfinska _ svenska _ engelska
linkkiVanda stad :
information om hemvårdsstödets kommuntilläggfinska _ svenska _ engelska
öppna daghem och invånarparker
öppna daghem ( avoin päiväkoti ) är avsedda för barn under skolåldern och de föräldrar och vårdare som tar hand om dem .
invånarparker ( asukaspuistot ) är avsedda för barn i alla åldrar och deras föräldrar eller vårdare .
små barn kan delta i verksamheten tillsammans med sin förälder eller vårdare .
verksamheten i öppna daghem och invånarparker är kostnadsfri och du behöver inte anmäla dig på förhand .
i verksamheten ingår lek och ledda aktiviteter , till exempel musik , motion och utflykter .
linkkiVanda stad :
Parker för invånare och öppna daghemfinska _ svenska _ engelska
klubbar
Vanda stad ordnar även klubbar ( kerho ) för 2,5 @-@ 5 @-@ åriga barn som vårdas i hemmet .
Klubbarna är avgiftsfria .
i klubben lär sig barnet tala finska , fungera i en grupp och där kan barnet träffa andra barn .
till klubben ansöker du om plats med samma ansökan om småbarnsfostran ( varhaiskasvatushakemus ) , med vilken du även ansöker om dagvårdsplats .
linkkiVanda stad :
Klubbverksamhetfinska _ svenska _ engelska
Barnpassningsservice för barn
om du vårdar ditt barn i hemmet och behöver tillfälligt en vårdplats för barnet , till exempel när du ska sköta ärenden , kan du kontakta barnpassningsservicen ( hoitoapupalvelu ) .
Barnpassningen är avgiftsbelagd .
linkkiVanda stad :
Barnpassningsservice för barnfinska _ engelska
tillfällig barnpassning
om du behöver tillfällig barnpassning i hemmet , kan du kontakta Mannerheims Barnskyddsförbund eller Väestöliitto .
den tillfälliga barnpassningshjälpen är avgiftsbelagd .
Läs mer : vård av barnet
linkkiMannerheims barnskyddsförbund :
Barnvaktshjälpfinska _ engelska
linkkiVanda stad :
hjälp i hemmet för barnfamiljer ( pdf , 500 kb ) finska _ engelska
problem i familjen
om du misstänker att ditt barn eller din ungdom behöver barnskyddets ( lastensuojelu ) hjälp , ska du kontakta en socialarbetare .
tfn växeln 09.83.911
mån @-@ fre kl . 8.15 @-@ 16.00
kvällar och helger
social- och krisjouren
tfn 09.8392.4005
linkkiVanda stad :
Barnskyddsanmälanfinska _ engelska
på InfoFinlands sida Problematiska situationer i Vanda hittar du information om var någonstans i Vanda det finns hjälp att få till barns och ungas problem .
information om barns och ungas problem finns även på InfoFinlands sidor Barns och ungas problem och Barnskydd .
på InfoFinlands sida Problem i äktenskap och parförhållande finns information om var man kan få hjälp med problem i parförhållanden .
äktenskap
skilsmässa
barnets födelse
vård av barn
problem i familjen
äldre människor
äktenskap
före äktenskapet ska du skriftligt begära hindersprövning ( avioliiton esteiden tutkiminen ) .
Hindersprövningen görs på magistraten ( maistraatti ) .
du kan begära hindersprövning på vilken magistrat som helst .
mer information hittar du på magistratens webbplats .
också borgerliga vigslar förrättas på magistraten .
Konvaljvägen 15 , PB 112
01301 Vanda
Läs mer : äktenskap .
Anhållan om prövning av hinder mot äktenskapfinska _ svenska
Ingående av äktenskapfinska _ svenska _ engelska
linkkiVanda församlingar :
information om kyrklig vigselfinska _ svenska _ engelska
linkkiHelsingfors ortodoxa församling :
information om ortodox vigselfinska _ ryska
skilsmässa
kvinnan eller mannen kan lämna in skilsmässoansökan i Vanda tingsrätts kansli .
makarna kan ansöka om skilsmässa tillsammans eller också kan den ena maken göra det ensam .
ansökan kan lämnas till tingsrättens kansli eller skickas dit per post , fax eller via e @-@ post .
tfn 029.56.45200
Läs mer : skilsmässa .
linkkiVanda stad :
information om skilsmässafinska _ engelska
att ansöka om skilsmässafinska _ svenska _ engelska
om du har barn och ska skilja dig tar du kontakt med barnatillsyningsmannen ( lastenvalvoja ) vid Vanda stad .
Socialväsendet bekräftar ett avtal om barnens boende , vårdnad , umgängesrätt och underhållsbidrag .
barnatillsyningsmännen ger även råd till föräldrar som ska skiljas .
kontaktuppgifterna till barnatillsyningsmannen hittar du på Vanda stads webbplats .
Läs mer :
barn vid skilsmässa .
linkkiVanda stad :
kontaktuppgifter till barnatillsyningsmännenfinska _ svenska _ engelska
barnets födelse
Uppgifterna om barnets födelse skickas från sjukhuset till befolkningsdataregistret i Finland .
du ska meddela barnets namn , modersmål och andra erforderliga uppgifter till magistraten ( Maistraatti ) med en separat blankett som skickas hem till dig .
du kan läsa mer om registrering av barnets födelse , faderskapserkännande och vårdnaden om barnet på InfoFinlands sida : när ett barn föds i Finland .
vård av barn
dagvård
på InfoFinlands sida Utbildning i Vanda hittar du information om dagvård för barn i Vanda .
hemvårdsstöd
om du tar hand om ett under treårigt barn , kan du få hemvårdsstöd ( kotihoidon tuki ) .
du ansöker om hemvårdsstödet hos FPA .
Vanda stad betalar dessutom ett kommuntillägg till hemvårdsstödet för barn till de familjer som vårdar ett under 1 ½ -årigt barn i hemmet .
du behöver inte ansöka separat om stödet , utan FPA betalar ut Vandatillägget ( Vantaa @-@ lisä ) med hemvårdsstödet .
information om hemvårdsstödfinska _ svenska _ engelska
linkkiVanda stad :
information om hemvårdsstödets kommuntilläggfinska _ svenska _ engelska
öppna daghem och invånarparker
öppna daghem ( avoin päiväkoti ) är avsedda för barn under skolåldern och de föräldrar och vårdare som tar hand om dem .
invånarparker ( asukaspuistot ) är avsedda för barn i alla åldrar och deras föräldrar eller vårdare .
små barn kan delta i verksamheten tillsammans med sin förälder eller vårdare .
verksamheten i öppna daghem och invånarparker är kostnadsfri och du behöver inte anmäla dig på förhand .
i verksamheten ingår lek och ledda aktiviteter , till exempel musik , motion och utflykter .
linkkiVanda stad :
Parker för invånare och öppna daghemfinska _ svenska _ engelska
klubbar
Vanda stad ordnar även klubbar ( kerho ) för 2,5 @-@ 5 @-@ åriga barn som vårdas i hemmet .
Klubbarna är avgiftsfria .
i klubben lär sig barnet tala finska , fungera i en grupp och där kan barnet träffa andra barn .
till klubben ansöker du om plats med samma ansökan om småbarnsfostran ( varhaiskasvatushakemus ) , med vilken du även ansöker om dagvårdsplats .
linkkiVanda stad :
Klubbverksamhetfinska _ svenska _ engelska
Barnpassningsservice för barn
om du vårdar ditt barn i hemmet och behöver tillfälligt en vårdplats för barnet , till exempel när du ska sköta ärenden , kan du kontakta barnpassningsservicen ( hoitoapupalvelu ) .
Barnpassningen är avgiftsbelagd .
linkkiVanda stad :
Barnpassningsservice för barnfinska _ engelska
tillfällig barnpassning
om du behöver tillfällig barnpassning i hemmet , kan du kontakta Mannerheims Barnskyddsförbund eller Väestöliitto .
den tillfälliga barnpassningshjälpen är avgiftsbelagd .
Läs mer : vård av barnet
linkkiMannerheims barnskyddsförbund :
Barnvaktshjälpfinska _ engelska
linkkiVanda stad :
hjälp i hemmet för barnfamiljer ( pdf , 500 kb ) finska _ engelska
problem i familjen
om du misstänker att ditt barn eller din ungdom behöver barnskyddets ( lastensuojelu ) hjälp , ska du kontakta en socialarbetare .
tfn växeln 09.83.911
mån @-@ fre kl . 8.15 @-@ 16.00
kvällar och helger
social- och krisjouren
tfn 09.8392.4005
linkkiVanda stad :
Barnskyddsanmälanfinska _ engelska
på InfoFinlands sida Problematiska situationer i Vanda hittar du information om var någonstans i Vanda det finns hjälp att få till barns och ungas problem .
information om barns och ungas problem finns även på InfoFinlands sidor Barns och ungas problem och Barnskydd .
på InfoFinlands sida Problem i äktenskap och parförhållande finns information om var man kan få hjälp med problem i parförhållanden .
äldre människor
i Vanda finns tjänster som är särskilt avsedda för äldre .
du får information om dem vid seniorrådgivningen .
seniorrådgivningen Tfn : 09.8392.4202
när du tar hand om en anhörig i hemmet
när en familjemedlem behöver kontinuerlig hjälp och vården är både bindande och krävande , finns det möjlighet att få stöd för närståendevård av kommunen .
seniorrådgivningen bedömer behovet av anhörigvård för en äldre person .
Läs mer : äldre människor .
linkkiVanda stad :
Seniorrådgivningenfinska _ svenska _ engelska
äktenskap
skilsmässa
barnets födelse
vård av barn
problem i familjen
äldre människor
äktenskap
före äktenskapet ska du skriftligt begära hindersprövning ( avioliiton esteiden tutkiminen ) .
Hindersprövningen görs på magistraten ( maistraatti ) .
du kan begära hindersprövning på vilken magistrat som helst .
mer information hittar du på magistratens webbplats .
också borgerliga vigslar förrättas på magistraten .
Konvaljvägen 15 , PB 112
01301 Vanda
Läs mer : äktenskap .
Anhållan om prövning av hinder mot äktenskapfinska _ svenska _ engelska
Ingående av äktenskapfinska _ svenska _ engelska
linkkiVanda församlingar :
information om kyrklig vigselfinska _ svenska _ engelska
linkkiHelsingfors ortodoxa församling :
information om ortodox vigselfinska _ ryska
skilsmässa
kvinnan eller mannen kan lämna in skilsmässoansökan i Vanda tingsrätts kansli .
makarna kan ansöka om skilsmässa tillsammans eller också kan den ena maken göra det ensam .
ansökan kan lämnas till tingsrättens kansli eller skickas dit per post , fax eller via e @-@ post .
tfn 029.56.45200
Läs mer : skilsmässa .
linkkiVanda stad :
information om skilsmässafinska _ engelska
att ansöka om skilsmässafinska _ svenska _ engelska
om du har barn och ska skilja dig tar du kontakt med barnatillsyningsmannen ( lastenvalvoja ) vid Vanda stad .
Socialväsendet bekräftar ett avtal om barnens boende , vårdnad , umgängesrätt och underhållsbidrag .
barnatillsyningsmännen ger även råd till föräldrar som ska skiljas .
kontaktuppgifterna till barnatillsyningsmannen hittar du på Vanda stads webbplats .
Läs mer :
barn vid skilsmässa .
linkkiVanda stad :
kontaktuppgifter till barnatillsyningsmännenfinska _ svenska _ engelska
barnets födelse
Uppgifterna om barnets födelse skickas från sjukhuset till befolkningsdataregistret i Finland .
du ska meddela barnets namn , modersmål och andra erforderliga uppgifter till magistraten ( Maistraatti ) med en separat blankett som skickas hem till dig .
du kan läsa mer om registrering av barnets födelse , faderskapserkännande och vårdnaden om barnet på InfoFinlands sida : när ett barn föds i Finland .
vård av barn
dagvård
på InfoFinlands sida Utbildning i Vanda hittar du information om dagvård för barn i Vanda .
hemvårdsstöd
om du tar hand om ett under treårigt barn , kan du få hemvårdsstöd ( kotihoidon tuki ) .
du ansöker om hemvårdsstödet hos FPA .
Vanda stad betalar dessutom ett kommuntillägg till hemvårdsstödet för barn till de familjer som vårdar ett under 1 ½ -årigt barn i hemmet .
du behöver inte ansöka separat om stödet , utan FPA betalar ut Vandatillägget ( Vantaa @-@ lisä ) med hemvårdsstödet .
information om hemvårdsstödfinska _ svenska _ engelska
linkkiVanda stad :
information om hemvårdsstödets kommuntilläggfinska _ svenska _ engelska
öppna daghem och invånarparker
öppna daghem ( avoin päiväkoti ) är avsedda för barn under skolåldern och de föräldrar och vårdare som tar hand om dem .
invånarparker ( asukaspuistot ) är avsedda för barn i alla åldrar och deras föräldrar eller vårdare .
små barn kan delta i verksamheten tillsammans med sin förälder eller vårdare .
verksamheten i öppna daghem och invånarparker är kostnadsfri och du behöver inte anmäla dig på förhand .
i verksamheten ingår lek och ledda aktiviteter , till exempel musik , motion och utflykter .
linkkiVanda stad :
Parker för invånare och öppna daghemfinska _ svenska _ engelska
klubbar
Vanda stad ordnar även klubbar ( kerho ) för 2,5 @-@ 5 @-@ åriga barn som vårdas i hemmet .
Klubbarna är avgiftsfria .
i klubben lär sig barnet tala finska , fungera i en grupp och där kan barnet träffa andra barn .
till klubben ansöker du om plats med samma ansökan om småbarnsfostran ( varhaiskasvatushakemus ) , med vilken du även ansöker om dagvårdsplats .
linkkiVanda stad :
Klubbverksamhetfinska _ svenska _ engelska
Barnpassningsservice för barn
om du vårdar ditt barn i hemmet och behöver tillfälligt en vårdplats för barnet , till exempel när du ska sköta ärenden , kan du kontakta barnpassningsservicen ( hoitoapupalvelu ) .
Barnpassningen är avgiftsbelagd .
linkkiVanda stad :
Barnpassningsservice för barnfinska _ engelska
tillfällig barnpassning
om du behöver tillfällig barnpassning i hemmet , kan du kontakta Mannerheims Barnskyddsförbund eller Väestöliitto .
den tillfälliga barnpassningshjälpen är avgiftsbelagd .
Läs mer : vård av barnet
linkkiMannerheims barnskyddsförbund :
Barnvaktshjälpfinska _ engelska
linkkiVanda stad :
hjälp i hemmet för barnfamiljer ( pdf , 500 kb ) finska _ engelska
problem i familjen
om du misstänker att ditt barn eller din ungdom behöver barnskyddets ( lastensuojelu ) hjälp , ska du kontakta en socialarbetare .
tfn växeln 09.83.911
mån @-@ fre kl . 8.15 @-@ 16.00
kvällar och helger
social- och krisjouren
tfn 09.8392.4005
linkkiVanda stad :
Barnskyddsanmälanfinska _ engelska
på InfoFinlands sida Problematiska situationer i Vanda hittar du information om var någonstans i Vanda det finns hjälp att få till barns och ungas problem .
information om barns och ungas problem finns även på InfoFinlands sidor Barns och ungas problem och Barnskydd .
på InfoFinlands sida Problem i äktenskap och parförhållande finns information om var man kan få hjälp med problem i parförhållanden .
äldre människor
i Vanda finns tjänster som är särskilt avsedda för äldre .
du får information om dem vid seniorrådgivningen .
seniorrådgivningen Tfn : 09.8392.4202
när du tar hand om en anhörig i hemmet
när en familjemedlem behöver kontinuerlig hjälp och vården är både bindande och krävande , finns det möjlighet att få stöd för närståendevård av kommunen .
seniorrådgivningen bedömer behovet av anhörigvård för en äldre person .
Läs mer : äldre människor .
linkkiVanda stad :
Seniorrådgivningenfinska _ svenska _ engelska
hälsotjänster i Vanda
privata hälsotjänster
barns hälsa
äldre människors hälsa
tandvård
mental hälsa
sexuell hälsa
när du väntar barn
handikappade
hälsotjänsterna i Vanda
om du behöver information om hälsotjänsterna , kan du ringa hälsorådgivningstelefonen : tfn ( 09 ) 839.10023 , mån @-@ fre kl . 8 @-@ 16 .
via tjänsten kan du också fråga om anvisningar för vård av sjukdomar .
du kan tala finska , svenska eller engelska .
Läs mer : hälsa .
linkkiVanda stad :
information om hälsorådgivningfinska _ svenska _ engelska
offentliga hälsovårdstjänster
om du har din hemkommun i Vanda , kan du utnyttja de offentliga hälsovårdstjänsterna .
offentliga hälsovårdstjänster tillhandahålls till exempel vid hälsostationer , tandkliniker , rådgivningsbyråer och sjukhus .
om du insjuknar plötsligt eller om du råkar ut för en olycka , får du akut sjukvård även om din hemkommun inte är Vanda .
i Vanda finns sju hälsostationer ( terveysasema ) som tillhandahåller offentliga hälsovårdstjänster .
hälsostationerna har öppet vardagar kl . 8.00 @-@ 16.00 .
hälsostationerna når du genom att ringa till respektive hälsostations eget telefonnummer eller hälsorådgivningens telefonnummer ( 09 ) 839.10023 och väljer din hälsostation med hjälpa av knappsatsen .
om du behöver akut vård samma dag , ska du ringa hälsostationen direkt då den öppnar .
hälsostationernas adresser :
Håkansböle hälsostation , Galoppbrinken 4
Korso hälsostation , Fjällrävsstigen 6
Västerkulla hälsostation , Kägelgränden 1
Myrbacka hälsostation , Jönsasvägen 4
Dickursby hälsostation , Konvaljvägen 11
närmare information hittar du på hälsostationernas egna webbplatser .
linkkiVanda stad :
Hälsostationernafinska _ svenska _ engelska
privata hälsotjänster
i Vanda finns flera läkarstationer som erbjuder privata hälsovårdstjänster .
du kan gå till en privat läkarstation även om du inte har rätt att använda den offentliga hälsovårdens tjänster i Finland .
på en privat läkarstation måste du betala samtliga kostnader själv .
i vissa fall ersätter Kela en liten del av kostnaderna för privat sjukvård .
privat läkarstationfinska _ svenska _ engelska
privat läkarstationfinska _ svenska _ engelska _ ryska
privat läkarstationfinska _ svenska _ engelska
linkkiAava :
privat läkarstationfinska _ svenska _ engelska
läkemedel
information om köp av läkemedel hittar du på InfoFinlands sida Läkemedel .
linkkiApotekareförbundet :
Apotekens kontaktuppgifterfinska
hälsovård för papperslösa
i Helsingfors finns Global Clinic , där personer som vistas i Finland utan tillstånd kan få primärhälsovård .
tjänsterna vid Global Clinic är avgiftsfria för kunderna .
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter .
för att skydda kunderna uppges inte klinikens adress eller öppettider offentligt .
telefonnumret till Helsingfors Global Clinicin är 044.948.1698 .
en sjuksköterska eller läkare svarar i telefonen .
Läs mer : hälsovårdstjänster i Finland .
hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
på kvällar , helger och storhelger är hälsostationerna stängda .
då vårdas akuta sjukfall och olycksfall på jourmottagningen ( päivystys ) .
jourmottagningen är öppen alla dagar dygnet runt
i Vanda finns jourmottagningen på Pejas sjukhus ( Peijaksen sairaala ) .
adress :
Sjukhusgatan 1
tfn 116.117
om du blir akut sjuk , kan du även besöka någon annan jourmottagning i huvudstadsregionen .
mer information om jourmottagningarna hittar du på Vanda stads webbplats om hälsovårdstjänster .
i nödsituationer ringer du det allmänna nödnumret 112 .
Läs mer : hälsovårdstjänster i Finland .
linkkiVanda stad :
Jourmottagningarfinska _ svenska _ engelska
barns hälsa
i hälsovården av barn under skolåldern får man hjälp av rådgivningsbyråerna ( neuvola ) .
där kan du fråga om råd och få stöd i föräldraskapet och fostran av barn .
på rådgivningsbyrån följs barnets hälsa , tillväxt och utveckling upp och där ges även vaccinationerna .
kontaktuppgifterna till rådgivningsbyråerna hittar du på Vanda webbplats .
via rådgivningsbyråernas telefontjänst kan du boka tid på rådgivningsbyrån och fråga hälsovårdaren om råd beträffande graviditet och barns hälsa .
numret till telefontjänsten är ( 09 ) 8392.5900 .
den är öppen mån @-@ tors kl . 8 @-@ 15 och fre kl . 8 @-@ 13 .
Skolhälsovården har hand om skolbarns hälsa .
mer information hittar du på Vanda stads webbplats .
om ett barn blir akut sjukt , ska du ta kontakt med hälsostationen eller jourmottagningen .
i nödsituationer ringer du det allmänna nödnumret 112 .
Läs mer : barns hälsa .
linkkiVanda stad :
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad :
tidsbokning och rådgivningfinska _ svenska _ engelska
linkkiVanda stad :
information om skolhälsovårdenfinska _ svenska _ engelska
linkkiVanda stad :
Hälsostationernafinska _ svenska _ engelska
linkkiVanda stad :
Jourmottagningarfinska _ svenska _ engelska
äldre människors hälsa
äldre människor använder samma hälsovårdstjänster som alla andra .
dessutom finns det i Vanda särskilda tjänster för äldre som du får information om via seniorrådgivningen ( seniorineuvonta ) .
tfn : ( 09 ) 8392.4202
mer information om tjänsterna för äldre hittar du på Vanda stads webbplats .
Läs mer : äldre människors hälsa och Äldre människor .
linkkiVanda stad :
Seniorrådgivningenfinska _ svenska _ engelska
linkkiVanda stad :
information om tjänster för äldrefinska _ svenska _ engelska
linkkiVanda stad :
Serviceguide för seniorer ( pdf , 1 MB ) finska
när du tar hand om en anhörig i hemmet
när en familjemedlem behöver kontinuerlig hjälp och vården är både bindande och krävande , finns det möjlighet att få stöd för närståendevård av kommunen .
behovet av närståendevård bedöms inom seniorrådgivningen .
tfn : ( 09 ) 8392.4202
behovet av närståendevård för personer under 65 år bedöms inom handikapprådgivningen .
tfn : ( 09 ) 8392.4682
linkkiVanda stad :
stöd för närståendevårdfinska _ svenska
tandvård
offentlig tandvård
Tidsbokningsnumret till Vanda tandvård ( hammashoito ) är ( 09 ) 8393.5300 .
tidsbokningen kan du ringa :
mån @-@ tors 7.30 @-@ 15
Fredagar och storhelgsaftnar 7.30 @-@ 14 .
om ditt ärende inte är brådskande , ring efter kl . 10.00 .
om tjänsten är hårt belastad , kan du lämna ett meddelande om att bli uppringd vid ett senare tillfälle .
om du behöver akut tandvård på en vardag , ska du ringa tidsbokningen så fort den öppnar .
linkkiVanda stad :
information om tandvårdenfinska _ svenska _ engelska
linkkiVanda stad :
Tandklinikerfinska _ svenska
Tandvårdens jourmottagning
under kvällar och veckoslut finns tandvårdsjouren ( hammashoidon päivystys ) vid Haartmanska sjukhuset i Helsingfors .
tfn ( 09 ) 310.49999 .
Tandvårdens nattjour ( hammashoidon yöpäivystys ) finns på Tölö sjukhus olycksfallsstation .
Tölö sjukhus olycksfallsstation , Oral och käkkirurgisk jourmottagning
tfn 040.621.5699
Tandvårdens jourmottagning kvällar och veckoslutfinska _ svenska _ engelska
barns tandvård
om tandvården för barn under skolåldern får du information på barnrådgivningen ( lastenneuvola ) och vid tandklinikerna ( hammashoitola ) .
barn under 17 år kallas till tandkliniken för undersökning med cirka två års mellanrum .
linkkiVanda stad :
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad :
information om tandvården för skolbarnfinska
privata tandvårdstjänster
i Vanda finns också privata tandläkare .
om du inte har rätt att använda de offentliga hälsovårdstjänsterna , kan du söka dig till en privat tandläkare .
hos en privat tandläkare måste du betala samtliga kostnader själv .
i vissa fall ersätter Kela en liten del av kostnaderna för privat tandvård .
Läs mer : tandvård .
Sök tandläkarefinska
mental hälsa
om du behöver psykisk hjälp eller stöd , ska du kontakta din hälsostation ( terveysasema ) .
på hälsostationen behandlas de vanligaste psykiska problemen .
från hälsostationen kan du remitteras vidare exempelvis till depressionsskötare .
om hälsostationen inte har öppet och situationen är akut , ska du kontakta samjouren vid Pejas sjukhus ( Peijaksen sairaalan yhteispäivystys ) .
Sjukhusgatan 1
tfn ( 09 ) 4716.7060
om du behöver omedelbar krishjälp , kan du också ta kontakt med social- och krisjouren .
den har öppet dygnet runt .
social- och krisjouren
tfn ( 09 ) 8392.4005
Läs mer : mental hälsa .
linkkiVanda stad :
information om mentalvårdstjänsternafinska _ svenska _ engelska
linkkiVanda stad :
Hälsostationernafinska _ svenska _ engelska
linkkiVanda stad :
Jourmottagningarfinska _ svenska _ engelska
linkkiVanda stad :
social- och krisjourenfinska _ svenska _ engelska
sexuell hälsa
om du vill har information om graviditetsprevention , abort , sexuell hälsa och könssjukdomar , kan du kontakta preventivmedels- och familjeplaneringsrådgivningen ( ehkäisy- ja perhesuunnitteluneuvola ) .
preventivmedels- och familjeplaneringsrådgivningarna betjänar kvinnor och män i alla åldrar .
du måste beställa tid vid rådgivningarna .
Besöken är avgiftsfria för kunderna .
information om kontaktuppgifter finns på Vanda stads webbplats .
boka en tid hos preventivmedelsrådgivningens läkare eller hälsovårdare om du behöver preventivmedel ( raskauden ehkäisy ) eller om du överväger abort ( abortti ) .
boka en tid hos hälsostationens allmänläkare om du till exempel har problem med blödningar eller smärtor i underlivet .
vid hälsostationerna vårdas även könssjukdomar ( sukupuolitauti ) .
Vandabor kan även besöka polikliniken för könssjukdomar i Helsingfors .
linkkiVanda stad :
rådgivningarna för familjeplaneringfinska _ svenska .
linkkiVanda stad :
Hälsostationernafinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS :
polikliniken för könssjukdomarfinska _ svenska _ engelska
när du väntar barn
vid mödrarådgivningen ( äitiysneuvola ) följs moderns , fostrets och hela familjens hälsotillstånd under graviditeten .
kontakta rådgivningsbyrån ( neuvola ) när du upptäcker att du är gravid .
Rådgivningarnas telefontjänst
mån @-@ tors kl . 8 @-@ 15 och fre kl . 8 @-@ 13
via rådgivningsbyråernas telefontjänst kan du boka tid på rådgivningsbyrån och fråga hälsovårdaren om råd beträffande graviditet och förlossning .
mer information om graviditet och förlossning hittar du på Vanda stads mödra- och barnrådgivning på Internet ( Nettineuvola ) .
Läs mer : när du väntar barn .
linkkiVanda stad :
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad :
rådgivningarna för familjeplaneringfinska _ svenska
linkkiVanda stad :
Förlossningen
Läs mer : förlossning .
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS :
Förlossningfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt :
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
handikappade
du kan få tjänster för handikappade ( vammaispalvelut ) om du eller en närstående till dig har en invaliditet eller en sjukdom som orsakar långvariga , betydande svårigheter att klara sig hemma och i livet utanför hemmet .
tjänster för handikappade är till exempel personlig assistans , serviceboende , färdtjänst och ombyggnadsarbeten i bostaden .
ta kontakt med handikapprådgivningen som utreder ditt behov av stöd , handledning och tjänster utifrån din situation .
Mån.-fre. kl . 9 @-@ 15
tfn : ( 09 ) 8392.4682
Läs mer : handikappade personer .
linkkiVanda stad :
information om handikapptjänsternafinska _ svenska _ engelska
hälsotjänster i Vanda
barns hälsa
tandvård
mental hälsa
sexuell hälsa och prevention
graviditet och förlossning
handikappade
hälsotjänsterna i Vanda
det allmänna nödnumret är 112 .
ring nödnumret endast om det handlar om ett nödfall , till exempel en akut sjukdomsattack .
om din hemkommun är Vanda kan du använda kommunens offentliga hälsovårdstjänster .
offentliga hälsovårdstjänster tillhandahålls till exempel vid hälsostationer , tandkliniker , rådgivningsbyråer och sjukhus .
om du insjuknar akut eller råkar ut för en olycka får du akut sjukvård även om din hemkommun inte är Vanda .
om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna , kan du boka tid på en privat läkarstation .
Läs mer : hälsovårdstjänster i Finland .
offentliga hälsovårdstjänster
telefonnumret till den gemensamma telefontjänsten för hälsostationerna i Vanda är 09.839.50.000 .
du kan ringa detta nummer om du behöver rådgivning i behandlingen av en sjukdom eller vill boka eller avboka en läkartid .
tjänsten har öppet måndag till fredag kl . 8 @-@ 16 .
i Vanda finns sju hälsostationer som tillhandahåller offentliga hälsovårdstjänster .
på hälsostationerna finns läkarens , sjukskötarens och hälsovårdarens mottagningar .
om du insjuknar akut kan du gå direkt till vilken som helst hälsostation .
det är bäst att gå till hälsostationen direkt på morgonen .
hälsostationerna har öppet vardagar kl . 8.00 @-@ 16.00 .
linkkiVanda stad :
information om hälsorådgivningfinska _ svenska _ engelska
linkkiVanda stad :
Hälsostationernafinska _ svenska _ engelska
privata hälsotjänster
i Vanda finns flera läkarstationer som erbjuder privata hälsovårdstjänster .
du kan gå till en privat läkarstation även om du inte har rätt att använda den offentliga hälsovårdens tjänster i Finland .
på en privat läkarstation måste du betala samtliga kostnader själv .
i vissa fall ersätter Kela en liten del av kostnaderna för privat sjukvård .
Läs mer : hälsovårdstjänster i Finland .
privat läkarstationfinska _ svenska _ engelska
privat läkarstationfinska _ svenska _ engelska _ ryska
privat läkarstationfinska _ svenska _ engelska
linkkiAava :
privat läkarstationfinska _ svenska _ engelska
läkemedel
information om köp av läkemedel hittar du på InfoFinlands sida Läkemedel .
linkkiApotekareförbundet :
Apotekens kontaktuppgifterfinska
hälsovård för papperslösa
i Helsingfors finns Global Clinic , där personer som vistas i Finland utan tillstånd kan få primärhälsovård .
tjänsterna vid Global Clinic är avgiftsfria för kunderna .
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter .
för att skydda kunderna uppges inte klinikens adress eller öppettider offentligt .
telefonnumret till Helsingfors Global Clinicin är 044.948.1698 .
en sjuksköterska eller läkare svarar i telefonen .
hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
på kvällar , helger och storhelger är hälsostationerna stängda .
om du insjuknar akut eller råkar ut för en olycka och inte kan vänta tills hälsostationen öppnar , kontakta jourmottagningen .
i Vanda finns jourmottagningen på Pejas sjukhus ( Peijaksen sairaala ) .
adress :
Sjukhusgatan 1
tfn 116.117
om du blir akut sjuk , kan du även besöka någon annan jourmottagning i huvudstadsregionen .
mer information om jourmottagningarna hittar du på Vanda stads webbplats om hälsovårdstjänster .
linkkiVanda stad :
Jourmottagningarfinska _ svenska _ engelska
barns hälsa
i hälsovården av barn under skolåldern får man hjälp av rådgivningsbyråerna ( neuvola ) .
telefonnumret till rådgivningsbyråerna i Vanda är 09.8392.5900 .
du kan boka en tid på rådgivningen eller fråga om råd om du har frågor kring barnets hälsa .
Skolhälsovården har hand om skolbarns hälsa .
mer information hittar du på Vanda stads webbplats .
om ett barn insjuknar akut , ska du kontakta hälsostationen .
hälsostationerna har öppet måndag till fredag kl . 8 @-@ 16 .
när hälsostationen har stängt ska du kontakta jourmottagningen vid Barnsjukhuset .
jourmottagningen tar endast hand om barn med brådskande hjälpbehov .
telefonnumret till jourmottagningen är 116.117 .
adress :
Barnsjukhuset
Stenbäcksgatan 9
du kan även ta barnet till en privat läkarstation .
i Vanda finns många privata läkarstationer som även tar hand om barn .
Läs mer : barns hälsa .
linkkiVanda stad :
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad :
tidsbokning och rådgivningfinska _ svenska _ engelska
linkkiVanda stad :
information om skolhälsovårdenfinska _ svenska _ engelska
linkkiVanda stad :
Hälsostationernafinska _ svenska _ engelska
linkkiVanda stad :
Jourmottagningarfinska _ svenska _ engelska
tandvård
offentlig tandvård
Tidsbokningsnumret till Vanda tandvård ( hammashoito ) är ( 09 ) 8393.5300 .
om du inte behöver brådskande tandvård , ring efter kl . 10.00 .
om du behöver brådskande tandvård , ska du ringa tidsbokningen så fort den öppnar kl . 7.30 .
mottagningen för brådskande vård finns vid Dickursby hälsostation måndag till fredag kl . 8 @-@ 14 .
linkkiVanda stad :
information om tandvårdenfinska _ svenska _ engelska
linkkiVanda stad :
Tandklinikerfinska _ svenska
Tandvårdens jourmottagning
under kvällar och veckoslut finns tandvårdsjouren ( hammashoidon päivystys ) vid Haartmanska sjukhuset i Helsingfors .
telefonnumret är 09.471.71110 .
tidsbokningen har öppet vardagar kl . 14 @-@ 21 och på veckoslut kl . 8 @-@ 21 .
Tandvårdens nattjour ( hammashoidon yöpäivystys ) finns på Tölö sjukhus olycksfallsstation .
Tölö sjukhus olycksfallsstation , Oral och käkkirurgisk jourmottagning
tfn 040.621.5699
Tandvårdens jourmottagning kvällar och veckoslutfinska _ svenska _ engelska
barns tandvård
om tandvården för barn under skolåldern får du information på barnrådgivningen ( lastenneuvola ) och vid tandklinikerna ( hammashoitola ) .
barn under 17 år kallas till tandkliniken för undersökning med cirka två års mellanrum .
linkkiVanda stad :
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad :
information om tandvården för skolbarnfinska
privata tandvårdstjänster
i Vanda finns också privata tandläkare .
om du inte har rätt att använda de offentliga hälsovårdstjänsterna , kan du söka dig till en privat tandläkare .
hos en privat tandläkare måste du betala samtliga kostnader själv .
i vissa fall ersätter Kela en liten del av kostnaderna för privat tandvård .
Läs mer : tandvård .
Sök tandläkarefinska
mental hälsa
om du behöver psykisk hjälp eller stöd , ska du kontakta din hälsostation ( terveysasema ) .
på hälsostationen behandlas de vanligaste psykiska problemen .
från hälsostationen kan du remitteras vidare exempelvis till depressionsskötare .
om hälsostationen inte har öppet och situationen är akut , ska du kontakta samjouren vid Pejas sjukhus ( Peijaksen sairaalan yhteispäivystys ) .
Sjukhusgatan 1
tfn 116.117
om du behöver omedelbar krishjälp , kan du också ta kontakt med social- och krisjouren .
den har öppet dygnet runt .
social- och krisjouren
tfn ( 09 ) 8392.4005
Läs mer : mental hälsa .
linkkiVanda stad :
information om mentalvårdstjänsternafinska _ svenska _ engelska
linkkiVanda stad :
Hälsostationernafinska _ svenska _ engelska
linkkiVanda stad :
Jourmottagningarfinska _ svenska _ engelska
linkkiVanda stad :
social- och krisjourenfinska _ svenska _ engelska
sexuell hälsa och prevention
om du behöver preventivmedel eller abort eller misstänker att du har en könssjukdom , kan du kontakta preventivmedels- och familjeplaneringsrådgivningen .
du kan boka tid per telefon .
numret är 09.839.50030 .
om du har en könssjukdom kan du även besöka polikliniken för könssjukdomar i Helsingfors eller en hälsostation .
Vanda erbjuder ungdomar under 20 år gratis preventivmedel .
även unga vuxna under 24 år kan få gratis preventivmedel om de använder långvariga preventivmedel såsom spiral eller p @-@ stav .
Läs mer : sexuell hälsa och prevention .
linkkiVanda stad :
rådgivningarna för familjeplaneringfinska _ svenska .
linkkiVanda stad :
Hälsostationernafinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS :
polikliniken för könssjukdomarfinska _ svenska _ engelska
graviditet och förlossning
vid mödrarådgivningen ( äitiysneuvola ) följs moderns , fostrets och hela familjens hälsotillstånd under graviditeten .
kontakta rådgivningsbyrån ( neuvola ) när du upptäcker att du är gravid .
Rådgivningarnas telefontjänst
via rådgivningsbyråernas telefontjänst kan du boka tid på rådgivningsbyrån och fråga hälsovårdaren om råd beträffande graviditet och förlossning .
Läs mer : graviditet och förlossning och När ett barn föds i Finland .
linkkiVanda stad :
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad :
rådgivningarna för familjeplaneringfinska _ svenska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS :
Förlossningfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt :
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
handikappade
du kan få tjänster för handikappade ( vammaispalvelut ) om du eller en närstående till dig har en invaliditet eller en sjukdom som orsakar långvariga , betydande svårigheter att klara sig hemma och i livet utanför hemmet .
tjänster för handikappade är till exempel personlig assistans , serviceboende , färdtjänst och ombyggnadsarbeten i bostaden .
ta kontakt med handikapprådgivningen som utreder ditt behov av stöd , handledning och tjänster utifrån din situation .
Mån.-fre. kl . 9 @-@ 15
tfn : ( 09 ) 8392.4682
Läs mer : handikappade personer .
linkkiVanda stad :
information om handikapptjänsternafinska _ svenska _ engelska
hälsotjänster i Vanda
barns hälsa
tandvård
mental hälsa
sexuell hälsa och prevention
graviditet och förlossning
handikappade
hälsotjänsterna i Vanda
det allmänna nödnumret är 112 .
ring nödnumret endast om det handlar om ett nödfall , till exempel en akut sjukdomsattack .
om din hemkommun är Vanda kan du använda kommunens offentliga hälsovårdstjänster .
offentliga hälsovårdstjänster tillhandahålls till exempel vid hälsostationer , tandkliniker , rådgivningsbyråer och sjukhus .
om du insjuknar akut eller råkar ut för en olycka får du akut sjukvård även om din hemkommun inte är Vanda .
om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna , kan du boka tid på en privat läkarstation .
Läs mer : hälsovårdstjänster i Finland .
offentliga hälsovårdstjänster
telefonnumret till den gemensamma telefontjänsten för hälsostationerna i Vanda är 09.839.50.000 .
du kan ringa detta nummer om du behöver rådgivning i behandlingen av en sjukdom eller vill boka eller avboka en läkartid .
tjänsten har öppet måndag till fredag kl . 8 @-@ 16 .
i Vanda finns sju hälsostationer som tillhandahåller offentliga hälsovårdstjänster .
på hälsostationerna finns läkarens , sjukskötarens och hälsovårdarens mottagningar .
om du insjuknar akut kan du gå direkt till vilken som helst hälsostation .
det är bäst att gå till hälsostationen direkt på morgonen .
hälsostationerna har öppet vardagar kl . 8.00 @-@ 16.00 .
linkkiVanda stad :
information om hälsorådgivningfinska _ svenska _ engelska
linkkiVanda stad :
Hälsostationernafinska _ svenska _ engelska
privata hälsotjänster
i Vanda finns flera läkarstationer som erbjuder privata hälsovårdstjänster .
du kan gå till en privat läkarstation även om du inte har rätt att använda den offentliga hälsovårdens tjänster i Finland .
på en privat läkarstation måste du betala samtliga kostnader själv .
i vissa fall ersätter Kela en liten del av kostnaderna för privat sjukvård .
Läs mer : hälsovårdstjänster i Finland .
privat läkarstationfinska _ svenska _ engelska
privat läkarstationfinska _ svenska _ engelska _ ryska
privat läkarstationfinska _ svenska _ engelska
linkkiAava :
privat läkarstationfinska _ svenska _ engelska
läkemedel
information om köp av läkemedel hittar du på InfoFinlands sida Läkemedel .
linkkiApotekareförbundet :
Apotekens kontaktuppgifterfinska
hälsovård för papperslösa
i Helsingfors finns Global Clinic , där personer som vistas i Finland utan tillstånd kan få primärhälsovård .
tjänsterna vid Global Clinic är avgiftsfria för kunderna .
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter .
för att skydda kunderna uppges inte klinikens adress eller öppettider offentligt .
telefonnumret till Helsingfors Global Clinicin är 044.948.1698 .
en sjuksköterska eller läkare svarar i telefonen .
hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
på kvällar , helger och storhelger är hälsostationerna stängda .
om du insjuknar akut eller råkar ut för en olycka och inte kan vänta tills hälsostationen öppnar , kontakta jourmottagningen .
i Vanda finns jourmottagningen på Pejas sjukhus ( Peijaksen sairaala ) .
adress :
Sjukhusgatan 1
tfn 116.117
om du blir akut sjuk , kan du även besöka någon annan jourmottagning i huvudstadsregionen .
mer information om jourmottagningarna hittar du på Vanda stads webbplats om hälsovårdstjänster .
linkkiVanda stad :
Jourmottagningarfinska _ svenska _ engelska
barns hälsa
i hälsovården av barn under skolåldern får man hjälp av rådgivningsbyråerna ( neuvola ) .
telefonnumret till rådgivningsbyråerna i Vanda är 09.8392.5900 .
du kan boka en tid på rådgivningen eller fråga om råd om du har frågor kring barnets hälsa .
Skolhälsovården har hand om skolbarns hälsa .
mer information hittar du på Vanda stads webbplats .
om ett barn insjuknar akut , ska du kontakta hälsostationen .
hälsostationerna har öppet måndag till fredag kl . 8 @-@ 16 .
när hälsostationen har stängt ska du kontakta jourmottagningen vid Barnsjukhuset .
jourmottagningen tar endast hand om barn med brådskande hjälpbehov .
telefonnumret till jourmottagningen är 116.117 .
adress :
Barnsjukhuset
Stenbäcksgatan 9
du kan även ta barnet till en privat läkarstation .
i Vanda finns många privata läkarstationer som även tar hand om barn .
Läs mer : barns hälsa .
linkkiVanda stad :
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad :
tidsbokning och rådgivningfinska _ svenska _ engelska
linkkiVanda stad :
information om skolhälsovårdenfinska _ svenska _ engelska
linkkiVanda stad :
Hälsostationernafinska _ svenska _ engelska
linkkiVanda stad :
Jourmottagningarfinska _ svenska _ engelska
tandvård
offentlig tandvård
Tidsbokningsnumret till Vanda tandvård ( hammashoito ) är ( 09 ) 8393.5300 .
om du inte behöver brådskande tandvård , ring efter kl . 10.00 .
om du behöver brådskande tandvård , ska du ringa tidsbokningen så fort den öppnar kl . 7.30 .
mottagningen för brådskande vård finns vid Dickursby hälsostation måndag till fredag kl . 8 @-@ 14 .
linkkiVanda stad :
information om tandvårdenfinska _ svenska _ engelska
linkkiVanda stad :
Tandklinikerfinska _ svenska
Tandvårdens jourmottagning
under kvällar och veckoslut finns tandvårdsjouren ( hammashoidon päivystys ) vid Haartmanska sjukhuset i Helsingfors .
telefonnumret är 09.471.71110 .
tidsbokningen har öppet vardagar kl . 14 @-@ 21 och på veckoslut kl . 8 @-@ 21 .
Tandvårdens nattjour ( hammashoidon yöpäivystys ) finns på Tölö sjukhus olycksfallsstation .
Tölö sjukhus olycksfallsstation , Oral och käkkirurgisk jourmottagning
tfn 040.621.5699
Tandvårdens jourmottagning kvällar och veckoslutfinska _ svenska _ engelska
barns tandvård
om tandvården för barn under skolåldern får du information på barnrådgivningen ( lastenneuvola ) och vid tandklinikerna ( hammashoitola ) .
barn under 17 år kallas till tandkliniken för undersökning med cirka två års mellanrum .
linkkiVanda stad :
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad :
information om tandvården för skolbarnfinska
privata tandvårdstjänster
i Vanda finns också privata tandläkare .
om du inte har rätt att använda de offentliga hälsovårdstjänsterna , kan du söka dig till en privat tandläkare .
hos en privat tandläkare måste du betala samtliga kostnader själv .
i vissa fall ersätter Kela en liten del av kostnaderna för privat tandvård .
Läs mer : tandvård .
Sök tandläkarefinska
mental hälsa
om du behöver psykisk hjälp eller stöd , ska du kontakta din hälsostation ( terveysasema ) .
på hälsostationen behandlas de vanligaste psykiska problemen .
från hälsostationen kan du remitteras vidare exempelvis till depressionsskötare .
om hälsostationen inte har öppet och situationen är akut , ska du kontakta samjouren vid Pejas sjukhus ( Peijaksen sairaalan yhteispäivystys ) .
Sjukhusgatan 1
tfn 116.117
om du behöver omedelbar krishjälp , kan du också ta kontakt med social- och krisjouren .
den har öppet dygnet runt .
social- och krisjouren
tfn ( 09 ) 8392.4005
Läs mer : mental hälsa .
linkkiVanda stad :
information om mentalvårdstjänsternafinska _ svenska _ engelska
linkkiVanda stad :
Hälsostationernafinska _ svenska _ engelska
linkkiVanda stad :
Jourmottagningarfinska _ svenska _ engelska
linkkiVanda stad :
social- och krisjourenfinska _ svenska _ engelska
sexuell hälsa och prevention
om du behöver preventivmedel eller abort eller misstänker att du har en könssjukdom , kan du kontakta preventivmedels- och familjeplaneringsrådgivningen .
du kan boka tid per telefon .
numret är 09.839.50030 .
om du har en könssjukdom kan du även besöka polikliniken för könssjukdomar i Helsingfors eller en hälsostation .
Vanda erbjuder ungdomar under 20 år gratis preventivmedel .
även unga vuxna under 24 år kan få gratis preventivmedel om de använder långvariga preventivmedel såsom spiral eller p @-@ stav .
Läs mer : sexuell hälsa och prevention .
linkkiVanda stad :
rådgivningarna för familjeplaneringfinska _ svenska .
linkkiVanda stad :
Hälsostationernafinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS :
polikliniken för könssjukdomarfinska _ svenska _ engelska
graviditet och förlossning
vid mödrarådgivningen ( äitiysneuvola ) följs moderns , fostrets och hela familjens hälsotillstånd under graviditeten .
kontakta rådgivningsbyrån ( neuvola ) när du upptäcker att du är gravid .
Rådgivningarnas telefontjänst
via rådgivningsbyråernas telefontjänst kan du boka tid på rådgivningsbyrån och fråga hälsovårdaren om råd beträffande graviditet och förlossning .
Läs mer : graviditet och förlossning och När ett barn föds i Finland .
linkkiVanda stad :
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad :
rådgivningarna för familjeplaneringfinska _ svenska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS :
Förlossningfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt :
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
handikappade
du kan få tjänster för handikappade ( vammaispalvelut ) om du eller en närstående till dig har en invaliditet eller en sjukdom som orsakar långvariga , betydande svårigheter att klara sig hemma och i livet utanför hemmet .
tjänster för handikappade är till exempel personlig assistans , serviceboende , färdtjänst och ombyggnadsarbeten i bostaden .
ta kontakt med handikapprådgivningen som utreder ditt behov av stöd , handledning och tjänster utifrån din situation .
Mån.-fre. kl . 9 @-@ 15
tfn : ( 09 ) 8392.4682
Läs mer : handikappade personer .
linkkiVanda stad :
information om handikapptjänsternafinska _ svenska _ engelska
dagvård
förskoleundervisning
grundläggande utbildning
yrkesutbildning
gymnasium
stöd och handledning för unga
Högskoleutbildning
övriga studiemöjligheter
dagvård
i Vanda finns både kommunala och privata daghem .
kommunen övervakar också den privata dagvården .
i Vanda ges dagvård på finska , svenska , ryska och engelska .
inom dagvården ges även undervisning i finska som andra språk .
dagvård ordnas också inom familjedagvården och i gruppfamiljedaghem .
man ska ansöka om dagvårdsplats för sitt barn minst fyra månader innan barnet ska börja i dagvården .
du kan ansöka om plats i den kommunala dagvården via Internet eller med en pappersblankett .
för en elektronisk ansökan behöver du egna nätbankskoder eller en elektronisk legitimation .
Pappersblanketter kan hämtas till exempel vid Vandainfo eller daghemmen .
privata dagvårdsplatser söks direkt på daghemmet .
frågor kring dagvård och ansökan om dagvårdsplats kan du ställa till daghemsföreståndaren eller skicka till adressen varhaiskasvatus ( at ) vantaa.fi .
vanligtvis ansöker man om dagvårdsplats i den egna kommunen .
om familjen bor nära gränsen till Helsingfors eller Esbo , kan du också söka dagvårdsplats i grannkommunen .
du ska ändå lämna in din ansökan i den egna kommunen .
mer information hittar du via tjänsten Helsingforsregionen.fi .
Läs mer : dagvård
linkkiVanda stad :
privat dagvårdfinska _ svenska _ engelska
linkkiVanda stad :
privat dagvårdfinska
linkkiVanda stad :
ansökan om dagvårdsplatsfinska _ svenska _ engelska
linkkiVanda stad :
elektronisk ansökningsblankett för dagvårdenfinska _ svenska _ engelska
information om dagvården finska _ svenska _ engelska
förskoleundervisning
förskoleundervisning ( esiopetus ) ordnas i både kommunala och privata daghem samt i förskoleenheter i skolornas lokaler .
i Vanda kan man få förskoleundervisning på finska , svenska och engelska .
du måste ansöka om plats i förskoleundervisningen .
ansökan kan göras elektroniskt via stadens webbplats eller med en pappersblankett .
ansökningstiden är i januari , men ansökan kan även lämnas in övriga tider , om familjen till exempel flyttar till Vanda mitt under året .
förberedande undervisning tillhandahålls för invandrarbarn som inte har tillräckliga kunskaper i finska för att klara sig i förskoleundervisningen .
den förberedande undervisningen är avsedd för 6 @-@ åriga barn med invandrarbakgrund .
den ordnas i daghemmens förskolegrupper .
daghemmet anvisar barnet till den förberedande undervisningen i samband med ansökningen till förskoleundervisningen .
du hittar mer information om förskoleundervisningen , ansökning till förskoleundervisningen och om undervisning som förbereder för förskoleundervisning på Vanda stads ( Vantaan kaupunki ) webbplats .
du kan även fråga om mer information på daghemmen .
Läs mer : förskoleundervisning
linkkiVanda stad :
ansökan till förskoleundervisningfinska _ svenska _ engelska
linkkiVanda stad :
information om den förberedande undervisningenfinska _ engelska
linkkiVanda stad :
elektronisk ansökningsblankett för förskoleundervisningenfinska _ svenska _ engelska
linkkiVanda stad :
daghem som ger förskoleundervisningfinska _ engelska
grundläggande utbildning
i Vanda finns finskspråkiga och svenskspråkiga grundskolor ( peruskoulu ) .
i Vanda finns även en internationell skola , där man kan avlägga grundskolan på engelska .
mer information om skolorna i Vanda hittar du på Vanda stads ( Vantaan kaupunki ) webbplats .
anmälan till grundskolan ska göras på förhand .
Anmälningstiden är vanligtvis i januari .
på stadens webbplats hittar du kontaktuppgifterna till skolorna och mer information om anmälan .
Läs mer : grundläggande utbildning
linkkiVanda stad :
anmälan till skolanfinska _ svenska _ engelska
linkkiVanda stad :
skolornas kontaktuppgifterfinska
Eftermiddagsverksamhetfinska _ svenska
förberedande utbildning inför grundskola
om barnets kunskaper i det finska språket inte är tillräckligt bra för studier i den finskspråkiga grundskolan , kan barnet få förberedande utbildning ( valmistava opetus ) .
i den förberedande utbildningen läser barnen det finska språket och grundskolans läroämnen .
undervisningen pågår vanligtvis i ett år .
om du har anlänt till Finland för en kort tid sedan och har barn under skolåldern ska du ta kontakt med områdeskoordinatorn för ditt bostadsområde ( aluekoordinaattori ) .
områdeskoordinatorn berättar om hur undervisningen ordnas och hjälper dig i frågor som rör barnets skolgång .
information om den förberedande undervisningenfinska
linkkiVanda stad :
Områdeskoordinatorerfinska
grundläggande utbildning för unga invandrare
vid Vanda vuxenutbildningsinstitut ( Vantaan aikuisopisto ) kan 17 @-@ 24 @-@ åriga invandrarungdomar avlägga grundskolans avgångsbetyg .
om man har hoppat av grundskolan , kan man avlägga grundskolans lärokurs också vid Eira vuxengymnasium ( Eiran aikuislukio ) .
grundläggande utbildning för invandrarefinska
linkkiEira vuxengymnasium :
grundundervisning för vuxnafinska
tionde klasserna
du kan ansöka till den grundläggande utbildningens tilläggsundervisning , det vill säga till en tionde klass ( kymppiluokka ) , om du fick grundskolans avgångsbetyg samma år eller året innan , men inte har fått en studieplats på andra stadiet .
på tionde klassen kan du höja dina betyg från grundskolan och du får en plan för fortsatta studier .
Tiondeklasserna i Vanda finns i östra och västra Vanda vid Varias verksamhetsställen och vid Lumo gymnasium ( Lumon lukio ) .
linkkiVanda stad :
Tiondeklasserfinska _ svenska
invandrare och grundläggande utbildning
i skolorna i Vanda ges hemspråksundervisning i flera olika språk .
i grundskolorna ges även utbildning i finska som andraspråk ( suomi toisena kielenä ) till elever som har ett annat modersmål än finska , svenska eller samiska , och vars kunskaper i det finska språket inte är i nivå med modersmålet .
när du anmäler dig till skolan , kan du samtidigt anmäla dig till hemspråksundervisning och undervisning i din egen religion .
du kan även anmäla dig till undervisningen genom att fylla i en blankett , som du får från din egen skola .
den ifyllda blanketten returneras till den egna skolan .
undervisning i den egna religionen kan ordnas om gruppen består av minst tre elever .
mer information om hemspråksundervisning och om undervisning i elevens egen religion hittar du på stadens webbplats och hos områdeskoordinatorerna ( aluekoordinaattori ) .
linkkiVanda stad :
information om hemspråksundervisningfinska
linkkiVanda stad :
undervisning i den egna religionenfinska
finska som andra språk i den grundläggande undervisningenfinska
linkkiVanda stad :
Områdeskoordinatorerfinska
yrkesutbildning
i Vanda ordnas yrkesutbildning vid yrkesinstitutet Vantaan ammattiopisto Varia , handelsläroanstalten MERCURIA samt TTS Arbetseffektivitetsföreningen rf:s verksamhetsställe i Vanda .
i Varia ordnas även engelskspråkig undervisning samt finskspråkiga yrkesutbildningar särskilt avsedda för invandrare .
Edupoli ordnar yrkesutbildning för vuxna .
i Vanda finns även Finavia Avia College som ger utbildning för olika luftfartsyrken .
Läs mer : yrkesutbildning .
linkkiVanda stad :
yrkesutbildningfinska _ svenska
linkkiYrkesläroanstalten Varia i Vanda :
yrkesutbildningfinska _ engelska
yrkesutbildningfinska _ engelska
linkkiTTS Arbetseffektivitetsföreningen rf:s verksamhetsställe i Vanda :
yrkesutbildningfinska
utbildning som handleder för yrkesutbildning ( VALMA )
utbildning som handleder för grundläggande yrkesutbildning ( Ammatilliseen peruskoulutukseen valmentava koulutus ) d.v.s. VALMA är avsedd för dem som vill avlägga en grundläggande yrkesutbildning .
under VALMA @-@ utbildningen får du kunskap och färdigheter som hjälper dig i dina senare yrkesinriktade studier .
du kan även förbättra din språkkunskap . du kan också höja dina grundskolebetyg .
i Vanda ordnas VALMA @-@ utbildning av Varia .
Läs mer om VALMA @-@ utbildningen på InfoFinlands sida Utbildning som handleder för yrkesutbildning .
linkkiVanda stad :
information om VALMA @-@ utbildningarfinska
linkkiYrkesläroanstalten Varia i Vanda :
i Vanda kan du studera på gymnasiet ( lukio ) på finska , svenska eller engelska .
undervisning på engelska erbjuds på IB @-@ linjen vid gymnasieskolan Tikkurilan lukio .
i Vanda finns även ett vuxengymnasium .
Läs mer : gymnasium .
linkkiVanda stad :
information om gymnasieutbildningfinska _ svenska
linkkiVanda stad :
gymnasierna och gymnasiernas hemsidorfinska
linkkiVanda stad :
Vuxengymnasiumfinska
linkkiVanda stad :
Distansgymnasiumfinska
linkkiVanda stad :
Steinergymnasietfinska
förberedande gymnasieutbildning ( LUVA )
om du vill förbättra dina kunskaper i finska eller svenska innan du söker till ett gymnasium , kan du söka till en förberedande gymnasieutbildning .
den är avsedd för invandrare .
i Vanda ordnas LUVA @-@ utbildning av Lumon lukio .
Läs mer om LUVA @-@ utbildningen på InfoFinlands sida Förberedande gymnasieutbildning .
linkkiVanda stad :
förberedande gymnasieutbildningfinska
stöd och handledning för unga
om du är under 30 år gammal kan du få råd och handledning via Ohjaamo @-@ tjänsten .
Ohjaamos personal hjälper dig om du inte har ett arbete eller en studieplats .
du kan även fråga om andra saker , som till exempel boende eller ekonomiska frågor .
linkkiOhjaamo :
stöd och handledning för ungafinska _ engelska
Vägledningscentret Kipinä
om du är under 29 år gammal , bor i Vanda och inte har ett jobb eller en studieplats , kan du få råd och handledning i Kipinä .
ring och boka en tid i förväg .
utan tidsbokning kan du besöka Kipinä på tisdagar och onsdagar kl . 12.00 @-@ 18.00 .
mer information hittar du på webbplatsen .
Kipinä
Banvägen 2 , Dickursby
tfn 050.312.4372
vägledning och stöd för ungafinska _ svenska
Högskoleutbildning
i Vanda finns två yrkeshögskolor ( ammattikorkeakoulu ) , Laurea och Metropolia .
de erbjuder utbildning inom många olika branscher .
mer information om utbildningsprogram och om ansökan hittar du på läroanstalternas webbplats .
också Helsingfors universitets öppna universitet ( avoin yliopisto ) har verksamhetsställen i Vanda . där ges undervisning på högskolenivå och fortbildning .
Läs mer : Högskoleutbildning .
linkkiVanda stad :
Högskoleutbildningfinska
yrkeshögskolafinska _ engelska
linkkiMetropolia :
yrkeshögskolafinska _ engelska
Ubildning vid öppna universitetet i Vandafinska _ svenska _ engelska
övriga studiemöjligheter
vid Vanda vuxenutbildningsinstitut ( Vantaan aikuisopisto ) kan du studera till exempel språk , handarbete och matlagning eller delta i ledd motion .
kurserna är avgiftsbelagda och de ordnas både dag- och kvällstid .
Vuxenutbildningsinstitutet ordnar även kurser för invandrare .
mer information hittar du på Vanda stads webbplats .
Läs mer : andra studiemöjligheter .
linkkiVanda vuxenutbildningsinstitut :
Studiehandbokfinska
linkkiVanda vuxenutbildningsinstitut :
kurser i finska och svenska språket för invandrarefinska
linkkiEdupoli :
Vuxenutbildningscenterfinska
dagvård
förskoleundervisning
grundläggande utbildning
yrkesutbildning
gymnasium
stöd och handledning för unga
Högskoleutbildning
övriga studiemöjligheter
dagvård
i Vanda finns både kommunala och privata daghem .
kommunen övervakar också den privata dagvården .
i Vanda ges dagvård på finska , svenska , ryska och engelska .
inom dagvården ges även undervisning i finska som andra språk .
dagvård ordnas också inom familjedagvården och i gruppfamiljedaghem .
man ska ansöka om dagvårdsplats för sitt barn minst fyra månader innan barnet ska börja i dagvården .
du kan ansöka om plats i den kommunala dagvården via Internet eller med en pappersblankett .
för en elektronisk ansökan behöver du egna nätbankskoder eller en elektronisk legitimation .
Pappersblanketter kan hämtas till exempel vid Vandainfo eller daghemmen .
privata dagvårdsplatser söks direkt på daghemmet .
frågor kring dagvård och ansökan om dagvårdsplats kan du ställa till daghemsföreståndaren eller skicka till adressen varhaiskasvatus ( at ) vantaa.fi .
vanligtvis ansöker man om dagvårdsplats i den egna kommunen .
om familjen bor nära gränsen till Helsingfors eller Esbo , kan du också söka dagvårdsplats i grannkommunen .
du ska ändå lämna in din ansökan i den egna kommunen .
mer information hittar du via tjänsten Helsingforsregionen.fi .
Läs mer : dagvård
linkkiVanda stad :
privat dagvårdfinska _ svenska _ engelska
linkkiVanda stad :
privat dagvårdfinska
linkkiVanda stad :
ansökan om dagvårdsplatsfinska _ svenska _ engelska
linkkiVanda stad :
elektronisk ansökningsblankett för dagvårdenfinska _ svenska _ engelska
information om dagvården finska _ svenska _ engelska
förskoleundervisning
förskoleundervisning ( esiopetus ) ordnas i både kommunala och privata daghem samt i förskoleenheter i skolornas lokaler .
i Vanda kan man få förskoleundervisning på finska , svenska och engelska .
du måste ansöka om plats i förskoleundervisningen .
ansökan kan göras elektroniskt via stadens webbplats eller med en pappersblankett .
ansökningstiden är i januari , men ansökan kan även lämnas in övriga tider , om familjen till exempel flyttar till Vanda mitt under året .
förberedande undervisning tillhandahålls för invandrarbarn som inte har tillräckliga kunskaper i finska för att klara sig i förskoleundervisningen .
den förberedande undervisningen är avsedd för 6 @-@ åriga barn med invandrarbakgrund .
den ordnas i daghemmens förskolegrupper .
daghemmet anvisar barnet till den förberedande undervisningen i samband med ansökningen till förskoleundervisningen .
du hittar mer information om förskoleundervisningen , ansökning till förskoleundervisningen och om undervisning som förbereder för förskoleundervisning på Vanda stads ( Vantaan kaupunki ) webbplats .
du kan även fråga om mer information på daghemmen .
Läs mer : förskoleundervisning
linkkiVanda stad :
ansökan till förskoleundervisningfinska _ svenska _ engelska
linkkiVanda stad :
information om den förberedande undervisningenfinska _ engelska
linkkiVanda stad :
elektronisk ansökningsblankett för förskoleundervisningenfinska _ svenska _ engelska
linkkiVanda stad :
daghem som ger förskoleundervisningfinska _ engelska
grundläggande utbildning
i Vanda finns finskspråkiga och svenskspråkiga grundskolor ( peruskoulu ) .
i Vanda finns även en internationell skola , där man kan avlägga grundskolan på engelska .
mer information om skolorna i Vanda hittar du på Vanda stads ( Vantaan kaupunki ) webbplats .
anmälan till grundskolan ska göras på förhand .
Anmälningstiden är vanligtvis i januari .
på stadens webbplats hittar du kontaktuppgifterna till skolorna och mer information om anmälan .
Läs mer : grundläggande utbildning
linkkiVanda stad :
anmälan till skolanfinska _ svenska _ engelska
linkkiVanda stad :
skolornas kontaktuppgifterfinska
Eftermiddagsverksamhetfinska _ svenska
förberedande utbildning inför grundskola
om barnets kunskaper i det finska språket inte är tillräckligt bra för studier i den finskspråkiga grundskolan , kan barnet få förberedande utbildning ( valmistava opetus ) .
i den förberedande utbildningen läser barnen det finska språket och grundskolans läroämnen .
undervisningen pågår vanligtvis i ett år .
om du har anlänt till Finland för en kort tid sedan och har barn under skolåldern ska du ta kontakt med områdeskoordinatorn för ditt bostadsområde ( aluekoordinaattori ) .
områdeskoordinatorn berättar om hur undervisningen ordnas och hjälper dig i frågor som rör barnets skolgång .
information om den förberedande undervisningenfinska
linkkiVanda stad :
Områdeskoordinatorerfinska
grundläggande utbildning för unga invandrare
vid Vanda vuxenutbildningsinstitut ( Vantaan aikuisopisto ) kan 17 @-@ 24 @-@ åriga invandrarungdomar avlägga grundskolans avgångsbetyg .
om man har hoppat av grundskolan , kan man avlägga grundskolans lärokurs också vid Eira vuxengymnasium ( Eiran aikuislukio ) .
grundläggande utbildning för invandrarefinska
linkkiEira vuxengymnasium :
grundundervisning för vuxnafinska
tionde klasserna
du kan ansöka till den grundläggande utbildningens tilläggsundervisning , det vill säga till en tionde klass ( kymppiluokka ) , om du fick grundskolans avgångsbetyg samma år eller året innan , men inte har fått en studieplats på andra stadiet .
på tionde klassen kan du höja dina betyg från grundskolan och du får en plan för fortsatta studier .
Tiondeklasserna i Vanda finns i östra och västra Vanda vid Varias verksamhetsställen och vid Lumo gymnasium ( Lumon lukio ) .
linkkiVanda stad :
Tiondeklasserfinska _ svenska
invandrare och grundläggande utbildning
i skolorna i Vanda ges hemspråksundervisning i flera olika språk .
i grundskolorna ges även utbildning i finska som andraspråk ( suomi toisena kielenä ) till elever som har ett annat modersmål än finska , svenska eller samiska , och vars kunskaper i det finska språket inte är i nivå med modersmålet .
när du anmäler dig till skolan , kan du samtidigt anmäla dig till hemspråksundervisning och undervisning i din egen religion .
du kan även anmäla dig till undervisningen genom att fylla i en blankett , som du får från din egen skola .
den ifyllda blanketten returneras till den egna skolan .
undervisning i den egna religionen kan ordnas om gruppen består av minst tre elever .
mer information om hemspråksundervisning och om undervisning i elevens egen religion hittar du på stadens webbplats och hos områdeskoordinatorerna ( aluekoordinaattori ) .
linkkiVanda stad :
information om hemspråksundervisningfinska
linkkiVanda stad :
undervisning i den egna religionenfinska
finska som andra språk i den grundläggande undervisningenfinska
linkkiVanda stad :
Områdeskoordinatorerfinska
yrkesutbildning
i Vanda ordnas yrkesutbildning vid yrkesinstitutet Vantaan ammattiopisto Varia , handelsläroanstalten MERCURIA samt TTS Arbetseffektivitetsföreningen rf:s verksamhetsställe i Vanda .
i Varia ordnas även engelskspråkig undervisning samt finskspråkiga yrkesutbildningar särskilt avsedda för invandrare .
Edupoli ordnar yrkesutbildning för vuxna .
i Vanda finns även Finavia Avia College som ger utbildning för olika luftfartsyrken .
Läs mer : yrkesutbildning .
linkkiVanda stad :
yrkesutbildningfinska _ svenska
linkkiYrkesläroanstalten Varia i Vanda :
yrkesutbildningfinska _ engelska
yrkesutbildningfinska _ engelska
linkkiTTS Arbetseffektivitetsföreningen rf:s verksamhetsställe i Vanda :
yrkesutbildningfinska
utbildning som handleder för yrkesutbildning ( VALMA )
utbildning som handleder för grundläggande yrkesutbildning ( Ammatilliseen peruskoulutukseen valmentava koulutus ) d.v.s. VALMA är avsedd för dem som vill avlägga en grundläggande yrkesutbildning .
under VALMA @-@ utbildningen får du kunskap och färdigheter som hjälper dig i dina senare yrkesinriktade studier .
du kan även förbättra din språkkunskap . du kan också höja dina grundskolebetyg .
i Vanda ordnas VALMA @-@ utbildning av Varia .
Läs mer om VALMA @-@ utbildningen på InfoFinlands sida Utbildning som handleder för yrkesutbildning .
linkkiVanda stad :
information om VALMA @-@ utbildningarfinska
linkkiYrkesläroanstalten Varia i Vanda :
i Vanda kan du studera på gymnasiet ( lukio ) på finska , svenska eller engelska .
undervisning på engelska erbjuds på IB @-@ linjen vid gymnasieskolan Tikkurilan lukio .
i Vanda finns även ett vuxengymnasium .
Läs mer : gymnasium .
linkkiVanda stad :
information om gymnasieutbildningfinska _ svenska
linkkiVanda stad :
gymnasierna och gymnasiernas hemsidorfinska
linkkiVanda stad :
Vuxengymnasiumfinska
linkkiVanda stad :
Distansgymnasiumfinska
linkkiVanda stad :
Steinergymnasietfinska
förberedande gymnasieutbildning ( LUVA )
om du vill förbättra dina kunskaper i finska eller svenska innan du söker till ett gymnasium , kan du söka till en förberedande gymnasieutbildning .
den är avsedd för invandrare .
i Vanda ordnas LUVA @-@ utbildning av Lumon lukio .
Läs mer om LUVA @-@ utbildningen på InfoFinlands sida Förberedande gymnasieutbildning .
linkkiVanda stad :
förberedande gymnasieutbildningfinska
stöd och handledning för unga
om du är under 30 år gammal kan du få råd och handledning via Ohjaamo @-@ tjänsten .
Ohjaamos personal hjälper dig om du inte har ett arbete eller en studieplats .
du kan även fråga om andra saker , som till exempel boende eller ekonomiska frågor .
linkkiOhjaamo :
stöd och handledning för ungafinska _ engelska
Vägledningscentret Kipinä
om du är under 29 år gammal , bor i Vanda och inte har ett jobb eller en studieplats , kan du få råd och handledning i Kipinä .
ring och boka en tid i förväg .
utan tidsbokning kan du besöka Kipinä på tisdagar och onsdagar kl . 12.00 @-@ 18.00 .
mer information hittar du på webbplatsen .
Kipinä
Banvägen 2 , Dickursby
tfn 050.312.4372
vägledning och stöd för ungafinska _ svenska
Högskoleutbildning
i Vanda finns två yrkeshögskolor ( ammattikorkeakoulu ) , Laurea och Metropolia .
de erbjuder utbildning inom många olika branscher .
mer information om utbildningsprogram och om ansökan hittar du på läroanstalternas webbplats .
också Helsingfors universitets öppna universitet ( avoin yliopisto ) har verksamhetsställen i Vanda . där ges undervisning på högskolenivå och fortbildning .
Läs mer : Högskoleutbildning .
linkkiVanda stad :
Högskoleutbildningfinska
yrkeshögskolafinska _ engelska
linkkiMetropolia :
yrkeshögskolafinska _ engelska
Ubildning vid öppna universitetet i Vandafinska _ svenska _ engelska
övriga studiemöjligheter
vid Vanda vuxenutbildningsinstitut ( Vantaan aikuisopisto ) kan du studera till exempel språk , handarbete och matlagning eller delta i ledd motion .
kurserna är avgiftsbelagda och de ordnas både dag- och kvällstid .
Vuxenutbildningsinstitutet ordnar även kurser för invandrare .
mer information hittar du på Vanda stads webbplats .
Läs mer : andra studiemöjligheter .
linkkiVanda vuxenutbildningsinstitut :
Studiehandbokfinska
linkkiVanda vuxenutbildningsinstitut :
kurser i finska och svenska språket för invandrarefinska
linkkiEdupoli :
Vuxenutbildningscenterfinska
dagvård
förskoleundervisning
grundläggande utbildning
yrkesutbildning
gymnasium
stöd och handledning för unga
Högskoleutbildning
övriga studiemöjligheter
dagvård
i Vanda finns både kommunala och privata daghem .
kommunen övervakar också den privata dagvården .
i Vanda ges dagvård på finska , svenska , ryska och engelska .
inom dagvården ges även undervisning i finska som andra språk .
dagvård ordnas också inom familjedagvården och i gruppfamiljedaghem .
man ska ansöka om dagvårdsplats för sitt barn minst fyra månader innan barnet ska börja i dagvården .
du kan ansöka om plats i den kommunala dagvården via Internet eller med en pappersblankett .
för en elektronisk ansökan behöver du egna nätbankskoder eller en elektronisk legitimation .
Pappersblanketter kan hämtas till exempel vid Vandainfo eller daghemmen .
privata dagvårdsplatser söks direkt på daghemmet .
frågor kring dagvård och ansökan om dagvårdsplats kan du ställa till daghemsföreståndaren eller skicka till adressen varhaiskasvatus ( at ) vantaa.fi .
vanligtvis ansöker man om dagvårdsplats i den egna kommunen .
om familjen bor nära gränsen till Helsingfors eller Esbo , kan du också söka dagvårdsplats i grannkommunen .
du ska ändå lämna in din ansökan i den egna kommunen .
mer information hittar du via tjänsten Helsingforsregionen.fi .
Läs mer : dagvård
linkkiVanda stad :
privat dagvårdfinska _ svenska _ engelska
linkkiVanda stad :
privat dagvårdfinska
linkkiVanda stad :
ansökan om dagvårdsplatsfinska _ svenska _ engelska
linkkiVanda stad :
elektronisk ansökningsblankett för dagvårdenfinska _ svenska _ engelska
information om dagvården finska _ svenska _ engelska
förskoleundervisning
förskoleundervisning ( esiopetus ) ordnas i både kommunala och privata daghem samt i förskoleenheter i skolornas lokaler .
i Vanda kan man få förskoleundervisning på finska , svenska och engelska .
du måste ansöka om plats i förskoleundervisningen .
ansökan kan göras elektroniskt via stadens webbplats eller med en pappersblankett .
ansökningstiden är i januari , men ansökan kan även lämnas in övriga tider , om familjen till exempel flyttar till Vanda mitt under året .
förberedande undervisning tillhandahålls för invandrarbarn som inte har tillräckliga kunskaper i finska för att klara sig i förskoleundervisningen .
den förberedande undervisningen är avsedd för 6 @-@ åriga barn med invandrarbakgrund .
den ordnas i daghemmens förskolegrupper .
daghemmet anvisar barnet till den förberedande undervisningen i samband med ansökningen till förskoleundervisningen .
du hittar mer information om förskoleundervisningen , ansökning till förskoleundervisningen och om undervisning som förbereder för förskoleundervisning på Vanda stads ( Vantaan kaupunki ) webbplats .
du kan även fråga om mer information på daghemmen .
Läs mer : förskoleundervisning
linkkiVanda stad :
ansökan till förskoleundervisningfinska _ svenska _ engelska
linkkiVanda stad :
information om den förberedande undervisningenfinska _ engelska
linkkiVanda stad :
elektronisk ansökningsblankett för förskoleundervisningenfinska _ svenska _ engelska
linkkiVanda stad :
daghem som ger förskoleundervisningfinska _ engelska
grundläggande utbildning
i Vanda finns finskspråkiga och svenskspråkiga grundskolor ( peruskoulu ) .
i Vanda finns även en internationell skola , där man kan avlägga grundskolan på engelska .
mer information om skolorna i Vanda hittar du på Vanda stads ( Vantaan kaupunki ) webbplats .
anmälan till grundskolan ska göras på förhand .
Anmälningstiden är vanligtvis i januari .
på stadens webbplats hittar du kontaktuppgifterna till skolorna och mer information om anmälan .
Läs mer : grundläggande utbildning
linkkiVanda stad :
anmälan till skolanfinska _ svenska _ engelska
linkkiVanda stad :
skolornas kontaktuppgifterfinska
Eftermiddagsverksamhetfinska _ svenska
förberedande utbildning inför grundskola
om barnets kunskaper i det finska språket inte är tillräckligt bra för studier i den finskspråkiga grundskolan , kan barnet få förberedande utbildning ( valmistava opetus ) .
i den förberedande utbildningen läser barnen det finska språket och grundskolans läroämnen .
undervisningen pågår vanligtvis i ett år .
om du har anlänt till Finland för en kort tid sedan och har barn under skolåldern ska du ta kontakt med områdeskoordinatorn för ditt bostadsområde ( aluekoordinaattori ) .
områdeskoordinatorn berättar om hur undervisningen ordnas och hjälper dig i frågor som rör barnets skolgång .
information om den förberedande undervisningenfinska
linkkiVanda stad :
Områdeskoordinatorerfinska
grundläggande utbildning för unga invandrare
vid Vanda vuxenutbildningsinstitut ( Vantaan aikuisopisto ) kan 17 @-@ 24 @-@ åriga invandrarungdomar avlägga grundskolans avgångsbetyg .
om man har hoppat av grundskolan , kan man avlägga grundskolans lärokurs också vid Eira vuxengymnasium ( Eiran aikuislukio ) .
grundläggande utbildning för invandrarefinska
linkkiEira vuxengymnasium :
grundundervisning för vuxnafinska
tionde klasserna
du kan ansöka till den grundläggande utbildningens tilläggsundervisning , det vill säga till en tionde klass ( kymppiluokka ) , om du fick grundskolans avgångsbetyg samma år eller året innan , men inte har fått en studieplats på andra stadiet .
på tionde klassen kan du höja dina betyg från grundskolan och du får en plan för fortsatta studier .
Tiondeklasserna i Vanda finns i östra och västra Vanda vid Varias verksamhetsställen och vid Lumo gymnasium ( Lumon lukio ) .
linkkiVanda stad :
Tiondeklasserfinska _ svenska
invandrare och grundläggande utbildning
i skolorna i Vanda ges hemspråksundervisning i flera olika språk .
i grundskolorna ges även utbildning i finska som andraspråk ( suomi toisena kielenä ) till elever som har ett annat modersmål än finska , svenska eller samiska , och vars kunskaper i det finska språket inte är i nivå med modersmålet .
när du anmäler dig till skolan , kan du samtidigt anmäla dig till hemspråksundervisning och undervisning i din egen religion .
du kan även anmäla dig till undervisningen genom att fylla i en blankett , som du får från din egen skola .
den ifyllda blanketten returneras till den egna skolan .
undervisning i den egna religionen kan ordnas om gruppen består av minst tre elever .
mer information om hemspråksundervisning och om undervisning i elevens egen religion hittar du på stadens webbplats och hos områdeskoordinatorerna ( aluekoordinaattori ) .
linkkiVanda stad :
information om hemspråksundervisningfinska
linkkiVanda stad :
undervisning i den egna religionenfinska
finska som andra språk i den grundläggande undervisningenfinska
linkkiVanda stad :
Områdeskoordinatorerfinska
yrkesutbildning
i Vanda ordnas yrkesutbildning vid yrkesinstitutet Vantaan ammattiopisto Varia , handelsläroanstalten MERCURIA samt TTS Arbetseffektivitetsföreningen rf:s verksamhetsställe i Vanda .
i Varia ordnas även engelskspråkig undervisning samt finskspråkiga yrkesutbildningar särskilt avsedda för invandrare .
Edupoli ordnar yrkesutbildning för vuxna .
i Vanda finns även Finavia Avia College som ger utbildning för olika luftfartsyrken .
Läs mer : yrkesutbildning .
linkkiVanda stad :
yrkesutbildningfinska _ svenska
linkkiYrkesläroanstalten Varia i Vanda :
yrkesutbildningfinska _ engelska
yrkesutbildningfinska _ engelska
linkkiTTS Arbetseffektivitetsföreningen rf:s verksamhetsställe i Vanda :
yrkesutbildningfinska
utbildning som handleder för yrkesutbildning ( VALMA )
utbildning som handleder för grundläggande yrkesutbildning ( Ammatilliseen peruskoulutukseen valmentava koulutus ) d.v.s. VALMA är avsedd för dem som vill avlägga en grundläggande yrkesutbildning .
under VALMA @-@ utbildningen får du kunskap och färdigheter som hjälper dig i dina senare yrkesinriktade studier .
du kan även förbättra din språkkunskap . du kan också höja dina grundskolebetyg .
i Vanda ordnas VALMA @-@ utbildning av Varia .
Läs mer om VALMA @-@ utbildningen på InfoFinlands sida Utbildning som handleder för yrkesutbildning .
linkkiVanda stad :
information om VALMA @-@ utbildningarfinska
linkkiYrkesläroanstalten Varia i Vanda :
i Vanda kan du studera på gymnasiet ( lukio ) på finska , svenska eller engelska .
undervisning på engelska erbjuds på IB @-@ linjen vid gymnasieskolan Tikkurilan lukio .
i Vanda finns även ett vuxengymnasium .
Läs mer : gymnasium .
linkkiVanda stad :
information om gymnasieutbildningfinska _ svenska
linkkiVanda stad :
gymnasierna och gymnasiernas hemsidorfinska
linkkiVanda stad :
Vuxengymnasiumfinska
linkkiVanda stad :
Distansgymnasiumfinska
linkkiVanda stad :
Steinergymnasietfinska
förberedande gymnasieutbildning ( LUVA )
om du vill förbättra dina kunskaper i finska eller svenska innan du söker till ett gymnasium , kan du söka till en förberedande gymnasieutbildning .
den är avsedd för invandrare .
i Vanda ordnas LUVA @-@ utbildning av Lumon lukio .
Läs mer om LUVA @-@ utbildningen på InfoFinlands sida Förberedande gymnasieutbildning .
linkkiVanda stad :
förberedande gymnasieutbildningfinska
stöd och handledning för unga
om du är under 30 år gammal kan du få råd och handledning via Ohjaamo @-@ tjänsten .
Ohjaamos personal hjälper dig om du inte har ett arbete eller en studieplats .
du kan även fråga om andra saker , som till exempel boende eller ekonomiska frågor .
linkkiOhjaamo :
stöd och handledning för ungafinska _ engelska
Vägledningscentret Kipinä
om du är under 29 år gammal , bor i Vanda och inte har ett jobb eller en studieplats , kan du få råd och handledning i Kipinä .
ring och boka en tid i förväg .
utan tidsbokning kan du besöka Kipinä på tisdagar och onsdagar kl . 12.00 @-@ 18.00 .
mer information hittar du på webbplatsen .
Kipinä
Banvägen 2 , Dickursby
tfn 050.312.4372
vägledning och stöd för ungafinska _ svenska
Högskoleutbildning
i Vanda finns två yrkeshögskolor ( ammattikorkeakoulu ) , Laurea och Metropolia .
de erbjuder utbildning inom många olika branscher .
mer information om utbildningsprogram och om ansökan hittar du på läroanstalternas webbplats .
också Helsingfors universitets öppna universitet ( avoin yliopisto ) har verksamhetsställen i Vanda . där ges undervisning på högskolenivå och fortbildning .
Läs mer : yrkeshögskolor , Universitet .
linkkiVanda stad :
Högskoleutbildningfinska
yrkeshögskolafinska _ engelska
linkkiMetropolia :
yrkeshögskolafinska _ engelska
Ubildning vid öppna universitetet i Vandafinska _ svenska _ engelska
övriga studiemöjligheter
vid Vanda vuxenutbildningsinstitut ( Vantaan aikuisopisto ) kan du studera till exempel språk , handarbete och matlagning eller delta i ledd motion .
kurserna är avgiftsbelagda och de ordnas både dag- och kvällstid .
Vuxenutbildningsinstitutet ordnar även kurser för invandrare .
mer information hittar du på Vanda stads webbplats .
Läs mer : studier som hobby .
linkkiVanda vuxenutbildningsinstitut :
Studiehandbokfinska
linkkiVanda vuxenutbildningsinstitut :
kurser i finska och svenska språket för invandrarefinska
linkkiEdupoli :
Vuxenutbildningscenterfinska
detta innehåll finns inte på det språk som du har valt .
Välj något annat språk .
finska
detta innehåll finns inte på det språk som du har valt .
Välj något annat språk .
finska
detta innehåll finns inte på det språk som du har valt .
Välj något annat språk .
finska
hyresbostad
boende i en krissituation
Bostadslöshet
Stöd- och serviceboende
Bostadens avfallshantering
hyresbostad
Hyresbostäderna är ofta dyra i huvudstadsregionen .
du är själv ansvarig för att skaffa bostad åt dig själv .
Varken staden eller andra hyresvärdar har skyldighet att erbjuda dig bostad .
Läs mer : hyresbostad .
privata hyresbostäder
i Vanda finns också många andra hyresvärdar , varav de största är VVO , Sato och Avara .
Därtill ägs hyresbostäder i Vanda av många försäkringsbolag , Kuntien eläkevakuutus och Kunta @-@ asunnot .
det kan gå snabbt att få bostad via en privat hyresvärd .
om du är studerande kan du ansöka om en hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS ( Helsingin seudun Opiskelija @-@ asuntosäätiö HOAS ) .
om du är yngre än 30 år , kan du söka bostad hos Förbundet för ungdomsbostäder ( Nuorisoasuntoliitto ) och stiftelsen Nuorisosäätiö ( Nuorisosäätiö ) .
linkkiSATO :
hyresbostäderfinska _ engelska
linkkiAvara :
hyresbostäderfinska
linkkiKommunbostäder :
hyresbostäderfinska _ svenska _ engelska
linkkiFörbundet för ungdomsbostäder :
hyresbostäder för personer under 30 årfinska _ engelska
hyresbostäder för ungafinska _ engelska
linkkiHOAS :
hyresbostäder för studerandefinska _ svenska _ engelska
stadens hyresbostäder
stadens hyresbostäder är vanligtvis förmånligare än de bostäder som hyrs ut av företag och privatpersoner .
Väntetiden för dessa bostäder kan dock vara lång och endast en liten del av de sökande får en bostad .
Vanda stads hyresbostäder ägs och hyrs ut av VAV Asunnot Oy .
Lokgränden 7
tfn 010.235.1450 ( kundtjänst )
du kan göra en bostadsansökan på VAV Asunnot Oy:s webbplats .
ansökan är giltig i fyra månader och måste sedan förnyas .
vid val av invånare till stadens hyresbostäder prioriteras de sökande som har ett akut bostadsbehov .
också sökandens inkomster beaktas , eftersom bostäderna främst är avsedda för personer med låga inkomster .
information om stadens hyresbostäderfinska _ engelska
ansökan om hyresbostad i stadenfinska _ engelska
boende i en krissituation
om din bostad har skadats till exempel till följd av brand eller vattenskada kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna .
kontakta ditt försäkringsbolag direkt när skadan har inträffat .
i krissituationer får man även hjälp vid Vanda stads social- och krisjour ( sosiaali- ja kriisipäivystys ) , som har öppet dygnet runt .
telefonnumret till social- och krisjouren är ( 09 ) 8392.4005
linkkiVanda stad :
social- och krisjourenfinska _ svenska _ engelska
skyddshem
om någon i din familj utövar våld mot dig eller hotar dig med våld , kan du kontakta ett skyddshem ( turvakoti ) .
Skyddshemmen har jourmottagning dygnet runt .
skyddshemmet Mona är ett skyddshem avsett för invandrarkvinnor och deras barn .
tfn 045.639.6274
du kan även gå till Vanda skyddshem eller huvudstadsregionens skyddshem .
tfn ( 09 ) 8392.0071
Steniusvägen 20
tfn ( 09 ) 4777.180
linkkiTurvakoti Mona :
skyddshemfinska
skyddshemfinska _ engelska
hjälp till offer för familjevåldfinska
hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
de ungas skyddshus
Finlands Röda Kors De ungas skyddshus ( Suomen Punaisen Ristin Nuorten turvatalo ) ger stöd och hjälp i krissituationer för 12 @-@ 19 @-@ åriga ungdomar .
skyddshuset har öppet kl . 17 @-@ 10 , telefonjouren betjänar dygnet runt .
Sjukhusgatan 3 ( Räckhals gård )
tfn ( 09 ) 871.4043
linkkiFinlands Röda Kors :
de ungas skyddshusfinska _ svenska _ engelska
Bostadslöshet
om du blir bostadslös ska du kontakta socialstationen ( sosiaaliasema ) för ditt eget område .
kontaktuppgifterna hittar du på Vanda stads webbplats .
om din hemkommun är Vanda , kan du få en bostad via Sininauha Oy eller Villenpirtti .
Läs mer : Bostadslöshet
linkkiVanda stad :
Socialtjänsterfinska _ svenska _ engelska
bostäder för bostadslösafinska
Stödboende för personer med psykisk ohälsa och missbruksproblemfinska
Stöd- och serviceboende
staden ordnar boendetjänster till exempel för åldringar och handikappade , som har svårt att klara av de dagliga sysslorna utan hjälp .
åldringar och handikappade som inte klarar av att bo självständigt , kan bo i servicehus ( palvelutalo ) eller på en vårdinrättning ( laitos ) .
mer information om dessa tjänster får du från enheten för socialt arbete ( sosiaalityön yksikkö ) i ditt bostadsområde .
Läs mer : Stöd- och serviceboende .
linkkiVanda stad :
information om hemvårdens stödtjänsterfinska
linkkiVanda stad :
information om stadens servicebostäderfinska
linkkiVanda stad :
privata servicehusfinska
linkkiVanda stad :
Socialtjänsterfinska _ svenska _ engelska
Bostadens avfallshantering
information om var din närmaste återvinningsstation ( kierrätyspiste ) ligger hittar du på webbplatsen kierrätys.info .
Läs mer : avfallshantering och återvinning .
linkkiAvfallsverksföreningen :
Återvinningsstationerfinska
linkkiHRM :
Återvinningsstationerfinska _ svenska _ engelska
hyresbostad
boende i en krissituation
Bostadslöshet
Stöd- och serviceboende
Bostadens avfallshantering
hyresbostad
Hyresbostäderna är ofta dyra i huvudstadsregionen .
du är själv ansvarig för att skaffa bostad åt dig själv .
Varken staden eller andra hyresvärdar har skyldighet att erbjuda dig bostad .
Läs mer : hyresbostad .
privata hyresbostäder
i Vanda finns också många andra hyresvärdar , varav de största är VVO , Sato och Avara .
Därtill ägs hyresbostäder i Vanda av många försäkringsbolag , Kuntien eläkevakuutus och Kunta @-@ asunnot .
det kan gå snabbt att få bostad via en privat hyresvärd .
om du är studerande kan du ansöka om en hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS ( Helsingin seudun Opiskelija @-@ asuntosäätiö HOAS ) .
om du är yngre än 30 år , kan du söka bostad hos Förbundet för ungdomsbostäder ( Nuorisoasuntoliitto ) och stiftelsen Nuorisosäätiö ( Nuorisosäätiö ) .
linkkiSATO :
hyresbostäderfinska _ engelska
linkkiAvara :
hyresbostäderfinska
linkkiKommunbostäder :
hyresbostäderfinska _ svenska _ engelska
linkkiFörbundet för ungdomsbostäder :
hyresbostäder för personer under 30 årfinska _ engelska
hyresbostäder för ungafinska _ engelska
linkkiHOAS :
hyresbostäder för studerandefinska _ svenska _ engelska
stadens hyresbostäder
stadens hyresbostäder är vanligtvis förmånligare än de bostäder som hyrs ut av företag och privatpersoner .
Väntetiden för dessa bostäder kan dock vara lång och endast en liten del av de sökande får en bostad .
Vanda stads hyresbostäder ägs och hyrs ut av VAV Asunnot Oy .
Lokgränden 7
tfn 010.235.1450 ( kundtjänst )
du kan göra en bostadsansökan på VAV Asunnot Oy:s webbplats .
ansökan är giltig i fyra månader och måste sedan förnyas .
vid val av invånare till stadens hyresbostäder prioriteras de sökande som har ett akut bostadsbehov .
också sökandens inkomster beaktas , eftersom bostäderna främst är avsedda för personer med låga inkomster .
information om stadens hyresbostäderfinska _ engelska
ansökan om hyresbostad i stadenfinska _ engelska
boende i en krissituation
om din bostad har skadats till exempel till följd av brand eller vattenskada kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna .
kontakta ditt försäkringsbolag direkt när skadan har inträffat .
i krissituationer får man även hjälp vid Vanda stads social- och krisjour ( sosiaali- ja kriisipäivystys ) , som har öppet dygnet runt .
telefonnumret till social- och krisjouren är ( 09 ) 8392.4005
linkkiVanda stad :
social- och krisjourenfinska _ svenska _ engelska
skyddshem
om någon i din familj utövar våld mot dig eller hotar dig med våld , kan du kontakta ett skyddshem ( turvakoti ) .
Skyddshemmen har jourmottagning dygnet runt .
skyddshemmet Mona är ett skyddshem avsett för invandrarkvinnor och deras barn .
tfn 045.639.6274
du kan även gå till Vanda skyddshem eller huvudstadsregionens skyddshem .
tfn ( 09 ) 8392.0071
Steniusvägen 20
tfn ( 09 ) 4777.180
linkkiTurvakoti Mona :
skyddshemfinska
skyddshemfinska _ engelska
hjälp till offer för familjevåldfinska
hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
de ungas skyddshus
Finlands Röda Kors De ungas skyddshus ( Suomen Punaisen Ristin Nuorten turvatalo ) ger stöd och hjälp i krissituationer för 12 @-@ 19 @-@ åriga ungdomar .
skyddshuset har öppet kl . 17 @-@ 10 , telefonjouren betjänar dygnet runt .
Sjukhusgatan 3 ( Räckhals gård )
tfn ( 09 ) 871.4043
linkkiFinlands Röda Kors :
de ungas skyddshusfinska _ svenska _ engelska
Bostadslöshet
om du blir bostadslös ska du kontakta socialstationen ( sosiaaliasema ) för ditt eget område .
kontaktuppgifterna hittar du på Vanda stads webbplats .
om din hemkommun är Vanda , kan du få en bostad via Sininauha Oy eller Villenpirtti .
Läs mer : Bostadslöshet
linkkiVanda stad :
Socialtjänsterfinska _ svenska _ engelska
bostäder för bostadslösafinska
Stödboende för personer med psykisk ohälsa och missbruksproblemfinska
Stöd- och serviceboende
staden ordnar boendetjänster till exempel för åldringar och handikappade , som har svårt att klara av de dagliga sysslorna utan hjälp .
åldringar och handikappade som inte klarar av att bo självständigt , kan bo i servicehus ( palvelutalo ) eller på en vårdinrättning ( laitos ) .
mer information om dessa tjänster får du från enheten för socialt arbete ( sosiaalityön yksikkö ) i ditt bostadsområde .
Läs mer : Stöd- och serviceboende .
linkkiVanda stad :
information om hemvårdens stödtjänsterfinska
linkkiVanda stad :
information om stadens servicebostäderfinska
linkkiVanda stad :
privata servicehusfinska
linkkiVanda stad :
Socialtjänsterfinska _ svenska _ engelska
Bostadens avfallshantering
information om var din närmaste återvinningsstation ( kierrätyspiste ) ligger hittar du på webbplatsen kierrätys.info .
Läs mer : avfallshantering och återvinning .
linkkiAvfallsverksföreningen :
Återvinningsstationerfinska
linkkiHRM :
Återvinningsstationerfinska _ svenska _ engelska
hyresbostad
boende i en krissituation
Bostadslöshet
Stöd- och serviceboende
Bostadens avfallshantering
hyresbostad
Hyresbostäderna är ofta dyra i huvudstadsregionen .
du är själv ansvarig för att skaffa bostad åt dig själv .
Varken staden eller andra hyresvärdar har skyldighet att erbjuda dig bostad .
Läs mer : hyresbostad .
privata hyresbostäder
i Vanda finns också många andra hyresvärdar , varav de största är VVO , Sato och Avara .
Därtill ägs hyresbostäder i Vanda av många försäkringsbolag , Kuntien eläkevakuutus och Kunta @-@ asunnot .
det kan gå snabbt att få bostad via en privat hyresvärd .
om du är studerande kan du ansöka om en hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS ( Helsingin seudun Opiskelija @-@ asuntosäätiö HOAS ) .
om du är yngre än 30 år , kan du söka bostad hos Förbundet för ungdomsbostäder ( Nuorisoasuntoliitto ) och stiftelsen Nuorisosäätiö ( Nuorisosäätiö ) .
linkkiSATO :
hyresbostäderfinska _ engelska
linkkiAvara :
hyresbostäderfinska
linkkiKommunbostäder :
hyresbostäderfinska _ svenska _ engelska
linkkiFörbundet för ungdomsbostäder :
hyresbostäder för personer under 30 årfinska _ engelska
hyresbostäder för ungafinska _ engelska
linkkiHOAS :
hyresbostäder för studerandefinska _ svenska _ engelska
stadens hyresbostäder
stadens hyresbostäder är vanligtvis förmånligare än de bostäder som hyrs ut av företag och privatpersoner .
Väntetiden för dessa bostäder kan dock vara lång och endast en liten del av de sökande får en bostad .
Vanda stads hyresbostäder ägs och hyrs ut av VAV Asunnot Oy .
Lokgränden 7
tfn 010.235.1450 ( kundtjänst )
du kan göra en bostadsansökan på VAV Asunnot Oy:s webbplats .
ansökan är giltig i fyra månader och måste sedan förnyas .
vid val av invånare till stadens hyresbostäder prioriteras de sökande som har ett akut bostadsbehov .
också sökandens inkomster beaktas , eftersom bostäderna främst är avsedda för personer med låga inkomster .
information om stadens hyresbostäderfinska _ engelska
ansökan om hyresbostad i stadenfinska _ engelska
boende i en krissituation
om din bostad har skadats till exempel till följd av brand eller vattenskada kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna .
kontakta ditt försäkringsbolag direkt när skadan har inträffat .
i krissituationer får man även hjälp vid Vanda stads social- och krisjour ( sosiaali- ja kriisipäivystys ) , som har öppet dygnet runt .
telefonnumret till social- och krisjouren är ( 09 ) 8392.4005
linkkiVanda stad :
social- och krisjourenfinska _ svenska _ engelska
skyddshem
om någon i din familj utövar våld mot dig eller hotar dig med våld , kan du kontakta ett skyddshem ( turvakoti ) .
Skyddshemmen har jourmottagning dygnet runt .
skyddshemmet Mona är ett skyddshem avsett för invandrarkvinnor och deras barn .
tfn 045.639.6274
du kan även gå till Vanda skyddshem eller huvudstadsregionens skyddshem .
tfn ( 09 ) 8392.0071
Steniusvägen 20
tfn ( 09 ) 4777.180
linkkiTurvakoti Mona :
skyddshemfinska
skyddshemfinska _ engelska
hjälp till offer för familjevåldfinska
hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
de ungas skyddshus
Finlands Röda Kors De ungas skyddshus ( Suomen Punaisen Ristin Nuorten turvatalo ) ger stöd och hjälp i krissituationer för 12 @-@ 19 @-@ åriga ungdomar .
skyddshuset har öppet kl . 17 @-@ 10 , telefonjouren betjänar dygnet runt .
Sjukhusgatan 3 ( Räckhals gård )
tfn ( 09 ) 871.4043
linkkiFinlands Röda Kors :
de ungas skyddshusfinska _ svenska _ engelska
Bostadslöshet
om du blir bostadslös ska du kontakta socialstationen ( sosiaaliasema ) för ditt eget område .
kontaktuppgifterna hittar du på Vanda stads webbplats .
om din hemkommun är Vanda , kan du få en bostad via Sininauha Oy eller Villenpirtti .
Läs mer : Bostadslöshet
linkkiVanda stad :
Socialtjänsterfinska _ svenska _ engelska
bostäder för bostadslösafinska
Stödboende för personer med psykisk ohälsa och missbruksproblemfinska
Stöd- och serviceboende
staden ordnar boendetjänster till exempel för åldringar och handikappade , som har svårt att klara av de dagliga sysslorna utan hjälp .
åldringar och handikappade som inte klarar av att bo självständigt , kan bo i servicehus ( palvelutalo ) eller på en vårdinrättning ( laitos ) .
mer information om dessa tjänster får du från enheten för socialt arbete ( sosiaalityön yksikkö ) i ditt bostadsområde .
Läs mer : Stöd- och serviceboende .
linkkiVanda stad :
information om hemvårdens stödtjänsterfinska
linkkiVanda stad :
information om stadens servicebostäderfinska
linkkiVanda stad :
privata servicehusfinska
linkkiVanda stad :
Socialtjänsterfinska _ svenska _ engelska
Bostadens avfallshantering
information om var din närmaste återvinningsstation ( kierrätyspiste ) ligger hittar du på webbplatsen kierrätys.info .
Läs mer : avfallshantering och återvinning .
linkkiAvfallsverksföreningen :
Återvinningsstationerfinska
linkkiHRM :
Återvinningsstationerfinska _ svenska _ engelska
möjligheter att studera det finska eller svenska språket
språkkurser
med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors , Vanda , Esbo eller Grankulla .
kurserna i svenska hittar du genom att klicka på länken på tjänstens startsida .
kurserna i tjänsten finnishcourses.fi är öppna för alla .
tjänsten omfattar inte arbets- och näringsbyråns kurser .
i Vanda anordnas kurser i finska och svenska språket för invandrare av Vanda vuxenutbildningsinstitut ( Vantaan aikuisopisto ) Kurserna vid institutet är öppna för alla .
Vuxenutbildningsinstitutet ligger i Dickursby , men kurser ordnas runtom i Vanda .
adress :
Näckrosvägen 5
tfn ( 09 ) 8392.4342
ytterligare information om kurser och anmälan hittar du på Vanda vuxenutbildningsinstituts webbplats och i studiehandboken .
du får studiehandboken till exempel på bibliotek eller Vandainfo samt i elektroniskt format på Vanda stads webbplats .
arbets- och näringsbyrån anvisar invandrare till kurser i finska språket som ingår i integrationsprocessen .
i samband med att en integrations- eller sysselsättningsplan upprättas för dig , kan du också få också en studieplats på en finskakurs reserverad eller också kan du ställas i kö för en studieplats .
mer information hittar du vid arbets- och näringsbyrån .
Läs mer : studier i finska och svenska
kurser i finska och svenska språketfinska _ engelska _ ryska
linkkiVanda vuxenutbildningsinstitut :
kurser i finska och svenska språket för invandrarefinska
linkkiArbets- och näringsministeriet :
utbildning i finska och svenska språketfinska _ svenska _ engelska
linkkiVanda vuxenutbildningsinstitut :
grundundervisning för vuxnafinska
samtal på finska
på Vanda stadsbibliotek anordnas språkcaféer ( kielikahvila ) , där man kan öva på att prata finska .
alla som vill lära sig tala finska är välkomna till caféerna .
på språkcaféerna talar vi finska , så det är bra om du redan kan lite finska .
språkcaféerna är avgiftsfria .
mer information om språkcaféerna får du från biblioteken .
i Vanda anordnas samtalsklubbar på finska också på Silkesportens verksamhetscenter ( Silkinportin toimintakeskus ) och Kafnettis och Myyrinkis boendeträffpunkter ( Kafnetin ja Myyringin asukastila ) .
Finskaklubbar avsedda för föräldrar som vårdar barn i hemmet anordnas i invånarparkerna ( asukaspuisto ) och i de öppna daghemmen ( avoin päiväkoti ) .
Klubbarna för att lära sig tala finska är avgiftsfria .
Läsundervisning
nätverket Vi läser tillsammans ( Luetaan yhdessä @-@ verkosto ) erbjuder undervisning i läsning och det finska språket för invandrarkvinnor .
flera olika Vi läser tillsammans @-@ nätverk är verksamma på olika håll i Vanda .
det är avgiftsfritt att delta i grupperna .
Språkkaféerfinska _ engelska _ ryska
linkkiVanda stad :
Invånarlokalfinska _ engelska
linkkiVanda stad :
Invånarlokalfinska _ engelska
linkkiVanda stad :
Parker för invånare och öppna daghemfinska _ svenska _ engelska
linkkiVi läser tillsammans @-@ nätverket :
Vi läser tillsammans i Vandafinska _ svenska _ engelska
allmän språkexamen
du kan avlägga allmän språkexamen i finska eller svenska språket .
på utbildningsstyrelsens ( Opetushallitus ) webbplats finns en sökmotor med vilken du kan kontrollera var och när du kan avlägga examen .
i Vanda ordnas språkexamina till exempel vid Vanda vuxenutbildningsinstitut ( Vantaan aikuisopisto ) .
Läs mer : Officiellt intyg på språkkunskaper .
linkkiUtbildningsstyrelsen :
att anmäla sig till en allmän språkexamen och examensavgifterfinska _ svenska _ engelska
linkkiVanda vuxenutbildningsinstitut :
allmän språkexamenfinska
linkkiUtbildningsstyrelsen :
Examenssökningfinska
möjligheter att studera det finska eller svenska språket
språkkurser
med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors , Vanda , Esbo eller Grankulla .
kurserna i svenska hittar du genom att klicka på länken på tjänstens startsida .
kurserna i tjänsten finnishcourses.fi är öppna för alla .
tjänsten omfattar inte arbets- och näringsbyråns kurser .
i Vanda anordnas kurser i finska och svenska språket för invandrare av Vanda vuxenutbildningsinstitut ( Vantaan aikuisopisto ) Kurserna vid institutet är öppna för alla .
Vuxenutbildningsinstitutet ligger i Dickursby , men kurser ordnas runtom i Vanda .
adress :
Näckrosvägen 5
tfn ( 09 ) 8392.4342
ytterligare information om kurser och anmälan hittar du på Vanda vuxenutbildningsinstituts webbplats och i studiehandboken .
du får studiehandboken till exempel på bibliotek eller Vandainfo samt i elektroniskt format på Vanda stads webbplats .
arbets- och näringsbyrån anvisar invandrare till kurser i finska språket som ingår i integrationsprocessen .
i samband med att en integrations- eller sysselsättningsplan upprättas för dig , kan du också få också en studieplats på en finskakurs reserverad eller också kan du ställas i kö för en studieplats .
mer information hittar du vid arbets- och näringsbyrån .
Läs mer : studier i finska och svenska
kurser i finska och svenska språketfinska _ engelska _ ryska
linkkiVanda vuxenutbildningsinstitut :
kurser i finska och svenska språket för invandrarefinska
linkkiArbets- och näringsministeriet :
utbildning i finska och svenska språketfinska _ svenska _ engelska
linkkiVanda vuxenutbildningsinstitut :
grundundervisning för vuxnafinska
samtal på finska
på Vanda stadsbibliotek anordnas språkcaféer ( kielikahvila ) , där man kan öva på att prata finska .
alla som vill lära sig tala finska är välkomna till caféerna .
på språkcaféerna talar vi finska , så det är bra om du redan kan lite finska .
språkcaféerna är avgiftsfria .
mer information om språkcaféerna får du från biblioteken .
i Vanda anordnas samtalsklubbar på finska också på Silkesportens verksamhetscenter ( Silkinportin toimintakeskus ) och Kafnettis och Myyrinkis boendeträffpunkter ( Kafnetin ja Myyringin asukastila ) .
Finskaklubbar avsedda för föräldrar som vårdar barn i hemmet anordnas i invånarparkerna ( asukaspuisto ) och i de öppna daghemmen ( avoin päiväkoti ) .
Klubbarna för att lära sig tala finska är avgiftsfria .
Läsundervisning
nätverket Vi läser tillsammans ( Luetaan yhdessä @-@ verkosto ) erbjuder undervisning i läsning och det finska språket för invandrarkvinnor .
flera olika Vi läser tillsammans @-@ nätverk är verksamma på olika håll i Vanda .
det är avgiftsfritt att delta i grupperna .
Språkkaféerfinska _ engelska _ ryska
linkkiVanda stad :
Invånarlokalfinska _ engelska
linkkiVanda stad :
Invånarlokalfinska _ engelska
linkkiVanda stad :
Parker för invånare och öppna daghemfinska _ svenska _ engelska
linkkiVi läser tillsammans @-@ nätverket :
Vi läser tillsammans i Vandafinska _ svenska _ engelska
allmän språkexamen
du kan avlägga allmän språkexamen i finska eller svenska språket .
på utbildningsstyrelsens ( Opetushallitus ) webbplats finns en sökmotor med vilken du kan kontrollera var och när du kan avlägga examen .
i Vanda ordnas språkexamina till exempel vid Vanda vuxenutbildningsinstitut ( Vantaan aikuisopisto ) .
Läs mer : Officiellt intyg på språkkunskaper .
linkkiUtbildningsstyrelsen :
att anmäla sig till en allmän språkexamen och examensavgifterfinska _ svenska _ engelska
linkkiVanda vuxenutbildningsinstitut :
allmän språkexamenfinska
linkkiUtbildningsstyrelsen :
Examenssökningfinska
möjligheter att studera det finska eller svenska språket
språkkurser
med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors , Vanda , Esbo eller Grankulla .
kurserna i svenska hittar du genom att klicka på länken på tjänstens startsida .
kurserna i tjänsten finnishcourses.fi är öppna för alla .
tjänsten omfattar inte arbets- och näringsbyråns kurser .
i Vanda anordnas kurser i finska och svenska språket för invandrare av Vanda vuxenutbildningsinstitut ( Vantaan aikuisopisto ) Kurserna vid institutet är öppna för alla .
Vuxenutbildningsinstitutet ligger i Dickursby , men kurser ordnas runtom i Vanda .
adress :
Näckrosvägen 5
tfn ( 09 ) 8392.4342
ytterligare information om kurser och anmälan hittar du på Vanda vuxenutbildningsinstituts webbplats och i studiehandboken .
du får studiehandboken till exempel på bibliotek eller Vandainfo samt i elektroniskt format på Vanda stads webbplats .
arbets- och näringsbyrån anvisar invandrare till kurser i finska språket som ingår i integrationsprocessen .
i samband med att en integrations- eller sysselsättningsplan upprättas för dig , kan du också få också en studieplats på en finskakurs reserverad eller också kan du ställas i kö för en studieplats .
mer information hittar du vid arbets- och näringsbyrån .
Läs mer : studier i finska och svenska
kurser i finska och svenska språketfinska _ engelska _ ryska
linkkiVanda vuxenutbildningsinstitut :
kurser i finska och svenska språket för invandrarefinska
linkkiArbets- och näringsministeriet :
utbildning i finska och svenska språketfinska _ svenska _ engelska
linkkiVanda vuxenutbildningsinstitut :
grundundervisning för vuxnafinska
samtal på finska
på Vanda stadsbibliotek anordnas språkcaféer ( kielikahvila ) , där man kan öva på att prata finska .
alla som vill lära sig tala finska är välkomna till caféerna .
på språkcaféerna talar vi finska , så det är bra om du redan kan lite finska .
språkcaféerna är avgiftsfria .
mer information om språkcaféerna får du från biblioteken .
i Vanda anordnas samtalsklubbar på finska också på Silkesportens verksamhetscenter ( Silkinportin toimintakeskus ) och Kafnettis och Myyrinkis boendeträffpunkter ( Kafnetin ja Myyringin asukastila ) .
Finskaklubbar avsedda för föräldrar som vårdar barn i hemmet anordnas i invånarparkerna ( asukaspuisto ) och i de öppna daghemmen ( avoin päiväkoti ) .
Klubbarna för att lära sig tala finska är avgiftsfria .
Läsundervisning
nätverket Vi läser tillsammans ( Luetaan yhdessä @-@ verkosto ) erbjuder undervisning i läsning och det finska språket för invandrarkvinnor .
flera olika Vi läser tillsammans @-@ nätverk är verksamma på olika håll i Vanda .
det är avgiftsfritt att delta i grupperna .
Språkkaféerfinska _ engelska _ ryska
linkkiVanda stad :
Invånarlokalfinska _ engelska
linkkiVanda stad :
Invånarlokalfinska _ engelska
linkkiVanda stad :
Parker för invånare och öppna daghemfinska _ svenska _ engelska
linkkiVi läser tillsammans @-@ nätverket :
Vi läser tillsammans i Vandafinska _ svenska _ engelska
allmän språkexamen
du kan avlägga allmän språkexamen i finska eller svenska språket .
på utbildningsstyrelsens ( Opetushallitus ) webbplats finns en sökmotor med vilken du kan kontrollera var och när du kan avlägga examen .
i Vanda ordnas språkexamina till exempel vid Vanda vuxenutbildningsinstitut ( Vantaan aikuisopisto ) .
Läs mer : Officiellt intyg på språkkunskaper .
linkkiUtbildningsstyrelsen :
att anmäla sig till en allmän språkexamen och examensavgifterfinska _ svenska _ engelska
linkkiVanda vuxenutbildningsinstitut :
allmän språkexamenfinska
linkkiUtbildningsstyrelsen :
Examenssökningfinska
var hittar jag jobb ?
hjälp med jobbsökningen
att starta ett företag
beskattning
var hittar jag jobb ?
TE @-@ byrån ( TE @-@ toimisto ) hjälper dig att söka arbete .
om du är arbetslös och söker efter arbete , ska du anmäla dig som arbetssökande hos TE @-@ byrån .
du kan anmäla dig antingen via nättjänsten eller personligen hos TE @-@ byrån .
medborgare i EU @-@ länderna , Island , Liechtenstein och Schweiz kan anmäla sig som arbetssökande via TE @-@ byråns nättjänst .
övriga länders medborgare måste anmäla sig personligen hos TE @-@ byrån .
ta med dig din legitimation och ditt uppehållstillstånd .
kontaktuppgifter :
information om TE @-@ byråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös .
information om att söka arbete i Finland hittar du på InfoFinlands sida : var hittar jag jobb ?
linkkiVanda arbets- och näringsbyrå :
kontaktuppgifter och tjänsterfinska _ svenska
linkkiArbets- och näringsministeriet :
lediga jobbfinska _ svenska
linkkiArbets- och näringsförvaltningen :
Länkar till jobbsajterfinska _ svenska _ engelska
linkkiVanda stad :
stöd för att hitta sysselsättningfinska _ svenska _ engelska
hjälp med jobbsökningen
stadens tjänster för arbetssökande
Vanda stad tillhandahåller olika tjänster för arbetslösa som hjälper dem att få kontakt med arbetslivet och hitta jobb .
i Vanda ordnas även många rekryteringsevenemang där arbetsgivarna söker arbetstagare .
du hittar mer information om stadens tjänster på Vanda stads webbplats .
linkkiVanda stad :
stadens tjänster för arbetssökandefinska _ svenska _ engelska
om du behöver hjälp med jobbsökningen eller med att hitta en studieplats kan du kontakta rådgivarna i Håkansböle internationella förenings Tsemppari @-@ projekt .
du hittar kontaktuppgifterna på Håkansböle internationella förenings webbplats .
Integrationscentret Kotoutumiskeskus Monika hjälper arbetslösa invandrarkvinnor att hitta jobb .
du kan få hjälp med att skriva din CV eller en jobbansökan , studera vardagsfinska och digitala färdigheter .
Luckan integration
Luckan Integration är en rådgivningstjänst , som erbjuder personlig rådgivning för invandrare och anordnar bland annat evenemang och grupper relaterade till jobbsökning .
språket som talas vid träffarna är engelska .
råd om jobbsökningfinska _ svenska _ engelska _ spanska
Väestöliittos karriärmentorskap är avsett för utbildade invandrare .
via programmet kan du få en mentor , som stödjer dig i sökningen efter arbete eller utbildningsplats eller i att starta eget företag .
verksamheten sker på finska .
Mentorskap i fråga om arbetskarriärfinska _ engelska
om du är under 30 år , kan du få råd och handledning via tjänsten Navigatorn .
Personalen vid Navigatorn hjälper dig om du inte har något arbete eller en studieplats .
Stödföreningen för unga invandrare R3 ( R3 Maahanmuuttajanuorten tuki ry ) hjälper ungdomar i frågor som rör utbildning och sysselsättning .
mer information hittar du på föreningens webbplats .
stöd för unga invandrarefinska
att starta ett företag
om du har ett företag i Vanda , kan du bli medlem i Vanda Företagare .
Vanda Företagare rf är företagarnas intressebevakningsorganisation som erbjuder sina medlemmar till exempel utbildning och rådgivning .
mer information hittar du på föreningens webbplats .
NewCo Helsinki erbjuder rådgivning och hjälp med att starta eget företag på finska , svenska , engelska , ryska , arabiska , estniska , tyska och italienska .
vid NewCo Helsinki ordnas informationsmöten om att starta eget för invandrare på finska , engelska , ryska , arabiska och estniska .
Infomötena är avgiftsfria .
NewCo Helsinki ordnar företagarutbildningar på finska , engelska och ryska .
en del av kurserna är avsedda för personer som ska starta eget företag och en del för dem som redan har eget företag .
kurser hålls på finska , engelska och ryska .
mer information och anmälan finns på NewCo Helsinki webbplats .
Nylands TE @-@ byrå ( TE @-@ toimisto ) erbjuder mångsidiga tjänster för personer som funderar på att starta eget och dem som är på väg att starta eget .
på Nylands TE @-@ byrå kan du till exempel delta i företagarutbildning och söka startpeng för att starta eget företag .
Läs mer : att grunda ett företag
tjänster för företagare med invandrarbakgrundfinska _ engelska
linkkiFöretagsFinland :
Företagsrådgivningfinska _ svenska _ engelska
Företagsrådgivningfinska _ engelska
företagarnas intressebevakningsorganisationfinska
beskattning
huvudstadsregionens skattebyrå betjänar kunderna i centrala Helsingfors .
kontaktuppgifter :
Alexandersgatan 9 ( Gloet )
tfn : 029.512.000
invandrare kan även sköta ärenden vid servicestället International House Helsinki .
på servicestället hjälper FPA:s och Skatteförvaltningens experter invandrare som kommer till Finland för att arbeta i frågor som rör beskattning och social trygghet
kontaktuppgifter till servicestället International House Helsinki :
Albertinkatu 25
Läs mer : beskattning
linkkiSkatteförvaltningen :
kontaktuppgifterfinska _ svenska _ engelska
rådgivning om social trygghet och beskattningfinska _ svenska _ engelska
IHH - serviceställe för dig som flyttar till Finland engelska
var hittar jag jobb ?
hjälp med jobbsökningen
att starta ett företag
beskattning
var hittar jag jobb ?
TE @-@ byrån ( TE @-@ toimisto ) hjälper dig att söka arbete .
om du är arbetslös och söker efter arbete , ska du anmäla dig som arbetssökande hos TE @-@ byrån .
du kan anmäla dig antingen via nättjänsten eller personligen hos TE @-@ byrån .
medborgare i EU @-@ länderna , Island , Liechtenstein och Schweiz kan anmäla sig som arbetssökande via TE @-@ byråns nättjänst .
övriga länders medborgare måste anmäla sig personligen hos TE @-@ byrån .
ta med dig din legitimation och ditt uppehållstillstånd .
kontaktuppgifter :
information om TE @-@ byråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös .
information om att söka arbete i Finland hittar du på InfoFinlands sida : var hittar jag jobb ?
linkkiVanda arbets- och näringsbyrå :
kontaktuppgifter och tjänsterfinska _ svenska
linkkiArbets- och näringsministeriet :
lediga jobbfinska _ svenska
linkkiArbets- och näringsförvaltningen :
Länkar till jobbsajterfinska _ svenska _ engelska
linkkiVanda stad :
stöd för att hitta sysselsättningfinska _ svenska _ engelska
hjälp med jobbsökningen
stadens tjänster för arbetssökande
Vanda stad tillhandahåller olika tjänster för arbetslösa som hjälper dem att få kontakt med arbetslivet och hitta jobb .
i Vanda ordnas även många rekryteringsevenemang där arbetsgivarna söker arbetstagare .
du hittar mer information om stadens tjänster på Vanda stads webbplats .
linkkiVanda stad :
stadens tjänster för arbetssökandefinska _ svenska _ engelska
om du behöver hjälp med jobbsökningen eller med att hitta en studieplats kan du kontakta rådgivarna i Håkansböle internationella förenings Tsemppari @-@ projekt .
du hittar kontaktuppgifterna på Håkansböle internationella förenings webbplats .
Integrationscentret Kotoutumiskeskus Monika hjälper arbetslösa invandrarkvinnor att hitta jobb .
du kan få hjälp med att skriva din CV eller en jobbansökan , studera vardagsfinska och digitala färdigheter .
Luckan integration
Luckan Integration är en rådgivningstjänst , som erbjuder personlig rådgivning för invandrare och anordnar bland annat evenemang och grupper relaterade till jobbsökning .
språket som talas vid träffarna är engelska .
råd om jobbsökningfinska _ svenska _ engelska _ spanska
Väestöliittos karriärmentorskap är avsett för utbildade invandrare .
via programmet kan du få en mentor , som stödjer dig i sökningen efter arbete eller utbildningsplats eller i att starta eget företag .
verksamheten sker på finska .
Mentorskap i fråga om arbetskarriärfinska _ engelska
om du är under 30 år , kan du få råd och handledning via tjänsten Navigatorn .
Personalen vid Navigatorn hjälper dig om du inte har något arbete eller en studieplats .
Stödföreningen för unga invandrare R3 ( R3 Maahanmuuttajanuorten tuki ry ) hjälper ungdomar i frågor som rör utbildning och sysselsättning .
mer information hittar du på föreningens webbplats .
stöd för unga invandrarefinska
att starta ett företag
om du har ett företag i Vanda , kan du bli medlem i Vanda Företagare .
Vanda Företagare rf är företagarnas intressebevakningsorganisation som erbjuder sina medlemmar till exempel utbildning och rådgivning .
mer information hittar du på föreningens webbplats .
NewCo Helsinki erbjuder rådgivning och hjälp med att starta eget företag på finska , svenska , engelska , ryska , arabiska , estniska , tyska och italienska .
vid NewCo Helsinki ordnas informationsmöten om att starta eget för invandrare på finska , engelska , ryska , arabiska och estniska .
Infomötena är avgiftsfria .
NewCo Helsinki ordnar företagarutbildningar på finska , engelska och ryska .
en del av kurserna är avsedda för personer som ska starta eget företag och en del för dem som redan har eget företag .
kurser hålls på finska , engelska och ryska .
mer information och anmälan finns på NewCo Helsinki webbplats .
Nylands TE @-@ byrå ( TE @-@ toimisto ) erbjuder mångsidiga tjänster för personer som funderar på att starta eget och dem som är på väg att starta eget .
på Nylands TE @-@ byrå kan du till exempel delta i företagarutbildning och söka startpeng för att starta eget företag .
Läs mer : att grunda ett företag
tjänster för företagare med invandrarbakgrundfinska _ engelska
linkkiFöretagsFinland :
Företagsrådgivningfinska _ svenska _ engelska
Företagsrådgivningfinska _ engelska
företagarnas intressebevakningsorganisationfinska
beskattning
huvudstadsregionens skattebyrå betjänar kunderna i centrala Helsingfors .
kontaktuppgifter :
Alexandersgatan 9 ( Gloet )
tfn : 029.512.000
invandrare kan även sköta ärenden vid servicestället International House Helsinki .
på servicestället hjälper FPA:s och Skatteförvaltningens experter invandrare som kommer till Finland för att arbeta i frågor som rör beskattning och social trygghet
kontaktuppgifter till servicestället International House Helsinki :
Albertinkatu 25
Läs mer : beskattning
linkkiSkatteförvaltningen :
kontaktuppgifterfinska _ svenska _ engelska
rådgivning om social trygghet och beskattningfinska _ svenska _ engelska
IHH - serviceställe för dig som flyttar till Finland engelska
var hittar jag jobb ?
hjälp med jobbsökningen
att starta ett företag
beskattning
var hittar jag jobb ?
TE @-@ byrån ( TE @-@ toimisto ) hjälper dig att söka arbete .
om du är arbetslös och söker efter arbete , ska du anmäla dig som arbetssökande hos TE @-@ byrån .
du kan anmäla dig antingen via nättjänsten eller personligen hos TE @-@ byrån .
medborgare i EU @-@ länderna , Island , Liechtenstein och Schweiz kan anmäla sig som arbetssökande via TE @-@ byråns nättjänst .
övriga länders medborgare måste anmäla sig personligen hos TE @-@ byrån .
ta med dig din legitimation och ditt uppehållstillstånd .
kontaktuppgifter :
information om TE @-@ byråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös .
information om att söka arbete i Finland hittar du på InfoFinlands sida : var hittar jag jobb ?
linkkiVanda arbets- och näringsbyrå :
kontaktuppgifter och tjänsterfinska _ svenska
linkkiArbets- och näringsministeriet :
lediga jobbfinska _ svenska
linkkiArbets- och näringsförvaltningen :
Länkar till jobbsajterfinska _ svenska _ engelska
linkkiVanda stad :
stöd för att hitta sysselsättningfinska _ svenska _ engelska
hjälp med jobbsökningen
stadens tjänster för arbetssökande
Vanda stad tillhandahåller olika tjänster för arbetslösa som hjälper dem att få kontakt med arbetslivet och hitta jobb .
i Vanda ordnas även många rekryteringsevenemang där arbetsgivarna söker arbetstagare .
du hittar mer information om stadens tjänster på Vanda stads webbplats .
linkkiVanda stad :
stadens tjänster för arbetssökandefinska _ svenska _ engelska
om du behöver hjälp med jobbsökningen eller med att hitta en studieplats kan du kontakta rådgivarna i Håkansböle internationella förenings Tsemppari @-@ projekt .
du hittar kontaktuppgifterna på Håkansböle internationella förenings webbplats .
Integrationscentret Kotoutumiskeskus Monika hjälper arbetslösa invandrarkvinnor att hitta jobb .
du kan få hjälp med att skriva din CV eller en jobbansökan , studera vardagsfinska och digitala färdigheter .
Luckan integration
Luckan Integration är en rådgivningstjänst , som erbjuder personlig rådgivning för invandrare och anordnar bland annat evenemang och grupper relaterade till jobbsökning .
språket som talas vid träffarna är engelska .
råd om jobbsökningfinska _ svenska _ engelska _ spanska
Väestöliittos karriärmentorskap är avsett för utbildade invandrare .
via programmet kan du få en mentor , som stödjer dig i sökningen efter arbete eller utbildningsplats eller i att starta eget företag .
verksamheten sker på finska .
Mentorskap i fråga om arbetskarriärfinska _ engelska
om du är under 30 år , kan du få råd och handledning via tjänsten Navigatorn .
Personalen vid Navigatorn hjälper dig om du inte har något arbete eller en studieplats .
Stödföreningen för unga invandrare R3 ( R3 Maahanmuuttajanuorten tuki ry ) hjälper ungdomar i frågor som rör utbildning och sysselsättning .
mer information hittar du på föreningens webbplats .
stöd för unga invandrarefinska
att starta ett företag
om du har ett företag i Vanda , kan du bli medlem i Vanda Företagare .
Vanda Företagare rf är företagarnas intressebevakningsorganisation som erbjuder sina medlemmar till exempel utbildning och rådgivning .
mer information hittar du på föreningens webbplats .
NewCo Helsinki erbjuder rådgivning och hjälp med att starta eget företag på finska , svenska , engelska , ryska , arabiska , estniska , tyska och italienska .
vid NewCo Helsinki ordnas informationsmöten om att starta eget för invandrare på finska , engelska , ryska , arabiska och estniska .
Infomötena är avgiftsfria .
NewCo Helsinki ordnar företagarutbildningar på finska , engelska och ryska .
en del av kurserna är avsedda för personer som ska starta eget företag och en del för dem som redan har eget företag .
kurser hålls på finska , engelska och ryska .
mer information och anmälan finns på NewCo Helsinki webbplats .
Nylands TE @-@ byrå ( TE @-@ toimisto ) erbjuder mångsidiga tjänster för personer som funderar på att starta eget och dem som är på väg att starta eget .
på Nylands TE @-@ byrå kan du till exempel delta i företagarutbildning och söka startpeng för att starta eget företag .
Läs mer : att grunda ett företag
tjänster för företagare med invandrarbakgrundfinska _ engelska
linkkiFöretagsFinland :
Företagsrådgivningfinska _ svenska _ engelska
Företagsrådgivningfinska _ engelska
företagarnas intressebevakningsorganisationfinska
beskattning
huvudstadsregionens skattebyrå betjänar kunderna i centrala Helsingfors .
kontaktuppgifter :
Alexandersgatan 9 ( Gloet )
tfn : 029.512.000
invandrare kan även sköta ärenden vid servicestället International House Helsinki .
på servicestället hjälper FPA:s och Skatteförvaltningens experter invandrare som kommer till Finland för att arbeta i frågor som rör beskattning och social trygghet
kontaktuppgifter till servicestället International House Helsinki :
Albertinkatu 25
Läs mer : beskattning
linkkiSkatteförvaltningen :
kontaktuppgifterfinska _ svenska _ engelska
rådgivning om social trygghet och beskattningfinska _ svenska _ engelska
IHH - serviceställe för dig som flyttar till Finland engelska
rådgivning för och integration av invandrare
inledande kartläggning
behöver du en tolk ?
rådgivning för och integration av invandrare
Invandrartjänster
Vanda stads tjänster för invandrare omfattar
mottagningstjänster för invandrare
integrationstjänster
Vanda stads tjänster för invandrare ( Vantaan maahanmuuttajapalvelut ) ger dig information om integration , social- och hälsovårdstjänster och om stadens och olika organisationers tjänster .
du kan bli klient om du flyttat till Finland på grund av familjeband , är flykting , offer för människohandel eller har rätt till en inledande kartläggning .
tfn ( 09 ) 839.21074 och ( 09 ) 839.32042
linkkiVanda stad :
Invandrartjänsterfinska _ engelska
Verksamhetscentret Silkesporten ( Silkinportin toimintakeskus ) ger rådgivning för invandrare och där ordnas många slags aktiviteter .
dickursbyvägen 44 F , vån .
tfn ( 09 ) 839.23651
linkkiSilkesportens verksamhetscenter :
rådgivning och verksamhet för invandrarefinska _ engelska
Vandainfo ger dig information om såväl Vandas stads som statens tjänster .
Vandainfon finns i Dickursby , Korso och Myrbacka .
Adresserna är :
Dixi , Banvägen 11 , 2:a vån .
tfn ( 09 ) 839.22133
tfn ( 09 ) 839.22133
tfn ( 09 ) 839.22133
kontaktuppgifterna och öppettiderna hittar du på Vanda stads webbplats .
linkkiVanda stad :
Vandainfofinska _ svenska _ engelska
den internationella föreningen i Håkansböle ( Hakunilan kansainvälinen yhdistys ) har en rådgivningspunkt som betjänar invandrare i Håkansböle , Björkby och andra områden i Vanda , som vill ha information om till exempel studier , språkkurser , arbete , hobbyverksamhet , krissituationer eller juridiska frågor .
Sporrgränden 2 A , vån . 3 ( Håkansböle )
tfn ( 09 ) 272.2775 och 040.501.3199 .
linkkiInternationella föreningen i Håkansböle :
rådgivning för invandrarefinska _ engelska _ ryska _ somaliska _ arabiska
på invandrarrådgivningen vid föreningen Vantaan Järjestörinki ry ( Vantaan Järjestörinki ry:n Maahanmuuttajien neuvontapiste ) kan du fråga om sådant som rör till exempel arbetslivet , social trygghet , hälsa , utbildning och uppehållstillstånd .
adress :
Ranunkelvägen 22
asukastila Myyrinki
Eldstadstorget 1 eller Kopparbergsvägen 10 B , vån .
Vanda Tfn ( 09 ) 839.35703 och 040.183.0930
Rautbergsgatan 3
tfn 045.134.1711
rådgivning för invandrarefinska
om du har flyttat till huvudstadsregionen nyligen , kan du vid International House Helsinki ( IHH ) få rådgivning och myndighetstjänster på ett och samma besök .
IHH - serviceställe för dig som flyttar till Finland engelska
inledande kartläggning
den inledande kartläggningen ( alkukartoitus ) hjälper dig att hitta lämpliga tjänster i din hemstad .
Vanda stad eller Nylands TE @-@ byrå ordnar en inledande kartläggning för varje ny invandrare i Vanda .
du har rätt att få en inledande kartläggning om
din hemkommun är Vanda
du har flyttat till Vanda från ett annat land eller en annan ort i Finland
någon inledande kartläggning inte har gjorts för dig tidigare
du har haft hemkommun i Finland i högst tre år .
i den inledande kartläggningen får du information om utbildning i finska eller svenska , arbetssökning , utbildning och tjänster i Vanda .
vid den inledande kartläggningen talas man vid med hjälp av tolk .
den inledande kartläggningen är avgiftsfri .
Begäran om inledande kartläggning
du kan begära en inledande kartläggning via e @-@ post eller så kan du boka en tid per telefon .
tfn 09.839.32622 , 09.839.27525 eller 09.839.31766
om du söker arbete , bör du anmäla dig till TE @-@ byrån .
TE @-@ byrån gör den inledande kartläggningen .
Läs mer om den inledande kartläggningen och integrationsplanen på InfoFinlands webbplats Integration i Finland
linkkiVanda stad :
inledande kartläggningfinska _ engelska
behöver du en tolk ?
om du måste sköta ärenden med myndigheter , men inte kan finska eller svenska och det inte heller finns något annat språk som både du och myndigheten talar , kan du använda en tolktjänst .
meddela alltid myndigheten i förväg om du behöver en tolk .
myndigheten bokar tolken och då får du tolkningstjänsten gratis .
om du själv bokar tolken och betalar kostnaderna , kan du anlita en tolk när som helst .
Läs mer : behöver du en tolk ?
linkkiVanda stad :
information om tolktjänsterfinska
linkkiFinlands översättar- och tolkförbund :
Sök tolk eller översättarefinska _ svenska _ engelska
rådgivning för och integration av invandrare
inledande kartläggning
behöver du en tolk ?
rådgivning för och integration av invandrare
Invandrartjänster
Vanda stads tjänster för invandrare omfattar
mottagningstjänster för invandrare
integrationstjänster
Vanda stads tjänster för invandrare ( Vantaan maahanmuuttajapalvelut ) ger dig information om integration , social- och hälsovårdstjänster och om stadens och olika organisationers tjänster .
du kan bli klient om du flyttat till Finland på grund av familjeband , är flykting , offer för människohandel eller har rätt till en inledande kartläggning .
tfn ( 09 ) 839.21074 och ( 09 ) 839.32042
linkkiVanda stad :
Invandrartjänsterfinska _ engelska
Verksamhetscentret Silkesporten ( Silkinportin toimintakeskus ) ger rådgivning för invandrare och där ordnas många slags aktiviteter .
dickursbyvägen 44 F , vån .
tfn ( 09 ) 839.23651
linkkiSilkesportens verksamhetscenter :
rådgivning och verksamhet för invandrarefinska _ engelska
Vandainfo ger dig information om såväl Vandas stads som statens tjänster .
Vandainfon finns i Dickursby , Korso och Myrbacka .
Adresserna är :
Dixi , Banvägen 11 , 2:a vån .
tfn ( 09 ) 839.22133
tfn ( 09 ) 839.22133
tfn ( 09 ) 839.22133
kontaktuppgifterna och öppettiderna hittar du på Vanda stads webbplats .
linkkiVanda stad :
Vandainfofinska _ svenska _ engelska
den internationella föreningen i Håkansböle ( Hakunilan kansainvälinen yhdistys ) har en rådgivningspunkt som betjänar invandrare i Håkansböle , Björkby och andra områden i Vanda , som vill ha information om till exempel studier , språkkurser , arbete , hobbyverksamhet , krissituationer eller juridiska frågor .
Sporrgränden 2 A , vån . 3 ( Håkansböle )
tfn ( 09 ) 272.2775 och 040.501.3199 .
linkkiInternationella föreningen i Håkansböle :
rådgivning för invandrarefinska _ engelska _ ryska _ somaliska _ arabiska
på invandrarrådgivningen vid föreningen Vantaan Järjestörinki ry ( Vantaan Järjestörinki ry:n Maahanmuuttajien neuvontapiste ) kan du fråga om sådant som rör till exempel arbetslivet , social trygghet , hälsa , utbildning och uppehållstillstånd .
adress :
Ranunkelvägen 22
asukastila Myyrinki
Eldstadstorget 1 eller Kopparbergsvägen 10 B , vån .
Vanda Tfn ( 09 ) 839.35703 och 040.183.0930
Rautbergsgatan 3
tfn 045.134.1711
rådgivning för invandrarefinska
om du har flyttat till huvudstadsregionen nyligen , kan du vid International House Helsinki ( IHH ) få rådgivning och myndighetstjänster på ett och samma besök .
IHH - serviceställe för dig som flyttar till Finland engelska
inledande kartläggning
den inledande kartläggningen ( alkukartoitus ) hjälper dig att hitta lämpliga tjänster i din hemstad .
Vanda stad eller Nylands TE @-@ byrå ordnar en inledande kartläggning för varje ny invandrare i Vanda .
du har rätt att få en inledande kartläggning om
din hemkommun är Vanda
du har flyttat till Vanda från ett annat land eller en annan ort i Finland
någon inledande kartläggning inte har gjorts för dig tidigare
du har haft hemkommun i Finland i högst tre år .
i den inledande kartläggningen får du information om utbildning i finska eller svenska , arbetssökning , utbildning och tjänster i Vanda .
vid den inledande kartläggningen talas man vid med hjälp av tolk .
den inledande kartläggningen är avgiftsfri .
Begäran om inledande kartläggning
du kan begära en inledande kartläggning via e @-@ post eller så kan du boka en tid per telefon .
tfn 09.839.32622 , 09.839.27525 eller 09.839.31766
om du söker arbete , bör du anmäla dig till TE @-@ byrån .
TE @-@ byrån gör den inledande kartläggningen .
Läs mer om den inledande kartläggningen och integrationsplanen på InfoFinlands webbplats Integration i Finland
linkkiVanda stad :
inledande kartläggningfinska _ engelska
behöver du en tolk ?
om du måste sköta ärenden med myndigheter , men inte kan finska eller svenska och det inte heller finns något annat språk som både du och myndigheten talar , kan du använda en tolktjänst .
meddela alltid myndigheten i förväg om du behöver en tolk .
myndigheten bokar tolken och då får du tolkningstjänsten gratis .
om du själv bokar tolken och betalar kostnaderna , kan du anlita en tolk när som helst .
Läs mer : behöver du en tolk ?
linkkiVanda stad :
information om tolktjänsterfinska
linkkiFinlands översättar- och tolkförbund :
Sök tolk eller översättarefinska _ svenska _ engelska
rådgivning för och integration av invandrare
inledande kartläggning
behöver du en tolk ?
rådgivning för och integration av invandrare
Invandrartjänster
Vanda stads tjänster för invandrare omfattar
mottagningstjänster för invandrare
integrationstjänster
Vanda stads tjänster för invandrare ( Vantaan maahanmuuttajapalvelut ) ger dig information om integration , social- och hälsovårdstjänster och om stadens och olika organisationers tjänster .
du kan bli klient om du flyttat till Finland på grund av familjeband , är flykting , offer för människohandel eller har rätt till en inledande kartläggning .
tfn ( 09 ) 839.21074 och ( 09 ) 839.32042
linkkiVanda stad :
Invandrartjänsterfinska _ engelska
Vandainfo ger dig information om såväl Vandas stads som statens tjänster .
Vandainfon finns i Dickursby , Korso och Myrbacka .
Adresserna är :
Dixi , Banvägen 11 , 2:a vån .
tfn ( 09 ) 839.22133
tfn ( 09 ) 839.22133
tfn ( 09 ) 839.22133
kontaktuppgifterna och öppettiderna hittar du på Vanda stads webbplats .
linkkiVanda stad :
Vandainfofinska _ svenska _ engelska
den internationella föreningen i Håkansböle ( Hakunilan kansainvälinen yhdistys ) har en rådgivningspunkt som betjänar invandrare i Håkansböle , Björkby och andra områden i Vanda , som vill ha information om till exempel studier , språkkurser , arbete , hobbyverksamhet , krissituationer eller juridiska frågor .
Sporrgränden 2 A , vån . 3 ( Håkansböle )
tfn ( 09 ) 272.2775 och 040.501.3199 .
linkkiInternationella föreningen i Håkansböle :
rådgivning för invandrarefinska _ engelska _ ryska _ somaliska _ arabiska
på invandrarrådgivningen vid föreningen Vantaan Järjestörinki ry ( Vantaan Järjestörinki ry:n Maahanmuuttajien neuvontapiste ) kan du fråga om sådant som rör till exempel arbetslivet , social trygghet , hälsa , utbildning och uppehållstillstånd .
adress :
Ranunkelvägen 22
asukastila Myyrinki
Eldstadstorget 1 eller Kopparbergsvägen 10 B , vån .
Vanda Tfn ( 09 ) 839.35703 och 040.183.0930
Rautbergsgatan 3
tfn 045.134.1711
rådgivning för invandrarefinska
om du har flyttat till huvudstadsregionen nyligen , kan du vid International House Helsinki ( IHH ) få rådgivning och myndighetstjänster på ett och samma besök .
IHH - serviceställe för dig som flyttar till Finland engelska
inledande kartläggning
den inledande kartläggningen ( alkukartoitus ) hjälper dig att hitta lämpliga tjänster i din hemstad .
Vanda stad eller Nylands TE @-@ byrå ordnar en inledande kartläggning för varje ny invandrare i Vanda .
du har rätt att få en inledande kartläggning om
din hemkommun är Vanda
du har flyttat till Vanda från ett annat land eller en annan ort i Finland
någon inledande kartläggning inte har gjorts för dig tidigare
du har haft hemkommun i Finland i högst tre år .
i den inledande kartläggningen får du information om utbildning i finska eller svenska , arbetssökning , utbildning och tjänster i Vanda .
vid den inledande kartläggningen talas man vid med hjälp av tolk .
den inledande kartläggningen är avgiftsfri .
Begäran om inledande kartläggning
du kan begära en inledande kartläggning via e @-@ post eller så kan du boka en tid per telefon .
tfn 09.839.32622 , 09.839.27525 eller 09.839.31766
om du söker arbete , bör du anmäla dig till TE @-@ byrån .
TE @-@ byrån gör den inledande kartläggningen .
Läs mer om den inledande kartläggningen och integrationsplanen på InfoFinlands webbplats Integration i Finland
linkkiVanda stad :
inledande kartläggningfinska _ engelska
behöver du en tolk ?
om du måste sköta ärenden med myndigheter , men inte kan finska eller svenska och det inte heller finns något annat språk som både du och myndigheten talar , kan du använda en tolktjänst .
meddela alltid myndigheten i förväg om du behöver en tolk .
myndigheten bokar tolken och då får du tolkningstjänsten gratis .
om du själv bokar tolken och betalar kostnaderna , kan du anlita en tolk när som helst .
Läs mer : behöver du en tolk ?
linkkiVanda stad :
information om tolktjänsterfinska
linkkiFinlands översättar- och tolkförbund :
Sök tolk eller översättarefinska _ svenska _ engelska
tillståndsärenden
på Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU @-@ medborgarens uppehållsrätt .
Migrationsverkets tjänsteställe i Helsingfors :
Göksgränd 3A
du kan också ansöka om många slags uppehållstillstånd och EU @-@ registrering på internet i tjänsten Enter Finland .
om du inte är van vid att använda en dator , fyll i en ansökan på papper och lämna in den på Migrationsverkets tjänsteställe .
Dät är alltid bra att boka en tid i förväg på tjänstestället .
du kan boka en tid på Migrationsverkets tidsbokningstjänst .
Observera att tjänstestället inte kan ge rådgivning om tillståndsärenden .
Läs mer : flytta till Finland .
linkkiEnterfinland.fi :
elektronisk ansökanfinska _ svenska _ engelska
elektronisk tidsbokningfinska _ svenska _ engelska
registrering som invånare
om du flyttar ditt stadigvarande boende till Vanda , ska du registrera dig som invånare i kommunen .
du kan registrera dig vid magistraten .
Albertsgatan 25
växel 029.55.39391
registrering av utlänningar 029.55.36.300
när du går till magistraten ska du ta med dig
legitimation ( till exempel pass )
uppehållstillstånd och uppehållskort ( om du behöver uppehållstillstånd i Finland )
registreringsintyget över uppehållsrätten ( oleskeluoikeuden rekisteröintitodistus ) om du är EU @-@ medborgare .
äktenskapsintyg
dina barns födelseattester .
Observera att utländska handlingar ska vara legaliserade .
du får mer information om att legalisera officiella handlingar vid magistraten eller beskickningen för ditt eget land i Finland .
Läs mer : registrering som invånare .
registrering av utlänningarfinska _ svenska _ engelska
om du har flyttat till huvudstadsregionen nyligen , kan du vid International House Helsinki ( IHH ) få rådgivning och myndighetstjänster på ett och samma besök .
du kan få :
kostnadsfri rådgivning och information kring att flytta på flera olika språk
en finländsk personbeteckning , registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1 @-@ intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare .
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket .
adress
Albertsgatan 25
IHH - serviceställe för dig som flyttar till Finland engelska
Webbappen IHH Service Advisor App engelska
tillståndsärenden
på Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU @-@ medborgarens uppehållsrätt .
Migrationsverkets tjänsteställe i Helsingfors :
Göksgränd 3A
du kan också ansöka om många slags uppehållstillstånd och EU @-@ registrering på internet i tjänsten Enter Finland .
om du inte är van vid att använda en dator , fyll i en ansökan på papper och lämna in den på Migrationsverkets tjänsteställe .
Dät är alltid bra att boka en tid i förväg på tjänstestället .
du kan boka en tid på Migrationsverkets tidsbokningstjänst .
Observera att tjänstestället inte kan ge rådgivning om tillståndsärenden .
Läs mer : flytta till Finland .
linkkiEnterfinland.fi :
elektronisk ansökanfinska _ svenska _ engelska
elektronisk tidsbokningfinska _ svenska _ engelska
registrering som invånare
om du flyttar ditt stadigvarande boende till Vanda , ska du registrera dig som invånare i kommunen .
du kan registrera dig vid magistraten .
Albertsgatan 25
växel 029.55.39391
registrering av utlänningar 029.55.36.300
när du går till magistraten ska du ta med dig
legitimation ( till exempel pass )
uppehållstillstånd och uppehållskort ( om du behöver uppehållstillstånd i Finland )
registreringsintyget över uppehållsrätten ( oleskeluoikeuden rekisteröintitodistus ) om du är EU @-@ medborgare .
äktenskapsintyg
dina barns födelseattester .
Observera att utländska handlingar ska vara legaliserade .
du får mer information om att legalisera officiella handlingar vid magistraten eller beskickningen för ditt eget land i Finland .
Läs mer : registrering som invånare .
registrering av utlänningarfinska _ svenska _ engelska
om du har flyttat till huvudstadsregionen nyligen , kan du vid International House Helsinki ( IHH ) få rådgivning och myndighetstjänster på ett och samma besök .
du kan få :
kostnadsfri rådgivning och information kring att flytta på flera olika språk
en finländsk personbeteckning , registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1 @-@ intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare .
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket .
adress
IHH - serviceställe för dig som flyttar till Finland engelska
Webbappen IHH Service Advisor App engelska
tillståndsärenden
på Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU @-@ medborgarens uppehållsrätt .
Migrationsverkets tjänsteställe i Helsingfors :
Göksgränd 3A
du kan också ansöka om många slags uppehållstillstånd och EU @-@ registrering på internet i tjänsten Enter Finland .
om du inte är van vid att använda en dator , fyll i en ansökan på papper och lämna in den på Migrationsverkets tjänsteställe .
Dät är alltid bra att boka en tid i förväg på tjänstestället .
du kan boka en tid på Migrationsverkets tidsbokningstjänst .
Observera att tjänstestället inte kan ge rådgivning om tillståndsärenden .
Läs mer : flytta till Finland .
linkkiEnterfinland.fi :
elektronisk ansökanfinska _ svenska _ engelska
elektronisk tidsbokningfinska _ svenska _ engelska
registrering som invånare
om du flyttar ditt stadigvarande boende till Vanda , ska du registrera dig som invånare i kommunen .
du kan registrera dig vid magistraten .
Albertsgatan 25
växel 029.55.39391
registrering av utlänningar 029.55.36.300
när du går till magistraten ska du ta med dig
legitimation ( till exempel pass )
uppehållstillstånd och uppehållskort ( om du behöver uppehållstillstånd i Finland )
registreringsintyget över uppehållsrätten ( oleskeluoikeuden rekisteröintitodistus ) om du är EU @-@ medborgare .
äktenskapsintyg
dina barns födelseattester .
Observera att utländska handlingar ska vara legaliserade .
du får mer information om att legalisera officiella handlingar vid magistraten eller beskickningen för ditt eget land i Finland .
Läs mer : registrering som invånare .
registrering av utlänningarfinska _ svenska _ engelska
om du har flyttat till huvudstadsregionen nyligen , kan du vid International House Helsinki ( IHH ) få rådgivning och myndighetstjänster på ett och samma besök .
du kan få :
kostnadsfri rådgivning och information kring att flytta på flera olika språk
en finländsk personbeteckning , registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1 @-@ intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare .
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket .
adress
IHH - serviceställe för dig som flyttar till Finland engelska
Webbappen IHH Service Advisor App engelska
trafik
beslutsfattande och påverkan
religion
grundläggande information
historia
trafik
kollektivtrafiken
Esbo och hela huvudstadsregionen har goda kollektivtrafikförbindelser .
i Esbo finns flera tåg- och metrostationer .
i staden finns flera busslinjer .
information och råd till resenärerfinska _ svenska _ engelska
Esbo tillhör samkommunen Helsingforsregionens trafik HRT ( HSL ) , som ordnar kollektivtrafiken i huvudstadsregionen .
du kan söka information om rutterna i reseplanerartjänsten ( Reittiopas ) .
tjänsten ger dig råd om olika kollektivtrafikförbindelser från ett ställe till ett annat .
Reseplanerarefinska _ svenska _ engelska _ ryska
i kollektivtrafiken kan du betala med kontanter eller resekort .
i närtågen måste du köpa biljetten i förväg .
mer information om resekorten och deras försäljningsställen i Esbo hittar du på HRT:s webbplats .
du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat .
Biljetter och priserfinska _ svenska _ engelska
att gå och cykla
om du vill gå eller cykla i Esbo kan du söka en lämplig rutt i reseplaneraren för cykling och gång .
Resplan för cycling och gångfinska _ svenska _ engelska _ ryska
Cykelkartor för Helsingfors , Vanda och Esbo delas ut vid samservicekontoren och idrottsverkens serviceställen .
Cykelkartorna är kostnadsfria .
Friluftskartafinska
bil och flyg
du kan parkera bilen på många järnvägsstationer och fortsätta färden med kollektivtrafiken .
Helsingfors @-@ Vanda flygplats ligger Esbos grannkommun Vanda .
Läs mer : trafik .
linkkiEsbo stad :
trafikfinska _ svenska _ engelska
linkkiEsbo stad :
Kartorfinska _ svenska _ engelska
beslutsfattande och påverkan
i Esbo beslutas ärenden av stadsfullmäktige .
i stadsfullmäktige sitter 75 ledamöter som representerar olika politiska grupper .
Fullmäktige väljs var fjärde år genom kommunalval .
invånarna i Esbo kan påverka beslutsfattandet och beredning av ärenden på många olika sätt .
du kan ge respons till beslutsfattarna och tjänstemännen till exempel via det elektroniska responssystemet .
du kan vara med i invånarverksamheten eller ta ett invånarinitiativ .
Läs mer om hur du kan påverka på Esbo stads webbplats .
i Esbo finns en delegation för mångkulturella frågor som utvecklar stadens mångkulturella politik .
i Esbo finns många politiska föreningar , invandrarföreningar och andra föreningar via vilka du också kan påverka beslutsfattandet .
Läs mer : beslutsfattande och påverkan
linkkiEsbo stad :
information om beslutsfattandefinska _ svenska _ engelska
linkkiEsbo stad :
information om påverkanfinska _ svenska _ engelska
linkkiEsbo stad :
elektroniskt responssystemfinska _ svenska _ engelska
linkkiEsbo stad :
mångkulturella ärendenfinska _ svenska _ engelska
religion
många religiösa samfund är verksamma i Esbo och Helsingfors .
via tjänsten Uskonnot Suomessa kan du söka information efter det religiösa samfundet och orten .
Läs mer : kulturer och religioner i Finland .
religiösa samfundfinska _ engelska
linkkiEsbo kyrkliga samfällighet :
evangelisk @-@ lutherska församlingarfinska _ svenska _ engelska
linkkiHelsingfors ortodoxa församling :
ortodoxa församlingenfinska _ ryska
grundläggande information
Esbo är en av huvudstadsregionens fyra kommuner .
det ligger bredvid Helsingfors , väster om staden .
Utöver dessa finns det flera mindre tätorter , landsbygd och skogar i Esbo .
Esbo har cirka 280.000 invånare .
de flesta invånarna är finskspråkiga .
ungefär 7 procent av invånarna är svenskspråkiga och 16 procent har andra modersmål .
Esbos areal är cirka 528 km2 , varav cirka 216 km2 är vatten .
linkkiEsbo stad :
information om Esbofinska _ svenska _ engelska
historia
Esboområdet var bebott redan för ungefär 8.000 år sedan .
då var södra Esbo fortfarande hav .
på 1200 @-@ talet flyttade många emigranter från Sverige till Esbo .
på 1400 @-@ talet blev Esbo en självständig socken med många byar .
i Esbo byggdes stora herrgårdar som hade stor betydelse för områdets utveckling .
när Finland blev en del av Ryssland blev Helsingfors huvudstad år 1812 .
även om Helsingfors växte snabbt , var Esbo ännu länge en fridfull landssocken .
Inflyttningen till Esbo blev livligare från och med 1940 @-@ talet .
år 1950 hade Esbo 25.000 invånare och 15 år senare redan 65.000 invånare .
Esbo blev en stad år 1972 .
linkkiEsbo stad :
historiafinska _ svenska
linkkiEsbo stad :
Museerfinska _ svenska _ engelska
trafik
beslutsfattande och påverkan
religion
grundläggande information
historia
trafik
kollektivtrafiken
Esbo och hela huvudstadsregionen har goda kollektivtrafikförbindelser .
i Esbo finns flera tåg- och metrostationer .
i staden finns flera busslinjer .
information och råd till resenärerfinska _ svenska _ engelska
Esbo tillhör samkommunen Helsingforsregionens trafik HRT ( HSL ) , som ordnar kollektivtrafiken i huvudstadsregionen .
du kan söka information om rutterna i reseplanerartjänsten ( Reittiopas ) .
tjänsten ger dig råd om olika kollektivtrafikförbindelser från ett ställe till ett annat .
Reseplanerarefinska _ svenska _ engelska _ ryska
i kollektivtrafiken kan du betala med kontanter eller resekort .
i närtågen måste du köpa biljetten i förväg .
mer information om resekorten och deras försäljningsställen i Esbo hittar du på HRT:s webbplats .
du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat .
Biljetter och priserfinska _ svenska _ engelska
att gå och cykla
om du vill gå eller cykla i Esbo kan du söka en lämplig rutt i reseplaneraren för cykling och gång .
Resplan för cycling och gångfinska _ svenska _ engelska _ ryska
Cykelkartor för Helsingfors , Vanda och Esbo delas ut vid samservicekontoren och idrottsverkens serviceställen .
Cykelkartorna är kostnadsfria .
Friluftskartafinska
bil och flyg
du kan parkera bilen på många järnvägsstationer och fortsätta färden med kollektivtrafiken .
Helsingfors @-@ Vanda flygplats ligger Esbos grannkommun Vanda .
Läs mer : trafik .
linkkiEsbo stad :
trafikfinska _ svenska _ engelska
linkkiEsbo stad :
Kartorfinska _ svenska _ engelska
beslutsfattande och påverkan
i Esbo beslutas ärenden av stadsfullmäktige .
i stadsfullmäktige sitter 75 ledamöter som representerar olika politiska grupper .
Fullmäktige väljs var fjärde år genom kommunalval .
invånarna i Esbo kan påverka beslutsfattandet och beredning av ärenden på många olika sätt .
du kan ge respons till beslutsfattarna och tjänstemännen till exempel via det elektroniska responssystemet .
du kan vara med i invånarverksamheten eller ta ett invånarinitiativ .
Läs mer om hur du kan påverka på Esbo stads webbplats .
i Esbo finns en delegation för mångkulturella frågor som utvecklar stadens mångkulturella politik .
i Esbo finns många politiska föreningar , invandrarföreningar och andra föreningar via vilka du också kan påverka beslutsfattandet .
Läs mer : beslutsfattande och påverkan
linkkiEsbo stad :
information om beslutsfattandefinska _ svenska _ engelska
linkkiEsbo stad :
information om påverkanfinska _ svenska _ engelska
linkkiEsbo stad :
elektroniskt responssystemfinska _ svenska _ engelska
linkkiEsbo stad :
mångkulturella ärendenfinska _ svenska _ engelska
religion
många religiösa samfund är verksamma i Esbo och Helsingfors .
via tjänsten Uskonnot Suomessa kan du söka information efter det religiösa samfundet och orten .
Läs mer : kulturer och religioner i Finland .
religiösa samfundfinska _ engelska
linkkiEsbo kyrkliga samfällighet :
evangelisk @-@ lutherska församlingarfinska _ svenska _ engelska
linkkiHelsingfors ortodoxa församling :
ortodoxa församlingenfinska _ ryska
grundläggande information
Esbo är en av huvudstadsregionens fyra kommuner .
det ligger bredvid Helsingfors , väster om staden .
Utöver dessa finns det flera mindre tätorter , landsbygd och skogar i Esbo .
Esbo har cirka 280.000 invånare .
de flesta invånarna är finskspråkiga .
ungefär 7 procent av invånarna är svenskspråkiga och 16 procent har andra modersmål .
Esbos areal är cirka 528 km2 , varav cirka 216 km2 är vatten .
linkkiEsbo stad :
information om Esbofinska _ svenska _ engelska
historia
Esboområdet var bebott redan för ungefär 8.000 år sedan .
då var södra Esbo fortfarande hav .
på 1200 @-@ talet flyttade många emigranter från Sverige till Esbo .
på 1400 @-@ talet blev Esbo en självständig socken med många byar .
i Esbo byggdes stora herrgårdar som hade stor betydelse för områdets utveckling .
när Finland blev en del av Ryssland blev Helsingfors huvudstad år 1812 .
även om Helsingfors växte snabbt , var Esbo ännu länge en fridfull landssocken .
Inflyttningen till Esbo blev livligare från och med 1940 @-@ talet .
år 1950 hade Esbo 25.000 invånare och 15 år senare redan 65.000 invånare .
Esbo blev en stad år 1972 .
linkkiEsbo stad :
historiafinska _ svenska
linkkiEsbo stad :
Museerfinska _ svenska _ engelska
trafik
beslutsfattande och påverkan
religion
grundläggande information
historia
trafik
kollektivtrafiken
Esbo och hela huvudstadsregionen har goda kollektivtrafikförbindelser .
i Esbo finns flera tåg- och metrostationer .
i staden finns flera busslinjer .
information och råd till resenärerfinska _ svenska _ engelska
Esbo tillhör samkommunen Helsingforsregionens trafik HRT ( HSL ) , som ordnar kollektivtrafiken i huvudstadsregionen .
du kan söka information om rutterna i reseplanerartjänsten ( Reittiopas ) .
tjänsten ger dig råd om olika kollektivtrafikförbindelser från ett ställe till ett annat .
Reseplanerarefinska _ svenska _ engelska
i kollektivtrafiken kan du betala med kontanter eller resekort .
i närtågen måste du köpa biljetten i förväg .
mer information om resekorten och deras försäljningsställen i Esbo hittar du på HRT:s webbplats .
du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat .
Biljetter och priserfinska _ svenska _ engelska
att gå och cykla
om du vill gå eller cykla i Esbo kan du söka en lämplig rutt i reseplaneraren för cykling och gång .
Resplan för cycling och gångfinska _ svenska _ engelska _ ryska
bil och flyg
du kan parkera bilen på många järnvägsstationer och fortsätta färden med kollektivtrafiken .
Helsingfors @-@ Vanda flygplats ligger Esbos grannkommun Vanda .
Läs mer : trafik .
linkkiEsbo stad :
trafikfinska _ svenska _ engelska
linkkiEsbo stad :
Kartorfinska _ svenska _ engelska
beslutsfattande och påverkan
i Esbo beslutas ärenden av stadsfullmäktige .
i stadsfullmäktige sitter 75 ledamöter som representerar olika politiska grupper .
Fullmäktige väljs var fjärde år genom kommunalval .
invånarna i Esbo kan påverka beslutsfattandet och beredning av ärenden på många olika sätt .
du kan ge respons till beslutsfattarna och tjänstemännen till exempel via det elektroniska responssystemet .
du kan vara med i invånarverksamheten eller ta ett invånarinitiativ .
Läs mer om hur du kan påverka på Esbo stads webbplats .
i Esbo finns en delegation för mångkulturella frågor som utvecklar stadens mångkulturella politik .
i Esbo finns många politiska föreningar , invandrarföreningar och andra föreningar via vilka du också kan påverka beslutsfattandet .
Läs mer : beslutsfattande och påverkan
linkkiEsbo stad :
information om beslutsfattandefinska _ svenska _ engelska
linkkiEsbo stad :
information om påverkanfinska _ svenska _ engelska
linkkiEsbo stad :
elektroniskt responssystemfinska _ svenska _ engelska
linkkiEsbo stad :
mångkulturella ärendenfinska _ svenska _ engelska
religion
många religiösa samfund är verksamma i Esbo och Helsingfors .
via tjänsten Uskonnot Suomessa kan du söka information efter det religiösa samfundet och orten .
Läs mer : kulturer och religioner i Finland .
religiösa samfundfinska _ engelska
linkkiEsbo kyrkliga samfällighet :
evangelisk @-@ lutherska församlingarfinska _ svenska _ engelska
linkkiHelsingfors ortodoxa församling :
ortodoxa församlingenfinska _ ryska
grundläggande information
Esbo är en av huvudstadsregionens fyra kommuner .
det ligger bredvid Helsingfors , väster om staden .
Utöver dessa finns det flera mindre tätorter , landsbygd och skogar i Esbo .
Esbo har cirka 280.000 invånare .
de flesta invånarna är finskspråkiga .
ungefär 7 procent av invånarna är svenskspråkiga och 16 procent har andra modersmål .
Esbos areal är cirka 528 km2 , varav cirka 216 km2 är vatten .
linkkiEsbo stad :
information om Esbofinska _ svenska _ engelska
historia
Esboområdet var bebott redan för ungefär 8.000 år sedan .
då var södra Esbo fortfarande hav .
på 1200 @-@ talet flyttade många emigranter från Sverige till Esbo .
på 1400 @-@ talet blev Esbo en självständig socken med många byar .
i Esbo byggdes stora herrgårdar som hade stor betydelse för områdets utveckling .
när Finland blev en del av Ryssland blev Helsingfors huvudstad år 1812 .
även om Helsingfors växte snabbt , var Esbo ännu länge en fridfull landssocken .
Inflyttningen till Esbo blev livligare från och med 1940 @-@ talet .
år 1950 hade Esbo 25.000 invånare och 15 år senare redan 65.000 invånare .
Esbo blev en stad år 1972 .
linkkiEsbo stad :
historiafinska _ svenska
linkkiEsbo stad :
Museerfinska _ svenska _ engelska
evenemang
bibliotek
motion
att röra sig i naturen
teater och film
museer
Fritidsverksamhet för barn och unga
föreningar
i Esbo finns många hobbymöjligheter .
invånarhusen Kivenkolo och Kylämaja är öppna för alla .
i invånarhusen kan områdets invånare vistas och samlas samt få anvisningar och råd .
Invånarhuset Kivenkolo
Sjöstöveln 1 A
linkkiEsbo stad :
Kivenkolo invånarhusfinska _ svenska _ engelska
Invånarhuset Kylämaja
Mattsgatan 7
linkkiEsbo stad :
Invånarhus Kylämajafinska
vid Esbo arbetarinstitut ( Espoon työväenopisto ) kan man till exempel skapa konst , handarbeten , laga mat , dansa eller idka motion .
där kan man även studera finska och andra språk .
linkkiEsbo stad :
Arbetarinstitutetfinska _ svenska _ engelska
i Esbo finns flera läroanstalter som ger grundundervisning i konstämnen speciellt för barn och unga .
olika konstarter är musik , bildkonst , dans , teater och cirkus .
linkkiEsbo stad :
konstundervisningfinska _ engelska .
Konsthuset Lilla Aurora ordnar kulturevenemang för barn .
linkkiEsbo stad :
kulturevenemang för barnfinska _ svenska _ engelska
Läs mer : Fritid .
evenemang
Evenemangfinska _ svenska _ engelska _ ryska _ kinesiska
linkkiEsbo stad :
Evenemangfinska
bibliotek
i Esbo finns flera bibliotek på olika håll i staden .
på biblioteket kan du låna böcker , tidningar , musik , filmer , spel och mycket annat .
biblioteken har böcker och annat material på flera olika språk .
i biblioteket kan du också använda dator .
ofta hålls också utställningar och evenemang på biblioteken .
linkkiEsbo stad :
Bibliotekfinska _ svenska _ engelska
Flerspråkiga biblioteket
Flerspråkiga biblioteket ligger i Böle i Helsingfors
här finns böcker , musik , tidningar och tidskrifter samt ljudböcker på flera olika språk .
du kan åka till Böle eller beställa material till ditt eget närbibliotek .
linkkiHelsingfors stadsbibliotek :
Flerspråkiga biblioteketfinska _ svenska _ engelska
huvudstadsregionens gemensamma bibliotekstjänstfinska _ svenska _ engelska _ somaliska _ persiska _ arabiska
Läs mer : bibliotek .
motion
i Esbo finns simhallar , flera idrottshallar , idrottsplaner och andra idrottsplatser för olika idrottsgrenar .
på motionsslingorna kan man springa på somrarna och åka skidor på vintrarna .
Läs mer : motion .
linkkiEsbo stad :
information om motionstjänsternafinska _ svenska _ engelska
linkkiEsbo stad :
Idrottsklubbarfinska _ svenska
att röra sig i naturen
i Esbo finns flera friluftsområden där man kan vandra i naturen .
till exempel Noux nationalpark ligger delvis på Esbos område .
linkkiEsbo stad :
Naturobjekt i Esbofinska _ svenska _ engelska
Webbsidorfinska _ svenska _ engelska _ ryska _ kinesiska
Hemstadsstigarfinska _ svenska _ engelska
i naturhuset Villa Elfvik ordnas utflykter , evenemang och utställningar .
naturhuset är öppet för alla och ligger vid sidan av Bredvikens naturskyddsområde .
linkkiVilla Elfvik :
Naturens husfinska _ svenska _ engelska
i Esbo finns motionsslingor och friluftsleder på olika håll i staden .
på vintern är många motionsslingor skidspår .
en del rutter är belysta .
linkkiEsbo stad :
Friluftslivfinska _ svenska _ engelska
linkkiEsbo stad :
friluftsområdenfinska _ svenska _ engelska
vid insjöarna och på havskusten finns många badstränder .
alla Esbobor får fritt fiska med metspö och pimpla .
om du använder andra fiskeredskap ska du ha ett fisketillstånd .
linkkiEsbo stad :
fiske och jaktfinska _ svenska _ engelska
Läs mer : att röra sig i naturen .
teater och film
i Esbo finns flera yrkes- och amatörteatrar .
i Esbo finns tre biografer .
mer information om filmerna hittar du på biografernas webbplatser .
Därtill ordnar Esbo stad filmvisningar .
Läs mer : teater och film .
linkkiFinnkino :
Filmerfinska _ engelska
Filmerfinska
Filmerfinska _ svenska _ engelska
linkkiEsbo stad :
Teatrar i Esbofinska _ svenska _ engelska
museer
i Esbo finns flera museer .
Esbo moderna konstmuseum EMMA är ett av Finlands största konstmuseer .
Läs mer : museer .
linkkiEsbo stad :
Museerfinska _ svenska _ engelska
linkkiEsbo stad :
Stadsmuseetfinska _ svenska _ engelska
linkkiEsbo stad :
museet för modern konst EMMAfinska _ svenska _ engelska _ ryska
Fritidsverksamhet för barn och unga
i Esbo finns flera läroanstalter som ger grundundervisning i konstämnen speciellt för barn och unga .
olika konstarter är musik , bildkonst , dans , teater och cirkuskonst .
i Esbo finns ungdomsgårdar med utbildade ledare som övervakar verksamheten .
ungdomsgårdarna är öppna för alla ungdomar i åldrarna 9 @-@ 17 .
på ungdomsgårdarna kan de unga vistas på fritiden .
där bedrivs det även hobbyklubbar och ordnas kurser och evenemang .
också föreningar och idrottsklubbar ordnar mycket verksamhet för ungdomar .
Läs mer : Fritidsverksamhet för barn och unga .
linkkiEsbo stad :
verksamhet för ungafinska _ svenska _ engelska
linkkiEsbo stad :
Ungdomsgårdarfinska _ svenska _ engelska
linkkiEsbo stad :
rådgivning för ungafinska _ svenska _ engelska
linkkiEsbo stad :
Idrottsklubbarfinska _ svenska
Hobbysökningfinska
föreningar
i Esbo finns många olika föreningar , till exempel kulturföreningar och idrottsklubbar .
Läs mer : föreningar .
linkkiEsbo stad :
Idrottsklubbarfinska _ svenska
Föreningsverksamhetfinska
linkkiEsbo stad :
föreningar för seniorerfinska _ svenska
evenemang
bibliotek
motion
att röra sig i naturen
teater och film
museer
Fritidsverksamhet för barn och unga
föreningar
i Esbo finns många hobbymöjligheter .
invånarhusen Kivenkolo och Kylämaja är öppna för alla .
i invånarhusen kan områdets invånare vistas och samlas samt få anvisningar och råd .
Invånarhuset Kivenkolo
Sjöstöveln 1 A
linkkiEsbo stad :
Kivenkolo invånarhusfinska _ svenska _ engelska
Invånarhuset Kylämaja
Mattsgatan 7
linkkiEsbo stad :
Invånarhus Kylämajafinska
vid Esbo arbetarinstitut ( Espoon työväenopisto ) kan man till exempel skapa konst , handarbeten , laga mat , dansa eller idka motion .
där kan man även studera finska och andra språk .
linkkiEsbo stad :
Arbetarinstitutetfinska _ svenska _ engelska
i Esbo finns flera läroanstalter som ger grundundervisning i konstämnen speciellt för barn och unga .
olika konstarter är musik , bildkonst , dans , teater och cirkus .
linkkiEsbo stad :
konstundervisningfinska _ engelska .
Konsthuset Lilla Aurora ordnar kulturevenemang för barn .
linkkiEsbo stad :
kulturevenemang för barnfinska _ svenska _ engelska
Läs mer : Fritid .
evenemang
Evenemangfinska _ svenska _ engelska _ ryska
linkkiEsbo stad :
Evenemangfinska
bibliotek
i Esbo finns flera bibliotek på olika håll i staden .
på biblioteket kan du låna böcker , tidningar , musik , filmer , spel och mycket annat .
biblioteken har böcker och annat material på flera olika språk .
i biblioteket kan du också använda dator .
ofta hålls också utställningar och evenemang på biblioteken .
linkkiEsbo stad :
Bibliotekfinska _ svenska _ engelska
Flerspråkiga biblioteket
Flerspråkiga biblioteket ligger i Böle i Helsingfors
här finns böcker , musik , tidningar och tidskrifter samt ljudböcker på flera olika språk .
du kan åka till Böle eller beställa material till ditt eget närbibliotek .
linkkiHelsingfors stadsbibliotek :
Flerspråkiga biblioteketfinska _ svenska _ engelska
huvudstadsregionens gemensamma bibliotekstjänstfinska _ svenska _ engelska _ somaliska _ persiska _ arabiska
Läs mer : bibliotek .
motion
i Esbo finns simhallar , flera idrottshallar , idrottsplaner och andra idrottsplatser för olika idrottsgrenar .
på motionsslingorna kan man springa på somrarna och åka skidor på vintrarna .
Läs mer : motion .
linkkiEsbo stad :
information om motionstjänsternafinska _ svenska _ engelska
linkkiEsbo stad :
Idrottsklubbarfinska _ svenska
att röra sig i naturen
i Esbo finns flera friluftsområden där man kan vandra i naturen .
till exempel Noux nationalpark ligger delvis på Esbos område .
linkkiEsbo stad :
Naturobjekt i Esbofinska _ svenska _ engelska
Webbsidorfinska _ svenska _ engelska _ ryska _ kinesiska
Hemstadsstigarfinska _ svenska _ engelska
i naturhuset Villa Elfvik ordnas utflykter , evenemang och utställningar .
naturhuset är öppet för alla och ligger vid sidan av Bredvikens naturskyddsområde .
linkkiVilla Elfvik :
Naturens husfinska _ svenska _ engelska
i Esbo finns motionsslingor och friluftsleder på olika håll i staden .
på vintern är många motionsslingor skidspår .
en del rutter är belysta .
linkkiEsbo stad :
Friluftslivfinska _ svenska _ engelska
linkkiEsbo stad :
friluftsområdenfinska _ svenska _ engelska
vid insjöarna och på havskusten finns många badstränder .
alla Esbobor får fritt fiska med metspö och pimpla .
om du använder andra fiskeredskap ska du ha ett fisketillstånd .
linkkiEsbo stad :
fiske och jaktfinska _ svenska _ engelska
Läs mer : att röra sig i naturen .
teater och film
i Esbo finns flera yrkes- och amatörteatrar .
i Esbo finns tre biografer .
mer information om filmerna hittar du på biografernas webbplatser .
Därtill ordnar Esbo stad filmvisningar .
Läs mer : teater och film .
linkkiFinnkino :
Filmerfinska _ engelska
Filmerfinska
Filmerfinska _ svenska _ engelska
linkkiEsbo stad :
Teatrar i Esbofinska _ svenska _ engelska
museer
i Esbo finns flera museer .
Esbo moderna konstmuseum EMMA är ett av Finlands största konstmuseer .
Läs mer : museer .
linkkiEsbo stad :
Museerfinska _ svenska _ engelska
linkkiEsbo stad :
Stadsmuseetfinska _ svenska _ engelska
linkkiEsbo stad :
museet för modern konst EMMAfinska _ svenska _ engelska _ ryska
Fritidsverksamhet för barn och unga
i Esbo finns flera läroanstalter som ger grundundervisning i konstämnen speciellt för barn och unga .
olika konstarter är musik , bildkonst , dans , teater och cirkuskonst .
i Esbo finns ungdomsgårdar med utbildade ledare som övervakar verksamheten .
ungdomsgårdarna är öppna för alla ungdomar i åldrarna 9 @-@ 17 .
på ungdomsgårdarna kan de unga vistas på fritiden .
där bedrivs det även hobbyklubbar och ordnas kurser och evenemang .
också föreningar och idrottsklubbar ordnar mycket verksamhet för ungdomar .
Läs mer : Fritidsverksamhet för barn och unga .
linkkiEsbo stad :
verksamhet för ungafinska _ svenska _ engelska
linkkiEsbo stad :
Ungdomsgårdarfinska _ svenska _ engelska
linkkiEsbo stad :
rådgivning för ungafinska _ svenska _ engelska
linkkiEsbo stad :
Idrottsklubbarfinska _ svenska
Hobbysökningfinska
föreningar
i Esbo finns många olika föreningar , till exempel kulturföreningar och idrottsklubbar .
Läs mer : föreningar .
linkkiEsbo stad :
Idrottsklubbarfinska _ svenska
Föreningsverksamhetfinska
linkkiEsbo stad :
föreningar för seniorerfinska _ svenska
evenemang
bibliotek
motion
att röra sig i naturen
teater och film
museer
Fritidsverksamhet för barn och unga
föreningar
i Esbo finns många hobbymöjligheter .
invånarhusen Kivenkolo och Kylämaja är öppna för alla .
i invånarhusen kan områdets invånare vistas och samlas samt få anvisningar och råd .
Invånarhuset Kivenkolo
Sjöstöveln 1 A
linkkiEsbo stad :
Kivenkolo invånarhusfinska _ svenska _ engelska
Invånarhuset Kylämaja
Mattsgatan 7
linkkiEsbo stad :
Invånarhus Kylämajafinska
vid Esbo arbetarinstitut ( Espoon työväenopisto ) kan man till exempel skapa konst , handarbeten , laga mat , dansa eller idka motion .
där kan man även studera finska och andra språk .
linkkiEsbo stad :
Arbetarinstitutetfinska _ svenska _ engelska
i Esbo finns flera läroanstalter som ger grundundervisning i konstämnen speciellt för barn och unga .
olika konstarter är musik , bildkonst , dans , teater och cirkus .
linkkiEsbo stad :
konstundervisningfinska _ engelska .
Konsthuset Lilla Aurora ordnar kulturevenemang för barn .
linkkiEsbo stad :
kulturevenemang för barnfinska _ svenska _ engelska
Läs mer : Fritid .
evenemang
Evenemangfinska _ svenska _ engelska _ ryska
linkkiEsbo stad :
Evenemangfinska
bibliotek
i Esbo finns flera bibliotek på olika håll i staden .
på biblioteket kan du låna böcker , tidningar , musik , filmer , spel och mycket annat .
biblioteken har böcker och annat material på flera olika språk .
i biblioteket kan du också använda dator .
ofta hålls också utställningar och evenemang på biblioteken .
linkkiEsbo stad :
Bibliotekfinska _ svenska _ engelska
Flerspråkiga biblioteket
Flerspråkiga biblioteket ligger i Böle i Helsingfors
här finns böcker , musik , tidningar och tidskrifter samt ljudböcker på flera olika språk .
du kan åka till Böle eller beställa material till ditt eget närbibliotek .
linkkiHelsingfors stadsbibliotek :
Flerspråkiga biblioteketfinska _ svenska _ engelska
huvudstadsregionens gemensamma bibliotekstjänstfinska _ svenska _ engelska _ somaliska _ persiska _ arabiska
Läs mer : bibliotek .
motion
i Esbo finns simhallar , flera idrottshallar , idrottsplaner och andra idrottsplatser för olika idrottsgrenar .
på motionsslingorna kan man springa på somrarna och åka skidor på vintrarna .
Läs mer : motion .
linkkiEsbo stad :
information om motionstjänsternafinska _ svenska _ engelska
linkkiEsbo stad :
Idrottsklubbarfinska _ svenska
att röra sig i naturen
i Esbo finns flera friluftsområden där man kan vandra i naturen .
till exempel Noux nationalpark ligger delvis på Esbos område .
linkkiEsbo stad :
Naturobjekt i Esbofinska _ svenska _ engelska
Webbsidorfinska _ svenska _ engelska _ ryska _ kinesiska
Hemstadsstigarfinska _ svenska _ engelska
i naturhuset Villa Elfvik ordnas utflykter , evenemang och utställningar .
naturhuset är öppet för alla och ligger vid sidan av Bredvikens naturskyddsområde .
linkkiVilla Elfvik :
Naturens husfinska _ svenska _ engelska
i Esbo finns motionsslingor och friluftsleder på olika håll i staden .
på vintern är många motionsslingor skidspår .
en del rutter är belysta .
linkkiEsbo stad :
Friluftslivfinska _ svenska _ engelska
linkkiEsbo stad :
friluftsområdenfinska _ svenska _ engelska
vid insjöarna och på havskusten finns många badstränder .
alla Esbobor får fritt fiska med metspö och pimpla .
om du använder andra fiskeredskap ska du ha ett fisketillstånd .
linkkiEsbo stad :
fiske och jaktfinska _ svenska _ engelska
Läs mer : att röra sig i naturen .
teater och film
i Esbo finns flera yrkes- och amatörteatrar .
i Esbo finns tre biografer .
mer information om filmerna hittar du på biografernas webbplatser .
Därtill ordnar Esbo stad filmvisningar .
Läs mer : teater och film .
linkkiFinnkino :
Filmerfinska _ engelska
Filmerfinska
Filmerfinska _ svenska _ engelska
linkkiEsbo stad :
Teatrar i Esbofinska _ svenska _ engelska
museer
i Esbo finns flera museer .
Esbo moderna konstmuseum EMMA är ett av Finlands största konstmuseer .
Läs mer : museer .
linkkiEsbo stad :
Museerfinska _ svenska _ engelska
linkkiEsbo stad :
Stadsmuseetfinska _ svenska _ engelska
linkkiEsbo stad :
museet för modern konst EMMAfinska _ svenska _ engelska _ ryska
Fritidsverksamhet för barn och unga
i Esbo finns flera läroanstalter som ger grundundervisning i konstämnen speciellt för barn och unga .
olika konstarter är musik , bildkonst , dans , teater och cirkuskonst .
i Esbo finns ungdomsgårdar med utbildade ledare som övervakar verksamheten .
ungdomsgårdarna är öppna för alla ungdomar i åldrarna 9 @-@ 17 .
på ungdomsgårdarna kan de unga vistas på fritiden .
där bedrivs det även hobbyklubbar och ordnas kurser och evenemang .
också föreningar och idrottsklubbar ordnar mycket verksamhet för ungdomar .
Läs mer : Fritidsverksamhet för barn och unga .
linkkiEsbo stad :
verksamhet för ungafinska _ svenska _ engelska
linkkiEsbo stad :
Ungdomsgårdarfinska _ svenska _ engelska
linkkiEsbo stad :
rådgivning för ungafinska _ svenska _ engelska
linkkiEsbo stad :
Idrottsklubbarfinska _ svenska
Hobbysökningfinska
föreningar
i Esbo finns många olika föreningar , till exempel kulturföreningar och idrottsklubbar .
Läs mer : föreningar .
linkkiEsbo stad :
Idrottsklubbarfinska _ svenska
Föreningsverksamhetfinska
linkkiEsbo stad :
föreningar för seniorerfinska _ svenska
problem med uppehållstillståndet
brott
behöver du en jurist ?
våld Problem i äktenskap eller parförhållande
barns och ungas problem
missbruksproblem
Dödsfall
ring nödnumret 112 om det är fråga om en nödsituation .
via nödnumret kan du tillkalla polis , ambulans eller brandkår .
ring inte nödnumret om det inte är en nödsituation .
Läs mer : nödsituationer
linkkiEsbo stad :
Jourmottagningarfinska _ svenska _ engelska
social- och krisjouren
social- och krisjouren ( sosiaali- ja kriisipäivystys ) hjälper dygnet runt om du eller din familj behöver hjälp i en akut krissituation .
Krisen kan till exempel ha med våld , parförhållandet eller barnens problem att göra .
du kan även kontakta social- och krisjouren om du har problem med din mentala hälsa , missbruksproblem eller om du råkat ut för en traumatisk händelse i livet .
social- och krisjouren
Jorvs sjukhus
Åbovägen 150
tfn ( 09 ) 816.42439
öppet varje dag dygnet runt .
linkkiEsbo stad :
social- och krisjourenfinska _ svenska _ engelska
föreningen för mental hälsa i Finland ( Suomen Mielenterveysseura ) har en krismottagning för invandrare .
Kontoret ligger i Böle i Helsingfors .
Krismottagningen ger dig hjälp och stöd i svåra situationer .
boka en tid per telefon på numret ( 09 ) 4135.0501 .
linkkiFöreningen för mental hälsa i Finland :
krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
problem med uppehållstillståndet
om du har problem eller oklarheter med uppehållstillståndet , ska du ta kontakt med migrationsverket .
Läs mer : problem med uppehållstillstånd
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
om du är flykting , asylsökande eller vistas i Finland av någon annan anledning kan du be om juridisk hjälp och rådgivning vid Flyktingrådgivningen rf .
Kontoret ligger i Helsingfors .
adress : Kaisaniemigatan 4 A
tfn 09.2313.9325
linkkiFlyktingrådgivningen r.f. :
rättshjälp till flyktingarfinska _ svenska _ engelska
brott
om du blir utsatt för ett brott , gör en brottsanmälan hos polisen .
du kan göra brottsanmälan på internet .
du kan även fylla i en blankett och lämna den till Esbo huvudpolisstation .
Esbo huvudpolisstation
Knektbrogränden 4
Läs mer : brott
kontaktuppgifterfinska _ svenska _ engelska
elektronisk polisanmälanfinska _ svenska _ engelska
behöver du en jurist ?
om du behöver juridisk hjälp , kan du kontakta Västra Nylands rättshjälpsbyrå .
Biskopsbron 9 B
tfn 029.56.61820
Läs mer : behöver du en jurist ?
linkkiVästra Nylands rättshjälpsbyrå :
rättshjälpfinska
våld
Omatila ( Omatila ) hjälper dig om du har blivit utsatt för närståendevåld eller våld inom familjen .
Omatila ordnar vid behov boende för dig och dina barn .
du kan ringa Omatila @-@ tjänsten dygnet runt . du behöver inte uppge ditt namn när du ringer .
du kan också komma utan tidsbokning för att prata om din situation , måndag till fredag kl . 9 @-@ 11 och onsdagar kl . 16 @-@ 20 .
Omatila
enheten för familjeärenden
Kamrersvägen 6 A
tfn 043.825.0535
Läs mer : våld
linkkiEsbo stad :
hjälp till offer för familjevåldfinska _ svenska _ engelska
Miehen Linja ( Miehen Linja ) är en tjänst som hjälper män , som har utsatt sina familjemedlemmar för våld . tjänsten är avsedd för invandrarmän .
Målargränden 3 B
tfn ( 09 ) 276.62899
hjälp för invandrarmänfinska _ engelska
problem i äktenskap eller parförhållande
om du har problem i ditt äktenskap eller parförhållande kan du kontakta familjerådgivningen .
familjerådgivningsbyråerna är i synnerhet avsedda för familjer med barn .
linkkiEsbo stad :
Familjerådgivningarfinska _ svenska _ engelska
Väestöliitto erbjuder rådgivning och terapi för par på finska och engelska .
linkkiBefolkningsförbundet :
rådgivning till invandrare telefonledes och via e @-@ postfinska _ svenska _ engelska
Familia Clubs projekt Duo erbjuder relationsrådgivning för par från två kulturer på finska och engelska .
rådgivningen är avgiftsbelagd .
relationsrådgivning för par från två kulturerfinska _ engelska
också kyrkans familjerådgivningscentral erbjuder familjerådgivning vid problem i parförhållandet .
kyrkans familjerådgivningfinska _ svenska _ engelska
Läs mer : problem i äktenskap och parförhållande
barns och ungas problem
hälsovårdaren vid barnrådgivningen ger råd i frågor som rör hälsan och utvecklingen av barn under skolåldern .
i Esbo finns flera rådgivningsbyråer runtom i staden .
rådgivningsbyråernas tidsbokning och rådgivning
tfn ( 09 ) 816.22800
linkkiEsbo stad :
rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
vid problem som berör barn i skolåldern hjälper till exempel skolans hälsovårdare .
linkkiEsbo stad :
information om hälsovården för skolbarnfinska _ svenska _ engelska
om du behöver råd i frågor kring barns psykiska utveckling , kan du boka en tid hos familjerådgivningen .
linkkiEsbo stad :
Familjerådgivningarfinska _ svenska _ engelska
Väestöliitto ger råd till invandrarfamiljer i frågor rörande barnfostran och familjens välmående .
rådgivningen på olika språk :
tfn 050.325.7173 ( ryska , engelska )
unga kan prata om sina problem med hälsovårdaren på den egna skolan eller läroanstalten .
det finns även andra ställen där man kan få hjälp .
en ung i åldern 13 @-@ 22 år kan få hjälp vid Ungdomspolikliniken Nupoli om hen har problem till exempel med den mentala hälsan , rusmedelsbruk , spelande eller fritidsaktiviteterna .
man kan ringa eller besöka Nupoli .
besök på Nupoli är kostnadsfria och konfidentiella .
tfn 09.816.31300
linkkiEsbo stad :
Nupoli - hjälp för ungafinska _ svenska
om den unga inte är trygg i sitt eget hem , kan hen kontakta Finlands Röda Kors De ungas skyddshus .
skyddshuset finns i Alberga .
de ungas skyddshus
tfn ( 09 ) 8195.5360
linkkiFinlands Röda Kors :
de ungas skyddshusfinska
Läs mer : barns och ungas problem
om du har ekonomiska problem kan du fråga om råd hos kommunens socialarbetare .
om du eller din familj inte har tillräckliga inkomster eller tillgångar för den nödvändiga dagliga försörjningen kan du söka grundläggande utkomststöd hos FPA .
information om utkomststödfinska _ svenska _ engelska _ ryska _ estniska
om du har problem med skulder , kontakta rättshjälpsbyråns ekonomi- och skuldrådgivning .
tjänsten är kostnadsfri .
linkkiRättshjälpsbyrå :
ekonomi- och skuldrådgivningfinska _ svenska _ engelska
missbruksproblem
kliniken för mental- och missbruksvård erbjuder vuxna Esbobor hjälp och vård vid problem med den mentala hälsan och missbruk .
Köpcentret Iso Omena
telefon : 09.816.31300
linkkiEsbo stad :
information om mentalvårdstjänsternafinska _ svenska _ engelska
unga i åldern 13 @-@ 22 med missbruksproblem kan få hjälp vid Ungdomspolikliniken Nupoli .
tfn 09.816.31300
linkkiEsbo stad :
Nupoli - hjälp för ungafinska _ svenska
Läs mer : missbruksproblem
Dödsfall
begravningsbyråer hjälper med de praktiska arrangemangen vid en begravning .
du kan söka begravningsbyråer till exempel på Finlands begravningsbyråers förbunds webbplats .
linkkiFinlands Begravningbyråers Förbund :
Begravningsbyråerfinska _ svenska _ engelska
i Esbo finns fem kristna begravningsplatser .
på Klockarmalmens begravningsplats finns ett gravområde för konfessionslösa .
där kan de avlidna begravas som hade en annan religionstillhörighet eller inte hörde till något religionssamfund .
linkkiEsbo församlingar :
Begravningsplatserfinska _ svenska _ engelska
om en närstående dör oväntat och du behöver stöd kan du kontakta social- och krisjouren i Esbo , telefon ( 09 ) 816.42439 .
Läs mer : Dödsfall
problem med uppehållstillståndet
brott
behöver du en jurist ?
våld Problem i äktenskap eller parförhållande
barns och ungas problem
missbruksproblem
Dödsfall
ring nödnumret 112 om det är fråga om en nödsituation .
via nödnumret kan du tillkalla polis , ambulans eller brandkår .
ring inte nödnumret om det inte är en nödsituation .
Läs mer : nödsituationer
linkkiEsbo stad :
Jourmottagningarfinska _ svenska _ engelska
social- och krisjouren
social- och krisjouren ( sosiaali- ja kriisipäivystys ) hjälper dygnet runt om du eller din familj behöver hjälp i en akut krissituation .
Krisen kan till exempel ha med våld , parförhållandet eller barnens problem att göra .
du kan även kontakta social- och krisjouren om du har problem med din mentala hälsa , missbruksproblem eller om du råkat ut för en traumatisk händelse i livet .
social- och krisjouren
Jorvs sjukhus
Åbovägen 150
tfn ( 09 ) 816.42439
öppet varje dag dygnet runt .
linkkiEsbo stad :
social- och krisjourenfinska _ svenska _ engelska
föreningen för mental hälsa i Finland ( Suomen Mielenterveysseura ) har en krismottagning för invandrare .
Kontoret ligger i Böle i Helsingfors .
Krismottagningen ger dig hjälp och stöd i svåra situationer .
boka en tid per telefon på numret ( 09 ) 4135.0501 .
linkkiFöreningen för mental hälsa i Finland :
krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
problem med uppehållstillståndet
om du har problem eller oklarheter med uppehållstillståndet , ska du ta kontakt med migrationsverket .
Läs mer : problem med uppehållstillstånd
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
om du är flykting , asylsökande eller vistas i Finland av någon annan anledning kan du be om juridisk hjälp och rådgivning vid Flyktingrådgivningen rf .
Kontoret ligger i Helsingfors .
adress : Kaisaniemigatan 4 A
tfn 09.2313.9325
linkkiFlyktingrådgivningen r.f. :
rättshjälp till flyktingarfinska _ svenska _ engelska
brott
om du blir utsatt för ett brott , gör en brottsanmälan hos polisen .
du kan göra brottsanmälan på internet .
du kan även fylla i en blankett och lämna den till Esbo huvudpolisstation .
Esbo huvudpolisstation
Knektbrogränden 4
Läs mer : brott
kontaktuppgifterfinska _ svenska _ engelska
elektronisk polisanmälanfinska _ svenska _ engelska
behöver du en jurist ?
om du behöver juridisk hjälp , kan du kontakta Västra Nylands rättshjälpsbyrå .
Biskopsbron 9 B
tfn 029.56.61820
Läs mer : behöver du en jurist ?
linkkiVästra Nylands rättshjälpsbyrå :
rättshjälpfinska
våld
Omatila ( Omatila ) hjälper dig om du har blivit utsatt för närståendevåld eller våld inom familjen .
Omatila ordnar vid behov boende för dig och dina barn .
du kan ringa Omatila @-@ tjänsten dygnet runt . du behöver inte uppge ditt namn när du ringer .
du kan också komma utan tidsbokning för att prata om din situation , måndag till fredag kl . 9 @-@ 11 och onsdagar kl . 16 @-@ 20 .
Omatila
enheten för familjeärenden
Kamrersvägen 6 A
tfn 043.825.0535
Läs mer : våld
linkkiEsbo stad :
hjälp till offer för familjevåldfinska _ svenska _ engelska
Miehen Linja ( Miehen Linja ) är en tjänst som hjälper män , som har utsatt sina familjemedlemmar för våld . tjänsten är avsedd för invandrarmän .
Målargränden 3 B
tfn ( 09 ) 276.62899
hjälp för invandrarmänfinska _ engelska
problem i äktenskap eller parförhållande
om du har problem i ditt äktenskap eller parförhållande kan du kontakta familjerådgivningen .
familjerådgivningsbyråerna är i synnerhet avsedda för familjer med barn .
linkkiEsbo stad :
Familjerådgivningarfinska _ svenska _ engelska
Väestöliitto erbjuder rådgivning och terapi för par på finska och engelska .
linkkiBefolkningsförbundet :
rådgivning till invandrare telefonledes och via e @-@ postfinska _ svenska _ engelska
Familia Clubs projekt Duo erbjuder relationsrådgivning för par från två kulturer på finska och engelska .
rådgivningen är avgiftsbelagd .
relationsrådgivning för par från två kulturerfinska _ engelska
också kyrkans familjerådgivningscentral erbjuder familjerådgivning vid problem i parförhållandet .
kyrkans familjerådgivningfinska _ svenska _ engelska
Läs mer : problem i äktenskap och parförhållande
barns och ungas problem
hälsovårdaren vid barnrådgivningen ger råd i frågor som rör hälsan och utvecklingen av barn under skolåldern .
i Esbo finns flera rådgivningsbyråer runtom i staden .
rådgivningsbyråernas tidsbokning och rådgivning
tfn ( 09 ) 816.22800
linkkiEsbo stad :
rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
vid problem som berör barn i skolåldern hjälper till exempel skolans hälsovårdare .
linkkiEsbo stad :
information om hälsovården för skolbarnfinska _ svenska _ engelska
om du behöver råd i frågor kring barns psykiska utveckling , kan du boka en tid hos familjerådgivningen .
linkkiEsbo stad :
Familjerådgivningarfinska _ svenska _ engelska
Väestöliitto ger råd till invandrarfamiljer i frågor rörande barnfostran och familjens välmående .
rådgivningen på olika språk :
tfn 050.325.7173 ( ryska , engelska )
unga kan prata om sina problem med hälsovårdaren på den egna skolan eller läroanstalten .
det finns även andra ställen där man kan få hjälp .
en ung i åldern 13 @-@ 22 år kan få hjälp vid Ungdomspolikliniken Nupoli om hen har problem till exempel med den mentala hälsan , rusmedelsbruk , spelande eller fritidsaktiviteterna .
man kan ringa eller besöka Nupoli .
besök på Nupoli är kostnadsfria och konfidentiella .
tfn 09.816.31300
linkkiEsbo stad :
Nupoli - hjälp för ungafinska _ svenska
om den unga inte är trygg i sitt eget hem , kan hen kontakta Finlands Röda Kors De ungas skyddshus .
skyddshuset finns i Alberga .
de ungas skyddshus
tfn ( 09 ) 8195.5360
linkkiFinlands Röda Kors :
de ungas skyddshusfinska
Läs mer : barns och ungas problem
om du har ekonomiska problem kan du fråga om råd hos kommunens socialarbetare .
om du eller din familj inte har tillräckliga inkomster eller tillgångar för den nödvändiga dagliga försörjningen kan du söka grundläggande utkomststöd hos FPA .
information om utkomststödfinska _ svenska _ engelska _ ryska _ estniska
om du har problem med skulder , kontakta rättshjälpsbyråns ekonomi- och skuldrådgivning .
tjänsten är kostnadsfri .
linkkiRättshjälpsbyrå :
ekonomi- och skuldrådgivningfinska _ svenska _ engelska
missbruksproblem
kliniken för mental- och missbruksvård erbjuder vuxna Esbobor hjälp och vård vid problem med den mentala hälsan och missbruk .
Köpcentret Iso Omena
telefon : 09.816.31300
linkkiEsbo stad :
information om mentalvårdstjänsternafinska _ svenska _ engelska
unga i åldern 13 @-@ 22 med missbruksproblem kan få hjälp vid Ungdomspolikliniken Nupoli .
tfn 09.816.31300
linkkiEsbo stad :
Nupoli - hjälp för ungafinska _ svenska
Läs mer : missbruksproblem
Dödsfall
begravningsbyråer hjälper med de praktiska arrangemangen vid en begravning .
du kan söka begravningsbyråer till exempel på Finlands begravningsbyråers förbunds webbplats .
linkkiFinlands Begravningbyråers Förbund :
Begravningsbyråerfinska
i Esbo finns fem kristna begravningsplatser .
på Klockarmalmens begravningsplats finns ett gravområde för konfessionslösa .
där kan de avlidna begravas som hade en annan religionstillhörighet eller inte hörde till något religionssamfund .
linkkiEsbo församlingar :
Begravningsplatserfinska _ svenska _ engelska
om en närstående dör oväntat och du behöver stöd kan du kontakta social- och krisjouren i Esbo , telefon ( 09 ) 816.42439 .
Läs mer : Dödsfall
problem med uppehållstillståndet
brott
behöver du en jurist ?
våld Problem i äktenskap eller parförhållande
barns och ungas problem
missbruksproblem
Dödsfall
ring nödnumret 112 om det är fråga om en nödsituation .
via nödnumret kan du tillkalla polis , ambulans eller brandkår .
ring inte nödnumret om det inte är en nödsituation .
Läs mer : nödsituationer
linkkiEsbo stad :
Jourmottagningarfinska _ svenska _ engelska
social- och krisjouren
social- och krisjouren ( sosiaali- ja kriisipäivystys ) hjälper dygnet runt om du eller din familj behöver hjälp i en akut krissituation .
Krisen kan till exempel ha med våld , parförhållandet eller barnens problem att göra .
du kan även kontakta social- och krisjouren om du har problem med din mentala hälsa , missbruksproblem eller om du råkat ut för en traumatisk händelse i livet .
social- och krisjouren
Jorvs sjukhus
Åbovägen 150
tfn ( 09 ) 816.42439
öppet varje dag dygnet runt .
linkkiEsbo stad :
social- och krisjourenfinska _ svenska _ engelska
föreningen för mental hälsa i Finland ( Suomen Mielenterveysseura ) har en krismottagning för invandrare .
Kontoret ligger i Böle i Helsingfors .
Krismottagningen ger dig hjälp och stöd i svåra situationer .
boka en tid per telefon på numret ( 09 ) 4135.0501 .
linkkiFöreningen för mental hälsa i Finland :
krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
problem med uppehållstillståndet
om du har problem eller oklarheter med uppehållstillståndet , ska du ta kontakt med migrationsverket .
Läs mer : problem med uppehållstillstånd
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
om du är flykting , asylsökande eller vistas i Finland av någon annan anledning kan du be om juridisk hjälp och rådgivning vid Flyktingrådgivningen rf .
Kontoret ligger i Helsingfors .
adress : Kaisaniemigatan 4 A
tfn 09.2313.9325
linkkiFlyktingrådgivningen r.f. :
rättshjälp till flyktingarfinska _ svenska _ engelska
brott
om du blir utsatt för ett brott , gör en brottsanmälan hos polisen .
du kan göra brottsanmälan på internet .
du kan även fylla i en blankett och lämna den till Esbo huvudpolisstation .
Esbo huvudpolisstation
Knektbrogränden 4
Läs mer : brott
kontaktuppgifterfinska _ svenska _ engelska
elektronisk polisanmälanfinska _ svenska _ engelska
behöver du en jurist ?
om du behöver juridisk hjälp , kan du kontakta Västra Nylands rättshjälpsbyrå .
Biskopsbron 9 B
tfn 029.56.61820
Läs mer : behöver du en jurist ?
linkkiVästra Nylands rättshjälpsbyrå :
rättshjälpfinska
våld
Omatila ( Omatila ) hjälper dig om du har blivit utsatt för närståendevåld eller våld inom familjen .
Omatila ordnar vid behov boende för dig och dina barn .
du kan ringa Omatila @-@ tjänsten dygnet runt . du behöver inte uppge ditt namn när du ringer .
du kan också komma utan tidsbokning för att prata om din situation , måndag till fredag kl . 9 @-@ 11 och onsdagar kl . 16 @-@ 20 .
Omatila
enheten för familjeärenden
Kamrersvägen 6 A
tfn 043.825.0535
Läs mer : våld
linkkiEsbo stad :
hjälp till offer för familjevåldfinska _ svenska _ engelska
Miehen Linja ( Miehen Linja ) är en tjänst som hjälper män , som har utsatt sina familjemedlemmar för våld . tjänsten är avsedd för invandrarmän .
Målargränden 3 B
tfn ( 09 ) 276.62899
hjälp för invandrarmänfinska _ engelska
problem i äktenskap eller parförhållande
om du har problem i ditt äktenskap eller parförhållande kan du kontakta familjerådgivningen .
familjerådgivningsbyråerna är i synnerhet avsedda för familjer med barn .
linkkiEsbo stad :
Familjerådgivningarfinska _ svenska _ engelska
Väestöliitto erbjuder rådgivning och terapi för par på finska och engelska .
linkkiBefolkningsförbundet :
rådgivning till invandrare telefonledes och via e @-@ postfinska _ svenska _ engelska
Familia Clubs projekt Duo erbjuder relationsrådgivning för par från två kulturer på finska och engelska .
rådgivningen är avgiftsbelagd .
relationsrådgivning för par från två kulturerfinska _ engelska
också kyrkans familjerådgivningscentral erbjuder familjerådgivning vid problem i parförhållandet .
kyrkans familjerådgivningfinska _ svenska _ engelska
Läs mer : problem i äktenskap och parförhållande
barns och ungas problem
hälsovårdaren vid barnrådgivningen ger råd i frågor som rör hälsan och utvecklingen av barn under skolåldern .
i Esbo finns flera rådgivningsbyråer runtom i staden .
rådgivningsbyråernas tidsbokning och rådgivning
tfn ( 09 ) 816.22800
linkkiEsbo stad :
rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
vid problem som berör barn i skolåldern hjälper till exempel skolans hälsovårdare .
linkkiEsbo stad :
information om hälsovården för skolbarnfinska _ svenska _ engelska
om du behöver råd i frågor kring barns psykiska utveckling , kan du boka en tid hos familjerådgivningen .
linkkiEsbo stad :
Familjerådgivningarfinska _ svenska _ engelska
Väestöliitto ger råd till invandrarfamiljer i frågor rörande barnfostran och familjens välmående .
rådgivningen på olika språk :
tfn 050.325.7173 ( ryska , engelska )
unga kan prata om sina problem med hälsovårdaren på den egna skolan eller läroanstalten .
det finns även andra ställen där man kan få hjälp .
en ung i åldern 13 @-@ 22 år kan få hjälp vid Ungdomspolikliniken Nupoli om hen har problem till exempel med den mentala hälsan , rusmedelsbruk , spelande eller fritidsaktiviteterna .
man kan ringa eller besöka Nupoli .
besök på Nupoli är kostnadsfria och konfidentiella .
tfn 09.816.31300
linkkiEsbo stad :
Nupoli - hjälp för ungafinska _ svenska
om den unga inte är trygg i sitt eget hem , kan hen kontakta Finlands Röda Kors De ungas skyddshus .
skyddshuset finns i Alberga .
de ungas skyddshus
tfn ( 09 ) 8195.5360
linkkiFinlands Röda Kors :
de ungas skyddshusfinska
Läs mer : barns och ungas problem
om du har ekonomiska problem kan du fråga om råd hos kommunens socialarbetare .
om du eller din familj inte har tillräckliga inkomster eller tillgångar för den nödvändiga dagliga försörjningen kan du söka grundläggande utkomststöd hos FPA .
information om utkomststödfinska _ svenska _ engelska _ ryska _ estniska
om du har problem med skulder , kontakta rättshjälpsbyråns ekonomi- och skuldrådgivning .
tjänsten är kostnadsfri .
linkkiRättshjälpsbyrå :
ekonomi- och skuldrådgivningfinska _ svenska _ engelska
missbruksproblem
kliniken för mental- och missbruksvård erbjuder vuxna Esbobor hjälp och vård vid problem med den mentala hälsan och missbruk .
Köpcentret Iso Omena
telefon : 09.816.31300
linkkiEsbo stad :
information om mentalvårdstjänsternafinska _ svenska _ engelska
unga i åldern 13 @-@ 22 med missbruksproblem kan få hjälp vid Ungdomspolikliniken Nupoli .
tfn 09.816.31300
linkkiEsbo stad :
Nupoli - hjälp för ungafinska _ svenska
Läs mer : missbruksproblem
Dödsfall
begravningsbyråer hjälper med de praktiska arrangemangen vid en begravning .
du kan söka begravningsbyråer till exempel på Finlands begravningsbyråers förbunds webbplats .
linkkiFinlands Begravningbyråers Förbund :
Begravningsbyråerfinska
i Esbo finns fem kristna begravningsplatser .
på Klockarmalmens begravningsplats finns ett gravområde för konfessionslösa .
där kan de avlidna begravas som hade en annan religionstillhörighet eller inte hörde till något religionssamfund .
linkkiEsbo församlingar :
Begravningsplatserfinska _ svenska _ engelska
om en närstående dör oväntat och du behöver stöd kan du kontakta social- och krisjouren i Esbo , telefon ( 09 ) 816.42439 .
Läs mer : Dödsfall
äktenskap
skilsmässa
Registrerat parförhållande
vård av barn Invånarparker och klubbar
problem i familjen
äktenskap
före äktenskapet ska du skriftligt begära hindersprövning ( avioliiton esteiden tutkiminen ) .
Hindersprövningen görs på magistraten ( maistraatti ) .
du kan begära hindersprövning på vilken magistrat som helst .
magistraten i Nyland , Esbo enhet
Miestentie 3
tfn 029.553.9391
Läs mer : äktenskap .
vigselfinska _ svenska _ engelska
Anhållan om prövning av hinder mot äktenskapfinska _ svenska
skilsmässa
kvinnan eller mannen kan lämna in skilsmässoansökan i Västra Nylands tingsrätts kansli .
du kan också söka skilsmässa ensam , utan din makes eller makas samtycke .
du kan skicka in ansökan till tingsrättens kansli per post , fax eller via e @-@ post .
tfn 029.564.4000
Läs mer : skilsmässa .
linkkiVästra Nylands tingsrätt :
kontaktuppgifterfinska _ svenska
barn vid skilsmässa
om du har barn under 13 år och överväger att skilja dig , ta kontakt med familjerådgivningen ( perheneuvola ) .
på familjerådgivningen kan du diskutera familjens situation med de anställda .
Familjerådgivningarnas kontaktuppgifter finns på Esbo stads webbplats .
om du planerar skilsmässa kan du också ta kontakt med barnatillsyningsmannen ( lastenvalvoja ) vid enheten för familjeärenden .
med barnatillsyningsmannen kan du diskutera skilsmässan och barnens framtid .
makarna ska ingå ett avtal om barnens boende , umgängesrätt och underhållsbidrag .
barnatillsyningsmännen bekräftar avtalet .
kontaktuppgifterna till barnatillsyningsmännen finns på Esbo stads webbplats .
Esbo stad har en rådgivningstelefon där man kan fråga om råd i frågor rörande barnen när föräldrarna skiljer sig .
tfn 046.877.3267
Läs mer : barn vid skilsmässa .
linkkiEsbo stad :
kontaktuppgifter till barnatillsyningsmännenfinska _ svenska
linkkiEsbo stad :
skilsmässa i en barnfamiljfinska _ svenska
vård av barn
information om dagvård av barn i Esbo finns på InfoFinlands sida Utbildning i Esbo .
tillfällig vård av barn
du kan föra barnet till en parktant för tillfällig vård .
det innebär kortvarig ( 2 @-@ 3 tim. per gång ) vård av småbarn ute i en lekpark .
du får närmare uppgifter av parktanterna per telefon .
du hittar telefonnumren på Esbo stads webbplats .
linkkiEsbo stad :
Parktanterfinska
om du behöver en tillfällig barnskötare hem , kan du kontakta Mannerheims Barnskyddsförbund eller Väestöliitto .
Barnavård och hemhjälpfinska
linkkiMannerheims Barnskyddsförbund :
Barnavårdfinska _ svenska _ engelska
Läs mer : dagvård .
hemvårdsstöd
om familjens yngsta barn är under tre år , kan barnets förälder få hemvårdsstöd ( kotihoidon tuki ) när han eller hon vårdar barnet i hemmet .
om du har rätt till hemvårdsstödet kan du ansöka om det hos FPA .
du kan fylla i ansökan på Internet eller posta den till FPA .
du kan också besöka FPA:s kontor .
Esbo stad betalar ett kommuntillägg till de familjer som vårdar ett under treårigt barn i hemmet .
man kan ansöka om Esbotillägget om en förälder tar hand om familjens alla barn under skolåldern i hemmet .
linkkiEsbo stad :
vård av barn i hemmetfinska _ svenska _ engelska
information om hemvårdsstödfinska _ svenska _ engelska
sköta ärenden på Internetfinska _ svenska _ engelska
kontaktuppgifter till FPAfinska _ svenska _ engelska
invånarparker och klubbar
Esbo stad ordnar mycket verksamhet för de föräldrar som vårdar barn i hemmet . det finns till exempel invånarparker , öppna daghem och klubbar .
Läs mer : stöd för vård av barn i hemmet
linkkiEsbo stad :
invånarparker och klubbarfinska _ engelska
problem i familjen
på InfoFinlands sida Problematiska situationer i Esbo hittar du uppgifter om vart du kan vända dig i Esbo för att få hjälp vid barns och ungas problem och problem i familjen .
du hittar uppgifter om barns och ungas problem också på InfoFinlands sida Barns och ungas problem och Var hittar jag hjälp när barn eller unga har problem ?
på InfoFinlands sida Problem i äktenskap och parförhållande finns uppgifter om vart du kan vända dig för att få hjälp vid problem i parförhållandet .
äktenskap
skilsmässa
Registrerat parförhållande
vård av barn Invånarparker och klubbar
problem i familjen
äktenskap
före äktenskapet ska du skriftligt begära hindersprövning ( avioliiton esteiden tutkiminen ) .
Hindersprövningen görs på magistraten ( maistraatti ) .
du kan begära hindersprövning på vilken magistrat som helst .
magistraten i Nyland , Esbo enhet
Miestentie 3
tfn 029.553.9391
Läs mer : äktenskap .
vigselfinska _ svenska _ engelska
Anhållan om prövning av hinder mot äktenskapfinska _ svenska
skilsmässa
kvinnan eller mannen kan lämna in skilsmässoansökan i Västra Nylands tingsrätts kansli .
du kan också söka skilsmässa ensam , utan din makes eller makas samtycke .
du kan skicka in ansökan till tingsrättens kansli per post , fax eller via e @-@ post .
tfn 029.564.4000
Läs mer : skilsmässa .
linkkiVästra Nylands tingsrätt :
kontaktuppgifterfinska _ svenska
barn vid skilsmässa
om du har barn under 13 år och överväger att skilja dig , ta kontakt med familjerådgivningen ( perheneuvola ) .
på familjerådgivningen kan du diskutera familjens situation med de anställda .
Familjerådgivningarnas kontaktuppgifter finns på Esbo stads webbplats .
om du planerar skilsmässa kan du också ta kontakt med barnatillsyningsmannen ( lastenvalvoja ) vid enheten för familjeärenden .
med barnatillsyningsmannen kan du diskutera skilsmässan och barnens framtid .
makarna ska ingå ett avtal om barnens boende , umgängesrätt och underhållsbidrag .
barnatillsyningsmännen bekräftar avtalet .
kontaktuppgifterna till barnatillsyningsmännen finns på Esbo stads webbplats .
Esbo stad har en rådgivningstelefon där man kan fråga om råd i frågor rörande barnen när föräldrarna skiljer sig .
tfn 046.877.3267
Läs mer : barn vid skilsmässa .
linkkiEsbo stad :
kontaktuppgifter till barnatillsyningsmännenfinska _ svenska
linkkiEsbo stad :
skilsmässa i en barnfamiljfinska _ svenska
vård av barn
information om dagvård av barn i Esbo finns på InfoFinlands sida Utbildning i Esbo .
tillfällig vård av barn
du kan föra barnet till en parktant för tillfällig vård .
det innebär kortvarig ( 2 @-@ 3 tim. per gång ) vård av småbarn ute i en lekpark .
du får närmare uppgifter av parktanterna per telefon .
du hittar telefonnumren på Esbo stads webbplats .
linkkiEsbo stad :
Parktanterfinska
om du behöver en tillfällig barnskötare hem , kan du kontakta Mannerheims Barnskyddsförbund eller Väestöliitto .
Barnavård och hemhjälpfinska
linkkiMannerheims Barnskyddsförbund :
Barnavårdfinska _ svenska _ engelska
Läs mer : dagvård .
hemvårdsstöd
om familjens yngsta barn är under tre år , kan barnets förälder få hemvårdsstöd ( kotihoidon tuki ) när han eller hon vårdar barnet i hemmet .
om du har rätt till hemvårdsstödet kan du ansöka om det hos FPA .
du kan fylla i ansökan på Internet eller posta den till FPA .
du kan också besöka FPA:s kontor .
Esbo stad betalar ett kommuntillägg till de familjer som vårdar ett under treårigt barn i hemmet .
man kan ansöka om Esbotillägget om en förälder tar hand om familjens alla barn under skolåldern i hemmet .
linkkiEsbo stad :
vård av barn i hemmetfinska _ svenska _ engelska
information om hemvårdsstödfinska _ svenska _ engelska
sköta ärenden på Internetfinska _ svenska _ engelska
kontaktuppgifter till FPAfinska _ svenska _ engelska
invånarparker och klubbar
Esbo stad ordnar mycket verksamhet för de föräldrar som vårdar barn i hemmet . det finns till exempel invånarparker , öppna daghem och klubbar .
Läs mer : stöd för vård av barn i hemmet
linkkiEsbo stad :
invånarparker och klubbarfinska _ engelska
äldre människor
åldringar kan använda tjänsterna vid de vanliga hälsostationerna .
dessutom erbjuds åldringar i Esbo egna tjänster , till exempel hemvårdens tjänster .
om du vill ha mer information om tjänster för äldre kan du kontakta seniorrådgivningen ( seniorineuvonta ) .
tfn ( 09 ) 816.33333
linkkiEsbo stad :
Seniorrådgivningenfinska _ svenska _ engelska
när du tar hand om en anhörig i hemmet
om du tar hand om en äldre , sjuk eller handikappad anhörig hemma så att hen ska kunna bo hemma , kan du ha rätt till stöd för närståendevård .
linkkiEsbo stad :
stöd för närståendevårdfinska _ svenska
äldre människor
problem i familjen
på InfoFinlands sida Problematiska situationer i Esbo hittar du uppgifter om vart du kan vända dig i Esbo för att få hjälp vid barns och ungas problem och problem i familjen .
du hittar uppgifter om barns och ungas problem också på InfoFinlands sida Barns och ungas problem och Var hittar jag hjälp när barn eller unga har problem ?
på InfoFinlands sida Problem i äktenskap och parförhållande finns uppgifter om vart du kan vända dig för att få hjälp vid problem i parförhållandet .
äktenskap
skilsmässa
Registrerat parförhållande
vård av barn Invånarparker och klubbar
problem i familjen
äktenskap
före äktenskapet ska du skriftligt begära hindersprövning ( avioliiton esteiden tutkiminen ) .
Hindersprövningen görs på magistraten ( maistraatti ) .
du kan begära hindersprövning på vilken magistrat som helst .
magistraten i Nyland , Esbo enhet
Miestentie 3
tfn 029.553.9391
Läs mer : äktenskap .
vigselfinska _ svenska _ engelska
Anhållan om prövning av hinder mot äktenskapfinska _ svenska
skilsmässa
kvinnan eller mannen kan lämna in skilsmässoansökan i Västra Nylands tingsrätts kansli .
du kan också söka skilsmässa ensam , utan din makes eller makas samtycke .
du kan skicka in ansökan till tingsrättens kansli per post , fax eller via e @-@ post .
tfn 029.564.4000
Läs mer : skilsmässa .
linkkiVästra Nylands tingsrätt :
kontaktuppgifterfinska _ svenska
barn vid skilsmässa
om du har barn under 13 år och överväger att skilja dig , ta kontakt med familjerådgivningen ( perheneuvola ) .
på familjerådgivningen kan du diskutera familjens situation med de anställda .
Familjerådgivningarnas kontaktuppgifter finns på Esbo stads webbplats .
om du planerar skilsmässa kan du också ta kontakt med barnatillsyningsmannen ( lastenvalvoja ) vid enheten för familjeärenden .
med barnatillsyningsmannen kan du diskutera skilsmässan och barnens framtid .
makarna ska ingå ett avtal om barnens boende , umgängesrätt och underhållsbidrag .
barnatillsyningsmännen bekräftar avtalet .
kontaktuppgifterna till barnatillsyningsmännen finns på Esbo stads webbplats .
Esbo stad har en rådgivningstelefon där man kan fråga om råd i frågor rörande barnen när föräldrarna skiljer sig .
tfn 046.877.3267
Läs mer : barn vid skilsmässa .
linkkiEsbo stad :
kontaktuppgifter till barnatillsyningsmännenfinska _ svenska
linkkiEsbo stad :
skilsmässa i en barnfamiljfinska _ svenska
vård av barn
information om dagvård av barn i Esbo finns på InfoFinlands sida Utbildning i Esbo .
tillfällig vård av barn
du kan föra barnet till en parktant för tillfällig vård .
det innebär kortvarig ( 2 @-@ 3 tim. per gång ) vård av småbarn ute i en lekpark .
du får närmare uppgifter av parktanterna per telefon .
du hittar telefonnumren på Esbo stads webbplats .
linkkiEsbo stad :
Parktanterfinska _ svenska
om du behöver en tillfällig barnskötare hem , kan du kontakta Mannerheims Barnskyddsförbund eller Väestöliitto .
Barnavård och hemhjälpfinska
linkkiMannerheims Barnskyddsförbund :
Barnavårdfinska _ svenska _ engelska
Läs mer : dagvård .
hemvårdsstöd
om familjens yngsta barn är under tre år , kan barnets förälder få hemvårdsstöd ( kotihoidon tuki ) när han eller hon vårdar barnet i hemmet .
om du har rätt till hemvårdsstödet kan du ansöka om det hos FPA .
du kan fylla i ansökan på Internet eller posta den till FPA .
du kan också besöka FPA:s kontor .
Esbo stad betalar ett kommuntillägg till de familjer som vårdar ett under treårigt barn i hemmet .
man kan ansöka om Esbotillägget om en förälder tar hand om familjens alla barn under skolåldern i hemmet .
linkkiEsbo stad :
vård av barn i hemmetfinska _ svenska _ engelska
information om hemvårdsstödfinska _ svenska _ engelska
sköta ärenden på Internetfinska _ svenska _ engelska
kontaktuppgifter till FPAfinska _ svenska _ engelska
invånarparker och klubbar
Esbo stad ordnar mycket verksamhet för de föräldrar som vårdar barn i hemmet . det finns till exempel invånarparker , öppna daghem och klubbar .
Läs mer : stöd för vård av barn i hemmet
linkkiEsbo stad :
invånarparker och klubbarfinska _ engelska
äldre människor
åldringar kan använda tjänsterna vid de vanliga hälsostationerna .
dessutom erbjuds åldringar i Esbo egna tjänster , till exempel hemvårdens tjänster .
om du vill ha mer information om tjänster för äldre kan du kontakta seniorrådgivningen ( seniorineuvonta ) .
tfn ( 09 ) 816.33333
linkkiEsbo stad :
Seniorrådgivningenfinska _ svenska _ engelska
när du tar hand om en anhörig i hemmet
om du tar hand om en äldre , sjuk eller handikappad anhörig hemma så att hen ska kunna bo hemma , kan du ha rätt till stöd för närståendevård .
linkkiEsbo stad :
stöd för närståendevårdfinska _ svenska
äldre människor
problem i familjen
på InfoFinlands sida Problematiska situationer i Esbo hittar du uppgifter om vart du kan vända dig i Esbo för att få hjälp vid barns och ungas problem och problem i familjen .
du hittar uppgifter om barns och ungas problem också på InfoFinlands sida Barns och ungas problem och Var hittar jag hjälp när barn eller unga har problem ?
på InfoFinlands sida Problem i äktenskap och parförhållande finns uppgifter om vart du kan vända dig för att få hjälp vid problem i parförhållandet .
hälsovårdstjänsterna i Esbo
äldre människors hälsa
tandvården
mental hälsa
sexuell hälsa
när du väntar barn
handikappade personer
ring nödnumret 112 om det är fråga om en brådskande nödsituation .
ring nödnumret till exempel vid en allvarlig olycka eller när någon drabbas av en sjukdomsattack .
ring inte nödnumret om det inte är en nödsituation .
om du har din hemkommun i Esbo kan du utnyttja de offentliga hälsovårdstjänsterna .
offentliga hälsovårdstjänster tillhandahålls vid hälsostationer , tandkliniker , rådgivningsbyråer och sjukhus .
om du inte har rätt till de offentliga hälsovårdstjänsterna , kan du söka hjälp på en privat läkarstation .
på en privat läkarstation måste du betala samtliga kostnader själv .
Läs mer : hälsa .
hälsovårdstjänsterna i Esbo
offentliga hälsovårdstjänster tillhandahålls av hälsostationerna ( terveysasema ) .
hälsostationerna har öppet vardagar klockan 8 @-@ 16 .
på hälsostationerna finns vanligtvis läkarens , sjukskötarens och hälsovårdarens mottagningar .
du kan boka tid på hälsostationen per telefon .
på Esbo stads webbplats finns kontaktuppgifterna och telefonnumren till hälsostationerna .
när du ringer hälsostationen , besvaras ditt samtal inte nödvändigtvis omedelbart .
ditt nummer sparas dock i en automat och du blir uppringd .
kom i tid till mottagningen .
om du inte kan komma till mottagningen , kom ihåg att avboka din tid senast föregående vardag före klockan 14 .
om du behöver första hjälpen snabbt , kan du komma till hälsostationen utan tidsbeställning .
linkkiEsbo stad :
Hälsostationernafinska _ svenska _ engelska
linkkiEsbo stad :
Hälsovårdscentralsavgifterfinska _ svenska
privata hälsovårdstjänster
Vem som helst kan gå till en privat hälsostation .
också de personer som inte har rätt till den offentliga hälsovården i Finland kan besöka privata hälsostationer .
på en privat hälsostation måste kunden själv betala samtliga kostnader .
i Esbo finns flera privata läkarstationer .
kontaktuppgifter till privata läkare hittar du till exempel på Internet .
linkkietsilaakari.fi :
privata hälsovårdstjänsterfinska
privat läkarstationfinska _ svenska _ engelska
privat läkarstationfinska _ svenska _ engelska
läkemedel
information om köp av läkemedel hittar du på InfoFinlands sida Läkemedel .
hälsovård för papperslösa
i Helsingfors finns Global Clinic , där personer som vistas i Finland utan tillstånd kan få primärhälsovård .
tjänsterna vid Global Clinic är avgiftsfria för kunderna .
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter .
för att skydda kunderna uppges inte klinikens adress eller öppettider offentligt .
telefonnumret till Global Clinic i Helsingfors är 044.977.4547 .
Samtalet besvaras av en sjukskötare eller en läkare .
hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Läs mer : hälsovårdstjänster i Finland
kvällstid och under veckoslut har hälsostationen stängt .
då vårdas akuta sjukfall och olycksfall på jourmottagningen ( päivystys ) .
den närmaste jourmottagningen för vuxna finns vid Jorv sjukhus .
ring den kostnadsfria Jourhjälpen på tfn 116.117 innan du kommer till jourmottagningen .
jourmottagningen vid Jorv sjukhus
Åbovägen 150
tfn ( 09 ) 4711
Jourmottagningar för barn under 16 år finns i Jorv och på Barnkliniken i Helsingfors .
du behöver inte boka tid på jourmottagningen .
linkkiEsbo stad :
Jourmottagningarfinska _ svenska _ engelska
Läs mer : hälsovårdstjänster i Finland
barns hälsa
i hälsovården av 1 @-@ 6 @-@ åriga barn får man hjälp av rådgivningsbyråns ( neuvola ) hälsovårdare och läkare .
dem kan du fråga om råd och få hjälp med fostran av barn .
på rådgivningsbyrån följs att barnet är friskt och växer som det ska .
i Esbo finns flera rådgivningsbyråer på olika håll i staden .
rådgivningsbyråernas kontaktuppgifter finns på Esbo stads webbplats .
du kan boka tid vid alla rådgivningsbyråer på samma nummer .
om ett barn blir sjukt och behöver snabbt vård , ta kontakt med hälsostationen ( terveysasema ) .
Skolhälsovårdaren har hand om skolbarns hälsa .
under kvällar och veckoslut finns jourmottagningen för barn under 16 år vid Jorv sjukhus och på Barnkliniken i Helsingfors .
du kan också ta ditt barn till en privat läkarstation .
Läs mer : barns hälsa .
linkkiEsbo stad :
Barnrådgivningsbyråernas tjänsterfinska _ svenska _ engelska
linkkiEsbo stad :
rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
linkkiEsbo stad :
Hälsostationernafinska _ svenska _ engelska
linkkiEsbo stad :
information om hälsovården för skolbarnfinska _ svenska _ engelska
linkkiEsbo stad :
Jourmottagningarfinska _ svenska _ engelska
äldre människors hälsa
åldringar kan använda tjänsterna vid de vanliga hälsostationerna .
dessutom erbjuds åldringar i Esbo egna tjänster , till exempel hemvårdens tjänster .
om du vill ha mer information om tjänster för äldre kan du kontakta seniorrådgivningen ( seniorineuvonta ) .
tfn ( 09 ) 816.33333
linkkiEsbo stad :
Seniorrådgivningenfinska _ svenska
när du tar hand om en anhörig i hemmet
om du tar hand om en äldre , sjuk eller handikappad anhörig hemma så att hen ska kunna bo hemma , kan du ha rätt till stöd för närståendevård .
linkkiEsbo stad :
stöd för närståendevårdfinska _ svenska
äldre människors hälsa , Äldre människor
tandvården
