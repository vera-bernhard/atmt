På InfoFinlands sida Avfallshantering och återvinning hittar du information om sopsortering.
linkkiHelsingforsregionens miljötjänster:
Sopsorteringsanvisningarfinska _ svenska _ engelska
linkkiHelsingforsregionens miljötjänster:
Återvinningsstationerfinska _ svenska _ engelska
Hyresbostad
Ägarbostad
Bostadsrättsbostad
Delägarbostad
Tillfälligt boende
Boende i en krissituation
Stöd- och serviceboende
Bostadslöshet
Avfallshantering och återvinning
Hyresbostad
I Esbo och huvudstadsregionen är hyrorna ofta högre än i resten av Finland.
Det kan vara svårt att hitta en bostad med lämplig hyra.
Det lönar sig att avsätta tid för bostadssökandet och undersöka olika alternativ.
Privata hyresbostäder
Hos en privat hyresvärd kan det gå snabbt att få en bostad, men hyran kan vara högre än i stadens hyresbostäder.
Du kan söka privata hyresbostäder i Esbo via hyresvärdarnas webbplatser:
Sökning av hyresbostäderfinska
Sökning av hyresbostäderfinska _ engelska
Hyresbostäder för ungafinska _ engelska
Hyresbostäder för ungafinska _ engelska
Om du är studerande kan du få en hyresbostad för studerande i Esbo.
Hyresbostäder för studerande erbjuds av Helsingforsregionens studentbostadsstiftelse HOAS och Aalto-universitets studentkår AUS.
linkkiHOAS:
Hyresbostäder för studerandefinska _ svenska _ engelska
Hyresbostäder för studerandefinska _ svenska _ engelska
Stadens hyresbostäder
Stadens hyresbostäder är ofta billigare än bostäder som man hyr av företag eller privatpersoner.
Det är dock många som ansöker om stadens bostäder och endast en liten del av de sökande får en bostad.
Störst är bristen på små bostäder.
Stadens hyresbostäder förvaltas av Espoon Asunnot Oy (Espoon Asunnot Oy).
Om du vill ansöka om en hyresbostad, fyll i en ansökningsblankett för hyresbostad på Espoon Asunnot Oy:s webbplats.
Du kan även fylla i ansökningsblanketten på Espoon Asunnot Oy:s kontor.
Du kan också få blanketten hemskickad per post.
Dina möjligheter att få en bostad påverkas av ditt bostadsbehov och dina tillgångar och inkomster.
För att kunna ansöka om en hyresbostad hos staden, måste du ha uppehållstillstånd för minst ett år.
Tfn (09) 816 5800
Ansökan är giltig i tre månader.
Efter det måste du förnya din ansökan om du fortfarande letar efter bostad.
Läs mer: Hyresbostad
linkkiEsbo Bostäder Ab:
Ansökan om hyresbostad i stadenfinska _ engelska
linkkiEsbo stad:
Stadens hyresbostäderfinska _ svenska _ engelska
linkkiEsbo stad:
Seniorbostäderfinska _ svenska
Ägarbostad
På internet finns många bostadsförsäljningsannonser.
Bostäderna i Esbo är tämligen dyra.
Information om köp av bostad hittar du på InfoFinlands sida Ägarbostad.
Bostadsrättsbostad
Om du ansöker om en bostadsrättsbostad, behöver du ett ordningsnummer. Du ansöker om ordningsnumret vid Esbo eller Helsingfors stad.
Läs mer: Bostadsrättsbostad.
linkkiEsbo stad:
Bostadsrättsbostäderfinska _ svenska _ engelska
Delägarbostad
Asuntosäätiö har delägarbostäder i Esbo.
Mer information hittar du på Asuntosäätiös webbplats.
Läs mer: Delägarbostad.
Delägarbostadfinska
Tillfälligt boende
I Esbo finns många olika hotell där man kan bo tillfälligt.
Läs mer: Tillfälligt boende.
linkkiVisitEspoo.fi:
Hotellfinska _ svenska _ engelska _ ryska
Brand eller vattenskada
Om din bostad har skadats till exempel till följd av brand eller vattenskada kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
Kontakta ditt försäkringsbolag direkt när skadan har inträffat.
Våld i hemmet
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta tjänsten Omatila (Omatila).
Omatila ordnar vid behov boende för dig och dina barn.
Omatila-tjänsten
Kamrersvägen 6 A
Tfn 043 825 0535
Öppet
Lördag-söndag kl. 9-16
Social- och krisjouren 24 h
Tfn 09 816 42439
linkkiEsbo stad:
Hjälp till offer för familjevåldfinska _ svenska _ engelska
Om du är ung och har problem hemma, kan du kontakta Finlands Röda Kors De ungas skyddshus.
Skyddshuset finns i Alberga.
De ungas skyddshus
Tfn (09) 8195 5360
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Stöd- och serviceboende
En del människor, till exempel åldringar och handikappade, har svårt att klara av de dagliga sysslorna utan hjälp.
Personer som har sin hemkommun i Esbo kan få hemvårdens stödtjänster av Esbo stad, till exempel måltidstjänster eller färdtjänst.
Dessa tjänster hjälper människorna att klara sig bättre hemma.
Åldringar och handikappade som inte klarar av att bo självständigt, kan bo i ett servicehus eller på en vårdinrättning.
Läs mer: Stöd- och serviceboende
Om du har frågor kring stödtjänsterna för handikappade, kontakta handikappservicen vid Esbo stad.
Esbo stads handikappservice
Telefonrådgivning: (09) 816 45285
linkkiEsbo stad:
Stödtjänster för handikappadefinska _ svenska _ engelska
Om du har frågor kring stödtjänsterna för äldre, kontakta Esbo stads rådgivning för seniorer.
Esbo stads rådgivning för seniorer
tfn (09) 816 33333
linkkiEsbo stad:
Stödtjänster för äldrefinska _ svenska _ engelska
linkkiEsbo stad:
Information om hemvårdens stödtjänsterfinska _ svenska
linkkiEsbo stad:
Information om boende i servicehusfinska _ svenska
Bostadslöshet
Om du blir bostadslös, kontakta Esbo stads verksamhetsställe för vuxensocialarbete.
linkkiEsbo stad:
Kontaktuppgifter till vuxensocialarbetetfinska _ svenska _ engelska
Om läget är akut, kan du även kontakta social- och krisjouren i Esbo.
Social- och krisjouren
Jorvs sjukhus
Åbovägen 150
Tfn (09) 816 42439
linkkiEsbo stad:
Social- och krisjourenfinska _ svenska _ engelska
Läs mer: Bostadslöshet
Avfallshantering och återvinning
På InfoFinlands sida Avfallshantering och återvinning hittar du information om sopsortering.
linkkiHelsingforsregionens miljötjänster:
Sopsorteringsanvisningarfinska _ svenska _ engelska
linkkiHelsingforsregionens miljötjänster:
Återvinningsstationerfinska _ svenska _ engelska
Hyresbostad
Ägarbostad
Bostadsrättsbostad
Delägarbostad
Tillfälligt boende
Boende i en krissituation
Stöd- och serviceboende
Bostadslöshet
Avfallshantering och återvinning
Hyresbostad
I Esbo och huvudstadsregionen är hyrorna ofta högre än i resten av Finland.
Det kan vara svårt att hitta en bostad med lämplig hyra.
Det lönar sig att avsätta tid för bostadssökandet och undersöka olika alternativ.
Privata hyresbostäder
Hos en privat hyresvärd kan det gå snabbt att få en bostad, men hyran kan vara högre än i stadens hyresbostäder.
Du kan söka privata hyresbostäder i Esbo via hyresvärdarnas webbplatser:
Sökning av hyresbostäderfinska
Sökning av hyresbostäderfinska _ engelska
Hyresbostäder för ungafinska _ engelska
Hyresbostäder för ungafinska _ engelska
Om du är studerande kan du få en hyresbostad för studerande i Esbo.
Hyresbostäder för studerande erbjuds av Helsingforsregionens studentbostadsstiftelse HOAS och Aalto-universitets studentkår AUS.
linkkiHOAS:
Hyresbostäder för studerandefinska _ svenska _ engelska
Hyresbostäder för studerandefinska _ svenska _ engelska
Stadens hyresbostäder
Stadens hyresbostäder är ofta billigare än bostäder som man hyr av företag eller privatpersoner.
Det är dock många som ansöker om stadens bostäder och endast en liten del av de sökande får en bostad.
Störst är bristen på små bostäder.
Stadens hyresbostäder förvaltas av Espoon Asunnot Oy (Espoon Asunnot Oy).
Om du vill ansöka om en hyresbostad, fyll i en ansökningsblankett för hyresbostad på Espoon Asunnot Oy:s webbplats.
Du kan även fylla i ansökningsblanketten på Espoon Asunnot Oy:s kontor.
Du kan också få blanketten hemskickad per post.
Dina möjligheter att få en bostad påverkas av ditt bostadsbehov och dina tillgångar och inkomster.
För att kunna ansöka om en hyresbostad hos staden, måste du ha uppehållstillstånd för minst ett år.
Tfn (09) 816 5800
Ansökan är giltig i tre månader.
Efter det måste du förnya din ansökan om du fortfarande letar efter bostad.
Läs mer: Hyresbostad
linkkiEsbo Bostäder Ab:
Ansökan om hyresbostad i stadenfinska _ engelska
linkkiEsbo stad:
Stadens hyresbostäderfinska _ svenska _ engelska
linkkiEsbo stad:
Seniorbostäderfinska _ svenska
Ägarbostad
På internet finns många bostadsförsäljningsannonser.
Bostäderna i Esbo är tämligen dyra.
Information om köp av bostad hittar du på InfoFinlands sida Ägarbostad.
Bostadsrättsbostad
Om du ansöker om en bostadsrättsbostad, behöver du ett ordningsnummer. Du ansöker om ordningsnumret vid Esbo eller Helsingfors stad.
Läs mer: Bostadsrättsbostad.
linkkiEsbo stad:
Bostadsrättsbostäderfinska _ svenska _ engelska
Delägarbostad
Asuntosäätiö har delägarbostäder i Esbo.
Mer information hittar du på Asuntosäätiös webbplats.
Läs mer: Delägarbostad.
Delägarbostadfinska
Tillfälligt boende
I Esbo finns många olika hotell där man kan bo tillfälligt.
Läs mer: Tillfälligt boende.
linkkiVisitEspoo.fi:
Hotellfinska _ svenska _ engelska _ ryska
Brand eller vattenskada
Om din bostad har skadats till exempel till följd av brand eller vattenskada kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
Kontakta ditt försäkringsbolag direkt när skadan har inträffat.
Våld i hemmet
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta tjänsten Omatila (Omatila).
Omatila ordnar vid behov boende för dig och dina barn.
Omatila-tjänsten
Kamrersvägen 6 A
Tfn 043 825 0535
Öppet
Lördag-söndag kl. 9-16
Social- och krisjouren 24 h
Tfn 09 816 42439
linkkiEsbo stad:
Hjälp till offer för familjevåldfinska _ svenska _ engelska
Om du är ung och har problem hemma, kan du kontakta Finlands Röda Kors De ungas skyddshus.
Skyddshuset finns i Alberga.
De ungas skyddshus
Tfn (09) 8195 5360
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Stöd- och serviceboende
En del människor, till exempel åldringar och handikappade, har svårt att klara av de dagliga sysslorna utan hjälp.
Personer som har sin hemkommun i Esbo kan få hemvårdens stödtjänster av Esbo stad, till exempel måltidstjänster eller färdtjänst.
Dessa tjänster hjälper människorna att klara sig bättre hemma.
Åldringar och handikappade som inte klarar av att bo självständigt, kan bo i ett servicehus eller på en vårdinrättning.
Läs mer: Stöd- och serviceboende
Om du har frågor kring stödtjänsterna för handikappade, kontakta handikappservicen vid Esbo stad.
Esbo stads handikappservice
Telefonrådgivning: (09) 816 45285
linkkiEsbo stad:
Stödtjänster för handikappadefinska _ svenska _ engelska
Om du har frågor kring stödtjänsterna för äldre, kontakta Esbo stads rådgivning för seniorer.
Esbo stads rådgivning för seniorer
tfn (09) 816 33333
linkkiEsbo stad:
Stödtjänster för äldrefinska _ svenska _ engelska
linkkiEsbo stad:
Information om hemvårdens stödtjänsterfinska _ svenska
linkkiEsbo stad:
Information om boende i servicehusfinska _ svenska
Bostadslöshet
Om du blir bostadslös, kontakta Esbo stads verksamhetsställe för vuxensocialarbete.
linkkiEsbo stad:
Kontaktuppgifter till vuxensocialarbetetfinska _ svenska _ engelska
Om läget är akut, kan du även kontakta social- och krisjouren i Esbo.
Social- och krisjouren
Jorvs sjukhus
Åbovägen 150
Tfn (09) 816 42439
linkkiEsbo stad:
Social- och krisjourenfinska _ svenska _ engelska
Läs mer: Bostadslöshet
Avfallshantering och återvinning
På InfoFinlands sida Avfallshantering och återvinning hittar du information om sopsortering.
linkkiHelsingforsregionens miljötjänster:
Sopsorteringsanvisningarfinska _ svenska _ engelska
linkkiHelsingforsregionens miljötjänster:
Återvinningsstationerfinska _ svenska _ engelska
Språkkurser
Med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors, Vanda, Esbo eller Grankulla.
I Esbo ordnas språkkurser i finska och svenska av Esbo arbetarinstitut, Esbo vuxengymnasium, Luksia och Axxell.
Kurser i finska och svenska språketfinska _ engelska _ ryska
Samtala på finska
På biblioteken i Esbo ordnas språkkaféer, där man kan öva sig i att prata finska.
På språkkaféerna samtalar man på finska, så det är bra om du redan kan lite finska.
Språkkaféerna är avgiftsfria.
Språkkaféer:
Entresse bibliotek, Iso Omena bibliotek, Stensvik bibliotek, Sello bibliotek och Hagalunds bibliotek.
Språkkaféerfinska _ engelska _ ryska
På den internationella träffpunkten Trapesa kan du delta i en samtals- och inlärningsgrupp på finska.
Gruppen är öppen för alla och den är avgiftsfri.
Diskussionsgrupp på finskafinska
Vi läser tillsammans för kvinnor
I Esbo finns även Vi läser tillsammans-grupper, där kvinnor kan studera finska språket.
linkkiVi läser tillsammans:
Finska för kvinnorfinska
Invånarlokalen i Kivenkolo
Man kan även träna sina finskakunskaper i invånarlokalen i Kivenkolo.
linkkiEsbo stad:
Kivenkolo invånarhusfinska _ svenska _ engelska
Om du är kund vid arbets- och näringsbyrån kan du fråga om språkkurser i finska och svenska vid arbets- och näringsbyrån.
Läs mer: Studier i finska och svenska
linkkiEsbo stad:
Kurser i finska och svenska språketfinska _ svenska _ engelska
linkkiEsbo stad:
Arbetarinstitutetfinska _ svenska _ engelska
linkkiEsbo stad:
Vuxengymnasietfinska
Kurser i finska och svenska språketfinska _ engelska
linkkiAxxell:
Kurser i finska och svenska språketfinska _ svenska
Allmän språkexamen
Du kan avlägga allmän språkexamen (yleinen kielitutkinto) i finska eller svenska i Esbo.
I Esbo ordnas språkexamina av Axxell och Esbo arbetarinstitut.
På utbildningsstyrelsens (opetushallitus) webbplats finns en sökmotor för språkexamina.
Med sökmotorn kan du kontrollera var och när du kan avlägga examen.
linkkiUtbildningsstyrelsen:
Examenssökningfinska
linkkiUtbildningsstyrelsen:
Allmänna språkexaminafinska _ svenska _ engelska
Språkkurser
Med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors, Vanda, Esbo eller Grankulla.
I Esbo ordnas språkkurser i finska och svenska av Esbo arbetarinstitut, Esbo vuxengymnasium, Luksia och Axxell.
Kurser i finska och svenska språketfinska _ engelska _ ryska
Samtala på finska
På biblioteken i Esbo ordnas språkkaféer, där man kan öva sig i att prata finska.
På språkkaféerna samtalar man på finska, så det är bra om du redan kan lite finska.
Språkkaféerna är avgiftsfria.
Språkkaféer:
Entresse bibliotek, Iso Omena bibliotek, Stensvik bibliotek, Sello bibliotek och Hagalunds bibliotek.
Språkkaféerfinska _ engelska _ ryska
På den internationella träffpunkten Trapesa kan du delta i en samtals- och inlärningsgrupp på finska.
Gruppen är öppen för alla och den är avgiftsfri.
Diskussionsgrupp på finskafinska
Vi läser tillsammans för kvinnor
I Esbo finns även Vi läser tillsammans-grupper, där kvinnor kan studera finska språket.
linkkiVi läser tillsammans:
Finska för kvinnorfinska
Invånarlokalen i Kivenkolo
Man kan även träna sina finskakunskaper i invånarlokalen i Kivenkolo.
linkkiEsbo stad:
Kivenkolo invånarhusfinska _ svenska _ engelska
Om du är kund vid arbets- och näringsbyrån kan du fråga om språkkurser i finska och svenska vid arbets- och näringsbyrån.
Läs mer: Studier i finska och svenska
linkkiEsbo stad:
Kurser i finska och svenska språketfinska _ svenska _ engelska
linkkiEsbo stad:
Arbetarinstitutetfinska _ svenska _ engelska
linkkiEsbo stad:
Vuxengymnasietfinska
Kurser i finska och svenska språketfinska _ engelska
linkkiAxxell:
Kurser i finska och svenska språketfinska _ svenska
Allmän språkexamen
Du kan avlägga allmän språkexamen (yleinen kielitutkinto) i finska eller svenska i Esbo.
I Esbo ordnas språkexamina av Axxell och Esbo arbetarinstitut.
På utbildningsstyrelsens (opetushallitus) webbplats finns en sökmotor för språkexamina.
Med sökmotorn kan du kontrollera var och när du kan avlägga examen.
linkkiUtbildningsstyrelsen:
Examenssökningfinska
linkkiUtbildningsstyrelsen:
Allmänna språkexaminafinska _ svenska _ engelska
Språkkurser
Med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors, Vanda, Esbo eller Grankulla.
I Esbo ordnas språkkurser i finska och svenska av Esbo arbetarinstitut, Esbo vuxengymnasium, Luksia och Axxell.
Kurser i finska och svenska språketfinska _ engelska _ ryska
Samtala på finska
På biblioteken i Esbo ordnas språkkaféer, där man kan öva sig i att prata finska.
På språkkaféerna samtalar man på finska, så det är bra om du redan kan lite finska.
Språkkaféerna är avgiftsfria.
Språkkaféer:
Entresse bibliotek, Iso Omena bibliotek, Stensvik bibliotek, Sello bibliotek och Hagalunds bibliotek.
Språkkaféerfinska _ engelska _ ryska
På den internationella träffpunkten Trapesa kan du delta i en samtals- och inlärningsgrupp på finska.
Gruppen är öppen för alla och den är avgiftsfri.
Diskussionsgrupp på finskafinska
Vi läser tillsammans för kvinnor
I Esbo finns även Vi läser tillsammans-grupper, där kvinnor kan studera finska språket.
linkkiVi läser tillsammans:
Finska för kvinnorfinska
Invånarlokalen i Kivenkolo
Man kan även träna sina finskakunskaper i invånarlokalen i Kivenkolo.
linkkiEsbo stad:
Kivenkolo invånarhusfinska _ svenska _ engelska
Om du är kund vid arbets- och näringsbyrån kan du fråga om språkkurser i finska och svenska vid arbets- och näringsbyrån.
Läs mer: Studier i finska och svenska
linkkiEsbo stad:
Kurser i finska och svenska språketfinska _ svenska _ engelska
linkkiEsbo stad:
Arbetarinstitutetfinska _ svenska _ engelska
linkkiEsbo stad:
Vuxengymnasietfinska
Kurser i finska och svenska språketfinska _ engelska
linkkiAxxell:
Kurser i finska och svenska språketfinska _ svenska
Allmän språkexamen
Du kan avlägga allmän språkexamen (yleinen kielitutkinto) i finska eller svenska i Esbo.
I Esbo ordnas språkexamina av Axxell och Esbo arbetarinstitut.
På utbildningsstyrelsens (opetushallitus) webbplats finns en sökmotor för språkexamina.
Med sökmotorn kan du kontrollera var och när du kan avlägga examen.
linkkiUtbildningsstyrelsen:
Examenssökningfinska
linkkiUtbildningsstyrelsen:
Allmänna språkexaminafinska _ svenska _ engelska
Var hittar jag jobb?
Hjälp med jobbsökningen
Att grunda ett företag
Beskattning
Var hittar jag jobb?
TE-byråns tjänster
Du kan få hjälp med jobbsökningen vid Nylands TE-byrå.
Verksamhetsstället i Esbo finns i Alberga.
linkkiArbets- och näringsministeriet:
Arbets- och näringsbyråerna i Nylandfinska _ svenska
TE-byrån betjänar på internet via sidan E-tjänster (Oma asiointi).
För att använda tjänsten behöver du nätbankskoder.
Medborgare i EU-länderna, Norge, Island, Liechtenstein och Schweiz kan anmäla sig som arbetssökande via TE-byråns E-tjänster.
Medborgare i andra länder måste anmäla sig personligen vid TE-byrån.
Ta med ett ID-kort och ditt uppehållstillstånd.
Information om TE-byråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös.
Information om jobbsökning i Finland hittar du på InfoFinlands sida Var hittar jag jobb?
linkkiTE-tjänster:
Anmälan utan nätbankskoderfinska _ svenska
linkkiArbets- och näringsministeriet:
Lediga jobbfinska _ svenska
linkkiArbets- och näringsförvaltningen:
Länkar till jobbsajterfinska _ svenska _ engelska
Lediga tjänster vid Esbo stad hittar du på stadens webbplats.
linkkiEsbo stad:
Arbetsplatser vid stadenfinska _ svenska _ engelska
Seure (Seure) är ett bemanningsbolag som erbjuder kortvariga jobb vid Helsingfors, Vanda, Esbo och Grankulla städer.
Jobben finns till exempel på skolor, daghem och sjukhus.
Arbetsplatser i kommunernafinska _ svenska
Hjälp med jobbsökningen
Råd om jobbsökningfinska _ svenska _ engelska _ spanska
Mentorskap i fråga om arbetskarriärfinska _ engelska
För unga under 30 år
linkkiEsbo stad:
Ohjaamofinska _ svenska _ engelska
Arbetslöshetsersättning
Information om att ansöka om arbetslöshetsersättning hittar du på InfoFinlands sida Arbetslöshetsförsäkring.
Att grunda ett företag
Om du vill grunda ett eget företag, kan du få hjälp vid FöretagsEsbo.
De hjälper dig att utveckla affärsidén och planera affärsverksamheten.
Tjänsterna är kostnadsfria.
linkkiFöretagsEsbo:
Företagsrådgivningfinska _ svenska _ engelska
Tjänster för företagarefinska _ svenska _ engelska
NewCo Yritys Helsinki erbjuder individuell rådgivning om grundande av företag samt ordnar informationsmöten och företagarutbildning på flera olika språk.
Tjänster för företagare med invandrarbakgrundfinska _ engelska
Guide om att grunda ett företagfinska _ engelska _ kinesiska
linkkiArbets- och näringsministeriet:
Tjänster för företagarefinska _ svenska _ engelska
Företagare i Esbo får även hjälp av Företagarna i Esbo rf.
Företagarna i Esbo rf är företagarnas egen organisation som erbjuder sina medlemmar till exempel utbildning, samarbete och rådgivning.
linkkiEsbo Företagare:
Företagarnas intressebevakningsorganisationfinska
Läs mer: Att grunda ett företag
Beskattning
Huvudstadsregionens skattebyrå ligger på Alexandersgatan 9 i Gloet i Helsingfors.
linkkiSkatteförvaltningen:
Kontaktuppgifter till skattebyråerfinska _ svenska _ engelska
Du kan även besöka servicestället In To Finland i Kampen i Helsingfors.
FPA:s och Skatteförvaltningens gemensamma rådgivning hjälper invandrare som har frågor om beskattningen eller den sociala tryggheten.
Här kan du hämta ett skattekort och ett inom byggbranschen obligatoriskt skattenummer.
Här kan dessutom utländska arbetstagare som ska arbeta i Finland tillfälligt få en finsk personbeteckning utan ett separat besök till magistraten.
Albertsgatan 25
Information om beskattningen hittar du på InfoFinlands sida Beskattning.
Var hittar jag jobb?
Hjälp med jobbsökningen
Att grunda ett företag
Beskattning
Var hittar jag jobb?
TE-byråns tjänster
Du kan få hjälp med jobbsökningen vid Nylands TE-byrå.
Verksamhetsstället i Esbo finns i Alberga.
linkkiArbets- och näringsministeriet:
Arbets- och näringsbyråerna i Nylandfinska _ svenska
TE-byrån betjänar på internet via sidan E-tjänster (Oma asiointi).
För att använda tjänsten behöver du nätbankskoder.
Medborgare i EU-länderna, Norge, Island, Liechtenstein och Schweiz kan anmäla sig som arbetssökande via TE-byråns E-tjänster.
Medborgare i andra länder måste anmäla sig personligen vid TE-byrån.
Ta med ett ID-kort och ditt uppehållstillstånd.
Information om TE-byråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös.
Information om jobbsökning i Finland hittar du på InfoFinlands sida Var hittar jag jobb?
linkkiTE-tjänster:
Anmälan utan nätbankskoderfinska _ svenska
linkkiArbets- och näringsministeriet:
Lediga jobbfinska _ svenska
linkkiArbets- och näringsförvaltningen:
Länkar till jobbsajterfinska _ svenska _ engelska
Lediga tjänster vid Esbo stad hittar du på stadens webbplats.
linkkiEsbo stad:
Arbetsplatser vid stadenfinska _ svenska _ engelska
Seure (Seure) är ett bemanningsbolag som erbjuder kortvariga jobb vid Helsingfors, Vanda, Esbo och Grankulla städer.
Jobben finns till exempel på skolor, daghem och sjukhus.
Arbetsplatser i kommunernafinska _ svenska
Hjälp med jobbsökningen
Råd om jobbsökningfinska _ svenska _ engelska _ spanska
Mentorskap i fråga om arbetskarriärfinska _ engelska
För unga under 30 år
linkkiEsbo stad:
Ohjaamofinska _ svenska _ engelska
Arbetslöshetsersättning
Information om att ansöka om arbetslöshetsersättning hittar du på InfoFinlands sida Arbetslöshetsförsäkring.
Att grunda ett företag
Om du vill grunda ett eget företag, kan du få hjälp vid FöretagsEsbo.
De hjälper dig att utveckla affärsidén och planera affärsverksamheten.
Tjänsterna är kostnadsfria.
linkkiFöretagsEsbo:
Företagsrådgivningfinska _ svenska _ engelska
Tjänster för företagarefinska _ svenska _ engelska
NewCo Yritys Helsinki erbjuder individuell rådgivning om grundande av företag samt ordnar informationsmöten och företagarutbildning på flera olika språk.
Tjänster för företagare med invandrarbakgrundfinska _ engelska
Guide om att grunda ett företagfinska _ engelska _ kinesiska
linkkiArbets- och näringsministeriet:
Tjänster för företagarefinska _ svenska _ engelska
Företagare i Esbo får även hjälp av Företagarna i Esbo rf.
Företagarna i Esbo rf är företagarnas egen organisation som erbjuder sina medlemmar till exempel utbildning, samarbete och rådgivning.
linkkiEsbo Företagare:
Företagarnas intressebevakningsorganisationfinska
Läs mer: Att grunda ett företag
Beskattning
Huvudstadsregionens skattebyrå ligger på Alexandersgatan 9 i Gloet i Helsingfors.
linkkiSkatteförvaltningen:
Kontaktuppgifter till skattebyråerfinska _ svenska _ engelska
Invandrare kan även sköta ärenden vid servicestället International House Helsinki.
På servicestället hjälper FPA:s och Skatteförvaltningens experter invandrare som kommer till Finland för att arbeta i frågor som rör beskattning och social trygghet.
Information om beskattningen hittar du på InfoFinlands sida Beskattning.
Var hittar jag jobb?
Hjälp med jobbsökningen
Att grunda ett företag
Beskattning
Var hittar jag jobb?
TE-byråns tjänster
Du kan få hjälp med jobbsökningen vid Nylands TE-byrå.
Verksamhetsstället i Esbo finns i Alberga.
linkkiArbets- och näringsministeriet:
Arbets- och näringsbyråerna i Nylandfinska _ svenska
TE-byrån betjänar på internet via sidan E-tjänster (Oma asiointi).
För att använda tjänsten behöver du nätbankskoder.
Medborgare i EU-länderna, Norge, Island, Liechtenstein och Schweiz kan anmäla sig som arbetssökande via TE-byråns E-tjänster.
Medborgare i andra länder måste anmäla sig personligen vid TE-byrån.
Ta med ett ID-kort och ditt uppehållstillstånd.
Information om TE-byråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös.
Information om jobbsökning i Finland hittar du på InfoFinlands sida Var hittar jag jobb?
linkkiTE-tjänster:
Anmälan utan nätbankskoderfinska _ svenska
linkkiArbets- och näringsministeriet:
Lediga jobbfinska _ svenska
linkkiArbets- och näringsförvaltningen:
Länkar till jobbsajterfinska _ svenska _ engelska
Lediga tjänster vid Esbo stad hittar du på stadens webbplats.
linkkiEsbo stad:
Arbetsplatser vid stadenfinska _ svenska _ engelska
Seure (Seure) är ett bemanningsbolag som erbjuder kortvariga jobb vid Helsingfors, Vanda, Esbo och Grankulla städer.
Jobben finns till exempel på skolor, daghem och sjukhus.
Arbetsplatser i kommunernafinska _ svenska _ engelska
Hjälp med jobbsökningen
Råd om jobbsökningfinska _ svenska _ engelska _ spanska
Mentorskap i fråga om arbetskarriärfinska _ engelska
För unga under 30 år
linkkiEsbo stad:
Ohjaamofinska _ svenska _ engelska
Arbetslöshetsersättning
Information om att ansöka om arbetslöshetsersättning hittar du på InfoFinlands sida Arbetslöshetsförsäkring.
Att grunda ett företag
Om du vill grunda ett eget företag, kan du få hjälp vid FöretagsEsbo.
De hjälper dig att utveckla affärsidén och planera affärsverksamheten.
Tjänsterna är kostnadsfria.
linkkiFöretagsEsbo:
Företagsrådgivningfinska _ svenska _ engelska
Tjänster för företagarefinska _ svenska _ engelska
NewCo Yritys Helsinki erbjuder individuell rådgivning om grundande av företag samt ordnar informationsmöten och företagarutbildning på flera olika språk.
Tjänster för företagare med invandrarbakgrundfinska _ engelska
Guide om att grunda ett företagfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ turkiska _ kinesiska _ arabiska
linkkiArbets- och näringsministeriet:
Tjänster för företagarefinska _ svenska _ engelska
Företagare i Esbo får även hjälp av Företagarna i Esbo rf.
Företagarna i Esbo rf är företagarnas egen organisation som erbjuder sina medlemmar till exempel utbildning, samarbete och rådgivning.
linkkiEsbo Företagare:
Företagarnas intressebevakningsorganisationfinska
Läs mer: Att grunda ett företag
Beskattning
Huvudstadsregionens skattebyrå ligger på Alexandersgatan 9 i Gloet i Helsingfors.
linkkiSkatteförvaltningen:
Kontaktuppgifter till skattebyråerfinska _ svenska _ engelska
Invandrare kan även sköta ärenden vid servicestället International House Helsinki.
På servicestället hjälper FPA:s och Skatteförvaltningens experter invandrare som kommer till Finland för att arbeta i frågor som rör beskattning och social trygghet.
Information om beskattningen hittar du på InfoFinlands sida Beskattning.
Rådgivning för och integration av invandrare
Inledande kartläggning och integrationsplan
Behöver du en tolk?
Rådgivning för och integration av invandrare
Servicepunkt
Vid Esbo stads servicepunkter (asiointipiste) får du mer information om stadens tjänster.
Servicepunkter finns på olika håll i staden.
Närmare kontaktuppgifter finns på Esbo stads webbplats.
Det gemensamma telefonnumret till servicepunkterna är (09) 816 57070 och e-postadressen är info(at)espoo.fi.
linkkiEsbo stad:
Servicepunktfinska _ svenska _ engelska
Kivenkolo
Invånarhuset Kivenkolo är ett öppet vardagsum där du kan få rådgivning och handledning på olika språk.
Kivenkolo
Sjöstöveln 1 A
Tfn 050 300 6093
linkkiEsbo stad:
Kivenkolo invånarhusfinska _ svenska _ engelska
Startpunkt för unga vuxna
Navigatorns Startpunkter erbjuder handledning och rådgivning utan tidsbokning till unga under 30 år.
Fågelbergavägen 2 A
Startpunkten i Iso Omena
linkkiEsbo stad:
Rådgivning för ungafinska _ svenska _ engelska
Den internationella mötesplatsen Trapesa erbjuder rådgivningstjänster.
Boka en tid i förväg.
Föreningen har även ett öppet vardagsrum, samtalsgrupper på finska och olika slags evenemang.
Stationsbron i Esbo
Tfn 010 583 7971
Invandrartjänster
Flyktingar kan även kontakta Esbo stads invandrartjänster (Maahanmuuttajapalvelut).
Vid servicerådgivningen får du råd och handledning utan tidsbeställning.
Rådgivningen ges på många olika språk.
Invandrartjänsterna
Fångstvägen 3
Tfn (09) 81621
linkkiEsbo stad:
Invandrartjänsterfinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
Du kan få:
kostnadsfri rådgivning och information kring att flytta på flera olika språk
en finländsk personbeteckning, registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1-intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
I tjänsten medverkar Helsingfors-info, magistraten i Nyland, skatteförvaltningens och FPA:s tjänst In To Finland, NTM-centralen i Nyland, Pensionsskyddscentralen och Helsingforsregionens handelskammare.
Adress
Albertsgatan 25
IHH – serviceställe för dig som flyttar till Finland engelska
Inledande kartläggning och integrationsplan
Inledande kartläggningar görs vid Esbo stads invandrartjänster eller enheten för vuxensocialarbete.
Invandrartjänsterna hjälper invandrare även i frågor som rör livet i Finland.
linkkiEsbo stad:
Invandrartjänsterfinska _ svenska _ engelska
linkkiEsbo stad:
Kontaktuppgifter till vuxensocialarbetetfinska _ svenska _ engelska
En anställd vid arbets- och näringsbyrån gör en inledande kartläggning tillsammans med dig, när du registrerar dig som arbetssökande.
Byrån i Esbo finns i Alberga.
Arbets- och näringsbyrån i Esbo
linkkiArbets- och näringsministeriet:
Arbets- och näringsbyråerna i Nylandfinska _ svenska
Behöver du en tolk?
Om du inte kan finska eller svenska kan du anlita en tolk när du sköter ärenden med myndigheter.
I vissa fall får du tolken via myndigheten.
Då är tolkningen kostnadsfri för dig.
Med myndigheter avses till exempel polisen, FPA, arbets- och näringsbyrån eller tjänstemän vid Esbo stad.
Myndigheten betalar dock inte alltid för en tolk.
Du ska alltså på förhand fråga om myndigheten betalar för tolktjänsterna.
Du kan använda en tolk när du vill, ifall du betalar och beställer tolken själv.
Du kan fråga om tolktjänsterna närmare till exempel vid Esbo stads invandrartjänster.
Läs mer: Behöver du en tolk?
linkkiEsbo stad:
Invandrartjänsterfinska _ svenska _ engelska
linkkiFinlands översättar- och tolkförbund:
Sök tolk eller översättarefinska _ svenska _ engelska
Rådgivning för och integration av invandrare
Inledande kartläggning och integrationsplan
Behöver du en tolk?
Rådgivning för och integration av invandrare
Servicepunkt
Vid Esbo stads servicepunkter (asiointipiste) får du mer information om stadens tjänster.
Servicepunkter finns på olika håll i staden.
Närmare kontaktuppgifter finns på Esbo stads webbplats.
Det gemensamma telefonnumret till servicepunkterna är (09) 816 57070 och e-postadressen är info(at)espoo.fi.
linkkiEsbo stad:
Servicepunktfinska _ svenska _ engelska
Kivenkolo
Invånarhuset Kivenkolo är ett öppet vardagsum där du kan få rådgivning och handledning på olika språk.
Kivenkolo
Sjöstöveln 1 A
Tfn 050 300 6093
linkkiEsbo stad:
Kivenkolo invånarhusfinska _ svenska _ engelska
Startpunkt för unga vuxna
Navigatorns Startpunkter erbjuder handledning och rådgivning utan tidsbokning till unga under 30 år.
Fågelbergavägen 2 A
Startpunkten i Iso Omena
linkkiEsbo stad:
Rådgivning för ungafinska _ svenska _ engelska
Den internationella mötesplatsen Trapesa erbjuder rådgivningstjänster.
Boka en tid i förväg.
Föreningen har även ett öppet vardagsrum, samtalsgrupper på finska och olika slags evenemang.
Stationsbron i Esbo
Tfn 010 583 7971
Invandrartjänster
Flyktingar kan även kontakta Esbo stads invandrartjänster (Maahanmuuttajapalvelut).
Vid servicerådgivningen får du råd och handledning utan tidsbeställning.
Rådgivningen ges på många olika språk.
Invandrartjänsterna
Fångstvägen 3
Tfn (09) 81621
linkkiEsbo stad:
Invandrartjänsterfinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
Du kan få:
kostnadsfri rådgivning och information kring att flytta på flera olika språk
en finländsk personbeteckning, registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1-intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
I tjänsten medverkar Helsingfors-info, magistraten i Nyland, skatteförvaltningens och FPA:s tjänst In To Finland, NTM-centralen i Nyland, Pensionsskyddscentralen och Helsingforsregionens handelskammare.
Adress
IHH – serviceställe för dig som flyttar till Finland engelska
Inledande kartläggning och integrationsplan
Inledande kartläggningar görs vid Esbo stads invandrartjänster eller enheten för vuxensocialarbete.
Invandrartjänsterna hjälper invandrare även i frågor som rör livet i Finland.
linkkiEsbo stad:
Invandrartjänsterfinska _ svenska _ engelska
linkkiEsbo stad:
Kontaktuppgifter till vuxensocialarbetetfinska _ svenska _ engelska
En anställd vid arbets- och näringsbyrån gör en inledande kartläggning tillsammans med dig, när du registrerar dig som arbetssökande.
Byrån i Esbo finns i Alberga.
Arbets- och näringsbyrån i Esbo
linkkiArbets- och näringsministeriet:
Arbets- och näringsbyråerna i Nylandfinska _ svenska
Behöver du en tolk?
Om du inte kan finska eller svenska kan du anlita en tolk när du sköter ärenden med myndigheter.
I vissa fall får du tolken via myndigheten.
Då är tolkningen kostnadsfri för dig.
Med myndigheter avses till exempel polisen, FPA, arbets- och näringsbyrån eller tjänstemän vid Esbo stad.
Myndigheten betalar dock inte alltid för en tolk.
Du ska alltså på förhand fråga om myndigheten betalar för tolktjänsterna.
Du kan använda en tolk när du vill, ifall du betalar och beställer tolken själv.
Du kan fråga om tolktjänsterna närmare till exempel vid Esbo stads invandrartjänster.
Läs mer: Behöver du en tolk?
linkkiEsbo stad:
Invandrartjänsterfinska _ svenska _ engelska
linkkiFinlands översättar- och tolkförbund:
Sök tolk eller översättarefinska _ svenska _ engelska
Rådgivning för och integration av invandrare
Inledande kartläggning och integrationsplan
Behöver du en tolk?
Rådgivning för och integration av invandrare
Servicepunkt
Vid Esbo stads servicepunkter (asiointipiste) får du mer information om stadens tjänster.
Servicepunkter finns på olika håll i staden.
Närmare kontaktuppgifter finns på Esbo stads webbplats.
Det gemensamma telefonnumret till servicepunkterna är (09) 816 57070 och e-postadressen är info(at)espoo.fi.
linkkiEsbo stad:
Servicepunktfinska _ svenska _ engelska
Kivenkolo
Invånarhuset Kivenkolo är ett öppet vardagsum där du kan få rådgivning och handledning på olika språk.
Kivenkolo
Sjöstöveln 1 A
Tfn 050 300 6093
linkkiEsbo stad:
Kivenkolo invånarhusfinska _ svenska _ engelska
Startpunkt för unga vuxna
Navigatorns Startpunkter erbjuder handledning och rådgivning utan tidsbokning till unga under 30 år.
Fågelbergavägen 2 A
Startpunkten i Iso Omena
linkkiEsbo stad:
Rådgivning för ungafinska _ svenska _ engelska
Den internationella mötesplatsen Trapesa erbjuder rådgivningstjänster.
Boka en tid i förväg.
Föreningen har även ett öppet vardagsrum, samtalsgrupper på finska och olika slags evenemang.
Stationsbron i Esbo
Tfn 010 583 7971
Invandrartjänster
Flyktingar kan även kontakta Esbo stads invandrartjänster (Maahanmuuttajapalvelut).
Vid servicerådgivningen får du råd och handledning utan tidsbeställning.
Rådgivningen ges på många olika språk.
Invandrartjänsterna
Fångstvägen 3
Tfn (09) 81621
linkkiEsbo stad:
Invandrartjänsterfinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
Du kan få:
kostnadsfri rådgivning och information kring att flytta på flera olika språk
en finländsk personbeteckning, registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1-intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
I tjänsten medverkar Helsingfors-info, Esbo stad, magistraten i Nyland, Migrationsverket, Skatteförvaltningen, FPA, NTM-centralen i Nyland, Pensionsskyddscentralen, Helsingforsregionens handelskammare och Finlands Fackförbunds Centralorganisation FFC.
Adress
IHH – serviceställe för dig som flyttar till Finland engelska
Inledande kartläggning och integrationsplan
Inledande kartläggningar görs vid Esbo stads invandrartjänster eller enheten för vuxensocialarbete.
Invandrartjänsterna hjälper invandrare även i frågor som rör livet i Finland.
linkkiEsbo stad:
Invandrartjänsterfinska _ svenska _ engelska
linkkiEsbo stad:
Kontaktuppgifter till vuxensocialarbetetfinska _ svenska _ engelska
En anställd vid arbets- och näringsbyrån gör en inledande kartläggning tillsammans med dig, när du registrerar dig som arbetssökande.
Byrån i Esbo finns i Alberga.
Arbets- och näringsbyrån i Esbo
linkkiArbets- och näringsministeriet:
Arbets- och näringsbyråerna i Nylandfinska _ svenska
Behöver du en tolk?
Om du inte kan finska eller svenska kan du anlita en tolk när du sköter ärenden med myndigheter.
I vissa fall får du tolken via myndigheten.
Då är tolkningen kostnadsfri för dig.
Med myndigheter avses till exempel polisen, FPA, arbets- och näringsbyrån eller tjänstemän vid Esbo stad.
Myndigheten betalar dock inte alltid för en tolk.
Du ska alltså på förhand fråga om myndigheten betalar för tolktjänsterna.
Du kan använda en tolk när du vill, ifall du betalar och beställer tolken själv.
Du kan fråga om tolktjänsterna närmare till exempel vid Esbo stads invandrartjänster.
Läs mer: Behöver du en tolk?
linkkiEsbo stad:
Invandrartjänsterfinska _ svenska _ engelska
linkkiFinlands översättar- och tolkförbund:
Sök tolk eller översättarefinska _ svenska _ engelska
Tillståndsärenden
På Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU-medborgarens uppehållsrätt.
Migrationsverkets tjänsteställe i Helsingfors :
Göksgränd 3A
Du kan också ansöka om många slags uppehållstillstånd och EU-registrering på internet i tjänsten Enter Finland.
Om du inte är van vid att använda en dator, fyll i en ansökan på papper och lämna in den på Migrationsverkets tjänsteställe.
Dät är alltid bra att boka en tid i förväg på tjänstestället.
Du kan boka en tid på Migrationsverkets tidsbokningstjänst.
Observera att tjänstestället inte kan ge rådgivning om tillståndsärenden.
Läs mer: Flytta till Finland.
Elektronisk tidsbokningfinska _ svenska _ engelska
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Registrering som invånare
Om du flyttar ditt stadigvarande boende till Esbo, ska du registrera dig som invånare i kommunen.
Du kan registrera dig vid magistraten i Nyland, Helsingfors enhet.
Magistraten i Nyland Helsingfors enhet
Albertsgatan 25
Tfn 029 55 39391
När du går till magistraten ska du ta med dig
legitimation (till exempel pass)
uppehållstillstånd och uppehållskort (om du behöver uppehållstillstånd i Finland)
registreringsintyget över uppehållsrätten (oleskeluoikeuden rekisteröintitodistus) om du är EU-medborgare.
äktenskapsintyg
dina barns födelseattester.
Observera att utländska handlingar ska vara legaliserade och översatta till finska, svenska eller engelska.
Du kan också ansöka om personbeteckning från magistraten.
Läs mer: Registrering som invånare, Hemkommun i Finland.
Registrering av utlänningarfinska _ svenska _ engelska
Kontaktuppgifter till magistratfinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
Du kan få:
kostnadsfri rådgivning och information kring att flytta på flera olika språk
en finländsk personbeteckning, registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1-intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
I tjänsten medverkar Helsingfors-info, magistraten i Nyland, skatteförvaltningens och FPA:s tjänst In To Finland, NTM-centralen i Nyland, Pensionsskyddscentralen och Helsingforsregionens handelskammare.
Adress
Albertsgatan 25
IHH – serviceställe för dig som flyttar till Finland engelska
Tillståndsärenden
På Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU-medborgarens uppehållsrätt.
Migrationsverkets tjänsteställe i Helsingfors :
Göksgränd 3A
Du kan också ansöka om många slags uppehållstillstånd och EU-registrering på internet i tjänsten Enter Finland.
Om du inte är van vid att använda en dator, fyll i en ansökan på papper och lämna in den på Migrationsverkets tjänsteställe.
Dät är alltid bra att boka en tid i förväg på tjänstestället.
Du kan boka en tid på Migrationsverkets tidsbokningstjänst.
Observera att tjänstestället inte kan ge rådgivning om tillståndsärenden.
Läs mer: Flytta till Finland.
Elektronisk tidsbokningfinska _ svenska _ engelska
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Registrering som invånare
Om du flyttar ditt stadigvarande boende till Esbo, ska du registrera dig som invånare i kommunen.
Du kan registrera dig vid magistraten i Nyland, Helsingfors enhet.
Magistraten i Nyland Helsingfors enhet
Tfn 029 55 39391
När du går till magistraten ska du ta med dig
legitimation (till exempel pass)
uppehållstillstånd och uppehållskort (om du behöver uppehållstillstånd i Finland)
registreringsintyget över uppehållsrätten (oleskeluoikeuden rekisteröintitodistus) om du är EU-medborgare.
äktenskapsintyg
dina barns födelseattester.
Observera att utländska handlingar ska vara legaliserade och översatta till finska, svenska eller engelska.
Du kan också ansöka om personbeteckning från magistraten.
Läs mer: Registrering som invånare, Hemkommun i Finland.
Registrering av utlänningarfinska _ svenska _ engelska
Kontaktuppgifter till magistratfinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
Du kan få:
kostnadsfri rådgivning och information kring att flytta på flera olika språk
en finländsk personbeteckning, registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1-intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
I tjänsten medverkar Helsingfors-info, magistraten i Nyland, skatteförvaltningens och FPA:s tjänst In To Finland, NTM-centralen i Nyland, Pensionsskyddscentralen och Helsingforsregionens handelskammare.
Adress
IHH – serviceställe för dig som flyttar till Finland engelska
Tillståndsärenden
På Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU-medborgarens uppehållsrätt.
Migrationsverkets tjänsteställe i Helsingfors :
Göksgränd 3A
Du kan också ansöka om många slags uppehållstillstånd och EU-registrering på internet i tjänsten Enter Finland.
Om du inte är van vid att använda en dator, fyll i en ansökan på papper och lämna in den på Migrationsverkets tjänsteställe.
Dät är alltid bra att boka en tid i förväg på tjänstestället.
Du kan boka en tid på Migrationsverkets tidsbokningstjänst.
Observera att tjänstestället inte kan ge rådgivning om tillståndsärenden.
Läs mer: Flytta till Finland.
Elektronisk tidsbokningfinska _ svenska _ engelska
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Registrering som invånare
Om du flyttar ditt stadigvarande boende till Esbo, ska du registrera dig som invånare i kommunen.
Du kan registrera dig vid magistraten i Nyland, Helsingfors enhet.
Magistraten i Nyland Helsingfors enhet
Tfn 029 55 39391
När du går till magistraten ska du ta med dig
legitimation (till exempel pass)
uppehållstillstånd och uppehållskort (om du behöver uppehållstillstånd i Finland)
registreringsintyget över uppehållsrätten (oleskeluoikeuden rekisteröintitodistus) om du är EU-medborgare.
äktenskapsintyg
dina barns födelseattester.
Observera att utländska handlingar ska vara legaliserade och översatta till finska, svenska eller engelska.
Du kan också ansöka om personbeteckning från magistraten.
Läs mer: Registrering som invånare, Hemkommun i Finland.
Registrering av utlänningarfinska _ svenska _ engelska
Kontaktuppgifter till magistratfinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
Du kan få:
kostnadsfri rådgivning och information kring att flytta på flera olika språk
en finländsk personbeteckning, registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1-intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
I tjänsten medverkar Helsingfors-info, magistraten i Nyland, skatteförvaltningens och FPA:s tjänst In To Finland, NTM-centralen i Nyland, Pensionsskyddscentralen och Helsingforsregionens handelskammare.
Adress
IHH – serviceställe för dig som flyttar till Finland engelska
Trafiken
Beslutsfattande och påverkan
Religion
Basfakta
Historia
Trafiken
Huvudstadsregionen har goda kollektivtrafikförbindelser.
I Helsingfors trafikerar tåg, bussar, spårvagnar, metron och Sveaborgsfärjorna.
Helsingfors är med i samkommunen Helsingforsregionens trafik (HRT) (Helsingin seudun liikenne -kuntayhtymä (HSL)) som sköter kollektivtrafiken i huvudstadsregionen.
I tjänsten Reseplaneraren (Reittiopas-palvelu) kan du söka information om kollektivtrafikens rutter i huvudstadsregionen.
Tjänsten ger dig förslag på olika kollektivtrafikförbindelser från ett ställe till ett annat.
I kollektivtrafikens färdmedel kan du betala med kontanter eller resekort (matkakortti).
Reseplanerarefinska _ svenska _ engelska _ ryska
Resekort
Med ett resekort (matkakortti) reser du förmånligare än med kontanter.
Resekortet gäller i lokaltrafikens bussar, närtågen, metron, spårvagnarna och Sveaborgsfärjorna.
Det finns två slags resekort.
Det är det billigaste sättet att resa.
Ett innehavarkort (haltijakohtainen kortti) kan användas av flera personer.
Innan du skaffar dig ett personligt kort ska du registrera dig som invånare i någon av kommunerna inom HRT-området.
Du kan köpa resekort vid HRT:s försäljningsställen (myyntipiste) eller serviceställen (palvelupiste).
De finns runtom i huvudstadsregionen.
Personligt resekort kan du köpa vid serviceställena.
Ta med dig identitetsbevis om du ska köpa personligt resekort.
Om du har finska nätbankskoder kan du även köpa personligt resekort på HRT:s webbplats.
Du kan resa med resekortet när du laddar kortet med period (kausi) eller värde (arvo).
En period betyder tid: till exempel en månad.
Värde betyder pengar.
Om du använder kollektivtrafiken ofta tjänar du på att ladda kortet med period.
Du kan ladda resekortet på vilket serviceställe för resekort (matkakortin latauspiste) som helst.
Du hittar mer information på HRT:s webbplats.
Ansökan om försäljningsplatserfinska _ svenska _ engelska
Information och råd till resenärerfinska _ svenska _ engelska
På cykel och till fots
I Helsingfors finns gott om cykelvägar.
I reseplaneraren för cykel- och gångtrafiken kan du söka en lämplig rutt om du vill gå eller cykla.
Bil och flyg
På många metrostationer kan du parkera din bil gratis för att fortsätta resan med kollektivtrafiken.
Helsingfors har goda landsvägsförbindelsermed resten av landet.
Den närmaste flygplatsen är Helsingfors-Vanda flygplats.
Läs mer: Trafiken.
Resplan för cycling och gångfinska _ svenska _ engelska _ ryska
linkkiVR:
Tågtidtabellerfinska _ svenska _ engelska _ ryska
Anslutningsparkeringfinska _ svenska _ engelska
Flygplatsenfinska _ svenska _ engelska _ ryska _ kinesiska
Beslutsfattande och påverkan
I Helsingfors beslutas ärenden av stadsfullmäktige.
Fullmäktigeledamöterna representerar olika politiska grupper.
Fullmäktige väljs vart fjärde år genom kommunalval.
Du kan följa fullmäktiges sammanträden och få mer information om beslutsfattandet på Helsingforskanalen eller på stadens webbplats.
Borgmästaren och stadens aktörer ordnar boendemöten runtom i Helsingfors för invånarna där man berättar om och diskuterar stadens ärenden.
Du kan även själv påverka beslutsfattande.
Att rösta i kommunalvalet är ett viktigt sätt att påverka.
Du kan även delta i utvecklingen av staden via olika slags elektroniska kanaler.
Till exempel på Helsingfors stads webbplats finns en färdig blankett, ett responssystem (palautejärjestelmä).
Via den kan du skicka frågor och förslag eller respons till staden.
I ditt bostadsområde arbetar dessutom stadens kontaktperson, stadslotsen (stadiluotsi), som kan hjälpa dig att föra vidare ditt förslag.
Stadslotsen har jour i områdets bibliotek vissa veckodagar och klockslag.
Mer information om stadslotsar och kontaktuppgifterna till dem hittar du på Helsingfors stads webbplats.
Stadsfullmäktigefinska _ svenska _ engelska
Stadsfullmäktiges sammanträden på Internetfinska _ svenska
Feedback till stadens ämbetsverk och inrättningarfinska _ svenska _ engelska
Delta och påverkafinska _ svenska _ engelska
Religion
I Helsingfors och Helsingforsregionen verkar många religiösa samfund.
I Helsingfors finns många olika religionssamfunds tempel och dessutom olika verksamhetscenter.
Via tjänsten Religionerna i Finland kan du söka information enligt religionssamfund och ort.
Läs mer: Kulturer och religioner i Finland.
Religiösa samfundfinska _ engelska
Basfakta
