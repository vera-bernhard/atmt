��&      ]�(�numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i4�����R�(K�<�NNNJ����J����K t�b�CTT                        Y           �     �
  '                 �t�bhhK ��h��R�(KK!��h�C��   �  D  '       �                           /                                             "        �t�bhhK ��h��R�(KK;��h�C�T      %   �     �              �     %                     �     
                 t           �     �   �     u  �         C   1
  �     %      �	  [        �        �     A           �t�bhhK ��h��R�(KK��h�C`      ^           �               T      �       "        #     �  r   "     �t�bhhK ��h��R�(KK��h�C`�   J   �  �  �  �      `            %      �
           �   J      `            �t�bhhK ��h��R�(KK��h�CP%      �
     �     %      �
     �         <     �      �         �t�bhhK ��h��R�(KK$��h�C�   �            �         C                               2                                �      7   g   7         �t�bhhK ��h��R�(KK��h�CHT      %      �                           G
              �t�bhhK ��h��R�(KK��h�CD            �     �  �              �              �t�bhhK ��h��R�(KK��h�Cd�      �  v        
      #        �   �           7   v  �   �   "   �   �        �t�bhhK ��h��R�(KK��h�C4   %      �         �   I   t  C   �        �t�bhhK ��h��R�(KKB��h�B     *   %   �      9   �               �  �                �  :                     �        �   �   :         �     q           �      %         �  %         �                  �   i   %         /                  �t�bhhK ��h��R�(KK��h�C@               }              �                �t�bhhK ��h��R�(KK��h�Ct      �        C               �  �     #     �            �        �   �   9      �         �t�bhhK ��h��R�(KK&��h�C�%   �     b                              "  �  '     �	                    �     �  '     �        �   H   7   r   "     �t�bhhK ��h��R�(KK��h�C|                              I                     #                                         �t�bhhK ��h��R�(KKG��h�B              �  ,           2   �  �                             �  �      %                "           �  �        �  �
  �        �                                          P           �            C           "        �t�bhhK ��h��R�(KK7��h�C�   *   2   �                                 "     �         �  �   �     �  �   c   "        %      �                              C        �     %   �         !
              �t�bhhK ��h��R�(KK+��h�C�            
      �     �      �                  I   �  �  �            �  �              C            I      �  �     C   Y           �t�bhhK ��h��R�(KK��h�C|                                 �  �                 
      �  �     �      7                 �t�bhhK ��h��R�(KK	��h�C$   I                        �t�bhhK ��h��R�(KK��h�C8�        �                    �     �     �t�bhhK ��h��R�(KK,��h�C�   �  �  %               "     �       �      "  �  �  �  �       �   N         �          r                 �       �         r      �t�bhhK ��h��R�(KK��h�C\�      �     �  �        #        �                 v                 �t�bhhK ��h��R�(KK+��h�C�   %   A      �  �   w                  �      �                                  �           #  �      �     �      �        v	        �t�bhhK ��h��R�(KK'��h�C�'       �                                    C      �                  �       �	  �  %   A      %           �            �t�bhhK ��h��R�(KK��h�C@        �     
      �     �                   �t�bhhK ��h��R�(KK��h�CT      2         �         �  �      "  �            
      "        �t�bhhK ��h��R�(KK��h�CD`        J   �                     i   N         �     �t�bhhK ��h��R�(KK��h�Cx�              �   �         j      �        I         �  �   D  S   i   -         �     �  r      �t�bhhK ��h��R�(KK8��h�C�         6        4           �   �                 �          "  �      �  �   �  "             �                          �  I      6  V   ^  �              �              �t�bhhK ��h��R�(KK��h�CD�     �        �   �     /      I      �  �  {         �t�bhhK ��h��R�(KK��h�CD%            �             �           C           �t�bhhK ��h��R�(KK(��h�C�   �                    �                              �      �        �     �              C   "                  �        �t�bhhK ��h��R�(KK/��h�C��               �                  <  �                  
                     q              �           �        %      �  O  %                  �t�bhhK ��h��R�(KK��h�CPT         c   �   �   �      b              �            Q         �t�bhhK ��h��R�(KK��h�CT�         g
  [                             [     q              �t�bhhK ��h��R�(KK$��h�C�   �                     �  T   �  �      *           v     #  
                     �                           �t�bhhK ��h��R�(KK��h�Ch   �                                                                           �t�bhhK ��h��R�(KK(��h�C��     �       "        "        *   �   �     �         �                "  �  
      "     T      �   �   o     �     �   �         �t�bhhK ��h��R�(KK��h�C8      G
  q     �         �      %            �t�bhhK ��h��R�(KK��h�Cp   s   �  7      �   �  �        n      �   w   �           I            �    �   ~  �     �t�bhhK ��h��R�(KK��h�CPG   �                    G   �                 �               �t�bhhK ��h��R�(KK$��h�C�      �           
      �                                                   �  `           �        I         �t�bhhK ��h��R�(KK��h�C\�     �     S     �            �   �  �                  �   �            �t�bhhK ��h��R�(KK��h�CP�      Z     �   �        �   �           �      �               �t�bhhK ��h��R�(KK,��h�C�   �         0           ;      H   �     T   �  %      �               �                  �     #   �     Y  �       #   6  C               �t�bhhK ��h��R�(KK��h�C\                           �                  Q      �         C         �t�bhhK ��h��R�(KK��h�Cx*   �   J   �        T      C                        %   �	           �               
            �t�bhhK ��h��R�(KK��h�C<      W              �              Q         �t�bhhK ��h��R�(KK��h�CXT   �                   �   �   �                          �        �t�bhhK ��h��R�(KK,��h�C�               �  H         %                   "              "     �   �      �            �        �  �      S  %         �   �            �t�bhhK ��h��R�(KK#��h�C�   �                        �   �     Q            �      N            �      �     N            �               �t�bhhK ��h��R�(KK��h�C\   �         �            �      �	  "   �     V      �     V      �        �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�CLO
     �
     �      �      +                        �        �t�bhhK ��h��R�(KK$��h�C�   �           �
     �      �   c   �                 �     2         v  �
        �               %      �         �t�bhhK ��h��R�(KK��h�C|                 �               �            �  �      �   �            .                       �t�bhhK ��h��R�(KK&��h�C�T   �                     �  �   *  s                  �                 P           c                  %               �t�bhhK ��h��R�(KK#��h�C�   �  �                �      �            �        �   %      �  O        ,        %      O     �              �t�bhhK ��h��R�(KK��h�Cl�               �         �            �     �        �           �        C         �t�bhhK ��h��R�(KK,��h�C��      �
     �                 �  �              (      �                    �         "                             >   '     "        �t�bhhK ��h��R�(KK(��h�C�            �                     �      �     �              �                       �         �               I  �        �t�bhhK ��h��R�(KK��h�C4   A                              �     �t�bhhK ��h��R�(KK��h�C\                                       �   �  P     �  6  �  �        �t�bhhK ��h��R�(KK��h�C<      '              '              �        �t�bhhK ��h��R�(KK��h�C<   �           �	  
   �  L      7   g   7         �t�bhhK ��h��R�(KK��h�CH�  %   �     C            %      �                        �t�bhhK ��h��R�(KK��h�C\]   �     �        �        q                 ^  �     �     �         �t�bhhK ��h��R�(KK"��h�C�               �   a        �         �   �   ;   6  ^                    �  �   %       
       �            �t�bhhK ��h��R�(KK)��h�C�      5                       ;               u     �      +        �     
               �        A   �  �     
   �   �        �t�bhhK ��h��R�(KK	��h�C$                           �t�bhhK ��h��R�(KK��h�Cp*     ]        �  �     �  �                 �               �           C           �t�bhhK ��h��R�(KK��h�Cx�        �                                 ]      W     C                  �                 �t�bhhK ��h��R�(KK,��h�C��   �        #  �   (   �        N            �             �              j   %      �   �        �     �        �              2        �t�bhhK ��h��R�(KK'��h�C�      /     �              �        ]                                :         �                                       �t�bhhK ��h��R�(KK��h�Cl                     �                 �  �        �   �   �                       �t�bhhK ��h��R�(KK(��h�C�*     _  �  �      �        T   �                             �         �                    �      �  ;         
            �t�bhhK ��h��R�(KK!��h�C�T      C                     Y              �                  "     +                 #     �  "     �t�bhhK ��h��R�(KK*��h�C�   �      �   �            �     u     
         �        �      �  %   I      �  %   �    #   N   s   �       #   N         s            �t�bhhK ��h��R�(KK!��h�C�               c   �            �               �         �           �           �                   �t�bhhK ��h��R�(KK(��h�C�   I   E  �  I   P     �                    �           �   �  %            I            �           �                        �t�bhhK ��h��R�(KK#��h�C�      �     �      
               �     :  '  C  7   W     S           C                                    �t�bhhK ��h��R�(KK��h�CD  +     �  �     +               _  �
  `            �t�bhhK ��h��R�(KK#��h�C�   �        A      �      9   �     _                        �                     �     
  #     �            �t�bhhK ��h��R�(KK!��h�C��         �     D  0         T                  �
  r   Y        Y     "         Y  �      �               �t�bhhK ��h��R�(KK/��h�C�T      �      �          "              V            "   T     o        
         �      �        �        �     "     �      T         �  
            �t�bhhK ��h��R�(KK��h�CD   x     �                    :   �  T     �
        �t�bhhK ��h��R�(KK��h�Cl            �               I   �                  �  �            �      �            �t�bhhK ��h��R�(KK��h�C`                     �            �  �                 �                  �t�bhhK ��h��R�(KK��h�C0   +        C            +           �t�bhhK ��h��R�(KK��h�Cp�      '  T   �   "   �        '   
       '        [        �   �  '     '        �     �t�bhhK ��h��R�(KK��h�C`T      �                        �  �
     �  �     �  �     I      C         �t�bhhK ��h��R�(KK.��h�C�   �        C   �      �     %   �           �  �            %            �  �            �      C   q     �         �      �   0      
   I   �        �t�bhhK ��h��R�(KK3��h�C̥          
      *              <              �           (             T      ]   �                 �           T            �                �  "        �t�bhhK ��h��R�(KK3��h�C̴  �  �      +     O                 ^                    �  ,      "                 �            *   %   �   h           �                �         �  "     �t�bhhK ��h��R�(KK��h�C0�      �
             �	  `            �t�bhhK ��h��R�(KK��h�CxG   +        q  �         �            6  �   �              C                                 �t�bhhK ��h��R�(KK��h�CX         �                 �        "                    "        �t�bhhK ��h��R�(KK��h�Cl   �  �               �            �   �     �  
   +  �              �     "        �t�bhhK ��h��R�(KK��h�Cd�  8   <              �         8              �  $      �      �	              �t�bhhK ��h��R�(KK&��h�C�           o        
         [           T               c         P   g                 �  2         
      "        �t�bhhK ��h��R�(KK-��h�C�   k                    H         �     %   �     
         �  �         2                  2                        �     �   H               �t�bhhK ��h��R�(KK��h�C`�              �  P     �                 w      �      �                  �t�bhhK ��h��R�(KK��h�CT   ]      �                  �     ^     �                       �t�bhhK ��h��R�(KK1��h�C�          "     �               `               �         6                            �     �      J                                    $      "        �t�bhhK ��h��R�(KK(��h�C�   �      �      �   �                 
         q  [                                        P     �     0                 �t�bhhK ��h��R�(KK��h�Cp*     �                  +            �  +   
         �  +         �     �               �t�bhhK ��h��R�(KK'��h�C�                  _           V                 V   D        N         �           �   A      �     I      �     �        �t�bhhK ��h��R�(KK��h�C<T               *   C                          �t�bhhK ��h��R�(KK:��h�C�     �  �     �  T      �  �         �            �                           +            $                      N            o  �        �           N         �   o  �     "        �t�bhhK ��h��R�(KK��h�C\'     +               '     +      8   <        �  �  2      `   9         �t�bhhK ��h��R�(KK��h�CX�     �   C         �            �        �     P        �   �        �t�bhhK ��h��R�(KK��h�CP          "           ;   �  �        �  �   �  8      "        �t�bhhK ��h��R�(KK��h�CP�      �                     �                 �              �t�bhhK ��h��R�(KK!��h�C��               �     #  �        +   �  �        �  ]            �   $            #  �      +   "        �t�bhhK ��h��R�(KK7��h�C�   �            �            %   �                 �         �     �  c   �           �          "           %   A      0    
  ]   "     �     �            C         �   �        �t�bhhK ��h��R�(KK��h�Ct   '       �     �        *   �         r   �     �            #  �   �                    �t�bhhK ��h��R�(KK%��h�C��     %   �     (        �  :            �            �                  �     %         �  �  #     �     �         �t�bhhK ��h��R�(KK,��h�C�   2      ^  P        P        P        �      P                                   �     �                           ]   
               �t�bhhK ��h��R�(KK��h�Cl         �                                      �                    �           �t�bhhK ��h��R�(KK��h�CX                  ]           S        �                          �t�bhhK ��h��R�(KK��h�C`]  $        %                     �      �	           �     
      "        �t�bhhK ��h��R�(KK��h�Cp�              �   
                  �  �      �                        Q               �t�bhhK ��h��R�(KK��h�CD                       q           �               �t�bhhK ��h��R�(KK)��h�C�   �         +   �               �   �        �                 T                  +      �        V           �      $            �t�bhhK ��h��R�(KK��h�CTT         �  �      b  g   7  �                    �     v	        �t�bhhK ��h��R�(KK��h�Ch�   *        �              +                      �         6       "        �t�bhhK ��h��R�(KK*��h�C�      �      
   �            �               {   �  -   �                       {      g               �        �  �     �            �t�bhhK ��h��R�(KK��h�C@�                        �            �           �t�bhhK ��h��R�(KK��h�Cl�                           "              �
        "                             �t�bhhK ��h��R�(KK��h�C@�      C         �     �              A            �t�bhhK ��h��R�(KK��h�C@        �   �              v                    �t�bhhK ��h��R�(KK ��h�C��   �  
   �       �   %      �
     �        �           4     �  %      C   �           �            �t�bhhK ��h��R�(KK��h�C                     �t�bhhK ��h��R�(KK'��h�C�         $               �         +      �                          0      �      
                    C      $   �        �t�bhhK ��h��R�(KK&��h�C�   �              ^     �         C   �   �                        �              C   �         �      C   �  Y           �t�bhhK ��h��R�(KK ��h�C�               P        �     �        �      �  �   �           �  #  �      �	  �      P  �         �t�bhhK ��h��R�(KK"��h�C�      �   5     W	        �  g   �        W	              W	           T      �            S        "        �t�bhhK ��h��R�(KK��h�C`   �   �        �     #         �              �                  "        �t�bhhK ��h��R�(KK��h�CtT      �   �      "        �            �   +         �  �              �                    �t�bhhK ��h��R�(KK3��h�C�
  �            �               �                          �     �     �     %         o        �  �
        �                                   +   "        �t�bhhK ��h��R�(KK#��h�C�`           �  �      �   C        A      C      
                 ~  �                     �   �   �           �t�bhhK ��h��R�(KK��h�CX�                     �     �             #     �      
   �	        �t�bhhK ��h��R�(KK��h�Cp   �        $         �     
      �     �         
         �         $      D  -        �t�bhhK ��h��R�(KK,��h�C�T            Y           �                                  "           �     �  �   +            *              �
     �   o     �         �t�bhhK ��h��R�(KK��h�Cx   �            �                  _  6              �      S           �   D  w              �t�bhhK ��h��R�(KK9��h�C�      2   i         /         #     H   7      �        P        i   �   H      �   P             C         P  [           �   �      j        T   �  �          i   �                     �t�bhhK ��h��R�(KK��h�CL                        �        �         %               �t�bhhK ��h��R�(KK��h�C,      �                  �	        �t�bhhK ��h��R�(KK+��h�C�   �                     �         t              �     �      ^  �           s            �     w         �        �   �      "        �t�bhhK ��h��R�(KK'��h�C�            �      "  8         �   8            $   �            Y  +                            �                     "     �t�bhhK ��h��R�(KK!��h�C�         �	  C   �                          �  �      �  �   �     �   �      �      %         9   �         �t�bhhK ��h��R�(KK&��h�C�           �      �            [        �
  �      +              
   �
        �
        �  +  �         �              �t�bhhK ��h��R�(KK(��h�C�                     �
  �        �   (         #     �   J                 �         �                    �                  �t�bhhK ��h��R�(KK��h�C4`                       `               �t�bhhK ��h��R�(KK��h�Cx               I   �   9   �     �  �                  �      �           /   c   �  �   Q         �t�bhhK ��h��R�(KK��h�C`   *   �     �      �   �   V   2      ~        �      #        ^              �t�bhhK ��h��R�(KK��h�Ct         �           �        �        �     %               <            <               �t�bhhK ��h��R�(KK��h�Ct�                      "  ]      N            �     �      �  0  �
     �     
      "        �t�bhhK ��h��R�(KK��h�Cd�   *      :         C   c            %           �     �        %   �          �t�bhhK ��h��R�(KK��h�CX�   �         *     �         Y        Y                             �t�bhhK ��h��R�(KK��h�C@�     �               -                           �t�bhhK ��h��R�(KK��h�CP   �     �  r           �   �        7                        �t�bhhK ��h��R�(KK/��h�C�         �    �     T         �        r        �     �          "  �        �  �
  "  r            �     �        �
         "  �         "  r      �t�bhhK ��h��R�(KK=��h�C��        +     6  �   +      �      %   �     ^  Y  +   �  %   �        +                  %         �     +   �              2      �  g
  `                  #        �     +            �        �t�bhhK ��h��R�(KK��h�CD            C            �         �   A              �t�bhhK ��h��R�(KK��h�C                     �t�bhhK ��h��R�(KK.��h�C��      �      N   R  
     �  �            
                        �            �                                   
                           �t�bhhK ��h��R�(KK��h�Cl*      �  a     q                            :            A            *           �t�bhhK ��h��R�(KK��h�C|'           �           2                  I         �              �                           �t�bhhK ��h��R�(KK��h�C|   �  �            I         �
  g   I          +  �        j   %               %   �              �t�bhhK ��h��R�(KK,��h�C�                           �     �            L               �                    L         �        �   �  �  �           P  <        �t�bhhK ��h��R�(KK"��h�C�         �                        �                 
      T  �     �         
   V  T        #           �t�bhhK ��h��R�(KK��h�Cx�     �              �           �                  S  �           {                       �t�bhhK ��h��R�(KK2��h�C�   *   %         %        �  �  �
           %   �
              m	     �                    %   �           �     �  '  �                 %      %            �t�bhhK ��h��R�(KK;��h�C�            �      "  ]         Q      �                                          �                $         �               �            +   *        `         �              �   "        �t�bhhK ��h��R�(KK)��h�C�*                              �        g   �  �     P  �               P                             �                        �t�bhhK ��h��R�(KK"��h�C�2   S        �            �         �  �     2            �         �  2      G   +   �         �               �t�bhhK ��h��R�(KK��h�CH      �  W     �
  �  �                         �          �t�bhhK ��h��R�(KK��h�C0   >   �   C                           �t�bhhK ��h��R�(KK"��h�C�j      �                       h   �                  V      �   <     �        �  P      �        6        �t�bhhK ��h��R�(KK,��h�C��             �      o    �     r   �         �     �
        �                       �     �     �                 �  �      �
        �t�bhhK ��h��R�(KK.��h�C�   �  T        %        �  0               r              U                      U  %           C         Y  !     %      �  �	  
           �t�bhhK ��h��R�(KK-��h�C�   �         �  �   C                                      �                                �     �           �            �   P           �t�bhhK ��h��R�(KK��h�CH   %         -   �        T   �  �        �     �         �t�bhhK ��h��R�(KK��h�C|      �  "  )     �   r   "               "  �                                         "        �t�bhhK ��h��R�(KK��h�Cd               �     �  �                        �        �  �               �t�bhhK ��h��R�(KK��h�Cx]                   ]                   ]       2      t      I      �                    �t�bhhK ��h��R�(KK��h�CL            �                     �        �     I         �t�bhhK ��h��R�(KK.��h�C�      �     C     �   
            g
        *         �        �        8         �           5  u        �   a  +                    "        �t�bhhK ��h��R�(KK��h�CPT      �      +            �         7    J   5     �
  r         �t�bhhK ��h��R�(KK��h�C@�  �     �        �     �      �                  �t�bhhK ��h��R�(KK��h�CTP           �      �           �           P        �           �t�bhhK ��h��R�(KK.��h�C��           O  
   �  �  T     �  �            v	  c      �         %      v	        v	     �     q     �  �  �   *         �         %   v	  6        �t�bhhK ��h��R�(KK/��h�C�"  �      %   �  :               �   �                 %  %   �  �                                   (                    �            �   �         �t�bhhK ��h��R�(KK��h�CH            �  �   �     r   *   �   �  C   g   8   �        �t�bhhK ��h��R�(KK��h�C<               �      #     �     �	  "        �t�bhhK ��h��R�(KK(��h�C�         W  �                       �                 *   �      �  *                 �   �      �        �        C         �t�bhhK ��h��R�(KK��h�C\I   �         c                     v           �  A   `  �   v           �t�bhhK ��h��R�(KK+��h�C�         �     �     �   �  G   C      C               �  V      %   *           �     �      Y           �         �   I     �           �t�bhhK ��h��R�(KK��h�Cp   �      ]        U  �     �     U              U  �               �         �         �t�bhhK ��h��R�(KK-��h�C�      N                    �  �  P                         �  �  P           %                        �   #   �  %     �      P     �     �t�bhhK ��h��R�(KK"��h�C��  �     �         �     �         g   8   �     �      "             <             J            �   "     �t�bhhK ��h��R�(KK��h�Cd�     %   ^     �            "     +               �  "        �  
            �t�bhhK ��h��R�(KK-��h�C�   �        I        V   2         t  �                        =                          �   �                       �                     �t�bhhK ��h��R�(KK��h�C|�     I   A   �     '           �      <     �   '                          <     �               �t�bhhK ��h��R�(KK��h�CX*         ]         %   C             "           �            r   "     �t�bhhK ��h��R�(KK.��h�C�                  �     ^        �            $                  �   �  �  �                    <        �  %   s  �  I         I      �        �t�bhhK ��h��R�(KK��h�C@�   �      �                          �   ~  �      �t�bhhK ��h��R�(KK��h�C8"   C                    I                  �t�bhhK ��h��R�(KK��h�CD      �            7   v     *   �      
               �t�bhhK ��h��R�(KK��h�Cl   �         �     ^           �      "     +      g
     �        J      +   "        �t�bhhK ��h��R�(KK��h�CL   �      ^                 P        �   �  
               �t�bhhK ��h��R�(KK&��h�C�T            %      ^           �     C              �   �     �        �     �      "                I      r   "     �t�bhhK ��h��R�(KK,��h�C�S  �  �            �                    �     �               �                        �      �           :   �      �        �   �        �t�bhhK ��h��R�(KK��h�C\�      �   :                        C   w   �                              �t�bhhK ��h��R�(KK!��h�C��   �               :   A   T           �           �     Q         �      P        �  �      �           �t�bhhK ��h��R�(KK��h�C@      �     
   �   s                              �t�bhhK ��h��R�(KK&��h�C�T               �   �              �      �      "          �	  [        "     �     C   �     �  �  �   b   
   �        �t�bhhK ��h��R�(KK��h�CD          "        +                   �  "        �t�bhhK ��h��R�(KK ��h�C�T      �                        "  �  #              '  �   "              (                       �t�bhhK ��h��R�(KK��h�Cl      8   �                 
         �         N                                    �t�bhhK ��h��R�(KK��h�CH   %            �     �               �     �            �t�bhhK ��h��R�(KK'��h�C�   �   J      ^                 �      �                           �     ^        )           �            �              �t�bhhK ��h��R�(KK)��h�C�
   �     �  �   �        /         �                  �      �         �  %      �         C      C  Q      V   %   �   �     �        �t�bhhK ��h��R�(KK<��h�C�                           �   /         %     �                 �           �     �     %                 Y  �            �   w      �         �                  �     �        �
        �t�bhhK ��h��R�(KK%��h�C�                 '     g   %      �            �     ]               �                 �   #  �        :            �t�bhhK ��h��R�(KK��h�CL�            �      
   �   �
     �            �             �t�bhhK ��h��R�(KK��h�C<   �                 �                        �t�bhhK ��h��R�(KK2��h�CȚ   V   �         �   I        �              j  �     *        �              �   �
        :      V      �            �      Y  �           �   �              �t�bhhK ��h��R�(KK!��h�C��   J   O  #                    *     �           �   �        �      �     %        �                 �t�bhhK ��h��R�(KK��h�C0               �                     �t�bhhK ��h��R�(KK��h�C|   T                 7        !  �   #  �       �      �      j         7     C   w      7        �t�bhhK ��h��R�(KK-��h�C�               �         "  +                                              �      �        �          ;              j                  �t�bhhK ��h��R�(KK&��h�C�T               �   �              �      �      "          �	  [        "     �     C   �     �  �  �   b   
   �        �t�bhhK ��h��R�(KK��h�CH               P           �   �           b     �     �t�bhhK ��h��R�(KK"��h�C�"           �  �                    �         �         j   �
  �   �   �   �     �                           �t�bhhK ��h��R�(KK��h�C\            0        �   �      ]  �  �     q     #      i               �t�bhhK ��h��R�(KK&��h�C�P     �                                                      g            �                                         �t�bhhK ��h��R�(KK��h�CD�      O  
   �            �                           �t�bhhK ��h��R�(KK2��h�C�                            �   �                 /         C                         �                                                                    �t�bhhK ��h��R�(KK)��h�C��     C  �        �   �                    %   �  
         ~              �   J     ]     �      *   C        �      �           �t�bhhK ��h��R�(KK0��h�C�   �     �  �        �     *               J   �   �                  �                                    �            �  �         +           "     �t�bhhK ��h��R�(KK��h�CH�   %               �            �      �   �  C     �     �t�bhhK ��h��R�(KK��h�C<                     �  i   H      �           �t�bhhK ��h��R�(KK��h�CT        �        I     j                        I              �t�bhhK ��h��R�(KK+��h�C�               �   g      �                                       �   �  6                   �         "   �     �                    �t�bhhK ��h��R�(KK1��h�C�         �   �           �       "                                      9      �        �               �      9         �   I         J  C   
      "        �t�bhhK ��h��R�(KK��h�CL`           �                 �                          �t�bhhK ��h��R�(KK��h�CX   �         �               ]   Q         Q                           �t�bhhK ��h��R�(KK��h�Ch         �  c         �      �   �           C   w            T   P           r      �t�bhhK ��h��R�(KK��h�C4�                  2            �        �t�bhhK ��h��R�(KK��h�Cd   #     >                        $                         �              �t�bhhK ��h��R�(KK��h�C4                  �  P                 �t�bhhK ��h��R�(KK$��h�C�   �        %                  �             �                                    ]   
                        �t�bhhK ��h��R�(KK��h�Ct         
         
   �     �              %   A            �         �                    �t�bhhK ��h��R�(KK��h�C\�           d        Q   �           �                    �           �t�bhhK ��h��R�(KK.��h�C�j         6        �           $                     �   <        V                        *   [    �     L   
   �     T         c   �           �t�bhhK ��h��R�(KK��h�CL      �   _      �  t     i                           �     �t�bhhK ��h��R�(KK��h�Cd   �  �      �  �  �         �         �     N               N   +               �t�bhhK ��h��R�(KK(��h�C�      �  
      �  �                    C   q              �            Y     �  �   "      L   T   [     �     �   �            �t�bhhK ��h��R�(KK��h�C\               �    �  �                        �            "        �t�bhhK ��h��R�(KK��h�CxT         �      "                             �  �         �  �  V   �         �      "        �t�bhhK ��h��R�(KK��h�CL                             Q        �   �              �t�bhhK ��h��R�(KK.��h�C�      �         �                     �                          �  �                          �  �               �   J      �     N            �t�bhhK ��h��R�(KK��h�CL   �   
   +        �   �  �     �     >   �      G   �        �t�bhhK ��h��R�(KK)��h�C�   �            C           �      2           t  �   �           �         �    �  �  �     �  �  �  2      �                  �t�bhhK ��h��R�(KK.��h�C�          "     �  �             Y  %  �      �        �           r   "               "  �     �                                   "        �t�bhhK ��h��R�(KK��h�C\�                     e     i      �        �   �  �         
   U        �t�bhhK ��h��R�(KK��h�C\      D        
           �
        �     �      w         �   C         �t�bhhK ��h��R�(KK��h�CX               �               �            �     �                 �t�bhhK ��h��R�(KK��h�CH               �      %   s         �                    �t�bhhK ��h��R�(KK#��h�C�V      �   C      �   �      *   �   �                       �      S        �      Y  �        �      �            �t�bhhK ��h��R�(KK��h�Cl                     %               �                                             �t�bhhK ��h��R�(KK��h�Cd         �                              �           �         �     0        �t�bhhK ��h��R�(KK��h�Ch          "  �      �  �         P                    g
  �     �  '              �t�bhhK ��h��R�(KK"��h�C�         �  �                                 �     �         �  *   �              �            ]         �t�bhhK ��h��R�(KK��h�Cd   %                "              �           *     %     �   s               �t�bhhK ��h��R�(KK��h�C,   �                               �t�bhhK ��h��R�(KK��h�C<   �                 �                        �t�bhhK ��h��R�(KK��h�CX                 T   2   J                  c   y     �              �t�bhhK ��h��R�(KK'��h�C�   �              a  g   $      7        7     �   �                      C      �                             "        �t�bhhK ��h��R�(KK��h�C@�                      �      �     �      r      �t�bhhK ��h��R�(KK ��h�C��   %            �         
   �   �     �           T      I                     �                    �t�bhhK ��h��R�(KK��h�CT   C        �                              �  %   6  V      �     �t�bhhK ��h��R�(KK��h�CX      �  8                           +   �   Y  �
     �   $   <         �t�bhhK ��h��R�(KK��h�Ct�                  �      �  �   �               2                     �   �  G               �t�bhhK ��h��R�(KK��h�CT      /                             �                        �     �t�bhhK ��h��R�(KK&��h�C��  �      
        2            k                 �        �   >   �  �      �  %               %      V         �        �t�bhhK ��h��R�(KK&��h�C�                           Y                       �           �  �         P  �                                   �t�bhhK ��h��R�(KK��h�Cl�      ]              %      �   �  
            �  �  P  ]  �     �        C         �t�bhhK ��h��R�(KK��h�Cp   �                  �   (   �                �      �                                �t�bhhK ��h��R�(KK+��h�C�         +         t     �      �   2         G   v	  �                  �     0   �      �                    �     0      �           �t�bhhK ��h��R�(KK.��h�C�   �                  �   �  �        �      +        +           b  �        �            A            �   �  �        %                        �t�bhhK ��h��R�(KK#��h�C�S        �         �        �   G
        �         �
     �     �              +      �           8   �        �t�bhhK ��h��R�(KK��h�CP�        �  �	           +        �           �               �t�bhhK ��h��R�(KK��h�C|         
           P           �                "     J   �      +               8   <  "        �t�bhhK ��h��R�(KK��h�C88               J   �         `               �t�bhhK ��h��R�(KK��h�Ch�            \                 �                                       "        �t�bhhK ��h��R�(KK��h�CH�   *   �      ]      �  �               �   �   �            �t�bhhK ��h��R�(KK��h�Cp#  �     �           ]            Q       "                    �              "  r      �t�bhhK ��h��R�(KK��h�CT               N              t                    �            �t�bhhK ��h��R�(KK��h�Cx   �   W  (                  "  �           v	  �     �     
   E
     �          V   "        �t�bhhK ��h��R�(KK2��h�C�           �
     I              �           �        �   \  �        �           
   o  b     �      �        -            �   �             �   �         �t�bhhK ��h��R�(KK��h�CX                                                                  �t�bhhK ��h��R�(KK��h�C8   
        �      "         V               �t�bhhK ��h��R�(KK��h�C\   �     J      C      �      �   �         �         �      a        �     �t�bhhK ��h��R�(KK"��h�C�         �          "        T                  +     r      -   �
     +     "              c               �t�bhhK ��h��R�(KK��h�CD      �                           �      �            �t�bhhK ��h��R�(KK.��h�C�T   �   �     0   �                            �   �  �        �                 �           �   �      �     �   �              �  �  �         �t�bhhK ��h��R�(KK��h�C\               C   �         �      �   �      �  �         �      �        �t�bhhK ��h��R�(KK��h�Cp   �   �                  "     G   �
  "     �   �   �	        �  �            W  c         �t�bhhK ��h��R�(KK3��h�C�T      �      �      "  S                   ,     �           �  �  +      *        [  �
  "        *   �      �   �  [  �     W        ~  �        �  �        �t�bhhK ��h��R�(KK��h�CT              8        s   �                 e        �        �t�bhhK ��h��R�(KK"��h�C�            V         ]         T       "     �         "     A          "     �                  �  "        �t�bhhK ��h��R�(KK��h�CP   �           C                  C      `                     �t�bhhK ��h��R�(KK"��h�C�]     C                              2            V         �            "  �  �            <      "        �t�bhhK ��h��R�(KK/��h�C��      I   �                          b  �     �     �                                   �                    j               �                 �t�bhhK ��h��R�(KK��h�Cx      +     
                  g   �   P        �      
            %   A               �
  �     �t�bhhK ��h��R�(KK/��h�C��   �      �   B  ~  +             G   +   �     �	  D  "      6     P              �   �  t              /      �      %   �        :                     �t�bhhK ��h��R�(KK5��h�C�T               �  #  �   �     
              �       "  #        �                    r     �     ]        �  9         �     >         +   :   �  q        r   "     �t�bhhK ��h��R�(KK��h�C,      �           �              �t�bhhK ��h��R�(KK��h�C<   C     �  �              �     �  r   "     �t�bhhK ��h��R�(KK��h�CL               G   �            P        �     g   �        �t�bhhK ��h��R�(KK*��h�C�            �  �                 o           r         �
                            $   L            G   �
        �        "     �t�bhhK ��h��R�(KK��h�Ct�      T                     \     P              9   P        �                �        �t�bhhK ��h��R�(KK��h�C|   �      I   �     �         �   �      �     �      �  #  �   �     �   �      �     �     "        �t�bhhK ��h��R�(KK2��h�C�   %   �  �     �                u     �                                    �                        9               "               %   #                 �t�bhhK ��h��R�(KK��h�CD�         :  j   7  �  �   *      W     �     �        �t�bhhK ��h��R�(KK��h�C\'     �                                       N               L         �t�bhhK ��h��R�(KK-��h�C�]      #              �              :         %         �     �                             �        �         �     g
  [                 �t�bhhK ��h��R�(KK��h�C|   �         �     �              "      
     2   q           "                  
   �   6         �t�bhhK ��h��R�(KK��h�C\*               :            -      :            I                       �t�bhhK ��h��R�(KK��h�C\   �
           �      �         �  s   �
     �      �         i            �t�bhhK ��h��R�(KK��h�Cl         �           �   �         "     �               �
     �        �   "        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CP         �   �           �           �  �     �   '           �t�bhhK ��h��R�(KK��h�CT     �                       �         >      c      Y  �
  r      �t�bhhK ��h��R�(KK ��h�C�     +            �      +           C   [  +      �      �     a  +                        Q         �t�bhhK ��h��R�(KK#��h�C�            �            "  #  J         �      �   +   r   "           �      "           �
  0   +     "        �t�bhhK ��h��R�(KK(��h�C�                     �  �   �                             �  �   �                               �                �     �t�bhhK ��h��R�(KK��h�Cd                  $            �  8               $               $   Z        �t�bhhK ��h��R�(KK��h�Ct            �          "           "        %                              V   
            �t�bhhK ��h��R�(KK-��h�C�      �      D     �                 �         j      5  �   �            �      �                 �            �  �         T   a  �          �t�bhhK ��h��R�(KK-��h�C�                  s   �   2           �  �            C      b     �      �         (   �  6  �            �      �   H  �  �         P  _        �t�bhhK ��h��R�(KK"��h�C�%                     �                                                                                 �t�bhhK ��h��R�(KK��h�CT      �  2                       �   ?                          �t�bhhK ��h��R�(KK%��h�C�   +                          V   ]   �                  �     �  I                  �   �   �                        �t�bhhK ��h��R�(KK1��h�C�*         �        �                  �   �  Y  I   �      �         Y        Y     /      Y        Y              Y     �     '  �      C      �   �         �t�bhhK ��h��R�(KK��h�Ct            *   �   �           7   v        2      �        �                              �t�bhhK ��h��R�(KK��h�Ch      C                              �   �   /      �                             �t�bhhK ��h��R�(KK��h�Ct%      C      �            %            %   �  t  c      �  %   �      "  �  �  *     r   "     �t�bhhK ��h��R�(KK��h�Cx   �      2                  2            �     /                                           �t�bhhK ��h��R�(KK��h�CX                                             �       C           �t�bhhK ��h��R�(KK ��h�C�      �            �  D  R     �                    �  T   �       �       �        �           �t�bhhK ��h��R�(KK!��h�C��  �           �       S                                *     �     �   �   �         �                 �t�bhhK ��h��R�(KK��h�C@               V         Q      �     �           �t�bhhK ��h��R�(KK��h�C<              �  #                          �t�bhhK ��h��R�(KK'��h�C�   *         �        %      �                "                          �   �        W  Q         �   H            "        �t�bhhK ��h��R�(KK*��h�C�*   %      ]         %            %         �      "     5                 H                     �              I      %      �        �t�bhhK ��h��R�(KK��h�C8   a        
            _  0     �        �t�bhhK ��h��R�(KK4��h�C�      �  ]   
  <     C      N   "     "     S                      �  "     "              �  �           "     ]     "                    �                 �t�bhhK ��h��R�(KK��h�CtT                         "  �         +         �            �     �      `      [  �
        �t�bhhK ��h��R�(KK��h�C4T            c   :            �           �t�bhhK ��h��R�(KK��h�CH               $               :                  �     �t�bhhK ��h��R�(KK+��h�C��   4     �  #                          �              0   #        I               �       �     �      %         '  �              �t�bhhK ��h��R�(KK��h�C<�   H                  �           �           �t�bhhK ��h��R�(KK=��h�C��   �           �           �                        �      %   *  �      �
        *  �  %               %   �  �	     g   �     �  2   �     g               �     �	  �     �  2      �            �t�bhhK ��h��R�(KK#��h�C�            �             "  �            �        �  �
     �                       j               "        �t�bhhK ��h��R�(KK��h�CL   �  [  �  P                             %              �t�bhhK ��h��R�(KK��h�CP                  r      �           r            -            �t�bhhK ��h��R�(KK��h�CX      �   �         �   �  �     �        �            
     �        �t�bhhK ��h��R�(KK.��h�C��         6  �        �           �  g      6  �  �     P        �   ]              �      �   �                                       "        �t�bhhK ��h��R�(KK��h�Cd   �     T                        �      "     %           �        "        �t�bhhK ��h��R�(KK��h�C<�   H                              �           �t�bhhK ��h��R�(KK��h�CL   q  �   :   P           �  :   P     �        :   �        �t�bhhK ��h��R�(KK��h�CLh   �         >   %            %   0                           �t�bhhK ��h��R�(KK��h�Cx      �     �          �        �      �   �  (                                             �t�bhhK ��h��R�(KK��h�C<   �   �              �  v	  ^  �  %            �t�bhhK ��h��R�(KK!��h�C�`     �              "     %         �      "  '                   '                 �  �   "        �t�bhhK ��h��R�(KK��h�C\   �         �            �      �	  "   �     V      �     V      �        �t�bhhK ��h��R�(KK%��h�C��                             �      2   �   T   *         �           
     �                              "        �t�bhhK ��h��R�(KK��h�C|         �                          �                           �           �                 �t�bhhK ��h��R�(KK��h�CP            P     �      �  P     �      �  P     �            �t�bhhK ��h��R�(KK��h�Cl   �     G   �         �   �  %   �           �  %                        "   �         �t�bhhK ��h��R�(KK2��h�Cȳ         o         "  *     �      �  �
  I           �               �                  �   �
        �      �  �                 o                 "        �t�bhhK ��h��R�(KK��h�C`�   *      W              �     �   Y  �        �   �     r                 �t�bhhK ��h��R�(KK#��h�C�T                  �        �        �     �                    $                           O              �t�bhhK ��h��R�(KK&��h�C��            �     �
                 �     �      b                          �      o  �     +           0            �t�bhhK ��h��R�(KK��h�CdV   �              "   <                                         I  �        �t�bhhK ��h��R�(KK��h�CP�     �
                             �
  
   �                 �t�bhhK ��h��R�(KK��h�CT   �  �      �   ]      T               S                         �t�bhhK ��h��R�(KK��h�C<   I   %                     %         /         �t�bhhK ��h��R�(KK'��h�C�   w            �                               +           +   
   +     6         �  �         `      +                     �t�bhhK ��h��R�(KK)��h�C�         ]            �         +   �     \     v        T            $                  [     �                                �t�bhhK ��h��R�(KK��h�C4               �     �  �                �t�bhhK ��h��R�(KK��h�Cp         ^     Y                                   �                 C               �t�bhhK ��h��R�(KK��h�CLT   *         �                     I      
                  �t�bhhK ��h��R�(KK��h�Cl      %  2                        �     I   %   Y           �  �     
      "        �t�bhhK ��h��R�(KK,��h�C�*   �   �           6  ^  g   �                       �                                   �   *   %   T      g   �        �                 �t�bhhK ��h��R�(KK��h�C8              '           �               �t�bhhK ��h��R�(KK��h�CH�           �  P     r   �     C   �   0  P     �  r      �t�bhhK ��h��R�(KK��h�CxV                        �        �      �  �     �                                 �        �t�bhhK ��h��R�(KK��h�Ch         
            *      �     �            g
     S       V   �  �            �t�bhhK ��h��R�(KK��h�CD   a                                               �t�bhhK ��h��R�(KK��h�CD                 [        �                       �t�bhhK ��h��R�(KK��h�Cd�               �        �         �              �           �               �t�bhhK ��h��R�(KK*��h�C��  �     �                   �        �   �      �  �           �         �  �        Y     �  ^  �            �   �      Y           �t�bhhK ��h��R�(KK��h�CH   �
     +        8               �        `            �t�bhhK ��h��R�(KK��h�Cd                                 /               A      T            �         �t�bhhK ��h��R�(KK+��h�C��  �              �               o  �           ~                     *   �      +               �      Y  +      �  2                  �t�bhhK ��h��R�(KK&��h�C�*   T      W  �                     �      "  �      �            "     '  �   �  �         r           �   I     "        �t�bhhK ��h��R�(KK+��h�C��        o  �           Q       "     T              r      
       #   V   r   "  �          %      �
     �            �   �     r      �t�bhhK ��h��R�(KK,��h�C�      $              �   �            %            $                 �   �        �   ]   �                       �                        �t�bhhK ��h��R�(KK��h�C0   2      9   �      I         u        �t�bhhK ��h��R�(KK#��h�C�             �     ]   �     �  �        �  C           �   �          O  +  ,     #     �  �  �        �t�bhhK ��h��R�(KK��h�CH         W  c               P              �   �  �     �t�bhhK ��h��R�(KK��h�C`         �                                                              �t�bhhK ��h��R�(KK��h�Cx   *      W  �   �            �       "  �      ;                              $      r   "     �t�bhhK ��h��R�(KK ��h�C�            �     +            J   N   P        �  �            +               J   �	  I   P     �     �t�bhhK ��h��R�(KK��h�C4�     �   C                              �t�bhhK ��h��R�(KK��h�C|        �               
   P           �            "  *              +         �   �            �t�bhhK ��h��R�(KK��h�C<                     *   �   �      7   v        �t�bhhK ��h��R�(KK!��h�C�P                             
                     *  �     �     *     �        �   �              �t�bhhK ��h��R�(KK��h�C<   C           �  �      �  C  �  Y  +         �t�bhhK ��h��R�(KK��h�Ct                              �            �            �           C      �     "        �t�bhhK ��h��R�(KK��h�C@      O  �   �     I           `     �            �t�bhhK ��h��R�(KK,��h�C�            �          "  �   �     �            *              �     �   :   ]   Q         Q      �                                 "        �t�bhhK ��h��R�(KK��h�C@                  %               %               �t�bhhK ��h��R�(KK��h�Ct�        �          "        +        G               �   �  �        �  :   P     �  "     �t�bhhK ��h��R�(KK��h�CD�            �   �               �
           �        �t�bhhK ��h��R�(KK*��h�C�U  _  �     P                    �         �      T   W        �                    o  �  %                "             �  "     �t�bhhK ��h��R�(KK��h�ClT         �  $          "  '                    �         �            c   �           �t�bhhK ��h��R�(KK��h�Ct�               �  *  �     V   �      "            
   �            "  -   �  �      �        �t�bhhK ��h��R�(KK��h�Cp      2            �      "        �            +   +                                   �t�bhhK ��h��R�(KK��h�Cx�            T               �   v	              �         %            �  (   6     �           �t�bhhK ��h��R�(KK��h�CD#  2           G               
        N            �t�bhhK ��h��R�(KK��h�CH+     J   �   �     [           +     J   �   �  ;         �t�bhhK ��h��R�(KK'��h�C�   �           �            #  v	     �  �   S  �                j      �
     �           c   �        �                 �t�bhhK ��h��R�(KK#��h�C�       �     �                    �  
            �           `         8   �     �        �   �   �            �t�bhhK ��h��R�(KK��h�Cp   �   W                       T      �               �           �  �   �              �t�b��      hhK ��h��R�(KK��h�C|T      �       "  *     $            (     �   �        �      �           (     �  $      "        �t�bhhK ��h��R�(KK��h�Ch   �        �        T         �  �   �  �                       �  �           �t�bhhK ��h��R�(KK%��h�C�             "              �   �                    %        *  �                    %      *  �        "        �t�bhhK ��h��R�(KK��h�C0   ]      �                           �t�bhhK ��h��R�(KK%��h�C�   �      �     (     P           �      0   6     
               �     
                     �   0      C            �t�bhhK ��h��R�(KK��h�C<      P           �           I   P  9         �t�bhhK ��h��R�(KK$��h�C�            �      *   �      H  �                           �   �     #           N                     C          �t�bhhK ��h��R�(KK��h�C<                  2   �         I   �            �t�bhhK ��h��R�(KK��h�C8%   �                             I        �t�bhhK ��h��R�(KK��h�Cl                                 I                       %            I           �t�bhhK ��h��R�(KK��h�CP*         ]         %   �  �              �     �              �t�bhhK ��h��R�(KK��h�C\   �   �        �                 �      %                  $   �         �t�bhhK ��h��R�(KK1��h�C�               �       "     �   i         �
  w      �   $  �   o           �   D     �      �        '  �     �  �   �          �   �         '  �           �t�bhhK ��h��R�(KK��h�C                         �t�bhhK ��h��R�(KK��h�CL�   �  �           2   0                                    �t�bhhK ��h��R�(KK��h�Cd   �              �         j         �     �  +   �   �      j            r      �t�bhhK ��h��R�(KK��h�CxT      �      �       "  :               :         W     "     �   9   �   _     %                 �t�bhhK ��h��R�(KK��h�C`         t     �        a                       C            �            �t�bhhK ��h��R�(KK
��h�C(                              �t�bhhK ��h��R�(KK$��h�C��         c            I               �      "  *   �              �                      �                 "     �t�bhhK ��h��R�(KK��h�C|   W  �                    �      I   �        �      �     �  �      �   �            
            �t�bhhK ��h��R�(KK#��h�C��                          �   �         /  �    �           =                 
     �   �         /        �t�bhhK ��h��R�(KK��h�CD�                    g
  �       �                     �t�bhhK ��h��R�(KKA��h�B                     "     �        �	  �      r   �            �        �   J     
     �      N      �         �  8               6     �   J      +                        P        �         �
        "        �t�bhhK ��h��R�(KK��h�CP   I                           �  �     %      C               �t�bhhK ��h��R�(KK��h�Ch%      T      ~  P  �        C   �     �         
      �     "   �  �      l         �t�bhhK ��h��R�(KK��h�C|         �   �              �   s            C              �         g   P                       �t�bhhK ��h��R�(KK&��h�C�*   �   �     �
        �                       #  D  %     �         �   g         S   i         2   �        �  r         �t�bhhK ��h��R�(KK��h�Ch   C  /                           %     I              �      %   A               �t�bhhK ��h��R�(KK��h�C    �      %                �t�bhhK ��h��R�(KK��h�Cx�      �  ^  �              �              �  �      �        �           �                 �t�bhhK ��h��R�(KK��h�CX*   %   �              �   �      %         �  I     �      �   �        �t�bhhK ��h��R�(KK��h�CX   �         0   }  �         %               �  �   �     �  �         �t�bhhK ��h��R�(KK#��h�C�            �     V   �                   "     �     �                                I                    �t�bhhK ��h��R�(KK��h�CX   �         �      "     �      6  `         $            +   "        �t�bhhK ��h��R�(KK��h�C4�               H	  �     j            �t�bhhK ��h��R�(KK'��h�C�   �            �                  ]         *   �   �                    �   �           �           P        �
  ]         �t�bhhK ��h��R�(KK ��h�C�         0   7               �      �      g   ]      C               v         C   g   1     �   7         �t�bhhK ��h��R�(KK��h�CTT      �      �
      6  �  �   J      +      �	  g
              "     �t�bhhK ��h��R�(KK��h�C<   %      C            C  �                    �t�bhhK ��h��R�(KK��h�C<                  �         �  �               �t�bhhK ��h��R�(KK��h�CP�        $   �   N      �   `               I   `            �     �t�bhhK ��h��R�(KK��h�C`   �         �       "  �                  ]                  o        �     �t�bhhK ��h��R�(KK!��h�C�   �  �           �  '                          �  �           �      �  �            ^     �        �t�bhhK ��h��R�(KK$��h�C�   *   �                  �      �               �               �
        �                  �   �     g
           �t�bhhK ��h��R�(KK��h�CL�        [     �     �     �                  9      �     �t�bhhK ��h��R�(KK��h�C`   I               /      �           %  %      ^           �     �  �     �t�bhhK ��h��R�(KK6��h�Cش  �           C            �      "  #        �  Y     �        �      �
  Y  +      S           �   �
     o              �   I     r   
                 Y  �
  "        �t�bhhK ��h��R�(KK=��h�C�   �   D     �  g   +  �                 #                    [     �     �            6  �  �     ]  A           _     *   �     #                    �      �     �  �            "        �t�bhhK ��h��R�(KK��h�CD   �                                               �t�bhhK ��h��R�(KK��h�CT�   �         g   o  �                 %   �  �  �                 �t�bhhK ��h��R�(KK��h�C4            I     �                      �t�bhhK ��h��R�(KK#��h�C�   %   �  �                          �              �   �             *  �           �   �                  �t�bhhK ��h��R�(KK��h�C`�     +        N   G   �         �      N   C           %   �  N   o  �        �t�bhhK ��h��R�(KK��h�Cd   *     %            g
  [  +   �     �        �                  :   +         �t�bhhK ��h��R�(KK��h�C8         �  ^  P              
   �         �t�bhhK ��h��R�(KK��h�Cx            2   �     �   �   �              #  �   �            �  �         "        "        �t�bhhK ��h��R�(KK'��h�C��   �                             v                   j                                    �     �  �   �  �            �t�be.