men Aron och hans söner ombesörjde offren på brännoffersaltaret och på rökelsealtaret , och skulle utföra all förrättning i det allraheligaste och bringa försoning för Israel , alldeles såsom Mose , Guds tjänare , hade bjudit .
och dessa voro Arons söner : hans son Eleasar , dennes son Pinehas , dennes son Abisua ,
dennes son Bucki , dennes son Ussi , dennes son Seraja ,
dennes son Merajot , dennes son Amarja , dennes son Ahitub ,
dennes son Sadok , dennes son Ahimaas .
och dessa voro deras boningsorter , efter deras tältläger inom deras område : åt Arons söner av kehatiternas släkt -- ty dem träffade nu lotten --
åt dem gav man Hebron i Juda land med dess utmarker runt omkring .
men åkerjorden och byarna som hörde till staden gav man åt Kaleb , Jefunnes son .
åt Arons söner gav man alltså fristäderna Hebron och Libna med dess utmarker , vidare Jattir och Estemoa med dess utmarker .
Hilen med dess utmarker , Debir med dess utmarker ,
Asan med dess utmarker och Bet @-@ Semes med dess utmarker ;
och ur Benjamins stam Geba med dess utmarker , Alemet med dess utmarker och Anatot med dess utmarker , så att deras städer tillsammans utgjorde tretton städer , efter deras släkter .
och Kehats övriga barn fingo ur en stamsläkt , nämligen den stamhalva som utgjorde ena hälften av Manasse stam , genom lottkastning tio städer .
Gersoms barn åter fingo , efter sina släkter , ur Isaskars stam , ur Asers stam , ur Naftali stam och ur Manasse stam i Basan tretton städer .
Meraris barn fingo , efter sina släkter , ur Rubens stam , ur Gads stam och ur Sebulons stam genom lottkastning tolv städer .
så gåvo Israels barn åt leviterna dessa städer med deras utmarker .
genom lottkastning gåvo de åt dem ur Juda barns stam , ur Simeons barns stam och ur Benjamins barns stam dessa städer , som de namngåvo .
och bland Kehats barns släkter fingo några följande städer ur Efraims stam såsom sitt område :
man gav dem fristäderna Sikem med dess utmarker i Efraims bergsbygd , Geser med dess utmarker ,
Jokmeam med dess utmarker , Bet @-@ Horon med dess utmarker ;
vidare Ajalon med dess utmarker och Gat @-@ Rimmon med dess utmarker ;
och ur ena hälften av Manasse stam Aner med dess utmarker och Bileam med dess utmarker . detta tillföll Kehats övriga barns släkt .
Gersoms barn fingo ur den släkt som utgjorde ena hälften av Manasse stam Golan i Basan med dess utmarker och Astarot med dess utmarker ;
och ur Isaskars stam Kedes med dess utmarker , Dobrat med dess utmarker ,
Ramot med dess utmarker och Anem med dess utmarker ;
och ur Asers stam Masal med dess utmarker , Abdon med dess utmarker ,
Hukok med dess utmarker och Rehob med dess utmarker ;
och ur Naftali stam Kedes i Galileen med dess utmarker , Hammon med dess utmarker och Kirjataim med dess utmarker .
Meraris övriga barn fingo ur Sebulons stam Rimmono med dess utmarker och Tabor med dess utmarker ,
och på andra sidan Jordan mitt emot Jeriko , öster om Jordan , ur Rubens stam Beser i öknen med dess utmarker , Jahas med dess utmarker ,
Kedemot med dess utmarker och Mefaat med dess utmarker ;
och ur Gads stam Ramot i Gilead med dess utmarker , Mahanaim med dess utmarker ,
Hesbon med dess utmarker och Jaeser med dess utmarker .
och Isaskars söner voro Tola och Pua , Jasib och Simron , tillsammans fyra .
Tolas söner voro Ussi , Refaja , Jeriel , Jamai , Jibsam och Samuel , huvudmän för sina familjer , ättlingar av Tola , tappra stridsmän , upptecknade efter sin ättföljd . i Davids tid var deras antal tjugutvå tusen sex hundra .
Ussis söner voro Jisraja , och Jisrajas söner voro Mikael , Obadja och Joel samt Jissia , tillhopa fem , allasammans huvudmän .
och med dem följde stridbara härskaror , trettiosex tusen man , efter sin ättföljd och sina familjer ; ty de hade många hustrur och barn .
och deras bröder i alla Isaskars släkter voro tappra stridsmän ; åttiosju tusen utgjorde tillsammans de som voro upptecknade i deras släktregister .
Benjamins söner voro Bela , Beker och Jediael , tillsammans tre .
Belas söner voro Esbon , Ussi , Ussiel , Jerimot och Iri , tillsammans fem , huvudmän för sina familjer , tappra stridsmän ; de som voro upptecknade i deras släktregister utgjorde tjugutvå tusen trettiofyra .
Bekers söner voro Semira , Joas , Elieser , Eljoenai , Omri , Jeremot , Abia , Anatot och Alemet . alla dessa voro Bekers söner .
de som voro upptecknade i deras släktregister , efter sin ättföljd , efter huvudmannen för sina familjer , tappra stridsmän , utgjorde tjugu tusen två hundra .
Jediaels söner voro Bilhan ; Bilhans söner voro Jeus , Benjamin , Ehud , Kenaana , Setan , Tarsis och Ahisahar .
alla dessa voro Jediaels söner , upptecknade efter huvudmännen för sina familjer , tappra stridsmän , sjutton tusen två hundra stridbara krigsmän .
och Suppim och Huppim voro Irs söner . -- Men Husim voro Ahers söner .
Naftalis söner voro Jahasiel , Guni , Jeser och Sallum , Bilhas söner .
Manasses söner voro Asriel , som kvinnan födde ; hans arameiska bihustru födde Makir , Gileads fader .
och Makir tog hustru åt Huppim och Suppim . hans syster hette Maaka . och den andre hette Selofhad . och Selofhad hade döttrar .
och Maaka , Makirs hustru , födde en son och gav honom namnet Peres , men hans broder hette Seres . hans söner voro Ulam och Rekem .
Ulams söner voro Bedan . dessa voro söner till Gilead , son till Makir , son till Manasse .
och hans syster var Hammoleket ; hon födde Is @-@ Hod , Abieser och Mahela .
och Semidas söner voro Ajan , Sekem , Likhi och Aniam .
och Efraims söner voro Sutela , dennes son Bered , dennes son Tahat , dennes son Eleada , dennes son Tahat ,
dennes son Sabad och dennes son Sutela , så ock Eser och Elead . och män från Gat , som voro födda där i landet , dräpte dem , därför att de hade dragit ned för att taga deras boskapshjordar .
då sörjde Efraim , deras fader , i lång tid , och hans bröder kommo för att trösta honom .
och han gick in till sin hustru , och hon blev havande och födde en son ; och han gav honom namnet Beria , därför att det hade skett under en olyckstid för hans hus .
hans dotter var Seera ; hon byggde Nedre och Övre Bet @-@ Horon , så ock Ussen @-@ Seera .
och hans son var Refa ; hans son var Resef , ävensom Tela ; hans son var Tahan .
hans son var Laedan ; hans son var Ammihud ; hans son var Elisama .
hans son var Non ; hans son var Josua .
och deras besittning och deras boningsorter voro Betel med underlydande orter , österut Naaran och västerut Geser med underlydande orter , vidare Sikem med underlydande orter , ända till Aja med underlydande orter .
men i Manasse barns ägo voro Bet @-@ Sean med underlydande orter , Taanak med underlydande orter , Megiddo med underlydande orter , Dor med underlydande orter . här bodde nu Josefs , Israels sons , barn .
Asers söner voro Jimna , Jisva , Jisvi och Beria ; och deras syster var Sera .
Berias söner voro Heber och Malkiel ; han var Birsaits fader .
och Heber födde Jaflet , Somer och Hotam , så ock Sua , deras syster .
och Jaflets söner voro Pasak , Bimhal och Asvat . dessa voro Jaflets söner .
Semers söner voro Ahi och Rohaga , Jaba och Aram .
hans broder Helems söner voro Sofa , Jimna , Seles och Amal .
Sofas söner voro Sua , Harnefer , Sual , Beri och Jimra ,
beser , Hod , Samma , Silsa , Jitran och Beera .
Jeters söner voro Jefunne , Pispa och Ara .
och Ullas söner voro Ara , Hanniel och Risja .
alla dessa voro Asers söner , huvudmän för sina familjer , utvalda tappra stridsmän , huvudmän bland hövdingarna ; och de som voro upptecknade i deras släktregister såsom dugliga till krigstjänst utgjorde ett antal av tjugusex tusen man .
och Benjamin födde Bela , sin förstfödde , Asbel , den andre , och Ahara , den tredje ,
Noha , den fjärde , och Rafa , den femte .
Bela hade följande söner : Addar , Gera , Abihud ,
Abisua , Naaman , Ahoa ,
gera , Sefufan och Huram .
och dessa voro Ehuds söner , och de voro familjehuvudmän för dem som bodde i Geba , och som blevo bortförda till Manahat ,
dit Gera jämte Naaman och Ahia förde bort dem : han födde Ussa och Ahihud .
och Saharaim födde barn i Moabs land , sedan han hade skilt sig från sina hustrur , Husim och Baara ;
med sin hustru Hodes födde han där Jobab , Sibja , Mesa , Malkam ,
Jeus , Sakeja och Mirma . dessa voro hans söner , huvudmän för familjer .
med Husim hade han fött Abitub och Elpaal .
och Elpaals söner voro Eber , Miseam och Semed . han var den som byggde Ono och Lod med underlydande orter .
Beria och Sema -- vilka voro familjehuvudmän för Ajalons invånare och förjagade Gats invånare --
så ock Ajo , Sasak och Jeremot .
och Sebadja , Arad , Eder ,
Mikael , Jispa och Joha voro Berias söner .
och Sebadja , Mesullam , Hiski , Heber ,
Jismerai , Jislia och Jobab voro Elpaals söner .
och Jakim , Sikri , Sabdi ,
Elienai , Silletai , Eliel ,
Adaja , Beraja och Simrat voro Simeis söner .
och Jispan , Eber , Eliel ,
Abdon , Sikri , Hanan ,
Hananja , Elam , Antotja ,
Jifdeja och Peniel voro Sasaks söner .
och Samserai , Seharja , Atalja ,
Jaaresja , Elia och Sikri voro Jerohams söner .
dessa vore huvudman för familjer , huvudmän efter sin ättföljd ; de bodde i Jerusalem .
i Gibeon bodde Gibeons fader , vilkens hustru hette Maaka .
och hans förstfödde son var Abdon ; vidare Sur , Kis , Baal , Nadab ,
Gedor , Ajo och Seker .
men Miklot födde Simea . också dessa bodde jämte sina bröder i Jerusalem , gent emot sina bröder .
och Ner födde Kis , Kis födde Saul , och Saul födde Jonatan , Malki @-@ Sua , Abinadab och Esbaal .
Jonatans son var Merib @-@ Baal , och Merib @-@ Baal födde Mika .
Mikas söner voro Piton , Melek , Taarea och Ahas .
Ahas födde Joadda , Joadda födde Alemet , Asmavet och Simri , och Simri födde Mosa .
Mosa födde Binea . hans son var Rafa ; hans son var Eleasa ; hans son var Asel .
och Asel hade sex söner , och dessa hette Asrikam , Bokeru , Ismael , Searja , Obadja och Hanan . alla dessa voro Asels söner .
och hans broder Eseks söner voro Ulam , hans förstfödde , Jeus , den andre , och Elifelet , den tredje .
och Ulams söner voro tappra stridsmän , som voro skickliga i att spänna båge ; och de hade många söner och sonsöner : ett hundra femtio . alla dessa voro av Benjamins barn
och hela Israel blev upptecknat i släktregister , och de finnas uppskrivna i boken om Israels konungar . och Juda fördes i fångenskap bort till Babel för sin otrohets skull .
men de förra invånarna som bodde där de hade sin arvsbesittning , i sina städer , utgjordes av vanliga israeliter , präster , leviter och tempelträlar .
i Jerusalem bodde en del av Juda barn , av Benjamins barn och av Efraims och Manasse barn , nämligen :
Utai , son till Ammihud , son till Omri , son till Imri , son till Bani , av Peres &apos; , Judas sons , barn ;
av siloniterna Asaja , den förstfödde , och hans söner ;
av Seras barn Jeguel och deras broder , sex hundra nittio ;
av Benjamins barn Sallu , son till Mesullam , son till Hodauja , son till Hassenua ,
vidare Jibneja , Jerohams son , och Ela , son till Ussi , son till Mikri , och Mesullam , son till Sefatja , son till Reguel , son till Jibneja ,
så ock deras bröder , efter deras ättföljd , nio hundra femtiosex . alla dessa män voro huvudmän för familjer , var och en för sin familj .
och av prästerna : Jedaja , Jojarib och Jakin ,
vidare Asarja , son till Hilkia , son till Mesullam , son till Sadok , son till Merajot , son till Ahitub , fursten i Guds hus ,
vidare Adaja , son till Jeroham , son till Pashur , son till Malkia , vidare Maasai , son till Adiel , son till Jasera , son till Mesullam , son till Mesillemit , son till Immer ,
så ock deras bröder , huvudmän för sina familjer , ett tusen sju hundra sextio , dugande män i de sysslor som hörde till tjänstgöringen i Guds hus .
och av leviterna : Semaja , som till Hassub , son till Asrikam , son till Hasabja , av Meraris barn ,
vidare Bakbackar , Heres och Galal , så ock Mattanja , son till Mika , son till Sikri , son till Asaf ,
vidare Obadja , son till Semaja , son till Galal , son till Jedutun , så ock Berekja , son till Asa , son till Elkana , som bodde i netofatiternas byar .
och dörrvaktarna : Sallum , Ackub , Talmon och Ahiman med sina bröder ; men Sallum var huvudmannen .
och ända till nu göra de tjänst vid Konungsporten , på östra sidan . dessa voro dörrvaktarna i Levi barns läger .
men Sallum , son till Kore , son till Ebjasaf , son till Kora , hade jämte sina bröder , dem som voro av hans familj , koraiterna , till tjänstgöringssyssla att hålla vakt vid tältets trösklar ; deras fäder hade nämligen i HERRENS läger hållit vakt vid ingången .
och Pinehas , Eleasars son , hade förut varit furste över dem -- med honom vare HERREN !
Sakarja , Meselemjas son , var dörrvaktare vid ingången till uppenbarelsetältet .
alla dessa voro utvalda till dörrvaktare vid trösklarna : två hundra tolv . de blevo i sina byar upptecknade i släktregistret . David och siaren Samuel hade tillsatt dem att tjäna på heder och tro .
de och deras söner stodo därför vid portarna till HERRENS hus , tälthuset , och höllo vakt .
efter de fyra väderstrecken hade dörrvaktarna sina platser : i öster , väster , norr och söder .
och deras bröder , de som fingo bo i sina byar , skulle var sjunde dag , alltid på samma timme , infinna sig hos dem .
ty på heder och tro voro dessa fyra anställda såsom förmän för dörrvaktarna . detta var nu leviterna . de hade ock uppsikten över kamrarna och förvaringsrummen i Guds hus .
och de vistades om natten runt omkring Guds hus , ty dem ålåg att hålla vakt , och de skulle öppna dörrarna var morgon .
somliga av dem hade uppsikten över de kärl som användes vid tjänstgöringen . de buro nämligen in dem , efter att hava räknat dem , och buro sedan ut dem , efter att åter hava räknat dem .
och somliga av dem voro förordnade till att hava uppsikten över de andra kärlen , över alla andra helgedomens kärl , så ock över det fina mjölet och vinet och oljan och rökelsen och de välluktande kryddorna .
men somliga av prästernas söner beredde salvan av de välluktande kryddorna .
och Mattitja , en av leviterna , koraiten Sallums förstfödde , hade på heder och tro uppsikten över bakverket .
och somliga av deras bröder , kehatiternas söner , hade uppsikten över skådebröden och skulle tillreda dem för var sabbat .
men de andra , nämligen sångarna , huvudmän för levitiska familjer , vistades i kamrarna , fria ifrån annan tjänstgöring , ty dag och natt voro de upptagna av sina egna sysslor .
dessa voro huvudmännen för de levitiska familjerna , huvudman efter sin ättföljd ; de bodde i Jerusalem .
i Gibeon bodde Gibeons fader Jeguel , vilkens hustru hette Maaka .
och hans förstfödde son var Abdon ; vidare Sur , Kis , Baal , Ner , Nadab
Gedor , Ajo , Sakarja och Miklot .
men Miklot födde Simeam . också de bodde jämte sina bröder i Jerusalem , gent emot sina bröder .
och Ner födde Kis , Kis födde Saul , och Saul födde Jonatan , Malki @-@ Sua , Abinadab och Esbaal .
Jonatans son var Merib @-@ Baal , och Merib @-@ Baal födde Mika .
Mikas söner voro Piton , Melek och Taharea .
Ahas födde Jaera , Jaera födde Alemet , Asmavet och Simri , och Simri födde Mosa .
Mosa födde Binea . hans son var Refaja ; hans son var Eleasa ; hans son var Asel .
och Asel hade sex söner , och dessa hette Asrikam , Bokeru , Ismael , Searja , Obadja och Hanan . dessa voro Asels söner
och filistéerna stridde mot Israel ; och Israels män flydde för filistéerna och föllo slagna på berget Gilboa .
och filistéerna ansatte ivrigt Saul och hans söner . och filistéerna dödade Jonatan , Abinadab och Malki @-@ Sua , Sauls söner .
när då Saul själv blev häftigt anfallen och bågskyttarna kommo över honom , greps han av förskräckelse för skyttarna .
och Saul sade till sin vapendragare : &quot; drag ut ditt svärd och genomborra mig därmed , så att icke dessa oomskurna komma och hantera mig skändligt &quot; . men hans vapendragare ville det icke , ty han fruktade storligen . då tog Saul själv svärdet och störtade sig därpå .
men när vapendragaren såg att Saul var död , störtade han sig ock på sitt svärd och dog .
så dogo då Saul och hans tre söner ; och alla som hörde till hans hus dogo på samma gång .
och när alla israeliterna i dalen förnummo att deras här hade flytt , och att Saul och hans söner voro döda , övergåvo de sina städer och flydde ; sedan kommo filistéerna och bosatte sig i dem .
dagen därefter kommo filistéerna för att plundra de slagna och funno då Saul och hans söner , där de lågo fallna på berget Gilboa .
och de plundrade honom och togo med sig hans huvud och hans vapen och sände dem omkring i filistéernas land och läto förkunna det glada budskapet för sina avgudar och för folket .
och de lade hans vapen i sitt gudahus , men hans huvudskål hängde de upp i Dagons tempel .
men när allt folket i Jabes i Gilead hörde allt vad filistéerna hade gjort med Saul ,
stodo de upp , alla stridbara män , och togo Sauls och hans söners lik och förde dem till Jabes ; och de begrovo deras ben under terebinten i Jabes och fastade så i sju dagar .
detta blev Sauls död , därför att han hade begått otrohet mot HERREN , i det att han icke hade hållit HERRENS ord , så ock därför att han hade frågat en ande och sökt svar hos en sådan .
han hade icke sökt svar hos HERREN ; därför dödade HERREN honom . och sedan överflyttade han konungadömet på David , Isais son .
då församlade sig hela Israel till David i Hebron och sade : &quot; vi äro ju ditt kött och ben .
redan för länge sedan , redan då Saul ännu var konung , var det du som var ledare och anförare för Israel . och till dig har HERREN , din Gud , sagt : du skall vara en herde för mitt folk Israel , ja , du skall vara en furste över mitt folk Israel &quot; .
när så alla de äldste i Israel kommo till konungen i Hebron , slöt David ett förbund med dem där i Hebron , inför HERREN ; och sedan smorde de David till konung över Israel , i enlighet med HERRENS ord genom Samuel .
och David drog med hela Israel till Jerusalem , det är Jebus ; där befunno sig jebuséerna , som ännu bodde kvar i landet .
och invånarna i Jebus sade till David : &quot; hitin kommer du icke &quot; . men David intog likväl Sions borg , det är Davids stad
och David sade : &quot; vemhelst som först slår ihjäl en jebusé , han skall bliva hövding och anförare &quot; . och Joab , Serujas son , kom först ditupp och blev så hövding .
sedan tog David sin boning i bergfästet ; därför kallade man det Davids stad .
och han uppförde befästningsverk runt omkring staden , från Millo och allt omkring ; och Joab återställde det övriga av staden .
och David blev allt mäktigare och mäktigare , och HERREN Sebaot var med honom
och dessa äro de förnämsta bland Davids hjältar , vilka gåvo honom kraftig hjälp att bliva konung , de jämte hela Israel , och så skaffade honom konungaväldet , enligt HERRENS ord angående Israel .
detta är förteckningen på Davids hjältar : Jasobeam , son till en hakmonit , den förnämste bland kämparna , han som svängde sitt spjut över tre hundra som hade blivit slagna på en gång .
och efter honom kom ahoaiten Eleasar , son till Dodo ; han var en av de tre hjältarna .
han var med David vid Pas @-@ Dammim , när filistéerna där hade församlat sig till strid . och där var ett åkerstycke , fullt med korn . och folket flydde för filistéerna .
då ställde de sig mitt på åkerstycket och försvarade det och slogo filistéerna ; och HERREN lät dem så vinna en stor seger .
en gång drogo tre av de trettio förnämsta männen ned över klippan till David vid Adullams grotta , medan en avdelning filistéer var lägrad i Refaimsdalen .
men David var då på borgen , under det att en filisteisk utpost fanns i Bet @-@ Lehem .
och David greps av lystnad och sade : &quot; Ack att någon ville giva mig vatten att dricka från brunnen vid Bet @-@ Lehems stadsport ! &quot;
då bröto de tre sig igenom filistéernas läger och hämtade vatten ur brunnen vid Bet @-@ Lehems stadsport och togo det och buro det till David . men David ville icke dricka det , utan göt ut det såsom ett drickoffer åt HERREN .
han sade nämligen : &quot; Gud låte det vara fjärran ifrån mig att jag skulle göra detta ! skulle jag dricka dessa mäns blod , som hava vågat sina liv ? ty med fara för sina liv hava de burit det hit &quot; . och han ville icke dricka det . sådana ting hade de tre hjältarna gjort .
Absai , Joabs broder , var den förnämste av tre andra ; han svängde en gång sitt spjut över tre hundra som hade blivit slagna . och han hade ett stort namn bland de tre .
han var dubbelt mer ansedd än någon annan i detta tretal , och han var deras hövitsman , men upp till de tre första kom han dock icke .
vidare Benaja , son till Jojada , som var son till en tapper , segerrik man från Kabseel ; han slog ned de två Arielerna i Moab , och det var han som en snövädersdag steg ned och slog ihjäl lejonet i brunnen .
han slog ock ned den egyptiske mannen som var så reslig : fem alnar lång . fastän egyptiern i handen hade ett spjut som liknade en vävbom , gick han ned mot honom , väpnad allenast med sin stav . och han ryckte spjutet ur egyptiern hand och dräpte honom med hans eget spjut .
sådana ting hade Benaja , Jojadas son , gjort . och han hade ett stort namn bland de tre hjältarna .
ja , han var mer ansedd än någon av de trettio , men upp till de tre första kom han icke . och David satte honom till anförare för sin livvakt .
de tappra hjältarna voro : Asael , Joabs broder , Elhanan , Dodos son , från Bet @-@ Lehem ;
haroriten Sammot ; peloniten Heles ;
tekoaiten Ira , Ickes &apos; son ; anatotiten Abieser ;
husatiten Sibbekai ; ahoaiten Ilai ;
netofatiten Maherai ; netofatiten Heled , Baanas son ;
Itai , Ribais son , från Gibea i Benjamins barns stam ; pirgatoniten Benaja ;
Hurai från Gaas &apos; dalar ; arabatiten Abiel ;
baharumiten Asmavet ; saalboniten Eljaba ;
gisoniten Bene @-@ Hasem ; harariten Jonatan , Sages son ;
harariten Ahiam , Sakars son ; Elifal , Urs son ;
mekeratiten Hefer ; peloniten Ahia ;
Hesro från Karmel ; Naarai , Esbais son ;
Joel , broder till Natan ; Mibhar , Hagris son ;
ammoniten Selek ; berotiten Naherai , vapendragare åt Joab , Serujas son ;
jeteriten Ira ; jeteriten Gareb ;
hetiten Uria ; Sabad , Alais son ;
rubeniten Adina , Sisas son , en huvudman bland rubeniterna , och jämte honom trettio andra ;
Hanan , Maakas son , och mitniten Josafat ;
astarotiten Ussia ; Sama och Jeguel , aroeriten Hotams söner ;
Jediael , Simris son , och hans broder Joha , tisiten ;
Eliel @-@ Hammahavim samt Jeribai och Josauja , Elnaams söner , och moabiten Jitma ;
slutligen Eliel , Obed och Jaasiel @-@ Hammesobaja .
och dessa voro de som kommo till David i Siklag , medan han ännu höll sig undan för Saul , Kis &apos; son ; de hörde till de hjältar som bistodo honom under kriget .
de voro väpnade med båge och skickliga i att , både med höger och med vänster hand , slunga stenar och avskjuta pilar från bågen . av Sauls stamfränder , benjaminiterna , kommo :
Ahieser , den förnämste , och Joas , gibeatiten Hassemaas söner ; Jesuel och Pelet , Asmavets söner ; Beraka ; anatotiten Jehu ;
gibeoniten Jismaja , en av de trettio hjältarna , anförare för de trettio ; Jeremia ; Jahasiel ; Johanan ; gederatiten Josabad ;
Eleusai ; Jerimot ; Bealja ; Semarja ; harufiten Sefatja ;
koraiterna Elkana , Jissia , Asarel , Joeser och Jasobeam ;
Joela och Sebadja , söner till Jeroham , av strövskaran .
och av gaditerna avföllo några och gingo till David i bergfästet i öknen , tappra män , krigsmän skickliga att strida , rustade med sköld och spjut ; de hade en uppsyn såsom lejon och voro snabba såsom gaseller på bergen :
Eser , den förnämste , Obadja , den andre , Eliab , den tredje ,
Masmanna , den fjärde , Jeremia , den femte ,
Attai , den sjätte , Eliel , den sjunde ,
Johanan , den åttonde , Elsabad , den nionde ,
Jeremia , den tionde , Makbannai , den elfte .
dessa hörde till Gads barn och till de förnämsta i hären ; den ringaste av dem var ensam så god som hundra , men den ypperste så god som tusen .
dessa voro de som i första månaden gingo över Jordan , när den var full över alla sina bräddar , och som förjagade alla dem som bodde i dalarna , åt öster och åt väster .
av Benjamins och Juda barn kommo några män till David ända till bergfästet .
då gick David ut emot dem och tog till orda och sade till dem : &quot; om I kommen till mig i fredlig avsikt och viljen bistå mig , så är mitt hjärta redo till förening med eder ; men om I kommen för att förråda mig åt mina ovänner , fastän ingen orätt är i mina händer , då må våra fäders Gud se därtill och straffa det &quot; .
men Amasai , den förnämste bland de trettio , hade blivit beklädd med andekraft , och han sade : &quot; dina äro vi , David , och med dig stå vi , du Isais son . frid vare med dig , frid , och frid vare med dem som bistå dig ty din Gud har bistått dig ! &quot; och David tog emot dem och gav dem plats bland de förnämsta i sin skara .
från Manasse gingo några över till David , när han med filistéerna drog ut i strid mot Saul , dock fingo de icke bistå dessa ; ty när filistéernas hövdingar hade rådplägat , skickade de bort honom , i det de sade : &quot; det gäller huvudet för oss , om han går över till sin herre Saul .
när han då drog till Siklag , gingo dessa från Manasse över till honom : Adna , Josabad , Jediael , Mikael , Josabad , Elihu och Silletai , huvudmän för de ätter som tillhörde Manasse .
dessa bistodo David mot strövskaran , ty de voro allasammans tappra stridsmän och blevo hövitsmän i hären .
dag efter dag kommo nämligen allt flera till David för att bistå honom , så att hans läger blev övermåttan stort .
detta är de tal som angiva summorna av det väpnade krigsfolk som kom till David i Hebron , för att efter HERRENS befallning flytta Sauls konungamakt över på honom :
Juda barn , som buro sköld och spjut , sex tusen åtta hundra , väpnade till strid ;
av Simeons barn tappra krigsmän , sju tusen ett hundra ;
av Levi barn fyra tusen sex hundra ;
därtill Jojada , fursten inom Arons släkt , och med honom tre tusen sju hundra ;
så ock Sadok , en tapper yngling , med sin familj , tjugutvå hövitsmän ;
av Benjamins barn , Sauls stamfränder , tre tusen ( ty ännu vid den tiden höllo de flesta av dem troget med Sauls hus ) ;
av Efraims barn tjugu tusen åtta hundra , tappra stridsmän , namnkunniga män i sina familjer ;
av ena hälften av Manasse stam aderton tusen namngivna män , som kommo för att göra David till konung ;
av Isaskars barn kommo män som väl förstodo tidstecknen och insågo vad Israel borde göra , två hundra huvudmän , därtill alla deras stamfränder under deras befäl ;
av Sebulon stridbara män , rustade till krig med alla slags vapen , femtio tusen , som samlades endräktigt ;
av Naftali ett tusen hövitsmän , och med dem trettiosju tusen , väpnade med sköld och spjut ;
av daniterna krigsrustade män , tjuguåtta tusen sex hundra ;
av Aser stridbara män , rustade till krig , fyrtio tusen ;
och från andra sidan Jordan , av rubeniterna , gaditerna och andra hälften av Manasse stam , ett hundra tjugu tusen , väpnade med alla slags vapen som brukas vid krigföring .
alla dessa krigsmän , ordnade till strid , kommo i sina hjärtans hängivenhet till Hebron för att göra David till konung över hela Israel . också hela det övriga Israel var enigt i att göra David till konung .
och de voro där hos David i tre dagar och åto och drucko , ty deras bröder hade försett dem med livsmedel .
de som bodde närmast dem , ända upp till Isaskar , Sebulon och Naftali , tillförde dem ock på åsnor , kameler , mulåsnor och oxar livsmedel i myckenhet till föda : mjöl , fikonkakor och russinkakor , vin och olja , fäkreatur och småboskap ; ty glädje rådde i Israel .
och David rådförde sig med över- och underhövitsmännen , med alla furstarna .
sedan sade David till Israels hela församling : &quot; om I så finnen för gott , och om detta är från HERREN , vår Gud , så låt oss sända bud åt alla håll till våra övriga bröder i alla Israels landsändar , och därjämte till prästerna och leviterna i de städer kring vilka de hava sina utmarker , att de må församla sig till oss ;
och låt oss flytta vår Guds ark till oss , ty i Sauls tid frågade vi icke efter den &quot; .
och hela församlingen svarade att man skulle göra så , ty förslaget behagade hela folket .
så församlade då David hela Israel , från Sihor i Egypten ända dit där vägen går till Hamat , för att hämta Guds ark från Kirjat @-@ Jearim .
och David drog med hela Israel upp till Baala , det är Kirjat @-@ Jearim , som hör till Juda , för att därifrån föra upp Guds , HERRENS , ark , hans som tronar på keruberna , och efter vilken den hade fått sitt namn .
och de satte Guds ark på en ny vagn och förde den bort ifrån Abinadabs hus ; och Ussa och Ajo körde vagnen .
och David och hela Israel fröjdade sig inför Gud av all makt , med sånger och med harpor , psaltare , pukor , cymbaler och trumpeter .
men när de kommo till Kidonslogen , räckte Ussa ut sin hand för att Fatta I arken , ty oxarna snavade .
då upptändes HERRENS vrede mot Ussa , och därför att han hade räckt ut sin hand mot arken , slog han honom , så att han föll ned död där inför Gud .
men det gick David hårt till sinnes att HERREN så hade brutit ned Ussa ; och han kallade det stället Peres @-@ Ussa , såsom det heter ännu i dag .
och David betogs av sådan fruktan för Gud på den dagen , att han sade : &quot; huru skulle jag töras låta föra Guds ark till mig ? &quot;
därför lät David icke flytta in arken till sig i Davids stad , utan lät sätta in den i gatiten Obed @-@ Edoms hus .
sedan blev Guds ark kvar vid Obed @-@ Edoms hus , där den stod i sitt eget hus , i tre månader ; men HERREN välsignade Obed @-@ Edoms hus och allt vad som hörde honom till .
och Hiram , konungen i Tyrus , skickade sändebud till David med cederträ , därjämte ock murare och timmermän , för att de skulle bygga honom ett hus .
och David märkte att HERREN hade befäst honom såsom konung över Israel ; ty han hade låtit hans rike bliva övermåttan upphöjt , för sitt folk Israels skull .
och David tog sig ännu flera hustrur i Jerusalem , och David födde ännu flera söner och döttrar .
dessa äro namnen på de söner som han fick i Jerusalem : Sammua , Sobab , Natan , Salomo ,
Jibhar , Elisua , Elpelet ,
noga , Nefeg , Jafia ,
Elisama , Beeljada och Elifelet .
men när filistéerna hörde att David hade blivit smord till konung över hela Israel , drogo de allasammans upp för att fånga David . när David hörde detta , drog han ut mot dem .
då nu filistéerna hade fallit in i Refaimsdalen och där företogo plundringståg ,
frågade David Gud : &quot; skall jag draga upp mot filistéerna ? vill du då giva dem i min hand ? &quot; HERREN svarade honom : &quot; drag upp ; jag vill giva dem i din hand &quot; .
och de drogo upp till Baal @-@ Perasim , och där slog David dem . då sade David : &quot; Gud har brutit ned mina fiender genom min hand , likasom en vattenflod bryter ned &quot; . därav fick det stället namnet Baal @-@ Perasim .
de lämnade där efter sig sina gudar ; och David befallde att dessa skulle brännas upp i eld .
men filistéerna företogo ännu en gång plundringståg i dalen .
när David då åter frågade Gud , svarade Gud honom : &quot; du skall icke draga upp efter dem ; du må kringgå dem på en omväg , så att du kommer över dem från det håll där bakaträden stå .
så snart du sedan hör ljudet av steg i bakaträdens toppar , drag då ut till strid , ty då har Gud dragit ut framför dig till att slå filistéernas här &quot; .
David gjorde såsom Gud hade bjudit honom ; och de slogo filistéernas här och förföljde dem från Gibeon ända till Geser .
och ryktet om David gick ut i alla länder , och HERREN lät fruktan för honom komma över alla folk .
och han uppförde åt sig hus i Davids stad ; sedan beredde han en plats åt Guds ark och slog upp ett tält åt den .
därvid befallde David : &quot; inga andra än leviterna må bära Guds ark ; ty dem har HERREN utvalt till att bära Guds ark och till att göra tjänst inför honom för evärdlig tid &quot; .
och David församlade hela Israel till Jerusalem för att hämta HERRENS ark upp till den plats som han hade berett åt den .
och David samlade tillhopa Arons barn och leviterna ;
av Kehats barn : Uriel , deras överste , och hans bröder , ett hundra tjugu ;
av Meraris barn : Asaja , deras överste , och hans bröder , två hundra tjugu ;
av Gersoms barn : Joel , deras överste , och hans bröder , ett hundra trettio ;
av Elisafans barn : Semaja , deras överste , och hans bröder , två hundra ;
av Hebrons barn : Eliel , deras överste , och hans bröder , åttio ;
av Ussiels barn : Amminadab , deras överste , och hans bröder , ett hundra tolv .
och David kallade till sig prästerna Sadok och Ebjatar jämte leviterna Uriel , Asaja , Joel , Semaja , Eliel och Amminadab .
och han sade till dem : &quot; i ären huvudmän för leviternas familjer . Helgen eder tillika med edra bröder , och hämten så HERRENS , Israels Guds , ark upp till den plats som jag har berett åt den .
ty därför att I förra gången icke voren tillstädes var det som HERREN , vår Gud , bröt ned en av oss , till straff för att vi icke sökte honom så , som tillbörligt var &quot; .
då helgade prästerna och leviterna sig till att hämta upp HERRENS , Israels Guds , ark .
och såsom Mose hade bjudit i enlighet med HERRENS ord , buro nu Levi barn Guds ark med stänger , som vilade på deras axlar .
och David sade till de översta bland leviterna att de skulle förordna sina bröder sångarna till tjänstgöring med musikinstrumenter , psaltare , harpor och cymbaler , som de skulle låta ljuda , under det att de höjde glädjesången .
leviterna förordnade då Heman , Joels son , och av hans bröder Asaf , Berekjas son , och av dessas bröder , Meraris barn , Etan , Kusajas son ,
och jämte dem deras bröder av andra ordningen Sakarja , Ben , Jaasiel , Semiramot , Jehiel , Unni , Eliab , Benaja , Maaseja , Mattitja , Elifalehu , Mikneja , Obed @-@ Edom och Jegiel , dörrvaktarna .
och sångarna , Heman , Asaf och Etan , skulle slå kopparcymbaler .
Sakarja , Asiel , Semiramot , Jehiel , Unni , Eliab , Maaseja och Benaja skulle spela på psaltare , till Alamót .
Mattitja , Elifalehu , Mikneja , Obed @-@ Edom , Jegiel och Asasja skulle leda sången med harpor , till Seminit .
Kenanja , leviternas anförare , när de buro , skulle undervisa i att bära , ty han var kunnig i sådant .
Berekja och Elkana skulle vara dörrvaktare vid arken .
Sebanja , Josafat , Netanel , Amasai , Sakarja , Benaja och Elieser , prästerna , skulle blåsa i trumpeter framför Guds ark . slutligen skulle Obed @-@ Edom och Jehia vara dörrvaktare vid arken .
så gingo då David och de äldste i Israel och överhövitsmännen åstad för att hämta HERRENS förbundsark upp ur Obed @-@ Edoms hus , under jubel .
och då Gud skyddade leviterna som buro HERRENS förbundsark , offrade man sju tjurar och sju vädurar .
därvid var David klädd i en kåpa av fint linne ; så voro ock alla leviterna som buro arken , så ock sångarna och Kenanja , som anförde sångarna , när de buro . och därjämte bar David en linne @-@ efod .
och hela Israel hämtade upp HERRENS förbundsark under jubel och basuners ljud ; och man blåste i trumpeter och slog cymbaler och lät psaltare och harpor ljuda .
när då HERRENS förbundsark kom till Davids stad , blickade Mikal , Sauls dotter , ut genom fönstret , och då hon såg konung David dansa och göra sig glad , fick hon förakt för honom i sitt hjärta .
sedan de hade fört Guds ark ditin , ställde de den i tältet som David hade slagit upp åt den , och framburo därefter brännoffer och tackoffer inför Guds ansikte .
när David hade offrat brännoffret och tackoffret , välsignade han folket i HERRENS namn .
och åt var och en av alla israeliterna , både man och kvinna , gav han en kaka bröd , ett stycke kött och en druvkaka .
och han förordnade vissa leviter till att göra tjänst inför HERRENS ark , för att de skulle prisa , tacka och lova HERREN , Israels Gud :
Asaf såsom anförare , näst efter honom Sakarja , och vidare Jegiel , Semiramot , Jehiel , Mattitja , Eliab , Benaja , Obed @-@ Edom och Jegiel med psaltare och harpor ; och Asaf skulle slå cymbaler .
men prästerna Benaja och Jahasiel skulle beständigt stå med sina trumpeter framför Guds förbundsark .
på den dagen var det som David först fastställde den ordningen att man genom Asaf och hans bröder skulle tacka HERREN på detta sätt :
&quot; Tacken HERREN , åkallen hans namn , gören hans gärningar kunniga bland folken .
sjungen till hans ära , lovsägen honom , talen om alla hans under .
Berömmen eder av hans heliga namn ; glädje sig av hjärtat de som söka HERREN .
frågen efter HERREN och hans makt , söken hans ansikte beständigt .
Tänken på de underbara verk som han har gjort , på hans under och hans muns domar ,
i Israels , hans tjänares , säd , I Jakobs barn , hans utvalda .
han är HERREN , vår Gud ; över hela jorden gå hans domar .
Tänken evinnerligen på hans förbund , intill tusen släkten på vad han har stadgat ,
på det förbund han slöt med Abraham och på hans ed till Isak .
han fastställde det för Jakob till en stadga , för Israel till ett evigt förbund ;
han sade : &apos; åt dig vill jag giva Kanaans land , det skall bliva eder arvedels lott . &apos;
då voren I ännu en liten hop , I voren ringa och främlingar därinne .
och de vandrade åstad ifrån folk till folk ifrån ett rike bort till ett annat .
han tillstadde ingen att göra dem skada , han straffade konungar för deras skull :
&apos; kommen icke vid mina smorda , och gören ej mina profeter något ont . &apos;
sjungen till HERRENS ära , alla länder , båden glädje var dag , förkunnen hans frälsning .
förtäljen bland hedningarna hans ära , bland alla folk hans under .
ty stor är HERREN och högt Lovad , och fruktansvärd är han mer än alla gudar .
ty folkens alla gudar äro avgudar , men HERREN är den som har gjort himmelen .
Majestät och härlighet äro inför hans ansikte , makt och fröjd i hans boning .
given åt HERREN , I folkens släkter , given åt HERREN ära och makt ;
given åt HERREN hans namns ära , bären fram skänker och kommen inför hans ansikte , tillbedjen HERREN i helig skrud .
Bäven för hans ansikte , alla länder ; se , jordkretsen står fast och vacklar icke .
himmelen vare glad , och jorden fröjde sig , och bland hedningarna säge man : &apos; HERREN är nu konung ! &apos;
havet bruse och allt vad däri är , marken glädje sig och allt som är därpå ;
ja , då juble skogens träd inför HERREN , ty han kommer för att döma jorden .
Tacken HERREN , ty han är god , ty hans nåd varar evinnerligen ,
och sägen : &apos; fräls oss , du vår frälsnings Gud , församla oss och rädda oss från hedningarna , så att vi få prisa ditt heliga namn och berömma oss av ditt lov . &apos;
Lovad vare HERREN , Israels Gud , från evighet till evighet ! &quot; och allt folket sade : &quot; Amen &quot; , och lovade HERREN .
och han gav där , inför HERRENS förbundsark , åt Asaf och hans bröder uppdraget att beständigt göra tjänst inför arken , var dag med de för den dagen bestämda sysslorna .
men Obed @-@ Edom och deras bröder voro sextioåtta ; och Obed @-@ Edom , Jedituns son , och Hosa gjorde han till dörrvaktare .
och prästen Sadok och hans bröder , prästerna , anställde han inför HERRENS tabernakel , på offerhöjden i Gibeon ,
för att de beständigt skulle offra åt HERREN brännoffer på brännoffersaltaret , morgon och afton , och göra allt vad som var föreskrivet i HERRENS lag , den som han hade givit åt Israel ;
och jämte dem Heman och Jedutun och de övriga namngivna utvalda , på det att de skulle tacka HERREN , därför att hans nåd varar evinnerligen .
och hos dessa , nämligen Heman och Jedutun , förvarades trumpeter och cymbaler åt dem som skulle spela , så ock andra instrumenter som hörde till gudstjänsten . och Jedutuns söner gjorde han till dörrvaktare .
sedan gick allt folket hem , var och en till sitt ; men David vände om för att hälsa sitt husfolk .
då nu David satt i sitt hus , sade han till profeten Natan : &quot; se , jag bor i ett hus av cederträ , under det att HERRENS förbundsark står under ett tält &quot; .
Natan sade till David : &quot; gör allt vad du har i sinnet ; ty Gud är med dig &quot; .
men om natten kom Guds ord till Natan ; han sade :
&quot; gå och säg till min tjänare David : så säger HERREN : icke du skall bygga mig det hus som jag skall bo i .
jag har ju icke bott i något hus , från den dag då jag förde Israel hitupp ända till denna dag , utan jag har flyttat ifrån tält till tält , ifrån tabernakel till tabernakel .
har jag då någonsin , varhelst jag flyttade omkring med hela Israel , talat och sagt så till någon enda av Israels domare , som jag har förordnat till herde för mitt folk : &apos; Varför haven I icke byggt mig ett hus av cederträ ? &apos;
och nu skall du säga så till min tjänare David : så säger HERREN Sebaot : från betesmarken , där du följde fåren , har jag hämtat dig , för att du skulle bliva en furste över mitt folk Israel .
och jag har varit med dig på alla dina vägar och utrotat alla dina fiender för dig . och jag vill göra dig ett namn , sådant som de störstes namn på jorden .
jag skall bereda en plats åt mitt folk Israel och plantera det , så att det får bo kvar där , utan att vidare bliva oroat . Orättfärdiga människor skola icke mer föröda det , såsom fordom skedde ,
och såsom det har varit allt ifrån den tid då jag förordnade domare över mitt folk Israel ; och jag skall kuva alla dina fiender . så förkunnar jag nu för dig att HERREN skall bygga ett hus åt dig .
ty det skall ske , att när din tid är ute och du går till dina fäder skall jag efter dig upphöja din son , en av dina avkomlingar ; och jag skall befästa hans konungamakt .
han skall bygga ett hus åt mig , och jag skall befästa hans tron för evig tid .
jag skall vara hans fader , och han skall vara min son ; och min nåd skall jag icke låta vika ifrån honom , såsom jag lät den vika ifrån din företrädare .
jag skall hålla honom vid makt i mitt hus och i mitt rike för evig tid , och hans tron skall vara befäst för evig tid &quot; .
alldeles i överensstämmelse med dessa ord och med denna syn talade nu Natan till David .
då gick konung David in och satte sig ned inför HERRENS ansikte och sade : &quot; vem är jag , HERRE Gud , och vad är mitt hus , eftersom du har låtit mig komma härtill ?
och detta har likväl synts dig vara för litet , o Gud ; du har talat angående din tjänares hus om det som ligger långt fram i tiden . ja , du har sett till mig på människosätt , for att upphöja mig , HERRE Gud .
vad skall nu David vidare säga till dig om den ära du har bevisat din tjänare ? du känner ju din tjänare .
herre , för din tjänares skull och efter ditt hjärta har du gjort allt detta stora och förkunnat alla dessa stora ting .
herre , ingen är dig lik , och ingen Gud finnes utom dig , efter allt vad vi hava hört med våra öron .
och var finnes på jorden något enda folk som är likt ditt folk Israel , vilket Gud själv har gått åstad att förlossa åt sig till ett folk -- för att så göra dig ett stort och fruktansvärt namn , i det att du förjagade hedningarna för ditt folk , det som du hade förlossat ifrån Egypten ?
och du har gjort ditt folk Israel till ett folk åt dig för evig tid , och du , HERRE , har blivit deras Gud
så må nu , HERRE , vad du har talat om din tjänare och om hans hus bliva fast för evig tid ; gör såsom du har talat .
då skall ditt namn anses fast och bliva stort till evig tid , så att man skall säga : &apos; HERREN Sebaot , Israels Gud , är Gud över Israel . &apos; och så skall din tjänare Davids hus bestå inför dig .
ty du , min Gud , har uppenbarat för din tjänare att du skall bygga honom ett hus ; därför har din tjänare dristat att bedja inför dig .
och nu , HERRE , du är Gud ; och då du har lovat din tjänare detta goda ,
så må du nu ock värdigas välsigna din tjänares hus , så att det förbliver evinnerligen inför dig . ty vad du , HERRE , välsignar , det är välsignat evinnerligen &quot; .
en tid härefter slog David filistéerna och kuvade dem . därvid tog han Gat med underlydande orter ur filistéernas hand .
han slog ock moabiterna ; så blevo moabiterna David underdåniga och förde till honom skänker .
likaledes slog David Hadareser , konungen i Soba , vid Hamat , när denne hade dragit åstad för att befästa sitt välde vid floden Frat .
och David tog ifrån honom ett tusen vagnar och tog till fånga sju tusen ryttare och tjugu tusen man fotfolk ; och David lät avskära fotsenorna på alla vagnshästarna , utom på ett hundra hästar , som han skonade .
när sedan araméerna från Damaskus kommo för att hjälpa Hadareser , konungen i Soba , nedgjorde David tjugutvå tusen man av dem .
och David insatte fogdar bland araméerna i Damaskus ; och araméerna blevo David underdåniga och förde till honom skänker . så gav HERREN seger åt David , varhelst han drog fram .
och David tog de gyllene sköldar som Hadaresers tjänare hade burit och förde dem till Jerusalem .
och från Hadaresers städer Tibhat och Kun tog David koppar i stor myckenhet ; därav gjorde sedan Salomo kopparhavet , pelarna och kopparkärlen .
då nu Tou , konungen i Hamat , hörde att David hade slagit Hadaresers , konungens i Soba , hela här ,
sände han sin son Hadoram till konung David för att hälsa honom och lyckönska honom , därför att han hade givit sig i strid med Hadareser och slagit honom ; ty Hadareser hade varit Tous fiende . han sände ock alla slags kärl av guld , silver och koppar .
också dessa helgade konung David åt HERREN , likasom han hade gjort med det silver och guld han hade hemfört från alla andra folk : från edoméerna , moabiterna , Ammons barn , filistéerna och amalekiterna .
och sedan Absai , Serujas son , hade slagit edoméerna i Saltdalen , aderton tusen man ,
insatte han fogdar i Edom ; och alla edoméer blevo David underdåniga . så gav HERREN seger åt David , varhelst han drog fram .
David regerade nu över hela Israel ; och han skipade lag och rätt åt allt sitt folk .
Joab , Serujas son , hade befälet över krigshären , och Josafat , Ahiluds son , var kansler .
Sadok , Ahitubs son , och Abimelek , Ebjatars son , voro präster , och Sausa var sekreterare .
Benaja , Jojadas son , hade befälet över keretéerna och peletéerna ; men Davids söner voro de förnämste vid konungens sida .
en tid härefter dog Nahas , Ammons barns konung , och hans son blev konung efter honom .
då sade David : &quot; jag vill bevisa Hanun , Nahas &apos; son , vänskap , eftersom hans fader bevisade mig vänskap &quot; . och David skickade sändebud för att trösta honom i hans sorg efter fadern . när så Davids tjänare kommo till Ammons barns land , till Hanun , för att trösta honom ,
sade Ammons barns furstar till Hanun : &quot; Menar du att David därmed att han sänder tröstare till dig vill visa dig att han ärar din fader ? Nej , för att undersöka och fördärva och bespeja landet hava hans tjänare kommit till dig &quot; .
då tog Hanun Davids tjänare och lät raka dem och skära av deras kläder mitt på , ända uppe vid sätet , och lät dem så gå .
och man kom och berättade för David vad som hade hänt männen ; då sände han bud emot dem , ty männen voro ju mycket vanärade . och konungen lät säga : &quot; stannen i Jeriko , till dess edert skägg hinner växa ut , och kommen så tillbaka &quot; .
då nu Ammons barn insågo att de hade gjort sig förhatliga för David , sände Hanun och Ammons barn ett tusen talenter silver för att leja sig vagnar och ryttare från Aram @-@ Naharaim , från Aram @-@ Maaka och från Soba .
de lejde sig trettiotvå tusen vagnar , ävensom hjälp av konungen i Maaka med hans folk ; dessa kommo och lägrade sig framför Medeba . Ammons barn församlade sig ock från sina städer och kommo för att strida .
när David hörde detta , sände han åstad Joab med hela hären , de tappraste krigarna .
och Ammons barn drogo ut och ställde upp sig till strid vid ingången till staden ; men de konungar som hade kommit dit ställde upp sig för sig själva på fältet .
då Joab nu såg att han hade fiender både framför sig och bakom sig , gjorde han ett urval bland allt Israels utvalda manskap och ställde sedan upp sig mot araméerna .
men det övriga folket överlämnade han åt sin broder Absai , och dessa fingo ställa upp sig mot Ammons barn .
och han sade : &quot; om araméerna bliva mig övermäktiga , så skall du komma mig till hjälp ; och om Ammons barn bliva dig övermäktiga , så vill jag hjälpa dig .
var nu vid gott mod ; ja , låt oss visa mod i striden för vårt folk och för vår Guds städer . sedan må HERREN göra vad honom täckes .
därefter ryckte Joab fram med sitt folk till strid mot araméerna , och de flydde för honom .
men när Ammons barn sågo att araméerna flydde , flydde också de för hans broder Absai och begåvo sig in i staden . då begav sig Joab till Jerusalem .
då alltså araméerna sågo att de hade blivit slagna av Israel , sände de bud att de araméer som bodde på andra sidan floden skulle rycka ut , anförda av Sofak , Hadaresers härhövitsman .
när detta blev berättat för David , församlade han hela Israel och gick över Jordan , och då han kom fram till dem , ställde han upp sig i slagordning mot dem ; och när David hade ställt upp sig till strid mot araméerna , gåvo dessa sig i strid med honom .
men araméerna flydde undan för Israel , och David dräpte av araméerna manskapet på sju tusen vagnar , så ock fyrtio tusen man fotfolk ; härhövitsmannen Sofak dödade han ock .
följande år , vid den tid då konungarna plägade draga i fält , tågade Joab ut med krigshären och härjade Ammons barns land , och kom så och belägrade Rabba , medan David stannade kvar i Jerusalem . och Joab intog Rabba och förstörde det .
och David tog deras konungs krona från hans huvud , den befanns väga en talent guld och var prydd med en dyrbar sten . den sattes nu på Davids huvud . och han förde ut byte från staden i stor myckenhet .
och folket därinne förde han ut och söndersargade dem med sågar och tröskvagnar av järn och med bilor . så gjorde David mot Ammons barns alla städer . sedan vände David med allt folket tillbaka till Jerusalem .
därefter uppstod en strid med filistéerna vid Geser ; husatiten Sibbekai slog då ned Sippai , en av rafaéernas avkomlingar ; så blevo de kuvade .
åter stod en strid med filistéerna ; Elhanan , Jaurs son , slog då ned Lami , gatiten Goljats broder , som hade ett spjut vars skaft liknade en vävbom .
åter stod en strid vid Gat . där var en reslig man som hade sex fingrar och sex tår , tillsammans tjugufyra ; han var ock en avkomling av rafaéerna .
denne smädade Israel ; då blev han nedgjord av Jonatan , son till Simea , Davids broder .
dessa voro avkomlingar av rafaéerna i Gat ; och de föllo för Davids och hans tjänares hand .
men Satan trädde upp mot Israel och uppeggade David till att räkna Israel .
då sade David till Joab och till folkets andra hövitsman : &quot; Gån åstad och räknen Israel , från Beer @-@ Seba ända till Dan , och given mig besked därom , så att jag får veta huru många de äro &quot; .
Joab svarade : &quot; må HERREN än vidare föröka sitt folk hundrafalt . äro de då icke , min herre konung , allasammans min herres tjänare ? Varför begär då min herre sådant ? Varför skulle man därmed draga skuld över Israel ?
likväl blev konungens befallning gällande , trots Joab . alltså drog Joab ut och for omkring i hela Israel , och kom så hem igen till Jerusalem .
och Joab uppgav för David vilken slutsumma folkräkningen utvisade : i Israel funnos tillsammans elva hundra tusen svärdbeväpnade män , och i Juda funnos fyra hundra sjuttio tusen svärdbeväpnade man .
men Levi och Benjamin hade han icke räknat jämte de andra , ty konungens befallning var en styggelse för Joab .
vad som hade skett misshagade Gud , och han hemsökte Israel .
då sade David till Gud : &quot; jag har syndat storligen däri att jag har gjort detta ; men tillgiv nu din tjänares missgärning , ty jag har handlat mycket dåraktigt &quot; .
men HERREN talade till Gad , Davids siare , och sade :
&quot; gå och tala till David och säg : så säger HERREN : tre ting lägger jag fram för dig ; välj bland dem ut åt dig ett som du vill att jag skall göra dig &quot; .
då gick Gad in till David och sade till honom : &quot; så säger HERREN :
tag vilketdera du vill : antingen hungersnöd i tre år , eller förödelse i tre månader genom dina ovänners anfall , utan att du kan undkomma dina fienders svärd , eller HERRENS svärd och pest i landet under tre dagar , i det att HERRENS ängel sprider fördärv inom hela Israels område . eftersinna nu vilket svar jag skall giva honom som har sänt mig &quot; .
David svarade Gad : &quot; jag är i stor vånda . men låt mig då falla i HERRENS hand , ty hans barmhärtighet är mycket stor ; i människohand vill jag icke falla &quot; .
så lät då HERREN pest komma i Israel , så att sjuttio tusen män av Israel föllo .
och Gud sände en ängel mot Jerusalem till att fördärva det . men när denne höll på att fördärva , såg HERREN därtill och ångrade det onda , så att han sade till ängeln , Fördärvaren : &quot; det är nog ; drag nu din hand tillbaka &quot; . och HERRENS ängel stod då vid jebuséen Ornans tröskplats .
när nu David lyfte upp sina ögon och fick se HERRENS ängel stående mellan jorden och himmelen med ett blottat svärd i sin hand , uträckt över Jerusalem , då föllo han och de äldste , höljda i sorgdräkt , ned på sina ansikten .
och David sade till Gud : &quot; det var ju jag som befallde att folket skulle räknas . det är då jag som har syndat och gjort vad ont är ; men dessa , min hjord , vad hava de gjort ? herre , min Gud , må din hand vända sig mot mig och min faders hus , men icke mot ditt folk , så att det bliver hemsökt &quot; .
men HERRENS ängel befallde Gad att säga till David att David skulle gå åstad och resa ett altare åt HERREN på jebuséen Ornans tröskplats .
och David gick åstad på grund av det ord som Gad hade talat i HERRENS namn .
då Ornan nu vände sig om , fick han se ängeln ; och hans fyra söner som voro med honom , gömde sig . men Ornan höll på att tröska vete .
och David kom till Ornan ; när då Ornan såg upp och fick se David , gick han fram ifrån tröskplatsen och föll ned till jorden på sitt ansikte för David .
och David sade till Ornan : &quot; Giv mig den plats där du tröskar din säd , så att jag där kan bygga ett altare åt HERREN ; giv mig den för full betalning ; och må så hemsökelsen upphöra bland folket &quot; .
då sade Ornan till David : &quot; tag den , och må sedan min herre konungen göra vad honom täckes . se , här giver jag dig fäkreaturen till brännoffer och tröskvagnarna till ved och vetet till spisoffer ; alltsammans giver jag &quot; .
men konung David svarade Ornan : &quot; Nej , jag vill köpa det för full betalning ; ty jag vill icke taga åt HERREN det som är ditt , och offra brännoffer som jag har fått för intet &quot; .
och David gav åt Ornan för platsen sex hundra siklar guld , i full vikt .
och David byggde där ett altare åt HERREN och offrade brännoffer och tackoffer . han ropade till HERREN , och han svarade honom med eld från himmelen på brännoffersaltaret .
och på HERRENS befallning stack ängeln sitt svärd tillbaka i skidan .
då , när David förnam att HERREN hade bönhört honom på jebuséen Ornans tröskplats , offrade han där .
men HERRENS tabernakel , som Mose hade låtit göra i öknen , stod jämte brännoffersaltaret , vid den tiden på offerhöjden i Gibeon .
dock vågade David icke komma inför Guds ansikte för att söka honom ; så förskräckt var han för HERRENS ängels svärd .
och David sade : &quot; här skall HERREN Guds hus stå , och här altaret för Israels brännoffer &quot; .
och David befallde att man skulle samla tillhopa de främlingar som funnos i Israels land ; och han anställde hantverkare , som skulle hugga ut stenar för att därmed bygga Guds hus .
och David anskaffade järn i myckenhet till spikar på dörrarna i portarna och till krampor , så ock koppar i sådan myckenhet att den icke kunde vägas ,
och cederbjälkar i otalig mängd ; ty sidonierna och tyrierna förde cederträ i myckenhet till David .
David tänkte nämligen : &quot; min son Salomo är ung och späd , men huset som skall byggas åt HERREN måste göras övermåttan stort , så att det bliver namnkunnigt och prisat i alla länder ; jag vill därför skaffa förråd åt honom &quot; . så skaffade David förråd i myckenhet före sin död .
och han kallade till sig sin son Salomo och bjöd honom att bygga ett hus åt HERREN , Israels Gud .
och David sade till sin son Salomo : &quot; jag hade själv i sinnet att bygga ett hus åt HERRENS , min Guds , namn .
men HERRENS ord kom till mig ; han sade : du har utgjutit blod i myckenhet och fört stora krig ; du skall icke bygga ett hus åt mitt namn , eftersom du har utgjutit så mycket blod på jorden , i min åsyn .
men se , åt dig skall födas en son ; han skall bliva en fridsäll man , och jag skall låta honom få fred med alla sina fiender runt omkring ; ty Salomo skall han heta , och frid och ro skall jag låta vila över Israel i hans dagar .
han skall bygga ett hus åt mitt namn ; han skall vara min son , och jag skall vara hans fader . och jag skall befästa hans konungatron över Israel för evig tid .
så vare nu HERREN med dig , min son ; må du bliva lyckosam och få bygga HERRENS , din Guds , hus , såsom han har lovat om dig .
må HERREN allenast giva dig klokhet och förstånd , när han sätter dig till härskare över Israel , och förhjälpa dig till att hålla HERRENS , din Guds , lag .
då skall du bliva lyckosam , om du håller och gör efter de stadgar och rätter som HERREN har bjudit Mose att ålägga Israel . var frimodig och oförfärad ; frukta icke och var icke försagd .
och se , trots mitt betryck har jag nu anskaffat till HERRENS hus ett hundra tusen talenter guld och tusen gånger tusen talenter silver , därtill av koppar och järn mer än som kan vägas , ty så mycket är det ; trävirke och sten har jag ock anskaffat , och mer må du själv anskaffa .
Arbetare har du ock i myckenhet hantverkare , stenhuggare och timmermän , och därtill allahanda folk som är kunnigt i allt slags annat arbete .
på guldet , silvret , kopparen och järnet kan ingen räkning hållas . upp då och gå till verket ; och vare HERREN med dig ! &quot;
därefter bjöd David alla Israels furstar att de skulle understödja hans son Salomo ; han sade :
&quot; HERREN , eder Gud , är ju med eder och har låtit eder få ro på alla sidor ; ty han har givit landets förra inbyggare i min hand , och landet har blivit HERREN och hans folk underdånigt .
så vänden nu edert hjärta och eder själ till att söka HERREN , eder Gud ; och stån upp och byggen HERREN Guds helgedom , så att man kan föra HERRENS förbundsark och vad annat som hör till Guds helgedom in i det hus som skall byggas åt HERRENS namn &quot; .
och när David blev gammal och levnadsmätt , gjorde han sin son Salomo till konung över Israel .
och han församlade alla Israels furstar , så ock prästerna och leviterna .
och leviterna blevo räknade , de nämligen som voro trettio år gamla eller därutöver ; och deras antal , antalet av alla personer av mankön , utgjorde trettioåtta tusen .
&quot; av dessa &quot; , sade han &quot; , skola tjugufyra tusen förestå sysslorna vid HERRENS hus , och sex tusen vara tillsyningsmän och domare ;
fyra tusen skola vara dörrvaktare och fyra tusen skola lovsjunga HERREN till de instrumenter som jag har låtit göra för lovsången &quot; .
och David delade dem i avdelningar efter Levis söner , Gerson Kehat och Merari .
till gersoniterna hörde Laedan och Simei .
Laedans söner voro Jehiel , huvudmannen , Setam och Joel , tillsammans tre .
Simeis söner voro Selomot , Hasiel och Haran , tillsammans tre . dessa voro huvudmän för Laedans familjer .
och Simeis söner voro Jahat , sina , Jeus och Beria . dessa voro Simeis söner , tillsammans fyra .
Jahat var huvudmannen , och Sisa var den andre . men Jeus och Beria hade icke många barn ; därför fingo de utgöra allenast en familj , en ordning .
Kehats söner voro Amram , Jishar , Hebron och Ussiel , tillsammans fyra .
Amrams söner voro Aron och Mose . och Aron blev jämte sina söner för evärdlig tid avskild till att helgas såsom höghelig , till att för evärdlig tid antända rökelse inför HERREN och göra tjänst inför honom och välsigna i hans namn .
men gudsmannen Moses söner räknades till Levi stam .
Moses söner voro Gersom och Elieser .
Gersoms söner voro Sebuel , huvudmannen .
och Eliesers söner voro Rehabja , huvudmannen . Elieser hade inga andra söner ; men Rehabjas söner voro övermåttan talrika .
Jishars söner voro Selomit , huvudmannen .
Hebrons söner voro Jeria , huvudmannen , Amarja , den andre , Jahasiel , den tredje , och Jekameam , den fjärde .
Ussiels söner voro Mika , huvudmannen , och Jissia , den andre .
