Men Aron och hans söner ombesörjde offren på brännoffersaltaret och på rökelsealtaret, och skulle utföra all förrättning i det allraheligaste och bringa försoning för Israel, alldeles såsom Mose, Guds tjänare, hade bjudit.
Och dessa voro Arons söner: hans son Eleasar, dennes son Pinehas, dennes son Abisua,
dennes son Bucki, dennes son Ussi, dennes son Seraja,
dennes son Merajot, dennes son Amarja, dennes son Ahitub,
dennes son Sadok, dennes son Ahimaas.
Och dessa voro deras boningsorter, efter deras tältläger inom deras område: Åt Arons söner av kehatiternas släkt -- ty dem träffade nu lotten --
åt dem gav man Hebron i Juda land med dess utmarker runt omkring.
Men åkerjorden och byarna som hörde till staden gav man åt Kaleb, Jefunnes son.
Åt Arons söner gav man alltså fristäderna Hebron och Libna med dess utmarker, vidare Jattir och Estemoa med dess utmarker.
Hilen med dess utmarker, Debir med dess utmarker,
Asan med dess utmarker och Bet-Semes med dess utmarker;
och ur Benjamins stam Geba med dess utmarker, Alemet med dess utmarker och Anatot med dess utmarker, så att deras städer tillsammans utgjorde tretton städer, efter deras släkter.
Och Kehats övriga barn fingo ur en stamsläkt, nämligen den stamhalva som utgjorde ena hälften av Manasse stam, genom lottkastning tio städer.
Gersoms barn åter fingo, efter sina släkter, ur Isaskars stam, ur Asers stam, ur Naftali stam och ur Manasse stam i Basan tretton städer.
Meraris barn fingo, efter sina släkter, ur Rubens stam, ur Gads stam och ur Sebulons stam genom lottkastning tolv städer.
Så gåvo Israels barn åt leviterna dessa städer med deras utmarker.
Genom lottkastning gåvo de åt dem ur Juda barns stam, ur Simeons barns stam och ur Benjamins barns stam dessa städer, som de namngåvo.
Och bland Kehats barns släkter fingo några följande städer ur Efraims stam såsom sitt område:
Man gav dem fristäderna Sikem med dess utmarker i Efraims bergsbygd, Geser med dess utmarker,
Jokmeam med dess utmarker, Bet-Horon med dess utmarker;
vidare Ajalon med dess utmarker och Gat-Rimmon med dess utmarker;
och ur ena hälften av Manasse stam Aner med dess utmarker och Bileam med dess utmarker. Detta tillföll Kehats övriga barns släkt.
Gersoms barn fingo ur den släkt som utgjorde ena hälften av Manasse stam Golan i Basan med dess utmarker och Astarot med dess utmarker;
och ur Isaskars stam Kedes med dess utmarker, Dobrat med dess utmarker,
Ramot med dess utmarker och Anem med dess utmarker;
och ur Asers stam Masal med dess utmarker, Abdon med dess utmarker,
Hukok med dess utmarker och Rehob med dess utmarker;
och ur Naftali stam Kedes i Galileen med dess utmarker, Hammon med dess utmarker och Kirjataim med dess utmarker.
Meraris övriga barn fingo ur Sebulons stam Rimmono med dess utmarker och Tabor med dess utmarker,
och på andra sidan Jordan mitt emot Jeriko, öster om Jordan, ur Rubens stam Beser i öknen med dess utmarker, Jahas med dess utmarker,
Kedemot med dess utmarker och Mefaat med dess utmarker;
och ur Gads stam Ramot i Gilead med dess utmarker, Mahanaim med dess utmarker,
Hesbon med dess utmarker och Jaeser med dess utmarker.
Och Isaskars söner voro Tola och Pua, Jasib och Simron, tillsammans fyra.
Tolas söner voro Ussi, Refaja, Jeriel, Jamai, Jibsam och Samuel, huvudmän för sina familjer, ättlingar av Tola, tappra stridsmän, upptecknade efter sin ättföljd. I Davids tid var deras antal tjugutvå tusen sex hundra.
Ussis söner voro Jisraja, och Jisrajas söner voro Mikael, Obadja och Joel samt Jissia, tillhopa fem, allasammans huvudmän.
Och med dem följde stridbara härskaror, trettiosex tusen man, efter sin ättföljd och sina familjer; ty de hade många hustrur och barn.
Och deras bröder i alla Isaskars släkter voro tappra stridsmän; åttiosju tusen utgjorde tillsammans de som voro upptecknade i deras släktregister.
Benjamins söner voro Bela, Beker och Jediael, tillsammans tre.
Belas söner voro Esbon, Ussi, Ussiel, Jerimot och Iri, tillsammans fem, huvudmän för sina familjer, tappra stridsmän; de som voro upptecknade i deras släktregister utgjorde tjugutvå tusen trettiofyra.
Bekers söner voro Semira, Joas, Elieser, Eljoenai, Omri, Jeremot, Abia, Anatot och Alemet. Alla dessa voro Bekers söner.
De som voro upptecknade i deras släktregister, efter sin ättföljd, efter huvudmannen för sina familjer, tappra stridsmän, utgjorde tjugu tusen två hundra.
Jediaels söner voro Bilhan; Bilhans söner voro Jeus, Benjamin, Ehud, Kenaana, Setan, Tarsis och Ahisahar.
Alla dessa voro Jediaels söner, upptecknade efter huvudmännen för sina familjer, tappra stridsmän, sjutton tusen två hundra stridbara krigsmän.
Och Suppim och Huppim voro Irs söner. -- Men Husim voro Ahers söner.
Naftalis söner voro Jahasiel, Guni, Jeser och Sallum, Bilhas söner.
Manasses söner voro Asriel, som kvinnan födde; hans arameiska bihustru födde Makir, Gileads fader.
Och Makir tog hustru åt Huppim och Suppim. Hans syster hette Maaka. Och den andre hette Selofhad. Och Selofhad hade döttrar.
Och Maaka, Makirs hustru, födde en son och gav honom namnet Peres, men hans broder hette Seres. Hans söner voro Ulam och Rekem.
Ulams söner voro Bedan. Dessa voro söner till Gilead, son till Makir, son till Manasse.
Och hans syster var Hammoleket; hon födde Is-Hod, Abieser och Mahela.
Och Semidas söner voro Ajan, Sekem, Likhi och Aniam.
Och Efraims söner voro Sutela, dennes son Bered, dennes son Tahat, dennes son Eleada, dennes son Tahat,
dennes son Sabad och dennes son Sutela, så ock Eser och Elead. Och män från Gat, som voro födda där i landet, dräpte dem, därför att de hade dragit ned för att taga deras boskapshjordar.
Då sörjde Efraim, deras fader, i lång tid, och hans bröder kommo för att trösta honom.
Och han gick in till sin hustru, och hon blev havande och födde en son; och han gav honom namnet Beria , därför att det hade skett under en olyckstid för hans hus.
Hans dotter var Seera; hon byggde Nedre och Övre Bet-Horon, så ock Ussen-Seera.
Och hans son var Refa; hans son var Resef, ävensom Tela; hans son var Tahan.
Hans son var Laedan; hans son var Ammihud; hans son var Elisama.
Hans son var Non; hans son var Josua.
Och deras besittning och deras boningsorter voro Betel med underlydande orter, österut Naaran och västerut Geser med underlydande orter, vidare Sikem med underlydande orter, ända till Aja med underlydande orter.
Men i Manasse barns ägo voro Bet-Sean med underlydande orter, Taanak med underlydande orter, Megiddo med underlydande orter, Dor med underlydande orter. Här bodde nu Josefs, Israels sons, barn.
Asers söner voro Jimna, Jisva, Jisvi och Beria; och deras syster var Sera.
Berias söner voro Heber och Malkiel; han var Birsaits fader.
Och Heber födde Jaflet, Somer och Hotam, så ock Sua, deras syster.
Och Jaflets söner voro Pasak, Bimhal och Asvat. Dessa voro Jaflets söner.
Semers söner voro Ahi och Rohaga, Jaba och Aram.
Hans broder Helems söner voro Sofa, Jimna, Seles och Amal.
Sofas söner voro Sua, Harnefer, Sual, Beri och Jimra,
Beser, Hod, Samma, Silsa, Jitran och Beera.
Jeters söner voro Jefunne, Pispa och Ara.
Och Ullas söner voro Ara, Hanniel och Risja.
Alla dessa voro Asers söner, huvudmän för sina familjer, utvalda tappra stridsmän, huvudmän bland hövdingarna; och de som voro upptecknade i deras släktregister såsom dugliga till krigstjänst utgjorde ett antal av tjugusex tusen man.
Och Benjamin födde Bela, sin förstfödde, Asbel, den andre, och Ahara, den tredje,
Noha, den fjärde, och Rafa, den femte.
Bela hade följande söner: Addar, Gera, Abihud,
Abisua, Naaman, Ahoa,
Gera, Sefufan och Huram.
Och dessa voro Ehuds söner, och de voro familjehuvudmän för dem som bodde i Geba, och som blevo bortförda till Manahat,
dit Gera jämte Naaman och Ahia förde bort dem: han födde Ussa och Ahihud.
Och Saharaim födde barn i Moabs land, sedan han hade skilt sig från sina hustrur, Husim och Baara;
med sin hustru Hodes födde han där Jobab, Sibja, Mesa, Malkam,
Jeus, Sakeja och Mirma. Dessa voro hans söner, huvudmän för familjer.
Med Husim hade han fött Abitub och Elpaal.
Och Elpaals söner voro Eber, Miseam och Semed. Han var den som byggde Ono och Lod med underlydande orter.
Beria och Sema -- vilka voro familjehuvudmän för Ajalons invånare och förjagade Gats invånare --
så ock Ajo, Sasak och Jeremot.
Och Sebadja, Arad, Eder,
Mikael, Jispa och Joha voro Berias söner.
Och Sebadja, Mesullam, Hiski, Heber,
Jismerai, Jislia och Jobab voro Elpaals söner.
Och Jakim, Sikri, Sabdi,
Elienai, Silletai, Eliel,
Adaja, Beraja och Simrat voro Simeis söner.
Och Jispan, Eber, Eliel,
Abdon, Sikri, Hanan,
Hananja, Elam, Antotja,
Jifdeja och Peniel voro Sasaks söner.
Och Samserai, Seharja, Atalja,
Jaaresja, Elia och Sikri voro Jerohams söner.
Dessa vore huvudman för familjer, huvudmän efter sin ättföljd; de bodde i Jerusalem.
I Gibeon bodde Gibeons fader, vilkens hustru hette Maaka.
Och hans förstfödde son var Abdon; vidare Sur, Kis, Baal, Nadab,
Gedor, Ajo och Seker.
Men Miklot födde Simea. Också dessa bodde jämte sina bröder i Jerusalem, gent emot sina bröder.
Och Ner födde Kis, Kis födde Saul, och Saul födde Jonatan, Malki-Sua, Abinadab och Esbaal.
Jonatans son var Merib-Baal, och Merib-Baal födde Mika.
Mikas söner voro Piton, Melek, Taarea och Ahas.
Ahas födde Joadda, Joadda födde Alemet, Asmavet och Simri, och Simri födde Mosa.
Mosa födde Binea. Hans son var Rafa; hans son var Eleasa; hans son var Asel.
Och Asel hade sex söner, och dessa hette Asrikam, Bokeru, Ismael, Searja, Obadja och Hanan. Alla dessa voro Asels söner.
Och hans broder Eseks söner voro Ulam, hans förstfödde, Jeus, den andre, och Elifelet, den tredje.
Och Ulams söner voro tappra stridsmän, som voro skickliga i att spänna båge; och de hade många söner och sonsöner: ett hundra femtio. Alla dessa voro av Benjamins barn
Och hela Israel blev upptecknat i släktregister, och de finnas uppskrivna i boken om Israels konungar. Och Juda fördes i fångenskap bort till Babel för sin otrohets skull.
Men de förra invånarna som bodde där de hade sin arvsbesittning, i sina städer, utgjordes av vanliga israeliter, präster, leviter och tempelträlar.
I Jerusalem bodde en del av Juda barn, av Benjamins barn och av Efraims och Manasse barn, nämligen:
Utai, son till Ammihud, son till Omri, son till Imri, son till Bani, av Peres', Judas sons, barn;
av siloniterna Asaja, den förstfödde, och hans söner;
av Seras barn Jeguel och deras broder, sex hundra nittio;
av Benjamins barn Sallu, son till Mesullam, son till Hodauja, son till Hassenua,
vidare Jibneja, Jerohams son, och Ela, son till Ussi, son till Mikri, och Mesullam, son till Sefatja, son till Reguel, son till Jibneja,
så ock deras bröder, efter deras ättföljd, nio hundra femtiosex. Alla dessa män voro huvudmän för familjer, var och en för sin familj.
Och av prästerna: Jedaja, Jojarib och Jakin,
vidare Asarja, son till Hilkia, son till Mesullam, son till Sadok, son till Merajot, son till Ahitub, fursten i Guds hus,
vidare Adaja, son till Jeroham, son till Pashur, son till Malkia, vidare Maasai, son till Adiel, son till Jasera, son till Mesullam, son till Mesillemit, son till Immer,
så ock deras bröder, huvudmän för sina familjer, ett tusen sju hundra sextio, dugande män i de sysslor som hörde till tjänstgöringen i Guds hus.
Och av leviterna: Semaja, som till Hassub, son till Asrikam, son till Hasabja, av Meraris barn,
vidare Bakbackar, Heres och Galal, så ock Mattanja, son till Mika, son till Sikri, son till Asaf,
vidare Obadja, son till Semaja, son till Galal, son till Jedutun, så ock Berekja, son till Asa, son till Elkana, som bodde i netofatiternas byar.
Och dörrvaktarna: Sallum, Ackub, Talmon och Ahiman med sina bröder; men Sallum var huvudmannen.
Och ända till nu göra de tjänst vid Konungsporten, på östra sidan. Dessa voro dörrvaktarna i Levi barns läger.
Men Sallum, son till Kore, son till Ebjasaf, son till Kora, hade jämte sina bröder, dem som voro av hans familj, koraiterna, till tjänstgöringssyssla att hålla vakt vid tältets trösklar; deras fäder hade nämligen i HERRENS läger hållit vakt vid ingången.
Och Pinehas, Eleasars son, hade förut varit furste över dem -- med honom vare HERREN!
Sakarja, Meselemjas son, var dörrvaktare vid ingången till uppenbarelsetältet.
Alla dessa voro utvalda till dörrvaktare vid trösklarna: två hundra tolv. De blevo i sina byar upptecknade i släktregistret. David och siaren Samuel hade tillsatt dem att tjäna på heder och tro.
De och deras söner stodo därför vid portarna till HERRENS hus, tälthuset, och höllo vakt.
Efter de fyra väderstrecken hade dörrvaktarna sina platser: i öster, väster, norr och söder.
Och deras bröder, de som fingo bo i sina byar, skulle var sjunde dag, alltid på samma timme, infinna sig hos dem.
Ty på heder och tro voro dessa fyra anställda såsom förmän för dörrvaktarna. Detta var nu leviterna. De hade ock uppsikten över kamrarna och förvaringsrummen i Guds hus.
Och de vistades om natten runt omkring Guds hus, ty dem ålåg att hålla vakt, och de skulle öppna dörrarna var morgon.
Somliga av dem hade uppsikten över de kärl som användes vid tjänstgöringen. De buro nämligen in dem, efter att hava räknat dem, och buro sedan ut dem, efter att åter hava räknat dem.
Och somliga av dem voro förordnade till att hava uppsikten över de andra kärlen, över alla andra helgedomens kärl, så ock över det fina mjölet och vinet och oljan och rökelsen och de välluktande kryddorna.
Men somliga av prästernas söner beredde salvan av de välluktande kryddorna.
Och Mattitja, en av leviterna, koraiten Sallums förstfödde, hade på heder och tro uppsikten över bakverket.
Och somliga av deras bröder, kehatiternas söner, hade uppsikten över skådebröden och skulle tillreda dem för var sabbat.
Men de andra, nämligen sångarna, huvudmän för levitiska familjer, vistades i kamrarna, fria ifrån annan tjänstgöring, ty dag och natt voro de upptagna av sina egna sysslor.
Dessa voro huvudmännen för de levitiska familjerna, huvudman efter sin ättföljd; de bodde i Jerusalem.
I Gibeon bodde Gibeons fader Jeguel, vilkens hustru hette Maaka.
Och hans förstfödde son var Abdon; vidare Sur, Kis, Baal, Ner, Nadab
Gedor, Ajo, Sakarja och Miklot.
Men Miklot födde Simeam. Också de bodde jämte sina bröder i Jerusalem, gent emot sina bröder.
Och Ner födde Kis, Kis födde Saul, och Saul födde Jonatan, Malki-Sua, Abinadab och Esbaal.
Jonatans son var Merib-Baal, och Merib-Baal födde Mika.
Mikas söner voro Piton, Melek och Taharea.
Ahas födde Jaera, Jaera födde Alemet, Asmavet och Simri, och Simri födde Mosa.
Mosa födde Binea. Hans son var Refaja; hans son var Eleasa; hans son var Asel.
Och Asel hade sex söner, och dessa hette Asrikam, Bokeru, Ismael, Searja, Obadja och Hanan. Dessa voro Asels söner
Och filistéerna stridde mot Israel; och Israels män flydde för filistéerna och föllo slagna på berget Gilboa.
Och filistéerna ansatte ivrigt Saul och hans söner. Och filistéerna dödade Jonatan, Abinadab och Malki-Sua, Sauls söner.
När då Saul själv blev häftigt anfallen och bågskyttarna kommo över honom, greps han av förskräckelse för skyttarna.
Och Saul sade till sin vapendragare: »Drag ut ditt svärd och genomborra mig därmed, så att icke dessa oomskurna komma och hantera mig skändligt.» Men hans vapendragare ville det icke, ty han fruktade storligen. Då tog Saul själv svärdet och störtade sig därpå.
Men när vapendragaren såg att Saul var död, störtade han sig ock på sitt svärd och dog.
Så dogo då Saul och hans tre söner; och alla som hörde till hans hus dogo på samma gång.
Och när alla israeliterna i dalen förnummo att deras här hade flytt, och att Saul och hans söner voro döda, övergåvo de sina städer och flydde; sedan kommo filistéerna och bosatte sig i dem.
Dagen därefter kommo filistéerna för att plundra de slagna och funno då Saul och hans söner, där de lågo fallna på berget Gilboa.
Och de plundrade honom och togo med sig hans huvud och hans vapen och sände dem omkring i filistéernas land och läto förkunna det glada budskapet för sina avgudar och för folket.
Och de lade hans vapen i sitt gudahus, men hans huvudskål hängde de upp i Dagons tempel.
Men när allt folket i Jabes i Gilead hörde allt vad filistéerna hade gjort med Saul,
stodo de upp, alla stridbara män, och togo Sauls och hans söners lik och förde dem till Jabes; och de begrovo deras ben under terebinten i Jabes och fastade så i sju dagar.
Detta blev Sauls död, därför att han hade begått otrohet mot HERREN, i det att han icke hade hållit HERRENS ord, så ock därför att han hade frågat en ande och sökt svar hos en sådan.
Han hade icke sökt svar hos HERREN; därför dödade HERREN honom. Och sedan överflyttade han konungadömet på David, Isais son.
Då församlade sig hela Israel till David i Hebron och sade: »Vi äro ju ditt kött och ben.
Redan för länge sedan, redan då Saul ännu var konung, var det du som var ledare och anförare för Israel. Och till dig har HERREN, din Gud, sagt: Du skall vara en herde för mitt folk Israel, ja, du skall vara en furste över mitt folk Israel.»
När så alla de äldste i Israel kommo till konungen i Hebron, slöt David ett förbund med dem där i Hebron, inför HERREN; och sedan smorde de David till konung över Israel, i enlighet med HERRENS ord genom Samuel.
Och David drog med hela Israel till Jerusalem, det är Jebus; där befunno sig jebuséerna, som ännu bodde kvar i landet.
Och invånarna i Jebus sade till David: »Hitin kommer du icke.» Men David intog likväl Sions borg, det är Davids stad
Och David sade: »Vemhelst som först slår ihjäl en jebusé, han skall bliva hövding och anförare.» Och Joab, Serujas son, kom först ditupp och blev så hövding.
Sedan tog David sin boning i bergfästet; därför kallade man det Davids stad.
Och han uppförde befästningsverk runt omkring staden, från Millo och allt omkring; och Joab återställde det övriga av staden.
Och David blev allt mäktigare och mäktigare, och HERREN Sebaot var med honom
Och dessa äro de förnämsta bland Davids hjältar, vilka gåvo honom kraftig hjälp att bliva konung, de jämte hela Israel, och så skaffade honom konungaväldet, enligt HERRENS ord angående Israel.
Detta är förteckningen på Davids hjältar: Jasobeam, son till en hakmonit, den förnämste bland kämparna, han som svängde sitt spjut över tre hundra som hade blivit slagna på en gång.
Och efter honom kom ahoaiten Eleasar, son till Dodo; han var en av de tre hjältarna.
Han var med David vid Pas-Dammim, när filistéerna där hade församlat sig till strid. Och där var ett åkerstycke, fullt med korn. Och folket flydde för filistéerna.
Då ställde de sig mitt på åkerstycket och försvarade det och slogo filistéerna; och HERREN lät dem så vinna en stor seger.
En gång drogo tre av de trettio förnämsta männen ned över klippan till David vid Adullams grotta, medan en avdelning filistéer var lägrad i Refaimsdalen.
Men David var då på borgen, under det att en filisteisk utpost fanns i Bet-Lehem.
Och David greps av lystnad och sade: »Ack att någon ville giva mig vatten att dricka från brunnen vid Bet-Lehems stadsport!»
Då bröto de tre sig igenom filistéernas läger och hämtade vatten ur brunnen vid Bet-Lehems stadsport och togo det och buro det till David. Men David ville icke dricka det, utan göt ut det såsom ett drickoffer åt HERREN.
Han sade nämligen: »Gud låte det vara fjärran ifrån mig att jag skulle göra detta! Skulle jag dricka dessa mäns blod, som hava vågat sina liv? Ty med fara för sina liv hava de burit det hit.» Och han ville icke dricka det. Sådana ting hade de tre hjältarna gjort.
Absai, Joabs broder, var den förnämste av tre andra; han svängde en gång sitt spjut över tre hundra som hade blivit slagna. Och han hade ett stort namn bland de tre.
Han var dubbelt mer ansedd än någon annan i detta tretal, och han var deras hövitsman, men upp till de tre första kom han dock icke.
Vidare Benaja, son till Jojada, som var son till en tapper, segerrik man från Kabseel; han slog ned de två Arielerna i Moab, och det var han som en snövädersdag steg ned och slog ihjäl lejonet i brunnen.
Han slog ock ned den egyptiske mannen som var så reslig: fem alnar lång. Fastän egyptiern i handen hade ett spjut som liknade en vävbom, gick han ned mot honom, väpnad allenast med sin stav. Och han ryckte spjutet ur egyptiern hand och dräpte honom med hans eget spjut.
Sådana ting hade Benaja, Jojadas son, gjort. Och han hade ett stort namn bland de tre hjältarna.
Ja, han var mer ansedd än någon av de trettio, men upp till de tre första kom han icke. Och David satte honom till anförare för sin livvakt.
De tappra hjältarna voro: Asael, Joabs broder, Elhanan, Dodos son, från Bet-Lehem;
haroriten Sammot; peloniten Heles;
tekoaiten Ira, Ickes' son; anatotiten Abieser;
husatiten Sibbekai; ahoaiten Ilai;
netofatiten Maherai; netofatiten Heled, Baanas son;
Itai, Ribais son, från Gibea i Benjamins barns stam; pirgatoniten Benaja;
Hurai från Gaas' dalar; arabatiten Abiel;
baharumiten Asmavet; saalboniten Eljaba;
gisoniten Bene-Hasem; harariten Jonatan, Sages son;
harariten Ahiam, Sakars son; Elifal, Urs son;
mekeratiten Hefer; peloniten Ahia;
Hesro från Karmel; Naarai, Esbais son;
Joel, broder till Natan; Mibhar, Hagris son;
ammoniten Selek; berotiten Naherai, vapendragare åt Joab, Serujas son;
jeteriten Ira; jeteriten Gareb;
hetiten Uria; Sabad, Alais son;
rubeniten Adina, Sisas son, en huvudman bland rubeniterna, och jämte honom trettio andra;
Hanan, Maakas son, och mitniten Josafat;
astarotiten Ussia; Sama och Jeguel, aroeriten Hotams söner;
Jediael, Simris son, och hans broder Joha, tisiten;
Eliel-Hammahavim samt Jeribai och Josauja, Elnaams söner, och moabiten Jitma;
slutligen Eliel, Obed och Jaasiel-Hammesobaja.
Och dessa voro de som kommo till David i Siklag, medan han ännu höll sig undan för Saul, Kis' son; de hörde till de hjältar som bistodo honom under kriget.
De voro väpnade med båge och skickliga i att, både med höger och med vänster hand, slunga stenar och avskjuta pilar från bågen. Av Sauls stamfränder, benjaminiterna, kommo:
Ahieser, den förnämste, och Joas, gibeatiten Hassemaas söner; Jesuel och Pelet, Asmavets söner; Beraka; anatotiten Jehu;
gibeoniten Jismaja, en av de trettio hjältarna, anförare för de trettio; Jeremia; Jahasiel; Johanan; gederatiten Josabad;
Eleusai; Jerimot; Bealja; Semarja; harufiten Sefatja;
koraiterna Elkana, Jissia, Asarel, Joeser och Jasobeam;
Joela och Sebadja, söner till Jeroham, av strövskaran.
Och av gaditerna avföllo några och gingo till David i bergfästet i öknen, tappra män, krigsmän skickliga att strida, rustade med sköld och spjut; de hade en uppsyn såsom lejon och voro snabba såsom gaseller på bergen:
Eser, den förnämste, Obadja, den andre, Eliab, den tredje,
Masmanna, den fjärde, Jeremia, den femte,
Attai, den sjätte, Eliel, den sjunde,
Johanan, den åttonde, Elsabad, den nionde,
Jeremia, den tionde, Makbannai, den elfte.
Dessa hörde till Gads barn och till de förnämsta i hären; den ringaste av dem var ensam så god som hundra, men den ypperste så god som tusen.
Dessa voro de som i första månaden gingo över Jordan, när den var full över alla sina bräddar, och som förjagade alla dem som bodde i dalarna, åt öster och åt väster.
Av Benjamins och Juda barn kommo några män till David ända till bergfästet.
Då gick David ut emot dem och tog till orda och sade till dem: »Om I kommen till mig i fredlig avsikt och viljen bistå mig, så är mitt hjärta redo till förening med eder; men om I kommen för att förråda mig åt mina ovänner, fastän ingen orätt är i mina händer, då må våra fäders Gud se därtill och straffa det.»
Men Amasai, den förnämste bland de trettio, hade blivit beklädd med andekraft, och han sade: »Dina äro vi, David, och med dig stå vi, du Isais son. Frid vare med dig, frid, och frid vare med dem som bistå dig ty din Gud har bistått dig!» Och David tog emot dem och gav dem plats bland de förnämsta i sin skara.
Från Manasse gingo några över till David, när han med filistéerna drog ut i strid mot Saul, dock fingo de icke bistå dessa; ty när filistéernas hövdingar hade rådplägat, skickade de bort honom, i det de sade: »Det gäller huvudet för oss, om han går över till sin herre Saul.
När han då drog till Siklag, gingo dessa från Manasse över till honom: Adna, Josabad, Jediael, Mikael, Josabad, Elihu och Silletai, huvudmän för de ätter som tillhörde Manasse.
Dessa bistodo David mot strövskaran, ty de voro allasammans tappra stridsmän och blevo hövitsmän i hären.
Dag efter dag kommo nämligen allt flera till David för att bistå honom, så att hans läger blev övermåttan stort.
Detta är de tal som angiva summorna av det väpnade krigsfolk som kom till David i Hebron, för att efter HERRENS befallning flytta Sauls konungamakt över på honom:
Juda barn, som buro sköld och spjut, sex tusen åtta hundra, väpnade till strid;
av Simeons barn tappra krigsmän, sju tusen ett hundra;
av Levi barn fyra tusen sex hundra;
därtill Jojada, fursten inom Arons släkt, och med honom tre tusen sju hundra;
så ock Sadok, en tapper yngling, med sin familj, tjugutvå hövitsmän;
av Benjamins barn, Sauls stamfränder, tre tusen (ty ännu vid den tiden höllo de flesta av dem troget med Sauls hus);
av Efraims barn tjugu tusen åtta hundra, tappra stridsmän, namnkunniga män i sina familjer;
av ena hälften av Manasse stam aderton tusen namngivna män, som kommo för att göra David till konung;
av Isaskars barn kommo män som väl förstodo tidstecknen och insågo vad Israel borde göra, två hundra huvudmän, därtill alla deras stamfränder under deras befäl;
av Sebulon stridbara män, rustade till krig med alla slags vapen, femtio tusen, som samlades endräktigt;
av Naftali ett tusen hövitsmän, och med dem trettiosju tusen, väpnade med sköld och spjut;
av daniterna krigsrustade män, tjuguåtta tusen sex hundra;
av Aser stridbara män, rustade till krig, fyrtio tusen;
och från andra sidan Jordan, av rubeniterna, gaditerna och andra hälften av Manasse stam, ett hundra tjugu tusen, väpnade med alla slags vapen som brukas vid krigföring.
Alla dessa krigsmän, ordnade till strid, kommo i sina hjärtans hängivenhet till Hebron för att göra David till konung över hela Israel. Också hela det övriga Israel var enigt i att göra David till konung.
Och de voro där hos David i tre dagar och åto och drucko, ty deras bröder hade försett dem med livsmedel.
De som bodde närmast dem, ända upp till Isaskar, Sebulon och Naftali, tillförde dem ock på åsnor, kameler, mulåsnor och oxar livsmedel i myckenhet till föda: mjöl, fikonkakor och russinkakor, vin och olja, fäkreatur och småboskap; ty glädje rådde i Israel.
Och David rådförde sig med över- och underhövitsmännen, med alla furstarna.
Sedan sade David till Israels hela församling: »Om I så finnen för gott, och om detta är från HERREN, vår Gud, så låt oss sända bud åt alla håll till våra övriga bröder i alla Israels landsändar, och därjämte till prästerna och leviterna i de städer kring vilka de hava sina utmarker, att de må församla sig till oss;
och låt oss flytta vår Guds ark till oss, ty i Sauls tid frågade vi icke efter den.»
Och hela församlingen svarade att man skulle göra så, ty förslaget behagade hela folket.
Så församlade då David hela Israel, från Sihor i Egypten ända dit där vägen går till Hamat, för att hämta Guds ark från Kirjat-Jearim.
Och David drog med hela Israel upp till Baala, det är Kirjat-Jearim, som hör till Juda, för att därifrån föra upp Guds, HERRENS, ark, hans som tronar på keruberna, och efter vilken den hade fått sitt namn.
Och de satte Guds ark på en ny vagn och förde den bort ifrån Abinadabs hus; och Ussa och Ajo körde vagnen.
Och David och hela Israel fröjdade sig inför Gud av all makt, med sånger och med harpor, psaltare, pukor, cymbaler och trumpeter.
Men när de kommo till Kidonslogen, räckte Ussa ut sin hand för att fatta I arken, ty oxarna snavade.
Då upptändes HERRENS vrede mot Ussa, och därför att han hade räckt ut sin hand mot arken, slog han honom, så att han föll ned död där inför Gud.
Men det gick David hårt till sinnes att HERREN så hade brutit ned Ussa ; och han kallade det stället Peres-Ussa , såsom det heter ännu i dag.
Och David betogs av sådan fruktan för Gud på den dagen, att han sade: »Huru skulle jag töras låta föra Guds ark till mig?»
Därför lät David icke flytta in arken till sig i Davids stad, utan lät sätta in den i gatiten Obed-Edoms hus.
Sedan blev Guds ark kvar vid Obed-Edoms hus, där den stod i sitt eget hus, i tre månader; men HERREN välsignade Obed-Edoms hus och allt vad som hörde honom till.
Och Hiram, konungen i Tyrus, skickade sändebud till David med cederträ, därjämte ock murare och timmermän, för att de skulle bygga honom ett hus.
Och David märkte att HERREN hade befäst honom såsom konung över Israel; ty han hade låtit hans rike bliva övermåttan upphöjt, för sitt folk Israels skull.
Och David tog sig ännu flera hustrur i Jerusalem, och David födde ännu flera söner och döttrar.
Dessa äro namnen på de söner som han fick i Jerusalem: Sammua, Sobab, Natan, Salomo,
Jibhar, Elisua, Elpelet,
Noga, Nefeg, Jafia,
Elisama, Beeljada och Elifelet.
Men när filistéerna hörde att David hade blivit smord till konung över hela Israel, drogo de allasammans upp för att fånga David. När David hörde detta, drog han ut mot dem.
Då nu filistéerna hade fallit in i Refaimsdalen och där företogo plundringståg,
frågade David Gud: »Skall jag draga upp mot filistéerna? Vill du då giva dem i min hand?» HERREN svarade honom: »Drag upp; jag vill giva dem i din hand.»
Och de drogo upp till Baal-Perasim, och där slog David dem. Då sade David: »Gud har brutit ned mina fiender genom min hand, likasom en vattenflod bryter ned.» Därav fick det stället namnet Baal-Perasim .
De lämnade där efter sig sina gudar; och David befallde att dessa skulle brännas upp i eld.
Men filistéerna företogo ännu en gång plundringståg i dalen.
När David då åter frågade Gud, svarade Gud honom: »Du skall icke draga upp efter dem; du må kringgå dem på en omväg, så att du kommer över dem från det håll där bakaträden stå.
Så snart du sedan hör ljudet av steg i bakaträdens toppar, drag då ut till strid, ty då har Gud dragit ut framför dig till att slå filistéernas här.»
David gjorde såsom Gud hade bjudit honom; och de slogo filistéernas här och förföljde dem från Gibeon ända till Geser.
Och ryktet om David gick ut i alla länder, och HERREN lät fruktan för honom komma över alla folk.
Och han uppförde åt sig hus i Davids stad; sedan beredde han en plats åt Guds ark och slog upp ett tält åt den.
Därvid befallde David: »Inga andra än leviterna må bära Guds ark; ty dem har HERREN utvalt till att bära Guds ark och till att göra tjänst inför honom för evärdlig tid.»
Och David församlade hela Israel till Jerusalem för att hämta HERRENS ark upp till den plats som han hade berett åt den.
Och David samlade tillhopa Arons barn och leviterna;
av Kehats barn: Uriel, deras överste, och hans bröder, ett hundra tjugu;
av Meraris barn: Asaja, deras överste, och hans bröder, två hundra tjugu;
av Gersoms barn: Joel, deras överste, och hans bröder, ett hundra trettio;
av Elisafans barn: Semaja, deras överste, och hans bröder, två hundra;
av Hebrons barn: Eliel, deras överste, och hans bröder, åttio;
av Ussiels barn: Amminadab, deras överste, och hans bröder, ett hundra tolv.
Och David kallade till sig prästerna Sadok och Ebjatar jämte leviterna Uriel, Asaja, Joel, Semaja, Eliel och Amminadab.
Och han sade till dem: »I ären huvudmän för leviternas familjer. Helgen eder tillika med edra bröder, och hämten så HERRENS, Israels Guds, ark upp till den plats som jag har berett åt den.
Ty därför att I förra gången icke voren tillstädes var det som HERREN, vår Gud, bröt ned en av oss, till straff för att vi icke sökte honom så, som tillbörligt var.»
Då helgade prästerna och leviterna sig till att hämta upp HERRENS, Israels Guds, ark.
Och såsom Mose hade bjudit i enlighet med HERRENS ord, buro nu Levi barn Guds ark med stänger, som vilade på deras axlar.
Och David sade till de översta bland leviterna att de skulle förordna sina bröder sångarna till tjänstgöring med musikinstrumenter, psaltare, harpor och cymbaler, som de skulle låta ljuda, under det att de höjde glädjesången.
Leviterna förordnade då Heman, Joels son, och av hans bröder Asaf, Berekjas son, och av dessas bröder, Meraris barn, Etan, Kusajas son,
och jämte dem deras bröder av andra ordningen Sakarja, Ben, Jaasiel, Semiramot, Jehiel, Unni, Eliab, Benaja, Maaseja, Mattitja, Elifalehu, Mikneja, Obed-Edom och Jegiel, dörrvaktarna.
Och sångarna, Heman, Asaf och Etan, skulle slå kopparcymbaler.
Sakarja, Asiel, Semiramot, Jehiel, Unni, Eliab, Maaseja och Benaja skulle spela på psaltare, till Alamót.
Mattitja, Elifalehu, Mikneja, Obed-Edom, Jegiel och Asasja skulle leda sången med harpor, till Seminit.
Kenanja, leviternas anförare, när de buro, skulle undervisa i att bära, ty han var kunnig i sådant.
Berekja och Elkana skulle vara dörrvaktare vid arken.
Sebanja, Josafat, Netanel, Amasai, Sakarja, Benaja och Elieser, prästerna, skulle blåsa i trumpeter framför Guds ark. Slutligen skulle Obed-Edom och Jehia vara dörrvaktare vid arken.
Så gingo då David och de äldste i Israel och överhövitsmännen åstad för att hämta HERRENS förbundsark upp ur Obed-Edoms hus, under jubel.
Och då Gud skyddade leviterna som buro HERRENS förbundsark, offrade man sju tjurar och sju vädurar.
Därvid var David klädd i en kåpa av fint linne; så voro ock alla leviterna som buro arken, så ock sångarna och Kenanja, som anförde sångarna, när de buro. Och därjämte bar David en linne-efod.
Och hela Israel hämtade upp HERRENS förbundsark under jubel och basuners ljud; och man blåste i trumpeter och slog cymbaler och lät psaltare och harpor ljuda.
När då HERRENS förbundsark kom till Davids stad, blickade Mikal, Sauls dotter, ut genom fönstret, och då hon såg konung David dansa och göra sig glad, fick hon förakt för honom i sitt hjärta.
Sedan de hade fört Guds ark ditin, ställde de den i tältet som David hade slagit upp åt den, och framburo därefter brännoffer och tackoffer inför Guds ansikte.
När David hade offrat brännoffret och tackoffret, välsignade han folket i HERRENS namn.
Och åt var och en av alla israeliterna, både man och kvinna, gav han en kaka bröd, ett stycke kött och en druvkaka.
Och han förordnade vissa leviter till att göra tjänst inför HERRENS ark, för att de skulle prisa, tacka och lova HERREN, Israels Gud:
Asaf såsom anförare, näst efter honom Sakarja, och vidare Jegiel, Semiramot, Jehiel, Mattitja, Eliab, Benaja, Obed-Edom och Jegiel med psaltare och harpor; och Asaf skulle slå cymbaler.
Men prästerna Benaja och Jahasiel skulle beständigt stå med sina trumpeter framför Guds förbundsark.
På den dagen var det som David först fastställde den ordningen att man genom Asaf och hans bröder skulle tacka HERREN på detta sätt:
»Tacken HERREN, åkallen hans namn, gören hans gärningar kunniga bland folken.
Sjungen till hans ära, lovsägen honom, talen om alla hans under.
Berömmen eder av hans heliga namn; glädje sig av hjärtat de som söka HERREN.
Frågen efter HERREN och hans makt, söken hans ansikte beständigt.
Tänken på de underbara verk som han har gjort, på hans under och hans muns domar,
I Israels, hans tjänares, säd, I Jakobs barn, hans utvalda.
Han är HERREN, vår Gud; över hela jorden gå hans domar.
Tänken evinnerligen på hans förbund, intill tusen släkten på vad han har stadgat,
på det förbund han slöt med Abraham och på hans ed till Isak.
Han fastställde det för Jakob till en stadga, för Israel till ett evigt förbund;
han sade: 'Åt dig vill jag giva Kanaans land, det skall bliva eder arvedels lott.'
Då voren I ännu en liten hop, I voren ringa och främlingar därinne.
Och de vandrade åstad ifrån folk till folk ifrån ett rike bort till ett annat.
Han tillstadde ingen att göra dem skada, han straffade konungar för deras skull:
'Kommen icke vid mina smorda, och gören ej mina profeter något ont.'
Sjungen till HERRENS ära, alla länder, båden glädje var dag, förkunnen hans frälsning.
Förtäljen bland hedningarna hans ära, bland alla folk hans under.
Ty stor är HERREN och högt lovad, och fruktansvärd är han mer än alla gudar.
Ty folkens alla gudar äro avgudar, men HERREN är den som har gjort himmelen.
Majestät och härlighet äro inför hans ansikte, makt och fröjd i hans boning.
Given åt HERREN, I folkens släkter, given åt HERREN ära och makt;
given åt HERREN hans namns ära, bären fram skänker och kommen inför hans ansikte, tillbedjen HERREN i helig skrud.
Bäven för hans ansikte, alla länder; se, jordkretsen står fast och vacklar icke.
Himmelen vare glad, och jorden fröjde sig, och bland hedningarna säge man: 'HERREN är nu konung!'
Havet bruse och allt vad däri är, marken glädje sig och allt som är därpå;
ja, då juble skogens träd inför HERREN, ty han kommer för att döma jorden.
Tacken HERREN, ty han är god, ty hans nåd varar evinnerligen,
och sägen: 'Fräls oss, du vår frälsnings Gud, församla oss och rädda oss från hedningarna, så att vi få prisa ditt heliga namn och berömma oss av ditt lov.'
Lovad vare HERREN, Israels Gud, från evighet till evighet!» Och allt folket sade: »Amen», och lovade HERREN.
Och han gav där, inför HERRENS förbundsark, åt Asaf och hans bröder uppdraget att beständigt göra tjänst inför arken, var dag med de för den dagen bestämda sysslorna.
Men Obed-Edom och deras bröder voro sextioåtta; och Obed-Edom, Jedituns son, och Hosa gjorde han till dörrvaktare.
Och prästen Sadok och hans bröder, prästerna, anställde han inför HERRENS tabernakel, på offerhöjden i Gibeon,
för att de beständigt skulle offra åt HERREN brännoffer på brännoffersaltaret, morgon och afton, och göra allt vad som var föreskrivet i HERRENS lag, den som han hade givit åt Israel;
och jämte dem Heman och Jedutun och de övriga namngivna utvalda, på det att de skulle tacka HERREN, därför att hans nåd varar evinnerligen.
Och hos dessa, nämligen Heman och Jedutun, förvarades trumpeter och cymbaler åt dem som skulle spela, så ock andra instrumenter som hörde till gudstjänsten. Och Jedutuns söner gjorde han till dörrvaktare.
Sedan gick allt folket hem, var och en till sitt; men David vände om för att hälsa sitt husfolk.
Då nu David satt i sitt hus, sade han till profeten Natan: »Se, jag bor i ett hus av cederträ, under det att HERRENS förbundsark står under ett tält.»
Natan sade till David: »Gör allt vad du har i sinnet; ty Gud är med dig.»
Men om natten kom Guds ord till Natan; han sade:
»Gå och säg till min tjänare David: Så säger HERREN: Icke du skall bygga mig det hus som jag skall bo i.
Jag har ju icke bott i något hus, från den dag då jag förde Israel hitupp ända till denna dag, utan jag har flyttat ifrån tält till tält, ifrån tabernakel till tabernakel.
Har jag då någonsin, varhelst jag flyttade omkring med hela Israel, talat och sagt så till någon enda av Israels domare, som jag har förordnat till herde för mitt folk: 'Varför haven I icke byggt mig ett hus av cederträ?'
Och nu skall du säga så till min tjänare David: Så säger HERREN Sebaot: Från betesmarken, där du följde fåren, har jag hämtat dig, för att du skulle bliva en furste över mitt folk Israel.
Och jag har varit med dig på alla dina vägar och utrotat alla dina fiender för dig. Och jag vill göra dig ett namn, sådant som de störstes namn på jorden.
Jag skall bereda en plats åt mitt folk Israel och plantera det, så att det får bo kvar där, utan att vidare bliva oroat. Orättfärdiga människor skola icke mer föröda det, såsom fordom skedde,
och såsom det har varit allt ifrån den tid då jag förordnade domare över mitt folk Israel; och jag skall kuva alla dina fiender. Så förkunnar jag nu för dig att HERREN skall bygga ett hus åt dig.
Ty det skall ske, att när din tid är ute och du går till dina fäder skall jag efter dig upphöja din son, en av dina avkomlingar; och jag skall befästa hans konungamakt.
Han skall bygga ett hus åt mig, och jag skall befästa hans tron för evig tid.
Jag skall vara hans fader, och han skall vara min son; och min nåd skall jag icke låta vika ifrån honom, såsom jag lät den vika ifrån din företrädare.
Jag skall hålla honom vid makt i mitt hus och i mitt rike för evig tid, och hans tron skall vara befäst för evig tid.»
Alldeles i överensstämmelse med dessa ord och med denna syn talade nu Natan till David.
Då gick konung David in och satte sig ned inför HERRENS ansikte och sade: »Vem är jag, HERRE Gud, och vad är mitt hus, eftersom du har låtit mig komma härtill?
Och detta har likväl synts dig vara för litet, o Gud; du har talat angående din tjänares hus om det som ligger långt fram i tiden. Ja, du har sett till mig på människosätt, for att upphöja mig, HERRE Gud.
Vad skall nu David vidare säga till dig om den ära du har bevisat din tjänare? Du känner ju din tjänare.
HERRE, för din tjänares skull och efter ditt hjärta har du gjort allt detta stora och förkunnat alla dessa stora ting.
HERRE, ingen är dig lik, och ingen Gud finnes utom dig, efter allt vad vi hava hört med våra öron.
Och var finnes på jorden något enda folk som är likt ditt folk Israel, vilket Gud själv har gått åstad att förlossa åt sig till ett folk -- för att så göra dig ett stort och fruktansvärt namn, i det att du förjagade hedningarna för ditt folk, det som du hade förlossat ifrån Egypten?
Och du har gjort ditt folk Israel till ett folk åt dig för evig tid, och du, HERRE, har blivit deras Gud
Så må nu, HERRE, vad du har talat om din tjänare och om hans hus bliva fast för evig tid; gör såsom du har talat.
Då skall ditt namn anses fast och bliva stort till evig tid, så att man skall säga: 'HERREN Sebaot, Israels Gud, är Gud över Israel.' Och så skall din tjänare Davids hus bestå inför dig.
Ty du, min Gud, har uppenbarat för din tjänare att du skall bygga honom ett hus; därför har din tjänare dristat att bedja inför dig.
Och nu, HERRE, du är Gud; och då du har lovat din tjänare detta goda,
så må du nu ock värdigas välsigna din tjänares hus, så att det förbliver evinnerligen inför dig. Ty vad du, HERRE, välsignar, det är välsignat evinnerligen.»
En tid härefter slog David filistéerna och kuvade dem. Därvid tog han Gat med underlydande orter ur filistéernas hand.
Han slog ock moabiterna; så blevo moabiterna David underdåniga och förde till honom skänker.
Likaledes slog David Hadareser, konungen i Soba, vid Hamat, när denne hade dragit åstad för att befästa sitt välde vid floden Frat.
Och David tog ifrån honom ett tusen vagnar och tog till fånga sju tusen ryttare och tjugu tusen man fotfolk; och David lät avskära fotsenorna på alla vagnshästarna, utom på ett hundra hästar, som han skonade.
När sedan araméerna från Damaskus kommo för att hjälpa Hadareser, konungen i Soba, nedgjorde David tjugutvå tusen man av dem.
Och David insatte fogdar bland araméerna i Damaskus; och araméerna blevo David underdåniga och förde till honom skänker. Så gav HERREN seger åt David, varhelst han drog fram.
Och David tog de gyllene sköldar som Hadaresers tjänare hade burit och förde dem till Jerusalem.
Och från Hadaresers städer Tibhat och Kun tog David koppar i stor myckenhet; därav gjorde sedan Salomo kopparhavet, pelarna och kopparkärlen.
Då nu Tou, konungen i Hamat, hörde att David hade slagit Hadaresers, konungens i Soba, hela här,
sände han sin son Hadoram till konung David för att hälsa honom och lyckönska honom, därför att han hade givit sig i strid med Hadareser och slagit honom; ty Hadareser hade varit Tous fiende. Han sände ock alla slags kärl av guld, silver och koppar.
Också dessa helgade konung David åt HERREN, likasom han hade gjort med det silver och guld han hade hemfört från alla andra folk: från edoméerna, moabiterna, Ammons barn, filistéerna och amalekiterna.
Och sedan Absai, Serujas son, hade slagit edoméerna i Saltdalen, aderton tusen man,
insatte han fogdar i Edom; och alla edoméer blevo David underdåniga. Så gav HERREN seger åt David, varhelst han drog fram.
David regerade nu över hela Israel; och han skipade lag och rätt åt allt sitt folk.
Joab, Serujas son, hade befälet över krigshären, och Josafat, Ahiluds son, var kansler.
Sadok, Ahitubs son, och Abimelek, Ebjatars son, voro präster, och Sausa var sekreterare.
Benaja, Jojadas son, hade befälet över keretéerna och peletéerna; men Davids söner voro de förnämste vid konungens sida.
En tid härefter dog Nahas, Ammons barns konung, och hans son blev konung efter honom.
Då sade David: »Jag vill bevisa Hanun, Nahas' son, vänskap, eftersom hans fader bevisade mig vänskap.» Och David skickade sändebud för att trösta honom i hans sorg efter fadern. När så Davids tjänare kommo till Ammons barns land, till Hanun, för att trösta honom,
sade Ammons barns furstar till Hanun: »Menar du att David därmed att han sänder tröstare till dig vill visa dig att han ärar din fader? Nej, för att undersöka och fördärva och bespeja landet hava hans tjänare kommit till dig.»
Då tog Hanun Davids tjänare och lät raka dem och skära av deras kläder mitt på, ända uppe vid sätet, och lät dem så gå.
Och man kom och berättade för David vad som hade hänt männen; då sände han bud emot dem, ty männen voro ju mycket vanärade. Och konungen lät säga: »Stannen i Jeriko, till dess edert skägg hinner växa ut, och kommen så tillbaka.»
Då nu Ammons barn insågo att de hade gjort sig förhatliga för David, sände Hanun och Ammons barn ett tusen talenter silver för att leja sig vagnar och ryttare från Aram-Naharaim, från Aram-Maaka och från Soba.
De lejde sig trettiotvå tusen vagnar, ävensom hjälp av konungen i Maaka med hans folk; dessa kommo och lägrade sig framför Medeba. Ammons barn församlade sig ock från sina städer och kommo för att strida.
När David hörde detta, sände han åstad Joab med hela hären, de tappraste krigarna.
Och Ammons barn drogo ut och ställde upp sig till strid vid ingången till staden; men de konungar som hade kommit dit ställde upp sig för sig själva på fältet.
Då Joab nu såg att han hade fiender både framför sig och bakom sig, gjorde han ett urval bland allt Israels utvalda manskap och ställde sedan upp sig mot araméerna.
Men det övriga folket överlämnade han åt sin broder Absai, och dessa fingo ställa upp sig mot Ammons barn.
Och han sade: »Om araméerna bliva mig övermäktiga, så skall du komma mig till hjälp; och om Ammons barn bliva dig övermäktiga, så vill jag hjälpa dig.
Var nu vid gott mod; ja, låt oss visa mod i striden för vårt folk och för vår Guds städer. Sedan må HERREN göra vad honom täckes.
Därefter ryckte Joab fram med sitt folk till strid mot araméerna, och de flydde för honom.
Men när Ammons barn sågo att araméerna flydde, flydde också de för hans broder Absai och begåvo sig in i staden. Då begav sig Joab till Jerusalem.
Då alltså araméerna sågo att de hade blivit slagna av Israel, sände de bud att de araméer som bodde på andra sidan floden skulle rycka ut, anförda av Sofak, Hadaresers härhövitsman.
När detta blev berättat för David, församlade han hela Israel och gick över Jordan, och då han kom fram till dem, ställde han upp sig i slagordning mot dem; och när David hade ställt upp sig till strid mot araméerna, gåvo dessa sig i strid med honom.
Men araméerna flydde undan för Israel, och David dräpte av araméerna manskapet på sju tusen vagnar, så ock fyrtio tusen man fotfolk; härhövitsmannen Sofak dödade han ock.
Följande år, vid den tid då konungarna plägade draga i fält, tågade Joab ut med krigshären och härjade Ammons barns land, och kom så och belägrade Rabba, medan David stannade kvar i Jerusalem. Och Joab intog Rabba och förstörde det.
Och David tog deras konungs krona från hans huvud, den befanns väga en talent guld och var prydd med en dyrbar sten. Den sattes nu på Davids huvud. Och han förde ut byte från staden i stor myckenhet.
Och folket därinne förde han ut och söndersargade dem med sågar och tröskvagnar av järn och med bilor. Så gjorde David mot Ammons barns alla städer. Sedan vände David med allt folket tillbaka till Jerusalem.
Därefter uppstod en strid med filistéerna vid Geser; husatiten Sibbekai slog då ned Sippai, en av rafaéernas avkomlingar; så blevo de kuvade.
Åter stod en strid med filistéerna; Elhanan, Jaurs son, slog då ned Lami, gatiten Goljats broder, som hade ett spjut vars skaft liknade en vävbom.
Åter stod en strid vid Gat. Där var en reslig man som hade sex fingrar och sex tår, tillsammans tjugufyra; han var ock en avkomling av rafaéerna.
Denne smädade Israel; då blev han nedgjord av Jonatan, son till Simea, Davids broder.
Dessa voro avkomlingar av rafaéerna i Gat; och de föllo för Davids och hans tjänares hand.
Men Satan trädde upp mot Israel och uppeggade David till att räkna Israel.
Då sade David till Joab och till folkets andra hövitsman: »Gån åstad och räknen Israel, från Beer-Seba ända till Dan, och given mig besked därom, så att jag får veta huru många de äro.»
Joab svarade: »Må HERREN än vidare föröka sitt folk hundrafalt. Äro de då icke, min herre konung, allasammans min herres tjänare? Varför begär då min herre sådant? Varför skulle man därmed draga skuld över Israel?
Likväl blev konungens befallning gällande, trots Joab. Alltså drog Joab ut och for omkring i hela Israel, och kom så hem igen till Jerusalem.
Och Joab uppgav för David vilken slutsumma folkräkningen utvisade: i Israel funnos tillsammans elva hundra tusen svärdbeväpnade män, och i Juda funnos fyra hundra sjuttio tusen svärdbeväpnade man.
Men Levi och Benjamin hade han icke räknat jämte de andra, ty konungens befallning var en styggelse för Joab.
Vad som hade skett misshagade Gud, och han hemsökte Israel.
Då sade David till Gud: »Jag har syndat storligen däri att jag har gjort detta; men tillgiv nu din tjänares missgärning, ty jag har handlat mycket dåraktigt.»
Men HERREN talade till Gad, Davids siare, och sade:
»Gå och tala till David och säg: Så säger HERREN: Tre ting lägger jag fram för dig; välj bland dem ut åt dig ett som du vill att jag skall göra dig.»
Då gick Gad in till David och sade till honom: »Så säger HERREN:
Tag vilketdera du vill: antingen hungersnöd i tre år, eller förödelse i tre månader genom dina ovänners anfall, utan att du kan undkomma dina fienders svärd, eller HERRENS svärd och pest i landet under tre dagar, i det att HERRENS ängel sprider fördärv inom hela Israels område. Eftersinna nu vilket svar jag skall giva honom som har sänt mig.»
David svarade Gad: »Jag är i stor vånda. Men låt mig då falla i HERRENS hand, ty hans barmhärtighet är mycket stor; i människohand vill jag icke falla.»
Så lät då HERREN pest komma i Israel, så att sjuttio tusen män av Israel föllo.
Och Gud sände en ängel mot Jerusalem till att fördärva det. Men när denne höll på att fördärva, såg HERREN därtill och ångrade det onda, så att han sade till ängeln, Fördärvaren: »Det är nog; drag nu din hand tillbaka.» Och HERRENS ängel stod då vid jebuséen Ornans tröskplats.
När nu David lyfte upp sina ögon och fick se HERRENS ängel stående mellan jorden och himmelen med ett blottat svärd i sin hand, uträckt över Jerusalem, då föllo han och de äldste, höljda i sorgdräkt, ned på sina ansikten.
Och David sade till Gud: »Det var ju jag som befallde att folket skulle räknas. Det är då jag som har syndat och gjort vad ont är; men dessa, min hjord, vad hava de gjort? HERRE, min Gud, må din hand vända sig mot mig och min faders hus, men icke mot ditt folk, så att det bliver hemsökt.»
Men HERRENS ängel befallde Gad att säga till David att David skulle gå åstad och resa ett altare åt HERREN på jebuséen Ornans tröskplats.
Och David gick åstad på grund av det ord som Gad hade talat i HERRENS namn.
Då Ornan nu vände sig om, fick han se ängeln; och hans fyra söner som voro med honom, gömde sig. Men Ornan höll på att tröska vete.
Och David kom till Ornan; när då Ornan såg upp och fick se David, gick han fram ifrån tröskplatsen och föll ned till jorden på sitt ansikte för David.
Och David sade till Ornan: »Giv mig den plats där du tröskar din säd, så att jag där kan bygga ett altare åt HERREN; giv mig den för full betalning; och må så hemsökelsen upphöra bland folket.»
Då sade Ornan till David: »Tag den, och må sedan min herre konungen göra vad honom täckes. Se, här giver jag dig fäkreaturen till brännoffer och tröskvagnarna till ved och vetet till spisoffer; alltsammans giver jag.»
Men konung David svarade Ornan: »Nej, jag vill köpa det för full betalning; ty jag vill icke taga åt HERREN det som är ditt, och offra brännoffer som jag har fått för intet.»
Och David gav åt Ornan för platsen sex hundra siklar guld, i full vikt.
Och David byggde där ett altare åt HERREN och offrade brännoffer och tackoffer. Han ropade till HERREN, och han svarade honom med eld från himmelen på brännoffersaltaret.
Och på HERRENS befallning stack ängeln sitt svärd tillbaka i skidan.
Då, när David förnam att HERREN hade bönhört honom på jebuséen Ornans tröskplats, offrade han där.
Men HERRENS tabernakel, som Mose hade låtit göra i öknen, stod jämte brännoffersaltaret, vid den tiden på offerhöjden i Gibeon.
Dock vågade David icke komma inför Guds ansikte för att söka honom; så förskräckt var han för HERRENS ängels svärd.
Och David sade: »Här skall HERREN Guds hus stå, och här altaret för Israels brännoffer.»
Och David befallde att man skulle samla tillhopa de främlingar som funnos i Israels land; och han anställde hantverkare, som skulle hugga ut stenar för att därmed bygga Guds hus.
Och David anskaffade järn i myckenhet till spikar på dörrarna i portarna och till krampor, så ock koppar i sådan myckenhet att den icke kunde vägas,
och cederbjälkar i otalig mängd; ty sidonierna och tyrierna förde cederträ i myckenhet till David.
David tänkte nämligen: »Min son Salomo är ung och späd, men huset som skall byggas åt HERREN måste göras övermåttan stort, så att det bliver namnkunnigt och prisat i alla länder; jag vill därför skaffa förråd åt honom.» Så skaffade David förråd i myckenhet före sin död.
Och han kallade till sig sin son Salomo och bjöd honom att bygga ett hus åt HERREN, Israels Gud.
Och David sade till sin son Salomo: »Jag hade själv i sinnet att bygga ett hus åt HERRENS, min Guds, namn.
Men HERRENS ord kom till mig; han sade: Du har utgjutit blod i myckenhet och fört stora krig; du skall icke bygga ett hus åt mitt namn, eftersom du har utgjutit så mycket blod på jorden, i min åsyn.
Men se, åt dig skall födas en son; han skall bliva en fridsäll man, och jag skall låta honom få fred med alla sina fiender runt omkring; ty Salomo skall han heta, och frid och ro skall jag låta vila över Israel i hans dagar.
Han skall bygga ett hus åt mitt namn; han skall vara min son, och jag skall vara hans fader. Och jag skall befästa hans konungatron över Israel för evig tid.
Så vare nu HERREN med dig, min son; må du bliva lyckosam och få bygga HERRENS, din Guds, hus, såsom han har lovat om dig.
Må HERREN allenast giva dig klokhet och förstånd, när han sätter dig till härskare över Israel, och förhjälpa dig till att hålla HERRENS, din Guds, lag.
Då skall du bliva lyckosam, om du håller och gör efter de stadgar och rätter som HERREN har bjudit Mose att ålägga Israel. Var frimodig och oförfärad; frukta icke och var icke försagd.
Och se, trots mitt betryck har jag nu anskaffat till HERRENS hus ett hundra tusen talenter guld och tusen gånger tusen talenter silver, därtill av koppar och järn mer än som kan vägas, ty så mycket är det; trävirke och sten har jag ock anskaffat, och mer må du själv anskaffa.
Arbetare har du ock i myckenhet hantverkare, stenhuggare och timmermän, och därtill allahanda folk som är kunnigt i allt slags annat arbete.
På guldet, silvret, kopparen och järnet kan ingen räkning hållas. Upp då och gå till verket; och vare HERREN med dig!»
Därefter bjöd David alla Israels furstar att de skulle understödja hans son Salomo; han sade:
»HERREN, eder Gud, är ju med eder och har låtit eder få ro på alla sidor; ty han har givit landets förra inbyggare i min hand, och landet har blivit HERREN och hans folk underdånigt.
Så vänden nu edert hjärta och eder själ till att söka HERREN, eder Gud; och stån upp och byggen HERREN Guds helgedom, så att man kan föra HERRENS förbundsark och vad annat som hör till Guds helgedom in i det hus som skall byggas åt HERRENS namn.»
Och när David blev gammal och levnadsmätt, gjorde han sin son Salomo till konung över Israel.
Och han församlade alla Israels furstar, så ock prästerna och leviterna.
Och leviterna blevo räknade, de nämligen som voro trettio år gamla eller därutöver; och deras antal, antalet av alla personer av mankön, utgjorde trettioåtta tusen.
»Av dessa», sade han, »skola tjugufyra tusen förestå sysslorna vid HERRENS hus, och sex tusen vara tillsyningsmän och domare;
fyra tusen skola vara dörrvaktare och fyra tusen skola lovsjunga HERREN till de instrumenter som jag har låtit göra för lovsången.»
Och David delade dem i avdelningar efter Levis söner, Gerson Kehat och Merari.
Till gersoniterna hörde Laedan och Simei.
Laedans söner voro Jehiel, huvudmannen, Setam och Joel, tillsammans tre.
Simeis söner voro Selomot, Hasiel och Haran, tillsammans tre. Dessa voro huvudmän för Laedans familjer.
Och Simeis söner voro Jahat, Sina, Jeus och Beria. Dessa voro Simeis söner, tillsammans fyra.
Jahat var huvudmannen, och Sisa var den andre. Men Jeus och Beria hade icke många barn; därför fingo de utgöra allenast en familj, en ordning.
Kehats söner voro Amram, Jishar, Hebron och Ussiel, tillsammans fyra.
Amrams söner voro Aron och Mose. Och Aron blev jämte sina söner för evärdlig tid avskild till att helgas såsom höghelig, till att för evärdlig tid antända rökelse inför HERREN och göra tjänst inför honom och välsigna i hans namn.
Men gudsmannen Moses söner räknades till Levi stam.
Moses söner voro Gersom och Elieser.
Gersoms söner voro Sebuel, huvudmannen.
Och Eliesers söner voro Rehabja, huvudmannen. Elieser hade inga andra söner; men Rehabjas söner voro övermåttan talrika.
Jishars söner voro Selomit, huvudmannen.
Hebrons söner voro Jeria, huvudmannen, Amarja, den andre, Jahasiel, den tredje, och Jekameam, den fjärde.
Ussiels söner voro Mika, huvudmannen, och Jissia, den andre.
