grundläggande information
historia
trafik
religion
beslutsfattande och påverkan
grundläggande information
Karleby finns i Mellersta Österbotten invid Bottniska viken .
Karleby stad är grundad 1620 och hette då Gamlakarleby .
senare blev Kokkola stadens finska namn .
vid Karleby centrum finns en av landets mest omfattande historiska trästadshelheter .
Stadsplanen är från 1650 @-@ talet .
den omfattar 12 kvarter med hundratals trähus och gårdsbyggnader .
de äldsta av dessa är från 1600 @-@ talet .
Karleby är en kulturstad med mycket att se och uppleva .
Karleby hamn ligger i stadsdelen Yxpila och är en av Finlands mest trafikerade godshamnar .
Grunden för näringslivet i Karleby är den internationella storindustrin .
i Karleby är den kemiska industrin och industri i anslutning till denna särskilt viktig .
Karleby är även en betydande handelsstad .
information om Karlebyfinska _ svenska _ engelska
historia
redan under medeltiden fanns det hamn , båtbygge och handelsplats i Karleby .
Landhöjningen har varit en central faktor i Karlebys historia .
den har format omgivningen i hög grad och bland annat påverkat utvecklingen av hamnverksamheten och handeln .
Handel bedrevs längs med Bottniska vikens kust och jordbruk , jakt , fiske och sälfångst var även viktiga näringar .
Exporten av tjära , som blev mycket viktig för Karlebys historia , inleddes redan på 1500 @-@ talet .
den sjunde september 1620 undertecknade Sveriges kung Gustav II Adolf en handling som gav den lilla jordbruks- och fiskebyn vid Ristrand status som stad .
Dagens stadssund var då en smal havsvik som sträckte sig ända till Kyrkbacken .
Sakta men säkert blev Karleby en viktig stad för sjöfart och skeppsbygge .
Skeppsvarv fanns bland annat i Kaustarviken , Svartskär och Soldatskär .
Inledningsvis seglade man endast till Åbo och Stockholm , eftersom Karleby som s.k. uppstad inte fick bedriva utrikeshandel .
år 1765 erhöll staden stapelrättigheter , dvs. rätt till fri utrikeshandel , främst tack vare den aktiva kyrkoherden och lantdagsmannen Anders Chydenius .
Karleby blev snabbt en förmögen stad i början av 1800 @-@ talet tack vare just handeln med tjära och rederiverksamheten .
stadens borgare köpte tjära av bönder och exporterade den , ofta till hamnar vid Medelhavet och i England .
Karleby handelsflotta var under perioder Finlands största .
den snabba ekonomiska utvecklingen avtog i mitten av 1800 @-@ talet , men tog ny fart i slutet av århundradet tack vare industrialiseringen .
Karleby blev en viktig industristad främst tack vare läder- och metallindustrin .
Karlebys historiafinska _ svenska _ engelska
trafik
Karleby har goda trafikförbindelser .
via Karleby löper riksväg 8 och 13 .
Järnvägsstationen finns i stadens centrum .
Restiden med tåg till Helsingfors är cirka fyra timmar .
Flygplatsen finns i Kronoby på endast 22 kilometers avstånd från Karleby centrum .
Stadsborna erbjuds även ett tryggt , omfattande , fungerande och trivsamt nätverk för den lätta trafiken .
Karleby har satsat på att förbättra förhållandena för cyklister .
Lokalbussarna trafikerar de olika delarna av staden på vardagar .
Läs mer : trafik .
Gator och trafikfinska _ svenska
Kollektivtrafikfinska _ svenska
linkkiVR :
Tågtidtabellerfinska _ svenska _ engelska _ ryska
Busstidtabellerfinska _ svenska _ engelska
flyg från Karleby @-@ Jakobstad flygplatsfinska _ svenska _ engelska
religion
i Karleby finns flera olika religiösa samfund .
i tjänsten Uskonnot Suomessa ( Religioner i Finland ) finns information om religiösa samfund enligt ort .
den evangelisk @-@ lutherska kyrkan har fyra finskspråkiga församlingar och en svenskspråkig församling i Karleby .
Läs mer på Karleby kyrkliga samfällighets webbplats .
i Karleby finns en ortodox kyrka .
mer information om den ortodoxa församlingens verksamhet i Karleby finns på Vasa ortodoxa församlings webbplats .
Läs mer : kulturer och religioner i Finland .
linkkiKarleby kyrkliga samfällighet :
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiVasa ortodoxa församling :
Vasa ortodoxa församlingfinska _ engelska _ ryska
beslutsfattande och påverkan
den högsta beslutsfattande makten i Karleby stad innehas av stadsfullmäktige .
Fullmäktigeledamöterna och deras suppleanter väljs vid kommunalval vart fjärde år .
på stadens webbplats finns information om stadsfullmäktige och dess beslut .
invånarna kan påverka stadens beslutsfattande redan då beslut bereds .
information om olika sätt att delta och påverka finns på stadens webbplats .
kommunens invånare har enligt kommunallagen rätt att lämna in motioner till kommunen i ärenden som gäller dess verksamhet .
i Karleby finns ungdomsfullmäktige , äldre- och handikappråd samt ett råd för kulturell mångfald .
Läs mer : Finlands förvaltning , Val och röstning i Finland
beslutsfattandefinska _ svenska _ engelska
grundläggande information
historia
trafik
religion
beslutsfattande och påverkan
grundläggande information
Karleby finns i Mellersta Österbotten invid Bottniska viken .
Karleby stad är grundad 1620 och hette då Gamlakarleby .
senare blev Kokkola stadens finska namn .
vid Karleby centrum finns en av landets mest omfattande historiska trästadshelheter .
Stadsplanen är från 1650 @-@ talet .
den omfattar 12 kvarter med hundratals trähus och gårdsbyggnader .
de äldsta av dessa är från 1600 @-@ talet .
Karleby är en kulturstad med mycket att se och uppleva .
Karleby hamn ligger i stadsdelen Yxpila och är en av Finlands mest trafikerade godshamnar .
Grunden för näringslivet i Karleby är den internationella storindustrin .
i Karleby är den kemiska industrin och industri i anslutning till denna särskilt viktig .
Karleby är även en betydande handelsstad .
information om Karlebyfinska _ svenska _ engelska
historia
redan under medeltiden fanns det hamn , båtbygge och handelsplats i Karleby .
Landhöjningen har varit en central faktor i Karlebys historia .
den har format omgivningen i hög grad och bland annat påverkat utvecklingen av hamnverksamheten och handeln .
Handel bedrevs längs med Bottniska vikens kust och jordbruk , jakt , fiske och sälfångst var även viktiga näringar .
Exporten av tjära , som blev mycket viktig för Karlebys historia , inleddes redan på 1500 @-@ talet .
den sjunde september 1620 undertecknade Sveriges kung Gustav II Adolf en handling som gav den lilla jordbruks- och fiskebyn vid Ristrand status som stad .
Dagens stadssund var då en smal havsvik som sträckte sig ända till Kyrkbacken .
Sakta men säkert blev Karleby en viktig stad för sjöfart och skeppsbygge .
Skeppsvarv fanns bland annat i Kaustarviken , Svartskär och Soldatskär .
Inledningsvis seglade man endast till Åbo och Stockholm , eftersom Karleby som s.k. uppstad inte fick bedriva utrikeshandel .
år 1765 erhöll staden stapelrättigheter , dvs. rätt till fri utrikeshandel , främst tack vare den aktiva kyrkoherden och lantdagsmannen Anders Chydenius .
Karleby blev snabbt en förmögen stad i början av 1800 @-@ talet tack vare just handeln med tjära och rederiverksamheten .
stadens borgare köpte tjära av bönder och exporterade den , ofta till hamnar vid Medelhavet och i England .
Karleby handelsflotta var under perioder Finlands största .
den snabba ekonomiska utvecklingen avtog i mitten av 1800 @-@ talet , men tog ny fart i slutet av århundradet tack vare industrialiseringen .
Karleby blev en viktig industristad främst tack vare läder- och metallindustrin .
Karlebys historiafinska _ svenska _ engelska
trafik
Karleby har goda trafikförbindelser .
via Karleby löper riksväg 8 och 13 .
Järnvägsstationen finns i stadens centrum .
Restiden med tåg till Helsingfors är cirka fyra timmar .
Flygplatsen finns i Kronoby på endast 22 kilometers avstånd från Karleby centrum .
Stadsborna erbjuds även ett tryggt , omfattande , fungerande och trivsamt nätverk för den lätta trafiken .
Karleby har satsat på att förbättra förhållandena för cyklister .
Lokalbussarna trafikerar de olika delarna av staden på vardagar .
Läs mer : trafik .
Gator och trafikfinska _ svenska
Kollektivtrafikfinska _ svenska
linkkiVR :
Tågtidtabellerfinska _ svenska _ engelska _ ryska
Busstidtabellerfinska _ svenska _ engelska
flyg från Karleby @-@ Jakobstad flygplatsfinska _ svenska _ engelska
religion
i Karleby finns flera olika religiösa samfund .
i tjänsten Uskonnot Suomessa ( Religioner i Finland ) finns information om religiösa samfund enligt ort .
den evangelisk @-@ lutherska kyrkan har fyra finskspråkiga församlingar och en svenskspråkig församling i Karleby .
Läs mer på Karleby kyrkliga samfällighets webbplats .
i Karleby finns en ortodox kyrka .
mer information om den ortodoxa församlingens verksamhet i Karleby finns på Vasa ortodoxa församlings webbplats .
Läs mer : kulturer och religioner i Finland .
linkkiKarleby kyrkliga samfällighet :
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiVasa ortodoxa församling :
Vasa ortodoxa församlingfinska _ engelska _ ryska
beslutsfattande och påverkan
den högsta beslutsfattande makten i Karleby stad innehas av stadsfullmäktige .
Fullmäktigeledamöterna och deras suppleanter väljs vid kommunalval vart fjärde år .
på stadens webbplats finns information om stadsfullmäktige och dess beslut .
invånarna kan påverka stadens beslutsfattande redan då beslut bereds .
information om olika sätt att delta och påverka finns på stadens webbplats .
kommunens invånare har enligt kommunallagen rätt att lämna in motioner till kommunen i ärenden som gäller dess verksamhet .
i Karleby finns ungdomsfullmäktige , äldre- och handikappråd samt ett råd för kulturell mångfald .
Läs mer : Finlands förvaltning , Val och röstning i Finland
beslutsfattandefinska _ svenska _ engelska
grundläggande information
historia
trafik
religion
beslutsfattande och påverkan
grundläggande information
Karleby finns i Mellersta Österbotten invid Bottniska viken .
Karleby stad är grundad 1620 och hette då Gamlakarleby .
senare blev Kokkola stadens finska namn .
vid Karleby centrum finns en av landets mest omfattande historiska trästadshelheter .
Stadsplanen är från 1650 @-@ talet .
den omfattar 12 kvarter med hundratals trähus och gårdsbyggnader .
de äldsta av dessa är från 1600 @-@ talet .
Karleby är en kulturstad med mycket att se och uppleva .
Karleby hamn ligger i stadsdelen Yxpila och är en av Finlands mest trafikerade godshamnar .
Grunden för näringslivet i Karleby är den internationella storindustrin .
i Karleby är den kemiska industrin och industri i anslutning till denna särskilt viktig .
Karleby är även en betydande handelsstad .
information om Karlebyfinska _ svenska _ engelska
historia
redan under medeltiden fanns det hamn , båtbygge och handelsplats i Karleby .
Landhöjningen har varit en central faktor i Karlebys historia .
den har format omgivningen i hög grad och bland annat påverkat utvecklingen av hamnverksamheten och handeln .
Handel bedrevs längs med Bottniska vikens kust och jordbruk , jakt , fiske och sälfångst var även viktiga näringar .
Exporten av tjära , som blev mycket viktig för Karlebys historia , inleddes redan på 1500 @-@ talet .
den sjunde september 1620 undertecknade Sveriges kung Gustav II Adolf en handling som gav den lilla jordbruks- och fiskebyn vid Ristrand status som stad .
Dagens stadssund var då en smal havsvik som sträckte sig ända till Kyrkbacken .
Sakta men säkert blev Karleby en viktig stad för sjöfart och skeppsbygge .
Skeppsvarv fanns bland annat i Kaustarviken , Svartskär och Soldatskär .
Inledningsvis seglade man endast till Åbo och Stockholm , eftersom Karleby som s.k. uppstad inte fick bedriva utrikeshandel .
år 1765 erhöll staden stapelrättigheter , dvs. rätt till fri utrikeshandel , främst tack vare den aktiva kyrkoherden och lantdagsmannen Anders Chydenius .
Karleby blev snabbt en förmögen stad i början av 1800 @-@ talet tack vare just handeln med tjära och rederiverksamheten .
stadens borgare köpte tjära av bönder och exporterade den , ofta till hamnar vid Medelhavet och i England .
Karleby handelsflotta var under perioder Finlands största .
den snabba ekonomiska utvecklingen avtog i mitten av 1800 @-@ talet , men tog ny fart i slutet av århundradet tack vare industrialiseringen .
Karleby blev en viktig industristad främst tack vare läder- och metallindustrin .
Karlebys historiafinska _ svenska _ engelska
trafik
Karleby har goda trafikförbindelser .
via Karleby löper riksväg 8 och 13 .
Järnvägsstationen finns i stadens centrum .
Restiden med tåg till Helsingfors är cirka fyra timmar .
Flygplatsen finns i Kronoby på endast 22 kilometers avstånd från Karleby centrum .
Stadsborna erbjuds även ett tryggt , omfattande , fungerande och trivsamt nätverk för den lätta trafiken .
Karleby har satsat på att förbättra förhållandena för cyklister .
Lokalbussarna trafikerar de olika delarna av staden på vardagar .
Läs mer : trafik .
Gator och trafikfinska _ svenska
Kollektivtrafikfinska _ svenska
linkkiVR :
Tågtidtabellerfinska _ svenska _ engelska _ ryska
Busstidtabellerfinska _ svenska _ engelska
flyg från Karleby @-@ Jakobstad flygplatsfinska _ svenska _ engelska
religion
i Karleby finns flera olika religiösa samfund .
i tjänsten Uskonnot Suomessa ( Religioner i Finland ) finns information om religiösa samfund enligt ort .
den evangelisk @-@ lutherska kyrkan har fyra finskspråkiga församlingar och en svenskspråkig församling i Karleby .
Läs mer på Karleby kyrkliga samfällighets webbplats .
i Karleby finns en ortodox kyrka .
mer information om den ortodoxa församlingens verksamhet i Karleby finns på Vasa ortodoxa församlings webbplats .
Läs mer : kulturer och religioner i Finland .
linkkiKarleby kyrkliga samfällighet :
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiVasa ortodoxa församling :
Vasa ortodoxa församlingfinska _ engelska _ ryska
beslutsfattande och påverkan
den högsta beslutsfattande makten i Karleby stad innehas av stadsfullmäktige .
Fullmäktigeledamöterna och deras suppleanter väljs vid kommunalval vart fjärde år .
på stadens webbplats finns information om stadsfullmäktige och dess beslut .
invånarna kan påverka stadens beslutsfattande redan då beslut bereds .
information om olika sätt att delta och påverka finns på stadens webbplats .
kommunens invånare har enligt kommunallagen rätt att lämna in motioner till kommunen i ärenden som gäller dess verksamhet .
i Karleby finns ungdomsfullmäktige , äldre- och handikappråd samt ett råd för kulturell mångfald .
Läs mer : Finlands förvaltning , Val och röstning i Finland
beslutsfattandefinska _ svenska _ engelska
detta innehåll finns inte på det språk som du har valt .
Välj något annat språk .
finska
detta innehåll finns inte på det språk som du har valt .
Välj något annat språk .
finska
detta innehåll finns inte på det språk som du har valt .
Välj något annat språk .
finska
bibliotek
motion
att röra sig i naturen
teater och film
museer
hobbyer för barn och unga
föreningar
Karleby är en gammal sjöstad som erbjuder mångsidiga möjligheter för utfärder och friluftsliv .
personer ntresserad av friluftsliv bör läsa mer om allemansrätten under rubriken &quot; Att röra sig i naturen &quot; i denna tjänst .
flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet .
föreningar och organisationer samt hobbygrupper och kommunala institut erbjuder kurser i idrott och kultur samt bl.a. språk och hantverk .
i Snellman @-@ salen och i stadens övriga kulturlokaler erbjuds kulturevenemang av varierande slag .
Årliga evenemang i Karleby är bland annat Veneziansk afton i slutet av sommaren , Kokkola Cup för fotbollsjuniorer , Stadsfestivalen Karleby sommarveckor , Lochteå kyrkomusikfest samt Vinterdans i Karleby och festivalen Karleby Vinterharmonika .
mer information om fritidstjänsterna i Karleby finns på Karleby stads webbplats .
på stadens webbplats finns även en länk till Evenemangskalendern med daglig information om stadens kultur- och motionsevenemang .
Läs mer : Fritid .
Evenemangskalenderfinska
Kulturtjänsterfinska _ svenska _ engelska
Idrottstjänsterfinska _ svenska _ engelska
bibliotek
Karleby stadsbibliotek finns i stadens centrum .
Närbiblioteken finns i Björkhagen , Kelviå , Lochteå samt Ullava kyrkby och Rahkonen .
information om bibliotekets öppettider och tjänster finns på dess webbplats .
biblioteket finns även på nätet .
där kan kunderna bläddra i bibliotekets samlingar , reservera material , förnya sina lån , beställa fjärrlån och låna e @-@ böcker under alla tider på dygnet .
tack vare det effektiva biblioteksnätverket i Finland är nästan alla finländska biblioteks samlingar tillgängliga för bibliotekskunderna i Karleby .
Karleby stadsbibliotek / huvudbiblioteket
Storgatan 3 , 67100 Karleby
telefon : 040.806.5124 , 040.806.5133
Läs mer : bibliotek .
Bibliotekstjänsterfinska _ svenska _ engelska
motion
i Karleby finns mångsidiga motionsmöjligheter året runt .
staden anordnar ledda aktiviteter i Simcentret VesiVeijari och motionshallarna .
dessutom finns det gym av flera olika slag .
gym anpassade för äldre finns i Furuåsens aktivitetscenter och Kuusikumpu servicehus .
staden underhåller cykelvägar , motionsrutter , joggingbanor , skidspår , badstränder , bollplaner och skridskobanor samt platser för närmotion .
i Karlebynejdens instituts nättjänst finns information om institutets mångsidiga motionsutbud .
i Karleby finns nära på hundra idrottsföreningar för olika grenar samt föreningar som arrangerar övrig motion .
mer information om motionsmöjligheter i Karleby finns på Karleby stads webbplats .
Läs mer :
motion .
Idrottstjänsterfinska _ svenska _ engelska
Motionsplatserfinska _ svenska
gym för äldrefinska
Karlebynejdens institutfinska _ svenska
att röra sig i naturen
att röra sig i naturen är en traditionell och populär form av avkoppling för finländarna under alla årstider .
i Finland kan man med stöd av allemansrätten plocka bär och svamp i skogen och röra sig till fots , med cykel eller skidor vintertid .
det är inte tillåtet att beträda folks gårdar utan lov .
för fiske krävs fiskelov , med undantag för mete och pilkning .
även jakt fordrar jakttillstånd .
allemansrätten ger inte rätt att skräpa ner i naturen , skada träd eller växter , störa eller skada fågelbon eller fågelungar , köra motorfordon utan markägarens tillstånd eller bygga ens tillfälliga byggen .
mer information om motionsrutterna , rastplatser , möjligheter till fiske och båtliv samt exempelvis fågeltorn i Karleby finns på stadens webbplats .
rutterna för camping , paddling , vandring , cykling och övriga rutter i Karleby finns i karttjänsten på nätet .
i karttjänsten visas även var största delen av motionsplatserna finns .
du kan köpa friluftskartor över Karleby hos Karleby Turism : Salutorget 5 , 67100 Karleby .
Läs mer : att röra sig i naturen .
linkkiMiljöförvaltningen :
Allemansrättenfinska _ svenska _ engelska _ ryska
Motionskarta över Karlebyfinska _ svenska
motionsrutter i Karlebyfinska _ svenska
teater och film
Karleby är en teaterstad med långa anor , som erbjuder scenkonst på hög nivå framförd av både proffs och amatörer .
Karleby stadsteater finns i det stämningsfulla Vartiolinna ( Torggatan 48 ) .
du kan läsa mer om amatörteatrarnas verksamhet på deras webbplats och i evenemangskalendern .
i Karleby finns biografen Bio Rex , vars två salar använder digital- och 3D @-@ teknik .
Bio Rex program finns under länken här intill .
Läs mer : teater och film .
Stadsteaternfinska
Biograffinska
teater och danskonst i Karlebyfinska _ svenska _ engelska
Evenemangskalenderfinska
museer
i hjärtat av staden , i det anrika Rooska gården , finns K.H.Renlunds museum .
Karleby stad grundade museet 1909 utgående från en testamentsgåva av affärsmannen Karl Herman Renlund ( 1850 @-@ 1908 ) .
på museet finns Renlunds samling av finländsk konst från guldåldern och tillfälliga utställningar i en kulturhistorisk miljö .
även i museikvarterens övriga byggnader finns utställningar om stadens kulturhistoria och utställningar med ITE @-@ konst .
på K.H.Renlunds museums webbplats finns mer information om museets tjänster , utställningar samt aktuell verksamhet .
Utöver K.H.Renlunds museum lönar det sig att besöka det naturhistoriska museet Kieppi ( Kieppi är stängt tills vidare på grund av brand ) samt de många hembygdsmuseerna och övriga de historiska resmålen i regionen .
exempelvis i Konst @-@ Vionoja @-@ centret presenteras konstnären Veikko Vionojas verk .
i Kelviå , ca 10 km norrut från Karleby , finns Toivonen djurpark och drängmuseum .
mer information om dessa museer finns under länkarna här intill .
Läs mer : museer .
museer och traditionsarbetefinska _ svenska _ engelska
K.H. Renlunds museum - Mellersta Österbottens landskapsmuseumfinska _ svenska _ engelska
Kieppi , Karleby naturvetenskapliga museumfinska _ svenska _ engelska
linkkiToivonens djurpark och drängmuseum :
Toivonens djurpark och drängmuseum finska _ svenska _ engelska
konst Vionojafinska
hobbyer för barn och unga
flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet .
flera olika föreningar samt kommunala institut ger unga möjlighet att studera idrott och kultur samt bl.a. språk och hantverk .
barn och unga kan delta i grundläggande undervisning i musik , dans , bildkonst och hantverk .
dessutom erbjuder stadens ungdomstjänster en rockskola .
stadens ungdomstjänster driver sju ungdomsgårdar runt om i Karleby .
de rusmedels- och rökfria ungdomslokalerna erbjuder handledd verksamhet för barn i årskurserna 3 @-@ 6 och unga i åldern 13 @-@ 17 år i olika delar av Karleby .
information om hobbyverksamheter för barn och unga finns på stadens webbplats .
rådgivningen vid Ungdomsgården Vinge ger aktuell information om bl.a. internationalisering , studier , arbetsliv , hälsa , hobbyverksamhet och boende .
Karlebynejdens institut erbjuder barn och unga olika former av hobbyverksamhet , exempelvis i konstämnen och musik .
kontrollera vilka kurser som är aktuella i institutets webbtjänst .
Karleby evangelisk @-@ lutherska församlingar erbjuder även hobbyverksamhet för barn och unga , såsom lekparksträffar , klubbar , musikverksamhet och läger .
mer information om verksamheten finns på Karleby församlingssammanslutnings webbplats .
ungdomsgården Vinge
67100 Karleby
Läs mer : hobbyer för barn och unga .
övrig undervisning i Karlebyfinska _ svenska
Ungdomstjänsterfinska _ svenska _ engelska
Karlebynejdens institutfinska _ svenska
linkkiKarleby kyrkliga samfällighet :
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
föreningar
Karleby har ett aktivt och mångsidigt föreningsliv för invånare i alla åldrar .
Läs mer : föreningar .
bibliotek
motion
att röra sig i naturen
teater och film
museer
hobbyer för barn och unga
föreningar
Karleby är en gammal sjöstad som erbjuder mångsidiga möjligheter för utfärder och friluftsliv .
personer ntresserad av friluftsliv bör läsa mer om allemansrätten under rubriken &quot; Att röra sig i naturen &quot; i denna tjänst .
flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet .
föreningar och organisationer samt hobbygrupper och kommunala institut erbjuder kurser i idrott och kultur samt bl.a. språk och hantverk .
i Snellman @-@ salen och i stadens övriga kulturlokaler erbjuds kulturevenemang av varierande slag .
Årliga evenemang i Karleby är bland annat Veneziansk afton i slutet av sommaren , Kokkola Cup för fotbollsjuniorer , Stadsfestivalen Karleby sommarveckor , Lochteå kyrkomusikfest samt Vinterdans i Karleby och festivalen Karleby Vinterharmonika .
mer information om fritidstjänsterna i Karleby finns på Karleby stads webbplats .
på stadens webbplats finns även en länk till Evenemangskalendern med daglig information om stadens kultur- och motionsevenemang .
Läs mer : Fritid .
Evenemangskalenderfinska
Kulturtjänsterfinska _ svenska _ engelska
Idrottstjänsterfinska _ svenska _ engelska
bibliotek
Karleby stadsbibliotek finns i stadens centrum .
Närbiblioteken finns i Björkhagen , Kelviå , Lochteå samt Ullava kyrkby och Rahkonen .
information om bibliotekets öppettider och tjänster finns på dess webbplats .
biblioteket finns även på nätet .
där kan kunderna bläddra i bibliotekets samlingar , reservera material , förnya sina lån , beställa fjärrlån och låna e @-@ böcker under alla tider på dygnet .
tack vare det effektiva biblioteksnätverket i Finland är nästan alla finländska biblioteks samlingar tillgängliga för bibliotekskunderna i Karleby .
Karleby stadsbibliotek / huvudbiblioteket
Storgatan 3 , 67100 Karleby
telefon : 040.806.5124 , 040.806.5133
Läs mer : bibliotek .
Bibliotekstjänsterfinska _ svenska _ engelska
motion
i Karleby finns mångsidiga motionsmöjligheter året runt .
staden anordnar ledda aktiviteter i Simcentret VesiVeijari och motionshallarna .
dessutom finns det gym av flera olika slag .
gym anpassade för äldre finns i Furuåsens aktivitetscenter och Kuusikumpu servicehus .
staden underhåller cykelvägar , motionsrutter , joggingbanor , skidspår , badstränder , bollplaner och skridskobanor samt platser för närmotion .
i Karlebynejdens instituts nättjänst finns information om institutets mångsidiga motionsutbud .
i Karleby finns nära på hundra idrottsföreningar för olika grenar samt föreningar som arrangerar övrig motion .
mer information om motionsmöjligheter i Karleby finns på Karleby stads webbplats .
Läs mer :
motion .
Idrottstjänsterfinska _ svenska _ engelska
Motionsplatserfinska _ svenska
gym för äldrefinska
Karlebynejdens institutfinska _ svenska
att röra sig i naturen
att röra sig i naturen är en traditionell och populär form av avkoppling för finländarna under alla årstider .
i Finland kan man med stöd av allemansrätten plocka bär och svamp i skogen och röra sig till fots , med cykel eller skidor vintertid .
det är inte tillåtet att beträda folks gårdar utan lov .
för fiske krävs fiskelov , med undantag för mete och pilkning .
även jakt fordrar jakttillstånd .
allemansrätten ger inte rätt att skräpa ner i naturen , skada träd eller växter , störa eller skada fågelbon eller fågelungar , köra motorfordon utan markägarens tillstånd eller bygga ens tillfälliga byggen .
mer information om motionsrutterna , rastplatser , möjligheter till fiske och båtliv samt exempelvis fågeltorn i Karleby finns på stadens webbplats .
rutterna för camping , paddling , vandring , cykling och övriga rutter i Karleby finns i karttjänsten på nätet .
i karttjänsten visas även var största delen av motionsplatserna finns .
du kan köpa friluftskartor över Karleby hos Karleby Turism : Salutorget 5 , 67100 Karleby .
Läs mer : att röra sig i naturen .
linkkiMiljöförvaltningen :
Allemansrättenfinska _ svenska _ engelska _ ryska
Motionskarta över Karlebyfinska _ svenska
motionsrutter i Karlebyfinska _ svenska
teater och film
Karleby är en teaterstad med långa anor , som erbjuder scenkonst på hög nivå framförd av både proffs och amatörer .
Karleby stadsteater finns i det stämningsfulla Vartiolinna ( Torggatan 48 ) .
du kan läsa mer om amatörteatrarnas verksamhet på deras webbplats och i evenemangskalendern .
i Karleby finns biografen Bio Rex , vars två salar använder digital- och 3D @-@ teknik .
Bio Rex program finns under länken här intill .
Läs mer : teater och film .
Stadsteaternfinska
Biograffinska
teater och danskonst i Karlebyfinska _ svenska _ engelska
Evenemangskalenderfinska
museer
i hjärtat av staden , i det anrika Rooska gården , finns K.H.Renlunds museum .
Karleby stad grundade museet 1909 utgående från en testamentsgåva av affärsmannen Karl Herman Renlund ( 1850 @-@ 1908 ) .
på museet finns Renlunds samling av finländsk konst från guldåldern och tillfälliga utställningar i en kulturhistorisk miljö .
även i museikvarterens övriga byggnader finns utställningar om stadens kulturhistoria och utställningar med ITE @-@ konst .
på K.H.Renlunds museums webbplats finns mer information om museets tjänster , utställningar samt aktuell verksamhet .
Utöver K.H.Renlunds museum lönar det sig att besöka det naturhistoriska museet Kieppi ( Kieppi är stängt tills vidare på grund av brand ) samt de många hembygdsmuseerna och övriga de historiska resmålen i regionen .
exempelvis i Konst @-@ Vionoja @-@ centret presenteras konstnären Veikko Vionojas verk .
i Kelviå , ca 10 km norrut från Karleby , finns Toivonen djurpark och drängmuseum .
mer information om dessa museer finns under länkarna här intill .
Läs mer : museer .
museer och traditionsarbetefinska _ svenska _ engelska
K.H. Renlunds museum - Mellersta Österbottens landskapsmuseumfinska _ svenska _ engelska
Kieppi , Karleby naturvetenskapliga museumfinska _ svenska _ engelska
linkkiToivonens djurpark och drängmuseum :
Toivonens djurpark och drängmuseum finska _ svenska _ engelska
konst Vionojafinska
hobbyer för barn och unga
flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet .
flera olika föreningar samt kommunala institut ger unga möjlighet att studera idrott och kultur samt bl.a. språk och hantverk .
barn och unga kan delta i grundläggande undervisning i musik , dans , bildkonst och hantverk .
dessutom erbjuder stadens ungdomstjänster en rockskola .
stadens ungdomstjänster driver sju ungdomsgårdar runt om i Karleby .
de rusmedels- och rökfria ungdomslokalerna erbjuder handledd verksamhet för barn i årskurserna 3 @-@ 6 och unga i åldern 13 @-@ 17 år i olika delar av Karleby .
information om hobbyverksamheter för barn och unga finns på stadens webbplats .
rådgivningen vid Ungdomsgården Vinge ger aktuell information om bl.a. internationalisering , studier , arbetsliv , hälsa , hobbyverksamhet och boende .
Karlebynejdens institut erbjuder barn och unga olika former av hobbyverksamhet , exempelvis i konstämnen och musik .
kontrollera vilka kurser som är aktuella i institutets webbtjänst .
Karleby evangelisk @-@ lutherska församlingar erbjuder även hobbyverksamhet för barn och unga , såsom lekparksträffar , klubbar , musikverksamhet och läger .
mer information om verksamheten finns på Karleby församlingssammanslutnings webbplats .
ungdomsgården Vinge
67100 Karleby
Läs mer : hobbyer för barn och unga .
övrig undervisning i Karlebyfinska _ svenska
Ungdomstjänsterfinska _ svenska _ engelska
Karlebynejdens institutfinska _ svenska
linkkiKarleby kyrkliga samfällighet :
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
föreningar
Karleby har ett aktivt och mångsidigt föreningsliv för invånare i alla åldrar .
Läs mer : föreningar .
bibliotek
motion
att röra sig i naturen
teater och film
museer
hobbyer för barn och unga
föreningar
Karleby är en gammal sjöstad som erbjuder mångsidiga möjligheter för utfärder och friluftsliv .
personer ntresserad av friluftsliv bör läsa mer om allemansrätten under rubriken &quot; Att röra sig i naturen &quot; i denna tjänst .
flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet .
föreningar och organisationer samt hobbygrupper och kommunala institut erbjuder kurser i idrott och kultur samt bl.a. språk och hantverk .
i Snellman @-@ salen och i stadens övriga kulturlokaler erbjuds kulturevenemang av varierande slag .
Årliga evenemang i Karleby är bland annat Veneziansk afton i slutet av sommaren , Kokkola Cup för fotbollsjuniorer , Stadsfestivalen Karleby sommarveckor , Lochteå kyrkomusikfest samt Vinterdans i Karleby och festivalen Karleby Vinterharmonika .
mer information om fritidstjänsterna i Karleby finns på Karleby stads webbplats .
på stadens webbplats finns även en länk till Evenemangskalendern med daglig information om stadens kultur- och motionsevenemang .
Läs mer : Fritid .
Evenemangskalenderfinska
Kulturtjänsterfinska _ svenska _ engelska
Idrottstjänsterfinska _ svenska _ engelska
bibliotek
Karleby stadsbibliotek finns i stadens centrum .
Närbiblioteken finns i Björkhagen , Kelviå , Lochteå samt Ullava kyrkby och Rahkonen .
information om bibliotekets öppettider och tjänster finns på dess webbplats .
biblioteket finns även på nätet .
där kan kunderna bläddra i bibliotekets samlingar , reservera material , förnya sina lån , beställa fjärrlån och låna e @-@ böcker under alla tider på dygnet .
tack vare det effektiva biblioteksnätverket i Finland är nästan alla finländska biblioteks samlingar tillgängliga för bibliotekskunderna i Karleby .
Karleby stadsbibliotek / huvudbiblioteket
Storgatan 3 , 67100 Karleby
telefon : 040.806.5124 , 040.806.5133
Läs mer : bibliotek .
Bibliotekstjänsterfinska _ svenska _ engelska
motion
i Karleby finns mångsidiga motionsmöjligheter året runt .
staden anordnar ledda aktiviteter i Simcentret VesiVeijari och motionshallarna .
dessutom finns det gym av flera olika slag .
gym anpassade för äldre finns i Furuåsens aktivitetscenter och Kuusikumpu servicehus .
staden underhåller cykelvägar , motionsrutter , joggingbanor , skidspår , badstränder , bollplaner och skridskobanor samt platser för närmotion .
i Karlebynejdens instituts nättjänst finns information om institutets mångsidiga motionsutbud .
i Karleby finns nära på hundra idrottsföreningar för olika grenar samt föreningar som arrangerar övrig motion .
mer information om motionsmöjligheter i Karleby finns på Karleby stads webbplats .
Läs mer :
motion .
Idrottstjänsterfinska _ svenska _ engelska
Motionsplatserfinska _ svenska
gym för äldrefinska
Karlebynejdens institutfinska _ svenska
att röra sig i naturen
att röra sig i naturen är en traditionell och populär form av avkoppling för finländarna under alla årstider .
i Finland kan man med stöd av allemansrätten plocka bär och svamp i skogen och röra sig till fots , med cykel eller skidor vintertid .
det är inte tillåtet att beträda folks gårdar utan lov .
för fiske krävs fiskelov , med undantag för mete och pilkning .
även jakt fordrar jakttillstånd .
allemansrätten ger inte rätt att skräpa ner i naturen , skada träd eller växter , störa eller skada fågelbon eller fågelungar , köra motorfordon utan markägarens tillstånd eller bygga ens tillfälliga byggen .
mer information om motionsrutterna , rastplatser , möjligheter till fiske och båtliv samt exempelvis fågeltorn i Karleby finns på stadens webbplats .
rutterna för camping , paddling , vandring , cykling och övriga rutter i Karleby finns i karttjänsten på nätet .
i karttjänsten visas även var största delen av motionsplatserna finns .
du kan köpa friluftskartor över Karleby hos Karleby Turism : Salutorget 5 , 67100 Karleby .
Läs mer : att röra sig i naturen .
linkkiMiljöförvaltningen :
Allemansrättenfinska _ svenska _ engelska _ ryska
Motionskarta över Karlebyfinska _ svenska
motionsrutter i Karlebyfinska _ svenska
teater och film
Karleby är en teaterstad med långa anor , som erbjuder scenkonst på hög nivå framförd av både proffs och amatörer .
Karleby stadsteater finns i det stämningsfulla Vartiolinna ( Torggatan 48 ) .
du kan läsa mer om amatörteatrarnas verksamhet på deras webbplats och i evenemangskalendern .
i Karleby finns biografen Bio Rex , vars två salar använder digital- och 3D @-@ teknik .
Bio Rex program finns under länken här intill .
Läs mer : teater och film .
Stadsteaternfinska
Biograffinska
teater och danskonst i Karlebyfinska _ svenska _ engelska
Evenemangskalenderfinska
museer
i hjärtat av staden , i det anrika Rooska gården , finns K.H.Renlunds museum .
Karleby stad grundade museet 1909 utgående från en testamentsgåva av affärsmannen Karl Herman Renlund ( 1850 @-@ 1908 ) .
på museet finns Renlunds samling av finländsk konst från guldåldern och tillfälliga utställningar i en kulturhistorisk miljö .
även i museikvarterens övriga byggnader finns utställningar om stadens kulturhistoria och utställningar med ITE @-@ konst .
på K.H.Renlunds museums webbplats finns mer information om museets tjänster , utställningar samt aktuell verksamhet .
Utöver K.H.Renlunds museum lönar det sig att besöka det naturhistoriska museet Kieppi ( Kieppi är stängt tills vidare på grund av brand ) samt de många hembygdsmuseerna och övriga de historiska resmålen i regionen .
exempelvis i Konst @-@ Vionoja @-@ centret presenteras konstnären Veikko Vionojas verk .
i Kelviå , ca 10 km norrut från Karleby , finns Toivonen djurpark och drängmuseum .
mer information om dessa museer finns under länkarna här intill .
Läs mer : museer .
museer och traditionsarbetefinska _ svenska _ engelska
K.H. Renlunds museum - Mellersta Österbottens landskapsmuseumfinska _ svenska _ engelska
Kieppi , Karleby naturvetenskapliga museumfinska _ svenska _ engelska
linkkiToivonens djurpark och drängmuseum :
Toivonens djurpark och drängmuseum finska _ svenska _ engelska
konst Vionojafinska
hobbyer för barn och unga
flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet .
flera olika föreningar samt kommunala institut ger unga möjlighet att studera idrott och kultur samt bl.a. språk och hantverk .
barn och unga kan delta i grundläggande undervisning i musik , dans , bildkonst och hantverk .
dessutom erbjuder stadens ungdomstjänster en rockskola .
stadens ungdomstjänster driver sju ungdomsgårdar runt om i Karleby .
de rusmedels- och rökfria ungdomslokalerna erbjuder handledd verksamhet för barn i årskurserna 3 @-@ 6 och unga i åldern 13 @-@ 17 år i olika delar av Karleby .
information om hobbyverksamheter för barn och unga finns på stadens webbplats .
rådgivningen vid Ungdomsgården Vinge ger aktuell information om bl.a. internationalisering , studier , arbetsliv , hälsa , hobbyverksamhet och boende .
Karlebynejdens institut erbjuder barn och unga olika former av hobbyverksamhet , exempelvis i konstämnen och musik .
kontrollera vilka kurser som är aktuella i institutets webbtjänst .
Karleby evangelisk @-@ lutherska församlingar erbjuder även hobbyverksamhet för barn och unga , såsom lekparksträffar , klubbar , musikverksamhet och läger .
mer information om verksamheten finns på Karleby församlingssammanslutnings webbplats .
ungdomsgården Vinge
67100 Karleby
Läs mer : hobbyer för barn och unga .
övrig undervisning i Karlebyfinska _ svenska
Ungdomstjänsterfinska _ svenska _ engelska
Karlebynejdens institutfinska _ svenska
linkkiKarleby kyrkliga samfällighet :
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
föreningar
Karleby har ett aktivt och mångsidigt föreningsliv för invånare i alla åldrar .
Läs mer : föreningar .
problem med uppehållstillstånd
brott
våld
diskriminering och rasism
behöver du en jurist ?
Död
problem i äktenskap eller parförhållande
skilsmässa
problem med den mentala hälsan
missbruksproblem
i en krissituation kan du ringa nödcentralen på numret 112 .
de slussar vid behov dig vidare till socialjouren .
du ska endast ringa nödcentralen i brådskande nödsituationer , där liv , egendom eller miljön är i fara .
problem med uppehållstillstånd
om du har problem eller oklarheter med ditt uppehållstillstånd kan du kontakta Migrationsverket .
Migrationsverket
Korsholmsesplanaden 45
Vasa
Läs mer : problem med uppehållstillstånd .
brott
om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112 .
ring inte nödnumret om det inte är fråga om en nödsituation .
du kan göra en polisanmälan på nätet .
mer information finns på Polisens webbplats .
du kan även skriva ut anmälningsblanketten på nätet och lämna in den till polisstationen .
Karleby polisstation
Karlebygatan 74
67100 Karleby
Läs mer : brott .
tidsbokningfinska _ svenska _ engelska
Polisamälanfinska _ svenska _ engelska
våld
om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112 .
Läs mer : våld .
diskriminering och rasism
om du misstänker att du blivit utsatt för diskriminering då du sökt arbete eller på arbetsplatsen ska du först ta upp detta på din arbetsplats .
om saken inte kan lösas på arbetsplatsen ska du kontakta arbetarskyddet vid Regionförvaltningsverket i Västra och Inre Finland .
Besöksadress :
Regionförvaltningsverket i Västra och Inre Finland
Wollfskavägen 35
65101 Vasa
telefon : 0295.018.450
om du utsätts för diskriminering kan du be om hjälp av Diskrimineringsombudsmannen .
om du fallit offer för ett rasistiskt motiverat brott kan du göra en polisanmälan på nätet eller polisstationen .
Läs mer : diskriminering och rasism .
linkkiRegionförvaltningsverket i Västra och Inre Finland :
Regionförvaltningsverket i Västra och Inre Finlandfinska _ svenska _ engelska
hjälp och information för personer som drabbats av etnisk diskrimineringfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
behöver du en jurist ?
juridiska tjänster är avgiftsbelagda men om du har små eller medelstora inkomster , kan du få helt eller delvis avgiftsfri rättshjälp från statens rättshjälpsbyrå .
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
Besöksadress : Ämbetshuset , Torggatan 40 , 67100 Karleby
telefon : 029.566.1270
information om enskilda jurister finns bland annat på Finlands Advokatförbunds webbplats .
Läs mer :
behöver du en jurist ?
linkkiFinlands advokatförbund :
Finlands advokatförbundfinska _ svenska _ engelska
Död
den evangelisk @-@ lutherska kyrkans församlingars begravningsplatser fungerar som allmänna begravningsplatser .
där kan även avlidna som inte är medlemmar i kyrkan begravas .
de är alltså avsedda för alla invånare i staden .
mer information finns på Karleby kyrkliga samfällighets webbplats .
om en närstående plötsligt dör kan du söka krishjälp vid din egen hälsostation , eller utanför tjänstetid vid samjouren för Mellersta Österbottens centralsjukhus .
de evangelisk @-@ lutherska församlingarna i Karlebynejden erbjuder även sorggrupper .
även församlingarnas diakonimottagningar erbjuder samtalshjälp för sorgearbetet .
Läs mer : Död .
linkkiKarleby kyrkliga samfällighet :
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Hälsostationernafinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
problem i äktenskap eller parförhållande
vid problem i äktenskap eller parförhållande får du hjälp av Mellersta Österbottens familjerådgivningscentral som underhålls av Karleby kyrkliga samfällighets och Mellersta Österbottens social- och hälsovårdssamkommun Soites familjerådgivning .
Familjerågivningscentralen
telefon : 050.3147.464 .
Karleby familjerådgivning
67100 Karleby
tel . 044.730.7640
Läs mer : problem i äktenskap eller parförhållande .
linkkiMellersta Österbottens Familjerådgivningscentral :
familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
familjerådgivningfinska _ svenska
skilsmässa
skilsmässa kan sökas av kvinnan , av mannen eller av båda makarna tillsammans .
man ansöker om skilsmässa i tingsrätten .
till att börja med görs en skriftlig skilsmässoansökan .
Österbottens tingsrätt Karleby kansli
Besöksadress : Karlebygatan 27 , 67100 Karleby
telefon : 029.56.49294
Läs mer : skilsmässa .
hälsovårdaren på barnrådgivningsbyrån ger råd i frågor som gäller små barns hälsa , tillväxt och utveckling .
barnrådgivningsbyrån ger information om platser som erbjuder hjälp vid behov .
vid problem hos unga i skolåldern hjälper exempelvis skolans hälsovårdare eller skolkuratorn .
Läs mer : barns och ungas problem .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Skolhälsovårdfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Barnrådgivningarfinska _ svenska
du kan ta upp problem med hälsovårdaren på skolan eller studieplatsen eller vuxna på ungdomsgården .
mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats .
föräldrar eller unga själva kan kontakta familjerådgivningen .
där kan man tala om problem och få hjälp och stöd .
mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats .
Familjerådgivningens telefonnummer : 044.730.7640 .
Läs mer : barns och ungas problem .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Studerandehälsovårdfinska _ svenska
ungdomsgårdar och -lokaler finska _ svenska
problem med den mentala hälsan
om du behöver hjälp och stöd för din mentala hälsa kan du boka en läkartid vid hälsostationen .
läkaren bedömer situationen .
vid behov skriver läkaren en remiss till psykiatrisk specialsjukvård .
Läs mer : mental hälsa .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Mentalvårdstjänsterfinska _ svenska
om du har ekonomiska problem kan du be om råd hos Mellersta Österbottens social- och hälsovårdssamkommun Soites enheter för socialarbete eller utkomststöd , tfn 040.806.5095 eller tjänstestyrningen , tfn 040.806.5093 .
om du har problem med skulder , kontakta rättshjälpsbyrån .
du kan anlita vilken som helst rättshjälpsbyrå oberoende av din hemkommun .
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
telefon : 029.566.1270
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Servicehandledningfinska _ svenska
missbruksproblem
om du har problem med alkohol , droger , läkemedel eller hasardspel kan du få vård och rehabilitering vid Porten , Mellersta Österbottens social- och hälsovårdssamkommun Soites center för missbruksproblem .
du kan ta upp problemet med proffs inom hälsovården eller företagshälsovården , som kan slussa dig vidare i vårdsystemet , eller direkt kontakta Soites missbrukstjänster , tfn 040.8068.101 .
för tillnyktrings- och avgiftningsvård debiteras en patientavgift liksom även för korttidsrehabilitering , öppen rehabilitering är gratis .
även Karleby evangelisk @-@ lutherska församlingssammanslutnings specialdiakoner erbjuder samtalshjälp vid missbruksproblem .
kontaktuppgifter
Hälsovägen 4
67200 Karleby
telefon : 040.806.8101
Läs mer : missbruksproblem .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Service för missbrukarefinska _ svenska
linkkiKarleby evangelisk @-@ lutherska församlingssammansutning :
Karleby evangelisk @-@ lutherska församlings arbete bland missbrukarefinska _ svenska
problem med uppehållstillstånd
brott
våld
diskriminering och rasism
behöver du en jurist ?
Död
problem i äktenskap eller parförhållande
skilsmässa
problem med den mentala hälsan
missbruksproblem
i en krissituation kan du ringa nödcentralen på numret 112 .
de slussar vid behov dig vidare till socialjouren .
du ska endast ringa nödcentralen i brådskande nödsituationer , där liv , egendom eller miljön är i fara .
problem med uppehållstillstånd
om du har problem eller oklarheter med ditt uppehållstillstånd kan du kontakta Migrationsverket .
Migrationsverket
Korsholmsesplanaden 45
Vasa
Läs mer : problem med uppehållstillstånd .
brott
om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112 .
ring inte nödnumret om det inte är fråga om en nödsituation .
du kan göra en polisanmälan på nätet .
mer information finns på Polisens webbplats .
du kan även skriva ut anmälningsblanketten på nätet och lämna in den till polisstationen .
Karleby polisstation
Karlebygatan 74
67100 Karleby
Läs mer : brott .
tidsbokningfinska _ svenska _ engelska
Polisamälanfinska _ svenska _ engelska
våld
om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112 .
Läs mer : våld .
diskriminering och rasism
om du misstänker att du blivit utsatt för diskriminering då du sökt arbete eller på arbetsplatsen ska du först ta upp detta på din arbetsplats .
om saken inte kan lösas på arbetsplatsen ska du kontakta arbetarskyddet vid Regionförvaltningsverket i Västra och Inre Finland .
Besöksadress :
Regionförvaltningsverket i Västra och Inre Finland
Wollfskavägen 35
65101 Vasa
telefon : 0295.018.450
om du utsätts för diskriminering kan du be om hjälp av Diskrimineringsombudsmannen .
om du fallit offer för ett rasistiskt motiverat brott kan du göra en polisanmälan på nätet eller polisstationen .
Läs mer : diskriminering och rasism .
linkkiRegionförvaltningsverket i Västra och Inre Finland :
Regionförvaltningsverket i Västra och Inre Finlandfinska _ svenska _ engelska
hjälp och information för personer som drabbats av etnisk diskrimineringfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
behöver du en jurist ?
juridiska tjänster är avgiftsbelagda men om du har små eller medelstora inkomster , kan du få helt eller delvis avgiftsfri rättshjälp från statens rättshjälpsbyrå .
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
Besöksadress : Ämbetshuset , Torggatan 40 , 67100 Karleby
telefon : 029.566.1270
information om enskilda jurister finns bland annat på Finlands Advokatförbunds webbplats .
Läs mer :
behöver du en jurist ?
linkkiFinlands advokatförbund :
Finlands advokatförbundfinska _ svenska _ engelska
Död
den evangelisk @-@ lutherska kyrkans församlingars begravningsplatser fungerar som allmänna begravningsplatser .
där kan även avlidna som inte är medlemmar i kyrkan begravas .
de är alltså avsedda för alla invånare i staden .
mer information finns på Karleby kyrkliga samfällighets webbplats .
om en närstående plötsligt dör kan du söka krishjälp vid din egen hälsostation , eller utanför tjänstetid vid samjouren för Mellersta Österbottens centralsjukhus .
de evangelisk @-@ lutherska församlingarna i Karlebynejden erbjuder även sorggrupper .
även församlingarnas diakonimottagningar erbjuder samtalshjälp för sorgearbetet .
Läs mer : Död .
linkkiKarleby kyrkliga samfällighet :
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Hälsostationernafinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
problem i äktenskap eller parförhållande
vid problem i äktenskap eller parförhållande får du hjälp av Mellersta Österbottens familjerådgivningscentral som underhålls av Karleby kyrkliga samfällighets och Mellersta Österbottens social- och hälsovårdssamkommun Soites familjerådgivning .
Familjerågivningscentralen
telefon : 050.3147.464 .
Karleby familjerådgivning
67100 Karleby
tel . 044.730.7640
Läs mer : problem i äktenskap eller parförhållande .
linkkiMellersta Österbottens Familjerådgivningscentral :
familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
familjerådgivningfinska _ svenska
skilsmässa
skilsmässa kan sökas av kvinnan , av mannen eller av båda makarna tillsammans .
man ansöker om skilsmässa i tingsrätten .
till att börja med görs en skriftlig skilsmässoansökan .
Österbottens tingsrätt Karleby kansli
Besöksadress : Karlebygatan 27 , 67100 Karleby
telefon : 029.56.49294
Läs mer : skilsmässa .
hälsovårdaren på barnrådgivningsbyrån ger råd i frågor som gäller små barns hälsa , tillväxt och utveckling .
barnrådgivningsbyrån ger information om platser som erbjuder hjälp vid behov .
vid problem hos unga i skolåldern hjälper exempelvis skolans hälsovårdare eller skolkuratorn .
Läs mer : barns och ungas problem .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Skolhälsovårdfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Barnrådgivningarfinska _ svenska
du kan ta upp problem med hälsovårdaren på skolan eller studieplatsen eller vuxna på ungdomsgården .
mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats .
föräldrar eller unga själva kan kontakta familjerådgivningen .
där kan man tala om problem och få hjälp och stöd .
mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats .
Familjerådgivningens telefonnummer : 044.730.7640 .
Läs mer : barns och ungas problem .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Studerandehälsovårdfinska _ svenska
ungdomsgårdar och -lokaler finska _ svenska
problem med den mentala hälsan
om du behöver hjälp och stöd för din mentala hälsa kan du boka en läkartid vid hälsostationen .
läkaren bedömer situationen .
vid behov skriver läkaren en remiss till psykiatrisk specialsjukvård .
Läs mer : mental hälsa .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Mentalvårdstjänsterfinska _ svenska
om du har ekonomiska problem kan du be om råd hos Mellersta Österbottens social- och hälsovårdssamkommun Soites enheter för socialarbete eller utkomststöd , tfn 040.806.5095 eller tjänstestyrningen , tfn 040.806.5093 .
om du har problem med skulder , kontakta rättshjälpsbyrån .
du kan anlita vilken som helst rättshjälpsbyrå oberoende av din hemkommun .
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
telefon : 029.566.1270
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Servicehandledningfinska _ svenska
missbruksproblem
om du har problem med alkohol , droger , läkemedel eller hasardspel kan du få vård och rehabilitering vid Porten , Mellersta Österbottens social- och hälsovårdssamkommun Soites center för missbruksproblem .
du kan ta upp problemet med proffs inom hälsovården eller företagshälsovården , som kan slussa dig vidare i vårdsystemet , eller direkt kontakta Soites missbrukstjänster , tfn 040.8068.101 .
för tillnyktrings- och avgiftningsvård debiteras en patientavgift liksom även för korttidsrehabilitering , öppen rehabilitering är gratis .
även Karleby evangelisk @-@ lutherska församlingssammanslutnings specialdiakoner erbjuder samtalshjälp vid missbruksproblem .
kontaktuppgifter
Hälsovägen 4
67200 Karleby
telefon : 040.806.8101
Läs mer : missbruksproblem .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Service för missbrukarefinska _ svenska
linkkiKarleby evangelisk @-@ lutherska församlingssammansutning :
Karleby evangelisk @-@ lutherska församlings arbete bland missbrukarefinska _ svenska
problem med uppehållstillstånd
brott
våld
diskriminering och rasism
behöver du en jurist ?
Död
problem i äktenskap eller parförhållande
skilsmässa
problem med den mentala hälsan
missbruksproblem
i en krissituation kan du ringa nödcentralen på numret 112 .
de slussar vid behov dig vidare till socialjouren .
du ska endast ringa nödcentralen i brådskande nödsituationer , där liv , egendom eller miljön är i fara .
problem med uppehållstillstånd
om du har problem eller oklarheter med ditt uppehållstillstånd kan du kontakta Migrationsverket .
Migrationsverket
Korsholmsesplanaden 45
Vasa
Läs mer : problem med uppehållstillstånd .
brott
om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112 .
ring inte nödnumret om det inte är fråga om en nödsituation .
du kan göra en polisanmälan på nätet .
mer information finns på Polisens webbplats .
du kan även skriva ut anmälningsblanketten på nätet och lämna in den till polisstationen .
Karleby polisstation
Karlebygatan 74
67100 Karleby
Läs mer : brott .
tidsbokningfinska _ svenska _ engelska
Polisamälanfinska _ svenska _ engelska
våld
om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112 .
Läs mer : våld .
diskriminering och rasism
om du misstänker att du blivit utsatt för diskriminering då du sökt arbete eller på arbetsplatsen ska du först ta upp detta på din arbetsplats .
om saken inte kan lösas på arbetsplatsen ska du kontakta arbetarskyddet vid Regionförvaltningsverket i Västra och Inre Finland .
Besöksadress :
Regionförvaltningsverket i Västra och Inre Finland
Wollfskavägen 35
65101 Vasa
telefon : 0295.018.450
om du utsätts för diskriminering kan du be om hjälp av Diskrimineringsombudsmannen .
om du fallit offer för ett rasistiskt motiverat brott kan du göra en polisanmälan på nätet eller polisstationen .
Läs mer : diskriminering och rasism .
linkkiRegionförvaltningsverket i Västra och Inre Finland :
Regionförvaltningsverket i Västra och Inre Finlandfinska _ svenska _ engelska
hjälp och information för personer som drabbats av etnisk diskrimineringfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
behöver du en jurist ?
juridiska tjänster är avgiftsbelagda men om du har små eller medelstora inkomster , kan du få helt eller delvis avgiftsfri rättshjälp från statens rättshjälpsbyrå .
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
Besöksadress : Ämbetshuset , Torggatan 40 , 67100 Karleby
telefon : 029.566.1270
information om enskilda jurister finns bland annat på Finlands Advokatförbunds webbplats .
Läs mer :
behöver du en jurist ?
linkkiFinlands advokatförbund :
Finlands advokatförbundfinska _ svenska _ engelska
Död
den evangelisk @-@ lutherska kyrkans församlingars begravningsplatser fungerar som allmänna begravningsplatser .
där kan även avlidna som inte är medlemmar i kyrkan begravas .
de är alltså avsedda för alla invånare i staden .
mer information finns på Karleby kyrkliga samfällighets webbplats .
om en närstående plötsligt dör kan du söka krishjälp vid din egen hälsostation , eller utanför tjänstetid vid samjouren för Mellersta Österbottens centralsjukhus .
de evangelisk @-@ lutherska församlingarna i Karlebynejden erbjuder även sorggrupper .
även församlingarnas diakonimottagningar erbjuder samtalshjälp för sorgearbetet .
Läs mer : Död .
linkkiKarleby kyrkliga samfällighet :
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Hälsostationernafinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
problem i äktenskap eller parförhållande
vid problem i äktenskap eller parförhållande får du hjälp av Mellersta Österbottens familjerådgivningscentral som underhålls av Karleby kyrkliga samfällighets och Mellersta Österbottens social- och hälsovårdssamkommun Soites familjerådgivning .
Familjerågivningscentralen
telefon : 050.3147.464 .
Karleby familjerådgivning
67100 Karleby
tel . 044.730.7640
Läs mer : problem i äktenskap eller parförhållande .
linkkiMellersta Österbottens Familjerådgivningscentral :
familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
familjerådgivningfinska _ svenska
skilsmässa
skilsmässa kan sökas av kvinnan , av mannen eller av båda makarna tillsammans .
man ansöker om skilsmässa i tingsrätten .
till att börja med görs en skriftlig skilsmässoansökan .
Österbottens tingsrätt Karleby kansli
Besöksadress : Karlebygatan 27 , 67100 Karleby
telefon : 029.56.49294
Läs mer : skilsmässa .
hälsovårdaren på barnrådgivningsbyrån ger råd i frågor som gäller små barns hälsa , tillväxt och utveckling .
barnrådgivningsbyrån ger information om platser som erbjuder hjälp vid behov .
vid problem hos unga i skolåldern hjälper exempelvis skolans hälsovårdare eller skolkuratorn .
Läs mer : barns och ungas problem .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Skolhälsovårdfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Barnrådgivningarfinska _ svenska
du kan ta upp problem med hälsovårdaren på skolan eller studieplatsen eller vuxna på ungdomsgården .
mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats .
föräldrar eller unga själva kan kontakta familjerådgivningen .
där kan man tala om problem och få hjälp och stöd .
mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats .
Familjerådgivningens telefonnummer : 044.730.7640 .
Läs mer : barns och ungas problem .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Studerandehälsovårdfinska _ svenska
ungdomsgårdar och -lokaler finska _ svenska
problem med den mentala hälsan
om du behöver hjälp och stöd för din mentala hälsa kan du boka en läkartid vid hälsostationen .
läkaren bedömer situationen .
vid behov skriver läkaren en remiss till psykiatrisk specialsjukvård .
Läs mer : mental hälsa .
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Mentalvårdstjänsterfinska _ svenska
om du har ekonomiska problem kan du be om råd hos Mellersta Österbottens social- och hälsovårdssamkommun Soites enheter för socialarbete eller utkomststöd , tfn 040.806.5095 eller tjänstestyrningen , tfn 040.806.5093 .
om du har problem med skulder , kontakta rättshjälpsbyrån .
du kan anlita vilken som helst rättshjälpsbyrå oberoende av din hemkommun .
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
telefon : 029.566.1270
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite :
Servicehandledningfinska _ svenska
missbruksproblem
om du har problem med alkohol , droger , läkemedel eller hasardspel kan du få vård och rehabilitering vid Porten , Mellersta Österbottens social- och hälsovårdssamkommun Soites center för missbruksproblem .
du kan ta upp problemet med proffs inom hälsovården eller företagshälsovården , som kan slussa dig vidare i vårdsystemet , eller direkt kontakta Soites missbrukstjänster , tfn 040.8068.101 .
för tillnyktrings- och avgiftningsvård debiteras en patientavgift liksom även för korttidsrehabilitering , öppen rehabilitering är gratis .
även Karleby evangelisk @-@ lutherska församlingssammanslutnings specialdiakoner erbjuder samtalshjälp vid missbruksproblem .
kontaktuppgifter
