����      ]�(�numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i4�����R�(K�<�NNNJ����J����K t�b�C,a  E   h   �   �   g                  �t�bhhK ��h��R�(KK��h�C4   �            
   �  �   �              �t�bhhK ��h��R�(KK��h�C8      �  �	     0            A   �	  �        �t�bhhK ��h��R�(KK��h�C0d  -   
            �                 �t�bhhK ��h��R�(KK��h�C�   T     �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C<�                    �     O                 �t�bhhK ��h��R�(KK��h�C   ?     �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   6   1     	        �t�bhhK ��h��R�(KK��h�CH      �      �        &      �                 l        �t�bhhK ��h��R�(KK��h�Cd      0  �   �  m     �   x      �      $     �     �   �      �      -           �t�bhhK ��h��R�(KK
��h�C(   �        2     �     D      �t�bhhK ��h��R�(KK��h�C,     �t�bhhK ��h��R�(KK��h�C
     �t�bhhK ��h��R�(KK��h�C,�     E      n     �     �        �t�bhhK ��h��R�(KK
��h�C(      4               v        �t�bhhK ��h��R�(KK��h�C4	   �  	   �	  	   �  	   �  	   �  	   �     �t�bhhK ��h��R�(KK��h�C<[     �     '      I   ?                       �t�bhhK ��h��R�(KK��h�C8�     �         �   ]  9   %   #             �t�bhhK ��h��R�(KK��h�CP�         I   l      ~            �              D              �t�bhhK ��h��R�(KK��h�Cd         .        �                       �                     8   S        �t�bhhK ��h��R�(KK��h�C@   �     .      �  9   �  7   �  �     .  �        �t�bhhK ��h��R�(KK��h�C8           D         z  �  �  �   �        �t�bhhK ��h��R�(KK��h�C   y     �t�bhhK ��h��R�(KK	��h�C$      �     �  
            �t�bhhK ��h��R�(KK	��h�C$�      '	     �  h           �t�bhhK ��h��R�(KK��h�C   �  	         �t�bhhK ��h��R�(KK��h�C8         �   ~        L      x              �t�bhhK ��h��R�(KK��h�CX*      �  )        H   �        S   &      F  �     �  +              �t�bhhK ��h��R�(KK��h�Ct      �              (      *  �      4   :   H     �        >      e  �                   �t�bhhK ��h��R�(KK��h�CP   E      4      m  &      �  I        $   �   �        r	        �t�bhhK ��h��R�(KK��h�CH   .   
   @   �   F   '                                   �t�bhhK ��h��R�(KK��h�C`   $   n      �	     .      H          �          f   �     %   I  �        �t�bhhK ��h��R�(KK��h�C4*   �   (        �     �       �        �t�bhhK ��h��R�(KK��h�C   9  �     �t�bhhK ��h��R�(KK
��h�C(   ?   �  
            F         �t�bhhK ��h��R�(KK ��h�C�m     �      �      �     �        t        �   l        ?   !   �     �   �   |  
   �   �             �t�bhhK ��h��R�(KK��h�Ch   (   <      +	  "   �           �     	                                        �t�bhhK ��h��R�(KK��h�C4      �   X     U   e   �   T              �t�bhhK ��h��R�(KK��h�CH.     &     B         �  �     �  �     C      �        �t�bhhK ��h��R�(KK��h�C@   X   '   q                s                     �t�bhhK ��h��R�(KK��h�C      |        �t�bhhK ��h��R�(KK��h�C4      N         D     *        �         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C[            �t�bhhK ��h��R�(KK��h�C<            7     F     �  �     �   �          �t�bhhK ��h��R�(KK��h�CL   `   �      �   �  �  
      6  c   &      =      �  4         �t�bhhK ��h��R�(KK	��h�C$!      �  
         	         �t�bhhK ��h��R�(KK��h�C          	      	         �t�bhhK ��h��R�(KK��h�C             �t�bhhK ��h��R�(KK��h�Ch*   $                  o  p           P      3     (     �  
   p                 �t�bhhK ��h��R�(KK��h�C8N  �      �     y      l  
      �  �         �t�bhhK ��h��R�(KK��h�CH   %                    [        D	     �     �        �t�bhhK ��h��R�(KK	��h�C$�   �  +      $        �      �t�bhhK ��h��R�(KK��h�C!         	         �t�bhhK ��h��R�(KK	��h�C$�  	              �         �t�bhhK ��h��R�(KK��h�CH#   !            �  ?      
   3   6   �
        1  r         �t�bhhK ��h��R�(KK��h�C8   	   �   	   I  	   U  	   /  	   s  	   �     �t�bhhK ��h��R�(KK��h�CL*      �      �  �  |      �                  #     +         �t�bhhK ��h��R�(KK��h�C@z  �  �               �   y   %   �  �               �t�bhhK ��h��R�(KK��h�C               �t�bhhK ��h��R�(KK��h�CH            ,         ,            -   d     �   &        �t�bhhK ��h��R�(KK��h�C4      P   B   j              �           �t�bhhK ��h��R�(KK��h�C4   r    �     U  �   A   �     |        �t�bhhK ��h��R�(KK!��h�C�   $   A                   $   ,   �        �   �         �  N      �        0         �     �           �t�bhhK ��h��R�(KK��h�C�      �     �t�bhhK ��h��R�(KK��h�CH         �      �	     �   �   8	  
   B        B           �t�bhhK ��h��R�(KK��h�C09   ,     0     �      r  j            �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�C   9     �t�bhhK ��h��R�(KK��h�C\�  {  *   D         �  �        �   �                 7   �  �  w        �t�bhhK ��h��R�(KK��h�CP�   >      �  �     C   w      �      >   %   �        �   �         �t�bhhK ��h��R�(KK��h�Ch      J                   +     +      &      �     �                         �t�bhhK ��h��R�(KK��h�C,�        }        	      	   U     �t�bhhK ��h��R�(KK��h�C       g  )               �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C@         o  �  Y          �  ;         �        �t�bhhK ��h��R�(KK��h�Ct            �  �     
   �        I   b        g      2            �     )     9  b        �t�bhhK ��h��R�(KK��h�C|      �	  (        +     :            +   �   0     �   s   7         �  �  3  T      �	     B        �t�bhhK ��h��R�(KK��h�C0]         �      R  *      d          �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C %   �           �         �t�bhhK ��h��R�(KK	��h�C$     �      2   0   �  r      �t�bhhK ��h��R�(KK��h�CB  ]      $   �         �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK	��h�C$�              0   <         �t�bhhK ��h��R�(KK��h�C4,   O            �     �         �         �t�bhhK ��h��R�(KK	��h�C$   .      (      o  �        �t�bhhK ��h��R�(KK��h�CD   &   -   a                        $   G              �t�bhhK ��h��R�(KK��h�CHV  $  �  �              %         �   �     9            �t�bhhK ��h��R�(KK��h�CHq   �                    �  0  �     �    �           �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C,�     ^    
      "      y        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�C [           a  	         �t�bhhK ��h��R�(KK��h�C�  Z     �t�bhhK ��h��R�(KK��h�C0�     �     �       x  d   S        �t�bhhK ��h��R�(KK��h�C       -   i  �  �        �t�bhhK ��h��R�(KK��h�C4   >   a         �       *               �t�bhhK ��h��R�(KK��h�Cb   #   
   $   N        �t�bhhK ��h��R�(KK��h�C`      G           #   i   #  �      &         w  v     
   $                 �t�bhhK ��h��R�(KK��h�CL*      �      �  C  �      (     	           #     +         �t�bhhK ��h��R�(KK��h�CP      D  =         +  G   4     >      a   4      �      7         �t�bhhK ��h��R�(KK��h�Cd!      �      �           "              '      .   
   �        F   
   ,         �t�bhhK ��h��R�(KK��h�C  p   �       �t�bhhK ��h��R�(KK��h�C         
   �         �t�bhhK ��h��R�(KK��h�Cl   V   �   +      �           (   <         �                    �           ;        �t�bhhK ��h��R�(KK��h�CPB              �     2      �           2   J   �     o         �t�bhhK ��h��R�(KK��h�C08     A     �  
   %  .	     �        �t�bhhK ��h��R�(KK��h�CZ            �t�bhhK ��h��R�(KK��h�CL   &   M      �         "  g              �  h              �t�bhhK ��h��R�(KK��h�Cl        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�CT      �        �  �     h   t        M   �      �                 �t�bhhK ��h��R�(KK��h�CX�                  ;        2   l  g      �     �   �        "        �t�bhhK ��h��R�(KK��h�C,1   S        �  :         D        �t�bhhK ��h��R�(KK��h�CT      �  R  4         D  l           �      �   ;      o           �t�bhhK ��h��R�(KK��h�C    �  �   �       �      �t�bhhK ��h��R�(KK��h�C`�        �  F         �  !      l      �     4              �  ~   ]        �t�bhhK ��h��R�(KK��h�C !      %   ^     	         �t�bhhK ��h��R�(KK��h�C0#   !      �  (      
   3   6            �t�bhhK ��h��R�(KK��h�Cl�      (     |      �      |      s	     �   +        �     !      u  �      �  �        �t�bhhK ��h��R�(KK��h�CP	  l      ;      #     I	  �        .   z      �      �          �t�bhhK ��h��R�(KK��h�CD      0   B  v  �  A              .   {      �         �t�bhhK ��h��R�(KK��h�C<            �   *      �               z          �t�bhhK ��h��R�(KK
��h�C(Z     L     �  	      	         �t�bhhK ��h��R�(KK��h�C8         �         �   �         U            �t�bhhK ��h��R�(KK ��h�C�         �           �     J      ,   K     x     `      &      M   �      �                          �t�bhhK ��h��R�(KK��h�C8�      (  ]       R     B   �     o         �t�bhhK ��h��R�(KK��h�C   :               �t�bhhK ��h��R�(KK	��h�C$      �                     �t�bhhK ��h��R�(KK��h�CX      J   �  +   �  �  
      �                 �   #        �        �t�bhhK ��h��R�(KK��h�C�
        �t�bhhK ��h��R�(KK��h�C8        $   �     s        
      F         �t�bhhK ��h��R�(KK	��h�C$      )   =      �   w         �t�bhhK ��h��R�(KK��h�C@M   -   �      3   �     [      �     �      D         �t�bhhK ��h��R�(KK��h�C@      '   m      �      D   w        �   	  V        �t�bhhK ��h��R�(KK��h�C4
   �   F   '   �  1     #   !      P        �t�bhhK ��h��R�(KK��h�Ce   �
     �t�bhhK ��h��R�(KK��h�C\                  j   �  \  @         �  �     �  �      �             �t�bhhK ��h��R�(KK��h�Ce   �   �
     �t�bhhK ��h��R�(KK��h�Ct   �     �  	      	      	   K   	   �   	   �   	     	   U  	   �   	   �  	   /  	   �  	        �t�bhhK ��h��R�(KK��h�CD|  $  I   /      ~           C  �     d             �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�C 1   #       �      �        �t�bhhK ��h��R�(KK��h�CX   5  _  D   �     �   f     _  C      ,   �              �  �        �t�bhhK ��h��R�(KK��h�C       �         �        �t�bhhK ��h��R�(KK!��h�C�                        �   S   Q   h   Q     >      F  $   �                 y      �      4      �         �t�bhhK ��h��R�(KK��h�C4�        �       �      �     9        �t�bhhK ��h��R�(KK��h�C4/   9     7   &   �   a      �      �        �t�bhhK ��h��R�(KK	��h�C$   �    
         >        �t�bhhK ��h��R�(KK��h�C ]      �                 �t�bhhK ��h��R�(KK��h�Ct   $   �  �   �     4         
   _      X  �     �           0   4         
   _      �        �t�bhhK ��h��R�(KK��h�C,6     �  
   �   y      �           �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C`     �	     �        �t�bhhK ��h��R�(KK��h�C@]   P     �  �  �
     d   �  )      �   ~   �         �t�bhhK ��h��R�(KK��h�C   �           �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C4   �  &                 �
     �         �t�bhhK ��h��R�(KK��h�C<%      �     �           �   �                  �t�bhhK ��h��R�(KK��h�C       w   D  l     �      �t�bhhK ��h��R�(KK	��h�C$   '   
         
           �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C1   #            �t�bhhK ��h��R�(KK ��h�C�                 �     �        V  �	     
   _                  U   @     �     �  �  �           �t�bhhK ��h��R�(KK
��h�C(      )   �         "   W         �t�bhhK ��h��R�(KK��h�C\      \     �   �  )               ;        R   h      �        �        �t�bhhK ��h��R�(KK��h�Cv     H
  
   7     �t�bhhK ��h��R�(KK��h�C.     �        �t�bhhK ��h��R�(KK��h�Cl         �         P      +        ;  �     �            �     0  "  i   A   *        �t�bhhK ��h��R�(KK,��h�C�         Y      O                     �   G      t  &      =      n     �     Y      O   
   _      �     �   �        
   �     �     �        �t�bhhK ��h��R�(KK��h�CX   �           .   �     	        �     �     %   �  !  j   <         �t�bhhK ��h��R�(KK��h�C8�  /      2     `  �      �   K              �t�bhhK ��h��R�(KK��h�C<      U      �  �      b      %      u  �         �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C`?     |     N   L  �     d     �      �
        ]  �     �     �  �        �t�bhhK ��h��R�(KK��h�C�       9     �t�bhhK ��h��R�(KK��h�C,�      L   "   �  �  
   �  F         �t�bhhK ��h��R�(KK��h�CH�     �   
      $                   .      �   D        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�CH   ?   #   !               
   3   6   �     �	              �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�CD#   !      ]   ?      
   3   6      �   4  o  4   r         �t�bhhK ��h��R�(KK��h�C0e                     q   .           �t�bhhK ��h��R�(KK��h�C06  �    
   �  �           @         �t�bhhK ��h��R�(KK��h�CH      �  d                                �  �	        �t�bhhK ��h��R�(KK��h�CX        �  q	                 �  m     �         �   �     �        �t�bhhK ��h��R�(KK��h�C,H   �  �   �  
         f           �t�bhhK ��h��R�(KK	��h�C$   >   T   v                  �t�bhhK ��h��R�(KK��h�C4   .      �   ^     �  �     4           �t�bhhK ��h��R�(KK��h�C,�         �   A         �        �t�bhhK ��h��R�(KK��h�C�   �           �      �t�bhhK ��h��R�(KK
��h�C("   >  �  �     �              �t�bhhK ��h��R�(KK
��h�C(n     !  
      	      	         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK"��h�C�#   !      4      �            Z     v        0   4   (      
   3   6   7  z            
   �     �     F         �t�bhhK ��h��R�(KK��h�C@/      p     z     "     �
     �  "              �t�bhhK ��h��R�(KK��h�C,      �            	      	         �t�bhhK ��h��R�(KK
��h�C(   ]   5      d   �  :   t         �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CD   (   #   !         =      �  4   
   3   6   �  4         �t�bhhK ��h��R�(KK
��h�C(!          �   �              �t�bhhK ��h��R�(KK
��h�C(A   O  �           �  �        �t�bhhK ��h��R�(KK��h�C<�      �         �  �  Q        	      	         �t�bhhK ��h��R�(KK��h�C�      P     �t�bhhK ��h��R�(KK��h�C4      J         g   �  P      �  �         �t�bhhK ��h��R�(KK	��h�C$   �   '   E     y  �        �t�bhhK ��h��R�(KK ��h�C��   |      �  �  8  �   �   V     l
           �      �     �  �   4        �      �     �  
   N        �t�bhhK ��h��R�(KK	��h�C$           j	  �  �        �t�bhhK ��h��R�(KK��h�C<      �	  f
  �        l            h            �t�bhhK ��h��R�(KK��h�C@         O      �   
  Q   5         4               �t�bhhK ��h��R�(KK��h�C\        +      �      �t�bhhK ��h��R�(KK	��h�C$         -   ^  �            �t�bhhK ��h��R�(KK
��h�C(1   #       �	     /      �         �t�bhhK ��h��R�(KK��h�C0#   !      �                         �t�bhhK ��h��R�(KK��h�C@   @   '      �  b
  B   j        .                  �t�bhhK ��h��R�(KK��h�C    ?   �  
              �t�bhhK ��h��R�(KK��h�C4�  <              "   \     
           �t�bhhK ��h��R�(KK
��h�C(             	      	         �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�CL   �  C      P      f   �  
   �  }         J  E      �        �t�bhhK ��h��R�(KK��h�Cd"   >  (      �      \      �         G   W      �     $   k         �      u         �t�bhhK ��h��R�(KK��h�Cb     �      �t�bhhK ��h��R�(KK��h�C@   �        �   	     �           K     C        �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C<   ?   �     �      .   
   q           F         �t�bhhK ��h��R�(KK��h�C,W  
         �  '      B            �t�bhhK ��h��R�(KK��h�C4      �  d   �     z   B   }      �         �t�bhhK ��h��R�(KK��h�C,,      A   }         �      	         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C+     �t�bhhK ��h��R�(KK��h�C,%   b           �  :   �     y     �t�bhhK ��h��R�(KK��h�CP      &   2   �   
   c  �        $  G   A      )   G   [          �t�bhhK ��h��R�(KK
��h�C(   P     F  2   �  -            �t�bhhK ��h��R�(KK
��h�C(   �        .      �   �          �t�bhhK ��h��R�(KK��h�CH      �   N   y     �  o     �        B   �   j            �t�bhhK ��h��R�(KK��h�C4%         �        �   n   
   A           �t�bhhK ��h��R�(KK	��h�C$�     �  �            �     �t�bhhK ��h��R�(KK
��h�C(H      �   �  :         M        �t�bhhK ��h��R�(KK��h�C@	     �     �  �      �t�bhhK ��h��R�(KK��h�C4�	        b            F     0	  u         �t�bhhK ��h��R�(KK��h�C4$   �           �     �      �   w         �t�bhhK ��h��R�(KK
��h�C(�     �   .  "   %   �  K        �t�bhhK ��h��R�(KK��h�C-   �  >   5  �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C�     z   ,            �t�bhhK ��h��R�(KK&��h�C�*      �   �         v     F  �        �     �        �      �   &   D  �   �     �   S           a   ;      [              �t�bhhK ��h��R�(KK��h�Ch   $   n      �	        .      H          �             f   �     %   I  �        �t�bhhK ��h��R�(KK��h�Cl4     5      4     
        Q         O           �            \   �     &   H        �t�bhhK ��h��R�(KK��h�C<     �     �  "         V                    �t�bhhK ��h��R�(KK��h�CD         �  �  :   \   �  `   b     W  �             �t�bhhK ��h��R�(KK��h�CT�  !      �      ,               ?      
   3   6   �        �         �t�bhhK ��h��R�(KK��h�C8#   !            ^
  ?      
   3   6   �	        �t�bhhK ��h��R�(KK	��h�C$            �     f        �t�bhhK ��h��R�(KK��h�CT*         �      $   �   �  �     .            �  �      l  �         �t�bhhK ��h��R�(KK��h�Cd         �         �  G     *  X    �   �     �   �   �  p      �     �         �t�bhhK ��h��R�(KK��h�CB   �     B   |        �t�bhhK ��h��R�(KK
��h�C(
   �        P      �          �t�bhhK ��h��R�(KK��h�C,t   C           0      k   "	        �t�bhhK ��h��R�(KK��h�CD               l     E  �   2   �     .     [        �t�bhhK ��h��R�(KK��h�C	  �  x     �t�bhhK ��h��R�(KK��h�C8D      ;      0   �      �   �   d     �         �t�bhhK ��h��R�(KK
��h�C(                             �t�bhhK ��h��R�(KK��h�Cl      '      7     8              �   &            
   �           �    
   �        �t�bhhK ��h��R�(KK��h�CZ   .     �t�bhhK ��h��R�(KK��h�C�  �   G   `     �t�bhhK ��h��R�(KK��h�C8      U   k  ^      �  �     �              �t�bhhK ��h��R�(KK��h�CX;     N           �         �     �   �  :   �        A   :            �t�bhhK ��h��R�(KK��h�C8�  �     W   v   c   �     �     �  b        �t�bhhK ��h��R�(KK��h�C\
   3   6         p   '   !      \      �      p   
   A   F     �              �t�bhhK ��h��R�(KK��h�C81   #   
   3   6        �      /      V        �t�bhhK ��h��R�(KK��h�C,   R     �      7  �     �        �t�bhhK ��h��R�(KK��h�CP                        �      V     v   :                 �t�bhhK ��h��R�(KK��h�C0w  l     E     P  &   �     {        �t�bhhK ��h��R�(KK
��h�C(!      1  '   
   X   �   F         �t�bhhK ��h��R�(KK��h�C             �           �t�bhhK ��h��R�(KK��h�CL_        �  �     �      �        h     %       �        �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK
��h�C(�        �     	      	         �t�bhhK ��h��R�(KK��h�CE         c  c     �t�bhhK ��h��R�(KK��h�C!            �t�bhhK ��h��R�(KK��h�CE       ,   I     �t�bhhK ��h��R�(KK��h�C<  �   �   B   R      	        .        
        �t�bhhK ��h��R�(KK��h�C0�  �     �        y  V      L        �t�bhhK ��h��R�(KK��h�C8      5   :  <         [         U           �t�bhhK ��h��R�(KK��h�C,�	        j         ?        �      �t�bhhK ��h��R�(KK��h�C4      �   ?        2     j  
            �t�bhhK ��h��R�(KK��h�Cp         $   8     �     B   _  z    �      .   9               �  _            4         �t�bhhK ��h��R�(KK��h�C4�     $   �        l                    �t�bhhK ��h��R�(KK��h�C   �              �t�bhhK ��h��R�(KK��h�C@      5   �           U   @   k     �  
           �t�bhhK ��h��R�(KK��h�C      R        �t�bhhK ��h��R�(KK��h�CL�     0     '   �     �                           g        �t�bhhK ��h��R�(KK��h�C4�     �     �  H   B   R      �           �t�bhhK ��h��R�(KK��h�C�   (   �   <   r      �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CT[      <      	  M  	      	      	   K   	     	   �  	   �   	   �     �t�bhhK ��h��R�(KK��h�C,�  >      	  %   R      %   5         �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�CX*   �      �       d   �      �     {     J     �  
   D
     A        �t�bhhK ��h��R�(KK��h�C      	           �t�bhhK ��h��R�(KK��h�C4   �                    w     �        �t�bhhK ��h��R�(KK��h�C8"   k    �           �    h  9   �        �t�bhhK ��h��R�(KK��h�CL   Q     |      �   '      �  V   2      +
  �   
   �   �         �t�bhhK ��h��R�(KK��h�C      '   -   �   �        �t�bhhK ��h��R�(KK��h�CD$   ;  \                P      
       E   (        �t�bhhK ��h��R�(KK��h�CX   @      M     �     e   (   /      u  `  �        �     h          �t�bhhK ��h��R�(KK��h�C�	  [   9        R     �t�bhhK ��h��R�(KK��h�CT   .   '      !      >     ,   �      @      �     M     �            �t�bhhK ��h��R�(KK��h�C�  �   G   �     �t�bhhK ��h��R�(KK��h�C0   e   '   �     
   B   �     4        �t�bhhK ��h��R�(KK��h�C�  �  
   w        �t�bhhK ��h��R�(KK��h�C \      2           r      �t�bhhK ��h��R�(KK��h�C,z  +      �     |      <  �        �t�bhhK ��h��R�(KK��h�CL      /   �   :     5     �      M   �           i           �t�bhhK ��h��R�(KK��h�C8H         j             �        �         �t�bhhK ��h��R�(KK��h�C8!      �  	      	   �   	   �  	   �   	   �     �t�bhhK ��h��R�(KK	��h�C$      �   �      ^   �        �t�bhhK ��h��R�(KK��h�C<      �      �  T               �   �  a        �t�bhhK ��h��R�(KK��h�C   �  B  �        �t�bhhK ��h��R�(KK��h�C_     �         �t�bhhK ��h��R�(KK��h�C�  �  
   �        �t�bhhK ��h��R�(KK��h�C4   ]      �            U   �     �        �t�bhhK ��h��R�(KK��h�CD�	     	  u      �           ,   	      	   K   	   �      �t�bhhK ��h��R�(KK��h�C4%   	              .            �
        �t�bhhK ��h��R�(KK��h�C4Q     F     �            k               �t�bhhK ��h��R�(KK��h�C                    �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�CD      ;     %   |     �        �  �   �     ,         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�CX      G  �   �        J   �  9      7      �   W   �   $   �     �        �t�bhhK ��h��R�(KK��h�C   z            �t�bhhK ��h��R�(KK��h�C8�     ;         �           �   $   "        �t�bhhK ��h��R�(KK��h�C0   �  �      �         �               �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C@K       :   �          �   �      �     9        �t�bhhK ��h��R�(KK��h�C<1     `	     d           �           �         �t�bhhK ��h��R�(KK��h�Cp      .   p                  �   �         �     $   L     �        c   �         :        �t�bhhK ��h��R�(KK��h�Ch      �  +           .         w      ]
  c                       �   �           �t�bhhK ��h��R�(KK��h�C4b   $   �      �  �  �   �        �         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK!��h�C�   $   �   �         +   �         �   x        8   4         )         G  �   
   _      �      �   s   7         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C�   �  �             �t�bhhK ��h��R�(KK��h�CX   �      /   9     7      �  �  &   �      �       �        �          �t�bhhK ��h��R�(KK��h�C        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK
��h�C(2           5   �     �        �t�bhhK ��h��R�(KK��h�C02     �           �     H  @         �t�bhhK ��h��R�(KK��h�C<E      )   �  �     �   T   �  �  
   �  �        �t�bhhK ��h��R�(KK��h�C8�      2   0   �   �  T   %   h  �     �        �t�bhhK ��h��R�(KK
��h�C(]   (      �  I  �     a	        �t�bhhK ��h��R�(KK��h�CX*      �      8     4               )           �  "	     q   i
        �t�bhhK ��h��R�(KK&��h�C�            4      m        $  {         ]  �         x  $   �     &      =         �  4      m        4   
   A   �        �t�bhhK ��h��R�(KK��h�CD      0   �  >      -              �   �               �t�bhhK ��h��R�(KK��h�CD   f   �         �     0   X	  )                       �t�bhhK ��h��R�(KK��h�C 1        	      	         �t�bhhK ��h��R�(KK1��h�C�      =      o  �   *         �    7           +           �  H   7                 8  �     ,            �  �     o        M     $   0     }           �t�bhhK ��h��R�(KK��h�C8                  
            :	  �        �t�bhhK ��h��R�(KK��h�C/      �t�bhhK ��h��R�(KK��h�C,     N  7               �   O      �t�bhhK ��h��R�(KK��h�C�         	     �t�bhhK ��h��R�(KK
��h�C(f	           Y    
   �         �t�bhhK ��h��R�(KK��h�C	  	         �t�bhhK ��h��R�(KK��h�CH      '   H         h  !      �              ]  \        �t�bhhK ��h��R�(KK��h�C4�     {     �     %   t	                 �t�bhhK ��h��R�(KK��h�C@v  �	        .   %      �     K     �     �        �t�bhhK ��h��R�(KK��h�C -   �  �        _         �t�bhhK ��h��R�(KK��h�C�	     �t�bhhK ��h��R�(KK��h�C<�    �      f   �        �      ,               �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CX           /      $   8     T      �  
     �   9   s   �  L            �t�bhhK ��h��R�(KK��h�CL      '   �     �   
      �  d  �   c            �  �         �t�bhhK ��h��R�(KK��h�C8"   >  �  �     �           �     +         �t�bhhK ��h��R�(KK
��h�C(      )   =           ^        �t�bhhK ��h��R�(KK	��h�C$1   #   
   3   6      p         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C         	      	         �t�bhhK ��h��R�(KK	��h�C$�        f  ^     �        �t�bhhK ��h��R�(KK��h�C�   =     �t�bhhK ��h��R�(KK��h�CD                        �  c      l      �   �        �t�bhhK ��h��R�(KK��h�C8      }     �  e  w      �      A   �        �t�bhhK ��h��R�(KK��h�CD   (         L   �  
      �   N  i   h      �   t        �t�bhhK ��h��R�(KK��h�C,      -   �   L   G      �   �        �t�bhhK ��h��R�(KK��h�C0Q  �   :   �             �   �         �t�bhhK ��h��R�(KK
��h�C(W  �     B  -      !  �        �t�bhhK ��h��R�(KK ��h�C�      �     L  �           "   �      (     �  |      �      |      s	                 �  
   �        �t�bhhK ��h��R�(KK��h�C@      ;      ,  %   �              k               �t�bhhK ��h��R�(KK��h�CD#   !      �   }   (      
              %   {
  �        �t�bhhK ��h��R�(KK��h�CX      �     P   �         D  \      �         E  �   �     o  �         �t�bhhK ��h��R�(KK��h�C8
   3   6   �       '   !      �     /         �t�bhhK ��h��R�(KK��h�C0      �  z     �           �        �t�bhhK ��h��R�(KK	��h�C$�      ]  �      �   �         �t�bhhK ��h��R�(KK��h�C�     C        �t�bhhK ��h��R�(KK��h�CX)      �     w        (
          �  �           D  ,               �t�bhhK ��h��R�(KK��h�C�             �t�bhhK ��h��R�(KK��h�CX            v   `         `  T   %         &      U                     �t�bhhK ��h��R�(KK
��h�C(      P   #     ^   �   *        �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C 1     v  �     5         �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�Ch      J   �  `   �     ,         y              9           P           �        �t�bhhK ��h��R�(KK*��h�C�<         	      	      	   K   	   �   	   �   	     	   I  	   �  	   U  	   �  	   �   	   �  	   �  	   /  	   �  	     	   s  	      	   )     �t�bhhK ��h��R�(KK��h�C0      �     i   u  
      �            �t�bhhK ��h��R�(KK��h�C�      L   
   �        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�Cz  +        ;        �t�bhhK ��h��R�(KK��h�C,   Z     �   �      �   \  ]         �t�bhhK ��h��R�(KK��h�CL      5   [      $   �     �     L     +   g      r  '        �t�bhhK ��h��R�(KK��h�CdV     l  �           :   M  &   N            �  �         ,                     �t�bhhK ��h��R�(KK��h�C!        �t�bhhK ��h��R�(KK	��h�C$�        �  i   h          �t�bhhK ��h��R�(KK��h�C        �t�bhhK ��h��R�(KK��h�C@�   q   7     �                    0  s           �t�bhhK ��h��R�(KK��h�C@
   �     2   )   �
        �   �     z   s  �        �t�bhhK ��h��R�(KK��h�CH   D         0   %     �   :   W      &   t  �      �        �t�bhhK ��h��R�(KK��h�C   �                 �t�bhhK ��h��R�(KK��h�C   /   �         �t�bhhK ��h��R�(KK��h�C<   �     �        V   @                       �t�bhhK ��h��R�(KK	��h�C$      )   z   �   
   &        �t�bhhK ��h��R�(KK
��h�C(�          
   ,               �t�bhhK ��h��R�(KK��h�CL               o  ~        8   �     Z     7      �        �t�bhhK ��h��R�(KK
��h�C(   
      �     �  $   
        �t�bhhK ��h��R�(KK��h�CP     S        �t�bhhK ��h��R�(KK��h�CB   	  �   B   R         �t�bhhK ��h��R�(KK	��h�C$   &   N         q            �t�bhhK ��h��R�(KK��h�C@!      ?        ?      
   3   6   )  ?   �   �   r      �t�bhhK ��h��R�(KK��h�CH#          '      #       ?           �   6  ?        �t�bhhK ��h��R�(KK��h�C<�        L      0     r     �   y   �   {        �t�bhhK ��h��R�(KK��h�C �     T  	      	         �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK��h�C89   �  �        �  �        
               �t�bhhK ��h��R�(KK��h�CT      J   M               �  �  &      �   a      �  W              �t�bhhK ��h��R�(KK��h�CL�  v           �  �      `   �            &   0      r
        �t�bhhK ��h��R�(KK��h�CDi     
   _          |  �                         �t�bhhK ��h��R�(KK	��h�C$4      �   :   A   Y      ?     �t�bhhK ��h��R�(KK
��h�C(B     �  
            7         �t�bhhK ��h��R�(KK��h�C0@      )      �  E                    �t�bhhK ��h��R�(KK��h�C0�  �     p      .      �             �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�Cp         8   ,
        ,               5      �      	        3     L           z	        �t�bhhK ��h��R�(KK	��h�C$�     �     z   "   �         �t�bhhK ��h��R�(KK
��h�C(!      R         	      	         �t�bhhK ��h��R�(KK��h�C8      �               .      �
     �
        �t�bhhK ��h��R�(KK��h�C8h        0  7     �              R         �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C   R       �t�bhhK ��h��R�(KK(��h�C�         $        �  
   _        >                   0   �   @        �     $   k            �  @        �                 �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�Cl      �               z         0         V      (   �   �   �     `   �         �        �t�bhhK ��h��R�(KK��h�C,w  �      �        R     �         �t�bhhK ��h��R�(KK��h�C�      /      �t�bhhK ��h��R�(KK��h�C       �     �            �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C�  �      �t�bhhK ��h��R�(KK��h�CD   �         �        #        i     "  �   n         �t�bhhK ��h��R�(KK��h�C@
   �  1  -   4  $   �         �        �	  o         �t�bhhK ��h��R�(KK��h�CX            [  L  y   �     b     �         -   �          �        �t�bhhK ��h��R�(KK��h�C\      ~      �  @         @         @      �  @   ?         "      y        �t�bhhK ��h��R�(KK
��h�C(   }         .   �      �        �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK	��h�C$            M              �t�bhhK ��h��R�(KK��h�C0@   �   �   �        �  �      p         �t�bhhK ��h��R�(KK��h�C"   �  �        �t�bhhK ��h��R�(KK��h�C<      �  c   8   �        o  �  
      �        �t�bhhK ��h��R�(KK��h�C`D      -   0        �      �         z   j   �               �   �  j   �         �t�bhhK ��h��R�(KK��h�C         w     �t�bhhK ��h��R�(KK��h�C       �     r  �  /      �t�bhhK ��h��R�(KK	��h�C$Q    e     %     R         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CU        B   �        �t�bhhK ��h��R�(KK��h�C       O         
  Q      �t�bhhK ��h��R�(KK��h�CT                    �        �      n	  
           �   D        �t�bhhK ��h��R�(KK��h�C;        �   �        �t�bhhK ��h��R�(KK��h�CHv        .   H         `     A         �                 �t�bhhK ��h��R�(KK��h�CX      w   �        J   M   c     �     �  �     �  
   $              �t�bhhK ��h��R�(KK��h�CP      5   #   !      t
     �     U   t      �     8   �   Q         �t�bhhK ��h��R�(KK��h�C\      0      r  �        &      )  +      �  ^   &  
   �                 �t�bhhK ��h��R�(KK��h�CH?
     J                   �	     2   �     �            �t�bhhK ��h��R�(KK��h�C@�   3        S   <     �     �                   �t�bhhK ��h��R�(KK��h�CL  i      z  �	  %            W     E     h       u        �t�bhhK ��h��R�(KK��h�CD   X     4	  q        :   �      '                     �t�bhhK ��h��R�(KK��h�Cz     	      	         �t�bhhK ��h��R�(KK��h�CH`     �   5     �     R        5      )  +   
   c        �t�bhhK ��h��R�(KK��h�C       �  d     L        �t�bhhK ��h��R�(KK	��h�C$1   �        
      �        �t�bhhK ��h��R�(KK��h�C|A   3  �              .      )                                                        	        �t�bhhK ��h��R�(KK��h�C,   =  �     +                     �t�bhhK ��h��R�(KK��h�Ch   &   �   )   D  *  8         K  3     #             `               �           �t�bhhK ��h��R�(KK��h�CT      3     �
  �     
   �   n              �   �  &   �            �t�bhhK ��h��R�(KK��h�Cw
        �t�bhhK ��h��R�(KK��h�CT      �      �      d     @      k  V   2   �           �   �         �t�bhhK ��h��R�(KK��h�C,�     �     z   "        .        �t�bhhK ��h��R�(KK��h�C   �  S        �t�bhhK ��h��R�(KK��h�C�                �t�bhhK ��h��R�(KK��h�C<      �      �t�be.