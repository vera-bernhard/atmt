����      ]�(�numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK&��h�dtype����i4�����R�(K�<�NNNJ����J����K t�b�C�!   �      '   l      ,
     G        N        �     �           �       �     S      �  8   J      �   h      $   �         �t�bhhK ��h��R�(KK��h�CL   `   p   �  l      '   ;   C     7  ;   �     7  ;            �t�bhhK ��h��R�(KK��h�C47  ;         7  ;         7  ;            �t�bhhK ��h��R�(KK��h�C47  ;         7  ;         7  ;            �t�bhhK ��h��R�(KK	��h�C$7  ;   �     7  ;   �        �t�bhhK ��h��R�(KK��h�Cl   `   p   P         =   P      �  P   �     +   �  l      �    �   7       k  1   ,  �      �t�bhhK ��h��R�(KK��h�C<+       �   9   2     �   I      w   �  =  �         �t�bhhK ��h��R�(KK��h�CD!            
        �   �   9   +        j  ;         �t�bhhK ��h��R�(KK��h�C\+   �  l   �   9   Q     2     `     w   �                   w   �        �t�bhhK ��h��R�(KK��h�C,      w   �     �     w   �        �t�bhhK ��h��R�(KK��h�C4      w   �     0  g   y     w   �        �t�bhhK ��h��R�(KK!��h�C�   n   =  �   �     w   �           w   �           w   �           P   �   �  �  *  �      =   P           �t�bhhK ��h��R�(KK��h�Ch   P  `  >   �  n            \        
   �  '  Q     �  �      �   �  (  �         �t�bhhK ��h��R�(KK��h�Cx   >      �     =   G        n   �  �      n   W  �      n   �  �      n   �  �      �  *  �         �t�bhhK ��h��R�(KK��h�Cd*  >   �     =   G        n   c  �      n   �  �      n   V  �   �   �  �  �         �t�bhhK ��h��R�(KK��h�C4   h  6   >   +   �  `   �      P   �        �t�bhhK ��h��R�(KK��h�Cp�   �  h     +       n   �   �   �      n     �   �      n   =  �   �   `   �      
               �t�bhhK ��h��R�(KK��h�CD   �   P  �     �  N  �  �   n   
  �   8   s   �        �t�bhhK ��h��R�(KK��h�CH9   �               w   �     
  -     h     w   �        �t�bhhK ��h��R�(KK��h�C4      w   �     0  g   �	     w   �        �t�bhhK ��h��R�(KK��h�C8  �     w   �     r  g   �     w   �        �t�bhhK ��h��R�(KK��h�Cd   n   '  Q     �  �         w   �           w   �     A   �	  P  `  �           �t�bhhK ��h��R�(KK��h�Ch   >   �  n        
   �  '  Q     �  �         �     w   �     �     w   �        �t�bhhK ��h��R�(KK��h�C<   n   �  �         w   �           w   �        �t�bhhK ��h��R�(KK��h�C,v     w   �           w   �        �t�bhhK ��h��R�(KK��h�C<   n   W  �         w   �           w   �        �t�bhhK ��h��R�(KK��h�C,      w   �     
     w   �        �t�bhhK ��h��R�(KK��h�CX   n   �  �               w   �           w   �           w   �        �t�bhhK ��h��R�(KK��h�CH*  `  >   �  n   V  �         w   �          w   �        �t�bhhK ��h��R�(KK��h�Ct      }   �   �      �   y     �  &   �      n   c  �              w   �           w   �        �t�bhhK ��h��R�(KK��h�C,      w   �           w   �        �t�bhhK ��h��R�(KK��h�CD   n   �  �   v     �     w   �     �     w   �        �t�bhhK ��h��R�(KK��h�C,�     w   �     �     w   �        �t�bhhK ��h��R�(KK��h�C@   �  l   p                     �     �  &        �t�bhhK ��h��R�(KK,��h�C�   l   p                                 	     ~     G   �                         �  =   /   o        1  �   ,   P   '  �  �   c  �         �t�bhhK ��h��R�(KK��h�C`   l   p               l   p         �
        �        k  �      m  ~        �t�bhhK ��h��R�(KK��h�Cl          �  -  +
        �   9      =   /   o     G   �     7      $   �       >         �t�bhhK ��h��R�(KK��h�C`   P   �      4   �    p              �   �  �     
   p   �     P            �t�bhhK ��h��R�(KK��h�C4=  l   p   �
                 �  �         �t�bhhK ��h��R�(KK%��h�C�   l   p                                 �  �      ~     G   �                
   p   �     P      �  �  �            �t�bhhK ��h��R�(KK��h�Cp   l   p         X                                              4   `   p      l         �t�bhhK ��h��R�(KK��h�Cp   
   p   �     P         =   /   o     =         G   �             �  v  �   z   �         �t�bhhK ��h��R�(KK��h�C\   l   p            l   p              �	                                �t�bhhK ��h��R�(KK��h�C`4   `   p      l      �  =   ]     G   �             �  �   z   �   -           �t�bhhK ��h��R�(KK��h�C@            p      l      �         p      l         �t�bhhK ��h��R�(KK��h�C<   l   p                              l         �t�bhhK ��h��R�(KK��h�CLJ  l   p         
   �       '          )     j  �         �t�bhhK ��h��R�(KK��h�Ch   )  �   �   +               '     �  8           �  �              $           �t�bhhK ��h��R�(KK��h�Ct   8     �  �           ;      �      �       !   '   �   �        '   l   p                  �t�bhhK ��h��R�(KK��h�CP   l   p         `   p   l      �     ;      )     ;      �        �t�bhhK ��h��R�(KK��h�CD   '     ,         R     r  g                        �t�bhhK ��h��R�(KK��h�C4      l   p                              �t�bhhK ��h��R�(KK��h�C\   
  l   p         7  ;         7  ;         7  ;         7  ;            �t�bhhK ��h��R�(KK*��h�C�7  ;         7  ;            e                  ~   3   r     
   p   ]  B      �      �         �         $   A  r         �   P            �t�bhhK ��h��R�(KK��h�CT   9  G     P   �         �  �         '   �   �         ;           �t�bhhK ��h��R�(KK%��h�C�   	   m   t      /   �         R   u   �          ;         	   �      �        �         $   �  �            '   ^         �t�bhhK ��h��R�(KK��h�CT'   �   ,         R   �           0  g   �	        e      g            �t�bhhK ��h��R�(KK��h�CP   '   ;   ,         '   ;   ,         �        '   ;   ,            �t�bhhK ��h��R�(KK��h�C@'   ;   ,         '   ;   ,         '   ;   ,   �        �t�bhhK ��h��R�(KK��h�C,'   ;   ,         '   ;   ,   �         �t�bhhK ��h��R�(KK#��h�C�   P   /     P      p   0     �  m     3        b  h     �  m            �  m     �            �  m        �t�bhhK ��h��R�(KK'��h�C�!      �  �   �  p   0  g   �     �  m          �  m          �  m     �     �  m     �     1        6   �     >         �t�bhhK ��h��R�(KK��h�CHW  l   p                              P     ,   �        �t�bhhK ��h��R�(KK��h�C4   l   p               	   ,      �         �t�bhhK ��h��R�(KK��h�CD                             e   �     P           �t�bhhK ��h��R�(KK��h�C@      l   p                     `   p      l         �t�bhhK ��h��R�(KK��h�C0   l   p                             �t�bhhK ��h��R�(KK��h�C8'   �      l   p                              �t�bhhK ��h��R�(KK��h�C8   l   p   �                                �t�bhhK ��h��R�(KK��h�C4�           
                          �t�bhhK ��h��R�(KK
��h�C(   l   p                        �t�bhhK ��h��R�(KK��h�C,      l   p                        �t�bhhK ��h��R�(KK(��h�C�4   `   p   W  l      ~     G   �     �          ~  �   h           
   p   �     P      8            �  2   '        �   9         �t�bhhK ��h��R�(KK��h�CP       �
     /   �              �                 �        �t�bhhK ��h��R�(KK��h�C0         �                 �        �t�bhhK ��h��R�(KK��h�C0�
  $   �  l                           �t�bhhK ��h��R�(KK��h�C      �              �t�bhhK ��h��R�(KK��h�Ce                    �t�bhhK ��h��R�(KK��h�Cd   `   p      l            p             
        �        
   K                 �t�bhhK ��h��R�(KK��h�CD�        �     �  �   �          	                   �t�bhhK ��h��R�(KK��h�CX        >      .  I      O   	   $   [  %   3   G                       �t�bhhK ��h��R�(KK��h�C@   /   �        	   B   P                          �t�bhhK ��h��R�(KK��h�C@                  `   p   '   l      ~     �        �t�bhhK ��h��R�(KK
��h�C(      $   	   "                 �t�bhhK ��h��R�(KK��h�C\      l   p   �	                 	   ,      
   �              �  m        �t�bhhK ��h��R�(KK��h�C@         �   9  p            -           -  �      �t�bhhK ��h��R�(KK	��h�C$   e                        �t�bhhK ��h��R�(KK��h�C                         �t�bhhK ��h��R�(KK
��h�C(               p      l         �t�bhhK ��h��R�(KK
��h�C(                              �t�bhhK ��h��R�(KK
��h�C(            P  p      l         �t�bhhK ��h��R�(KK��h�C                         �t�bhhK ��h��R�(KK��h�C                     �t�bhhK ��h��R�(KK
��h�C(               p      l         �t�bhhK ��h��R�(KK��h�C          �	              �t�bhhK ��h��R�(KK��h�C                     �t�bhhK ��h��R�(KK��h�C                     �t�bhhK ��h��R�(KK��h�C          p      l         �t�bhhK ��h��R�(KK��h�C                �
        �t�bhhK ��h��R�(KK
��h�C(      �        p      l         �t�bhhK ��h��R�(KK��h�CD`   �        �     ~  =   /   o             ~        �t�bhhK ��h��R�(KK��h�C0   �       �      �  �   �  8        �t�bhhK ��h��R�(KK��h�CD   '   �  ;   ,           �     �
     j     Q        �t�bhhK ��h��R�(KK��h�C                     �t�bhhK ��h��R�(KK��h�CP!              �   `       G   �      ~     c  �   G   �         �t�bhhK ��h��R�(KK��h�C\        �
     �
    �         �     {        g   �                    �t�bhhK ��h��R�(KK��h�C<�  ;   ,      g   j           g   j    ~        �t�bhhK ��h��R�(KK��h�C0  l   p                     �        �t�bhhK ��h��R�(KK��h�CH�                           �        �             �t�bhhK ��h��R�(KK��h�CP           '   ;   ,         '   ;   ,         '   ;   ,            �t�bhhK ��h��R�(KK��h�Cp      $   c  l         `   �              �           �
           4   `   p      l         �t�bhhK ��h��R�(KK��h�C\   '   �      l   p         '   �              �                 �        �t�bhhK ��h��R�(KK"��h�C�      l   p           
   p               �           $   �  l            2   �   �     4   `   p      =  >      �t�bhhK ��h��R�(KK ��h�C�   [   S   u   Z                 �           &   6   3        �   
     �  �            /      A        �t�bhhK ��h��R�(KK��h�Cp!        =  
     B      $   /   V        G   �      �       u     �                    �t�bhhK ��h��R�(KK��h�CX   ~       (     �   >         =  >         
     �  >      \        �t�bhhK ��h��R�(KK��h�Cp      ;            ;           ;            ;                 L      :  �     >         �t�bhhK ��h��R�(KK��h�C0               �        '   l         �t�bhhK ��h��R�(KK��h�C4      >         P   �      c  �            �t�bhhK ��h��R�(KK��h�CH   =  >         ;            ;            ;               �t�bhhK ��h��R�(KK!��h�C�           ;         �     ;            ;                     ;            ;      �     ;               �t�bhhK ��h��R�(KK��h�Ct   e   P   �      =   P   o     �  �         4   `   ~   p   ~     �     ,            /   t	        �t�bhhK ��h��R�(KK��h�C,      �                 �        �t�bhhK ��h��R�(KK��h�Ct  @     ;            ;            ;      �     ;            ;            %     �   ^         �t�bhhK ��h��R�(KK'��h�C�        ;            ;            ;                    ;            ;            ;            ;            ;               �t�bhhK ��h��R�(KK��h�Cx   e   P   �      ~     G   �     2   �   �   �   4     �  ~         �  
        x     �   ^         �t�bhhK ��h��R�(KK��h�C\      �           
            ;            ;               *  >         �t�bhhK ��h��R�(KK��h�C`                       e         ;      ~     ;            ;               �t�bhhK ��h��R�(KK"��h�C�  �
     ;            ;            ;               e         ;           ;      r     
           �        �t�bhhK ��h��R�(KK��h�CP                                 G   �      !      ,            �t�bhhK ��h��R�(KK��h�C\   �      1   T        ?            �  �      `   p         �  �   �        �t�bhhK ��h��R�(KK3��h�C�!         ;            ;            ;      <     $     G   �          
   p      '   t	                    �   �
  ?            P   �   $   \     @   �  �  �
  ?   �        �t�bhhK ��h��R�(KK��h�CL   �     �  ;      $   1  -  P  <       �         �      �      �t�bhhK ��h��R�(KK��h�C4         ;      ,      ?   �     *        �t�bhhK ��h��R�(KK%��h�C�4   `   p   �        ?         z   �   �        K     G   �  �           V         	  $             �           �        �t�bhhK ��h��R�(KK��h�CL      P   l   4  �   ?         @   ^               �  �
        �t�bhhK ��h��R�(KK��h�CL=      &     $      G   �        �           �     �        �t�bhhK ��h��R�(KK��h�Cp   P   �         
   �  4     G   �     �   ,   �  |      )     �            %   �             �t�bhhK ��h��R�(KK ��h�C�7            �  p   `   &     8               A   ,   1   �        $   e      <               �   ^         �t�bhhK ��h��R�(KK��h�Ch      
  &   Z  =  �   �   ^      7             �   �
           �   �  �	  ,   I        �t�bhhK ��h��R�(KK'��h�C�{         $      <      $  
   t  ?   x        e  \  t          =      X   o            e  O   F          =         X   o            �t�bhhK ��h��R�(KK'��h�C�   {         p            X      <      }   V     <   4   }      $        e   <         {     I     �     �        '           �t�bhhK ��h��R�(KK��h�C4!   {        l               '           �t�bhhK ��h��R�(KK��h�CT               �           �     $            �     <            �t�bhhK ��h��R�(KK��h�CX   {     P   �      �  l      $      <   n     �   �         ,   �        �t�bhhK ��h��R�(KK"��h�C�!      }      \        ~     �
  �     
           4  �   l  �     7   |      �  p            G   �  �        �t�bhhK ��h��R�(KK��h�CL`   p   ]        �
  �        =   /   o             ~        �t�bhhK ��h��R�(KK��h�C4   �       �         �  �   �  8        �t�bhhK ��h��R�(KK��h�CH   '   �  ;   ,           �     �
     j           Q     �t�bhhK ��h��R�(KK	��h�C$                           �t�bhhK ��h��R�(KK��h�CP!              �          G   �      ~     c  �   G   �         �t�bhhK ��h��R�(KK��h�C\        �
     �
    �         �     {        g   �                    �t�bhhK ��h��R�(KK��h�C<�  ;   ,      g   j           g   j    ~        �t�bhhK ��h��R�(KK
��h�C(  l   p                        �t�bhhK ��h��R�(KK��h�CH�                           �        �             �t�bhhK ��h��R�(KK��h�CP           '   ;   ,         '   ;   ,         '   ;   ,            �t�bhhK ��h��R�(KK��h�Ch      $   c  l         `   �              �           �
           `   p      l      �t�bhhK ��h��R�(KK��h�CP   #  /  K   S         6   ~   �     #       �     $  4        �t�bhhK ��h��R�(KK��h�C`   #  $     �      '   l         #    {              g   �     �  l         �t�bhhK ��h��R�(KK��h�CT*      �   �   u   
           �   <         �  	                    �t�bhhK ��h��R�(KK4��h�C�   �         /   z        �  F   �   �     "  (                 `   *
  �         (            !   '   z  k           7   	   �  �        �   �   �   N     7	  %   }        �t�bhhK ��h��R�(KK��h�CP!   *      �      �   ,   z     7	  	   %   e      s   �     �        �t�bhhK ��h��R�(KK��h�CX   #	     �      '   �   l         4   
        '   ^   #	     �   �        �t�bhhK ��h��R�(KK'��h�C�   *   4   �     �        P   �   $   �           �      '   l   p   H     �     G   �      �     O   �   #     �  %                �t�bhhK ��h��R�(KK��h�Ch�   �   �   #              �     �     �      '   l      B      R        $  4        �t�bhhK ��h��R�(KK"��h�C�      �        �     %   '        '   H     �       �      �  I      �  �     c        G   �        ]         �t�bhhK ��h��R�(KK��h�CP        '   H     s         !   '      ]     0        �        �t�bhhK ��h��R�(KK��h�CH!   *   C   ]           �    C   :   #  $   �      �         �t�bhhK ��h��R�(KK&��h�C�4     0      4   -  ~         �  �     '   �  �     �                       P     �   M          �
        �   �         �t�bhhK ��h��R�(KK)��h�C�A   u   �  z     �      	   $   +     K                  	      $   �  @   �         e   �      	   $         7        n  �      �        �t�bhhK ��h��R�(KK��h�Cd	   $         n  �         �                 O      	        V      x  ;         �t�bhhK ��h��R�(KK��h�CX     %   [   S      V      2              \   �   �   �   �             �t�bhhK ��h��R�(KK:��h�C�w     g  O      w     �   �   ,   k      ,         
   ,   �     �     S            "            )   5      �            N      "        a   S      �            N      P  <      a   S            �t�bhhK ��h��R�(KK-��h�C�*      4      8     S   �      U      2       V   2   _         B      2     o            O   7     V      k   <   S         s     @   �   �   	        �t�bhhK ��h��R�(KK��h�Ch   V   �      [   S      ~        #   �     B      %        
   �     �      �         �t�bhhK ��h��R�(KK��h�Cl   =     �        V         �  �               !   V   �  U              #   1  �     �t�bhhK ��h��R�(KK$��h�C�   V               
   	  
  �           	      �   �     �           T     2  ;      f   	  $     u      �        �t�bhhK ��h��R�(KK��h�C@O   �   V   /   �           �   �  9      1  �        �t�bhhK ��h��R�(KK��h�C\   	         =  �   �      3   �
     C   �         T        `     �         �t�bhhK ��h��R�(KK��h�C<   V   u   C   �     �           �  ,            �t�bhhK ��h��R�(KK$��h�C�   `   �      �
  �   1        9  h        /     �   k           [   S            9           �  @   �     S         �t�bhhK ��h��R�(KK$��h�C�A   #         1              ;                     �         	   
     s   |  <   �   �   
   $   �   �        �        �t�bhhK ��h��R�(KK��h�CP   =      f      C     ;            	   ,            �   j        �t�bhhK ��h��R�(KK#��h�C�	   ,      V   ?      g         *   #  B   $   �  %      �        B   ,   2   �
     I     U        ]   �     #        �t�bhhK ��h��R�(KK��h�Cd   �     %                          #           �                X  �        �t�bhhK ��h��R�(KK��h�Cp   �  2  �         �  �
  h  r   <   _     V   ?      0     �        �  ,         �        �t�bhhK ��h��R�(KK��h�CP!   V   ,              �               /  �     0  g   �        �t�bhhK ��h��R�(KK��h�Cp   V   �                    I     i   k  x   (   �      �  3   B  ?   0  g      �	  �         �t�bhhK ��h��R�(KK-��h�C�   m     �   %   �  �  �     �  �   n   B  ?   0  g      �	     �        e        V      !   V   k     �        �   �  F      8   2   b  +            �t�bhhK ��h��R�(KK<��h�C�	      \        5   b     N   �  �   (         �   T   A   �   �      �  `   �
  C     
   X      G   )  H   7      �     G   )  X      �     <           	   k     �        o  l  $      �   j  �         �t�bhhK ��h��R�(KK%��h�C�      �  �      ,            �   }      	        �  s   |  <   �   �   
   $   �   �        	   $   2   9  �   �      �         �t�bhhK ��h��R�(KK��h�Cx	   ,     �      �   i   l     A            	   ,   P   S     !   0         �   �  f   	   D           �t�bhhK ��h��R�(KK-��h�C�  �     ;      �     
   ,   ;                  9   3         	   +  r      z         �           ,   	   
           r      +  �  �
     B        �t�bhhK ��h��R�(KK8��h�C�	   +  e   r      @  �   
   ,            �   q  �     �  �       $   2   |  
              m   	   r   K            �      /   �        	   o  w  n   �  q      �        '   �  |        �t�bhhK ��h��R�(KK��h�CXo  l  $   �     �  ;      �         	   $   2   9  �   �      �   j        �t�bhhK ��h��R�(KK!��h�C��      	   ,   �      �   i         �     !   0         �   �  f   	            V   �         �     /            �t�bhhK ��h��R�(KK��h�CT     j  p      s     �  �               ;      3   0  g   �        �t�bhhK ��h��R�(KK��h�C                     �t�bhhK ��h��R�(KK��h�C,            L   ;                  �t�bhhK ��h��R�(KK��h�C                     �t�bhhK ��h��R�(KK
��h�C(                     ;         �t�bhhK ��h��R�(KK��h�C@         ;      3   �     =  �   �         �        �t�bhhK ��h��R�(KK
��h�C(   3      L                     �t�bhhK ��h��R�(KK��h�C                     �t�bhhK ��h��R�(KK��h�C0   �  g            {        ;         �t�bhhK ��h��R�(KK��h�C0            ;               ;         �t�bhhK ��h��R�(KK��h�C   �        �        �t�bhhK ��h��R�(KK
��h�C(   3   	              ;         �t�bhhK ��h��R�(KK��h�C0      �      1              ;         �t�bhhK ��h��R�(KK��h�C8                  z  +   T     2  ;         �t�bhhK ��h��R�(KK��h�C                     �t�bhhK ��h��R�(KK	��h�C$�  �              ;         �t�bhhK ��h��R�(KK��h�CH            ;            �   �
             �  }         �t�bhhK ��h��R�(KK
��h�C(         ;            �        �t�bhhK ��h��R�(KK��h�C0                           l         �t�bhhK ��h��R�(KK��h�C4         ;         '   �                  �t�bhhK ��h��R�(KK��h�C@   g      �                 l                     �t�bhhK ��h��R�(KK
��h�C(         �	        g            �t�bhhK ��h��R�(KK$��h�C�   `   p      
   �      V      i     �  	   �     %   b     �      �
  L   ;                    
         �   �        �t�bhhK ��h��R�(KK#��h�C�   p   �     �                 E     ]        �  q         B        �
  3   H        �              �         �t�bhhK ��h��R�(KK��h�Cd                  X           l                     l               m        �t�bhhK ��h��R�(KK��h�C`                  �  j     �        �                                   �t�bhhK ��h��R�(KK��h�C0                                    �t�bhhK ��h��R�(KK��h�C0   r                                �t�bhhK ��h��R�(KK��h�C0            l                        �t�bhhK ��h��R�(KK+��h�C�      �
     N     �      V                   ~               �                |        $         8   �     p      8                 �t�bhhK ��h��R�(KK��h�C@               �
        �     s	        �        �t�bhhK ��h��R�(KK��h�C,         �              �        �t�bhhK ��h��R�(KK��h�C,         �              �        �t�bhhK ��h��R�(KK��h�C,         �                       �t�bhhK ��h��R�(KK��h�C,         C                       �t�bhhK ��h��R�(KK ��h�C�`        �  >            �
     �                  ,   �     �  
   �      !            �  
   �         �t�bhhK ��h��R�(KK%��h�C�`   p      
      �  �  �   <   �      *      ,   E  <   4   G            
      4       
              +   �     +            �t�bhhK ��h��R�(KK��h�C<   =     �   >   �   N  ~      V   �               �t�bhhK ��h��R�(KKH��h�B      m   V   F   �          �      �                     &   .        (               �     (         #      !  �           -      !   &   .              (   +   �   '     �  �   �  #      �   �        M   �  �  5   _   G                    �t�bhhK ��h��R�(KKL��h�B0  !               �      �     $   �                  	            j   �   \      V            "   ,  \         x  ;        �      "                �          
      "   7   )   5         "   �         V   �   �          �         �      �
     /   �        �t�bhhK ��h��R�(KK<��h�C�3   �  �   N  <      V      *   	      #  �   F      �  K   �      D  �           `      7   *   �  S  $         �     �                              �  �     W      &   	   ;  <      /   �   �         �t�bhhK ��h��R�(KK&��h�C�*   	      �      i     �   `   3   �  <                                                      ~        �  
     �        �t�bhhK ��h��R�(KK��h�CL`      V   K         7      p   m          K       �        �t�bhhK ��h��R�(KK��h�C\|   =   |   �   \  C   c     V                        '   �  u   �  9        �t�bhhK ��h��R�(KK��h�C|A   #      �  
               �     
   f      V      2           =   @   �  �  �     <               �t�bhhK ��h��R�(KK��h�CL�   >      
   e       |     c  �   �  �      �     �        �t�bhhK ��h��R�(KK��h�C0     >           �   �   2   �         �t�bhhK ��h��R�(KK	��h�C$   �  >   &  �   c  �         �t�bhhK ��h��R�(KK��h�CDG  �     %  �  �                �   �   �   �         �t�bhhK ��h��R�(KK��h�C@   e   �           �	        /   t	     �          �t�bhhK ��h��R�(KK��h�Cl   =  >      �        �   �   p  7   �   ?      �  �                     �  ^   q        �t�bhhK ��h��R�(KK��h�CH   
  >   v  �   �  �                 ~      G   �        �t�bhhK ��h��R�(KK��h�CT   '  Q     �  �   �	  �      ~      
   �         T   V      k         �t�bhhK ��h��R�(KK��h�Ct   �  >   �   ~   
                 :   S      T      z   �   ~     G  4   P      �   P            �t�bhhK ��h��R�(KK��h�CT   �  -  ~            �     4     H     �  �      
               �t�bhhK ��h��R�(KK��h�CL   �  2   �                    �      �          |        �t�bhhK ��h��R�(KK��h�C,         ~         �   c  �         �t�bhhK ��h��R�(KK��h�C4     -  ~            �     �  �         �t�bhhK ��h��R�(KK!��h�C�   3   }   �   �         �
     �
     }   Q     �  �      2   �   v  �      �     4     H  
      ?            �t�bhhK ��h��R�(KK(��h�C�4   `               �     �      G            2        T   V      k   <   [   S      �   [      `  S   ,            T   V      k         �t�bhhK ��h��R�(KK��h�C`      p   B   �   V      �   �      d          7   P   �   $                     �t�bhhK ��h��R�(KK5��h�C�   
     �         �   0      O     �     �            e      �     �           �            D                      �     �               7     #     S         �t�bhhK ��h��R�(KK��h�C8   V      %      �
     �        4            �t�bhhK ��h��R�(KKD��h�B  O      V      6   [   �        &   .      n             &   A   #   3         �   5         �   W   i    +   4   f     �  `  �      4   6            M     �     �        �      9     X   G   �           M   �  %      W         �t�bhhK ��h��R�(KK��h�CX   �   W   �  �   �   �     W      7      �  �   F  \      =               �t�bhhK ��h��R�(KK��h�CD   [   e  c      9   �   T         7      C  [   ]         �t�bhhK ��h��R�(KK��h�Cx        V   [   S      3         �   �   �   B   B  ;     x	           �  �   �  3   �  g   �	        �t�bhhK ��h��R�(KK0��h�C�   V   �      [   S   0               #   �  g   �	     
   J     �            O    0   �      @      �     '   
         �        =   P     $   �  s   �         �t�bhhK ��h��R�(KK��h�Cd      �   �   �        ?  �     �      �   �      ^                    S        �t�bhhK ��h��R�(KK��h�Cp   V      [   S     %   o   5      �  h                             �                    �t�bhhK ��h��R�(KK��h�C\!   *      �            �    F   /   q            .   �     7               �t�bhhK ��h��R�(KK"��h�C�   S  @     K           �      	   $      F   /   q   K   �     +  	               	   �  r   z  B   o   5         �t�bhhK ��h��R�(KK ��h�C�!      m   V   T                 $   <  r           	   �     �    g        8      �  �      |         �t�bhhK ��h��R�(KK��h�Cx   V   �     �  �     5         �         	            �   �         �     �   �     (   H         �t�bhhK ��h��R�(KK��h�Ch�   �   V      �  t   �     %      1  �     �   �   Y  t         9  �	  g     ^         �t�bhhK ��h��R�(KK'��h�C�O   u   �   �  �   ?   �	  g     ^      B      �      s   �  ^         �   �     !      �  �	  g     ^      C   :   
                 �t�bhhK ��h��R�(KK��h�Cx   |     U      �
     �  �     V      y     M  e                        �        2   ^         �t�bhhK ��h��R�(KK��h�Cx   V   *        $   �     8   k   <   S      7   	   $   u  '   �  �   �  �        s   a   6   A        �t�bhhK ��h��R�(KK��h�CP   V   �   %   �   c       ~        V     �   c  l              �t�bhhK ��h��R�(KK��h�CT`   �           l   
   	   �      ~                 1             �t�bhhK ��h��R�(KK��h�C                     �t�bhhK ��h��R�(KK��h�Ca                    �t�bhhK ��h��R�(KK��h�C�                    �t�bhhK ��h��R�(KK$��h�C�!   *   #       V   $   �   d
     k   <   [   S      2     m  0         �  V      *   V     A      �   	   F   K             �t�bhhK ��h��R�(KK��h�C8   1   #  $   A  t      �     B               �t�bhhK ��h��R�(KK(��h�C�F  V   5                 0   K   #  H   d         x          D   q   H         c            �  0         d   x          )   q            �t�bhhK ��h��R�(KK/��h�C�      2  0      j  g            B   +  V                V         5      <  r   �   �  �   D   q      �        �  r         %  �      �  �  j  g            �t�bhhK ��h��R�(KK��h�CP   Q  B   =   %   G   d        V         `   �   V  0              �t�bhhK ��h��R�(KK��h�C,!   #     �      �        �        �t�bhhK ��h��R�(KK*��h�C�*   V         F  5      c   5                       0   =             M                               �   <       3      f  B      ,        �t�bhhK ��h��R�(KK"��h�C�   �     O   J                      �     F      �     7         5   A  F   �   "         �  �  �            �t�bhhK ��h��R�(KK��h�C\V   v   8   5   $   �                 �  �      �      3   �  �      h        �t�bhhK ��h��R�(KK��h�CX   f  &   V   m   F      4              �   �        �   <   4   a         �t�bhhK ��h��R�(KK��h�Cl   	      +   %   ^      1  �     O      	        +   �   �     +  0   2     +            �t�bhhK ��h��R�(KK%��h�C�J     V         Z  }   �   �  M   �   �   �     7             �        �   �   �           T     o         r  �            �t�bhhK ��h��R�(KK��h�C`   V     [   S      ~        �  @   �  0           
   	   $      +            �t�bhhK ��h��R�(KK
��h�C(   V   C  k  �  >      �        �t�bhhK ��h��R�(KK��h�CH   P  >            P   �        '   �      2   �   v        �t�bhhK ��h��R�(KK��h�CH   *  >            P   �        '   �      z   �   v        �t�bhhK ��h��R�(KK��h�CH      >            P   �        '   �      2   �   �        �t�bhhK ��h��R�(KK��h�CD      >            P   �        '   �      z   �         �t�bhhK ��h��R�(KK��h�C@      >            P   �        '   �      �        �t�bhhK ��h��R�(KK��h�CH      >            P   �        '   �      2   �   �        �t�bhhK ��h��R�(KK��h�C`   V   �     %   �  �     T    �                                         �t�bhhK ��h��R�(KK*��h�C�   	                      P  ~     �  �        -   �     �   �         O     @      6   �      �  0           
            +            �t�bhhK ��h��R�(KK'��h�C�7   �      .          �  +  ,      
         �   5      �  r         W                  \      `           
      ,            �t�bhhK ��h��R�(KK��h�CH   7  �     �  %         �  0   @      6   �      �        �t�bhhK ��h��R�(KK��h�Cl   8   J   $   �      s     @   �      e  1   �  >   �   �     �     
   �     P           �t�bhhK ��h��R�(KK(��h�C�   V               �   �        �      G   �         �                             
      �   �         �            �           �t�bhhK ��h��R�(KK��h�C|�                 ;            '   �            ;            &  �      *  >               ;         �t�bhhK ��h��R�(KK)��h�C�         P   �      }            �                             s	     �                             �	  g   �                    �t�bhhK ��h��R�(KK��h�C8                           �   �           �t�bhhK ��h��R�(KK��h�C`                              s	           �  �                           �t�bhhK ��h��R�(KK��h�C\                  �	  g   �              �                             �t�bhhK ��h��R�(KK��h�C\      �  �     *      e     �            �      7   	   ,         f        �t�bhhK ��h��R�(KK
��h�C(      r  �   N      ?   �        �t�bhhK ��h��R�(KK%��h�C�      �                       �           �     �   /	        �   �   �        �   �	  g   �        N      ?   �        �t�bhhK ��h��R�(KK��h�Cp   �      V         8     S         �         �  @   .  0   n   �	  g     ^      �   
        �t�bhhK ��h��R�(KK��h�CL      5      �  
   e  @   .     �  9   �   T     �   l        �t�bhhK ��h��R�(KK,��h�C�J  ,   V                 �  �        p   e   4   �  
   e  �        e               
            *      e        M  �  V      �  g   R	        �t�bhhK ��h��R�(KK��h�Ct   [   S   �  0   @   .  �   
                9               +        �                     �t�bhhK ��h��R�(KK)��h�C�*      @   .  f      1  �     �  1     �  �      F   �   {           R   �   k   V         T   %         �   R               s   !        �t�bhhK ��h��R�(KK ��h�C�O      $   n  �   �  <     �           �  
   V   $   _  0   +               �        �  o   �   �         �t�bhhK ��h��R�(KK��h�C@*   V   $   �  u     v     �  	   ]      @   �         �t�bhhK ��h��R�(KK��h�Cp   +   ,            4   �     E  9      ?     �   	      �  �     2   *  �                 �t�bhhK ��h��R�(KK��h�Cp   	                  T     o   @   �              �   �           3        6   5         �t�bhhK ��h��R�(KK(��h�C�   8   �     �  =                                         s	     �     �	  g   �                             �   �           �t�bhhK ��h��R�(KK��h�C@!   �  �        �     ,     G      �   �   .        �t�bhhK ��h��R�(KK��h�Ch      �   ,      
   V   	              9   �         '   �   �            A   :        �t�bhhK ��h��R�(KK��h�C@               '   �      _  '   (     �   �        �t�bhhK ��h��R�(KK��h�C<      '                 0	  &   4   '   �         �t�bhhK ��h��R�(KK��h�CD   -      '   �  �        %      U
     
               �t�bhhK ��h��R�(KK��h�C4   =         '   h        '   �           �t�bhhK ��h��R�(KK��h�CL              
   	      �         '   �      '               �t�bhhK ��h��R�(KK��h�C@   6      '   e     e     .   5  >      '   �        �t�bhhK ��h��R�(KK��h�C<	   #         �   5      <   [   �   b   '            �t�bhhK ��h��R�(KK��h�C@   �     '   _     �  �        :   	               �t�bhhK ��h��R�(KK��h�C<      _  	                '   S     x        �t�bhhK ��h��R�(KK��h�CD	            �         �        S      2   �  _        �t�bhhK ��h��R�(KK��h�CT	         L   +   "   d      x   �  I            �   -     |     L      �t�bhhK ��h��R�(KK��h�C@   �  .   �      �  �     .   �       �  �        �t�bhhK ��h��R�(KK��h�CD      �  �   �   a      a   �   2   �  �      2   �        �t�bhhK ��h��R�(KK��h�C@	   �  �      T       E	     	      3     P   A        �t�bhhK ��h��R�(KK��h�CDL        ?   �   �        _  W  �   �  y   @     L      �t�bhhK ��h��R�(KK��h�CH      @        4             ,   |         '   V        �t�bhhK ��h��R�(KK��h�C4   �   p	  '        �   4   a   '   �         �t�bhhK ��h��R�(KK��h�CH7   X  #         �             #   	   �   �   4   d        �t�bhhK ��h��R�(KK��h�CD7      4   d  �   �     !      #      
      �   U        �t�bhhK ��h��R�(KK��h�C@      I  �   o   '   �      h           '   �        �t�bhhK ��h��R�(KK��h�C@�  +         .           �  +           h        �t�bhhK ��h��R�(KK��h�C\�  +      '   �       �  Z   A       o   '   �      �        �           �t�bhhK ��h��R�(KK��h�CH      '   �      4        _         �  �                 �t�bhhK ��h��R�(KK��h�C\U  �            �      %         �   p	     9      L      #   1   k   �   L      �t�bhhK ��h��R�(KK��h�CH�        C   :   �  #      [    %      C   
   #   }        �t�bhhK ��h��R�(KK��h�CH�               }  o         7   	   �         �  �         �t�bhhK ��h��R�(KK��h�C<         7   	   #   �     7   '   �  �  �        �t�bhhK ��h��R�(KK%��h�C�   �     L      W         �      5      �  W        W   3   p	           \   �   �  �   �  �         W      �   e     L      �t�bhhK ��h��R�(KK��h�Cl  �         6   5      3            �         C   ]                       e           �t�bhhK ��h��R�(KK!��h�C�   	   �   B      o   @   .     +         '   �           T     o   �     ,   |               �   �           �t�bhhK ��h��R�(KK��h�Ch!   �	  g   �     P   �   p            �	  g   �        ;            v   	               �t�bhhK ��h��R�(KK��h�CT   �   �     '   �      �     �  	   o   @   �        �
     �        �t�bhhK ��h��R�(KK$��h�C�           �   �   +           G     I     �        T   C   :   
   ,        @   (        
   	   $   �   +   S         �t�bhhK ��h��R�(KK��h�Cp                        `     �                 �            �      '   �  �  �        �t�bhhK ��h��R�(KK%��h�C�   �   `      \                          +       
   �            e   }      
                    l   v   	               �t�bhhK ��h��R�(KK��h�C\O   m   C   ]        ,            s      !   V     &         �
  s           �t�bhhK ��h��R�(KK%��h�C�   1   V   �     s   ^         	      �  1        _         #     2   ^      y     �         @   .  �  �   2              �t�bhhK ��h��R�(KK��h�CX1        V         �   C   :                 7   5   #      "            �t�bhhK ��h��R�(KK��h�C4!   &   Z  f   �   �      1     	            �t�bhhK ��h��R�(KK��h�Cl   b      L     D   h   V         �                    (      ^   
         4           �t�bhhK ��h��R�(KK%��h�C�      �      �     y   ^      3      |         �   S   l  �      �   |      �            �             �   �     �        �t�bhhK ��h��R�(KK0��h�C�         6	     	     �
  �      [   S      j     �         i   Z     6   �     
               "        a      L     �   .      �  (   2   ^      y  H   L      �t�bhhK ��h��R�(KK*��h�C�   1         �         D   h   V         �      �     3         B      �  j           �  "               �   �      P  <      a   S         �t�bhhK ��h��R�(KK#��h�C�         -     "      4   j   �     �  4   j   �     "            d   T   "   2   �      f  
         �      �         �t�bhhK ��h��R�(KK(��h�C�             +      a   S                        �   4  �   B      �        �               Q      �            8   �  �        �t�bhhK ��h��R�(KK*��h�C�   8         -  C   �      �            �  <      a   S                  4   j   �              1      "              2   ^   +   "         �t�bhhK ��h��R�(KK&��h�C�7         �        *   )   �   #   �        ;     j   �         =   "   	  )   ;            j   f              z  '            �t�bhhK ��h��R�(KK��h�CL	        2   ^   +   (               z  '   �     �  �         �t�bhhK ��h��R�(KK"��h�C�      N   '   �         	      N   D   ;         D   �           �   �  �         8      �      �  �   )            �t�bhhK ��h��R�(KK��h�Ct      �      ?   h        ^            �     �  �         '   �     N   �     �  �            �t�bhhK ��h��R�(KK��h�CD�           `   �         �      �   1   1     V         �t�bhhK ��h��R�(KK&��h�C�   m   k   V   t      �   %   r   o   @   �               |  #         [  5         :   #      ^      �         u  (   �   �	  H      �t�bhhK ��h��R�(KK0��h�C�   A      U     "   N      F     K  5            j    )   e  ^   &      
   w  v  Z      �     �            5     (            )     	  (      [  5         �t�bhhK ��h��R�(KK��h�C`:      1   V     �      "   &                )   h   H      &  �   )   h         �t�bhhK ��h��R�(KK��h�C`�         )   e  A     =   �   !        �   C   A   V     �  4   `   V  l        �t�bhhK ��h��R�(KK��h�Cd�      �   #   "   �        �   5     �  "      =   C   :   \   X   E     �  �        �t�bhhK ��h��R�(KK;��h�C�   ,        �   y   Z  a   
   #   �  �   a   S      �  5   �      i  �         +   %      2   a   �            T   "   2   9        �                     p	     �   a         
      $   h  �   �   H      �t�bhhK ��h��R�(KK��h�Ch         �   �   a   S      2   a   +   "      �  �               [        �   P   5      �t�bhhK ��h��R�(KK��h�Cx   M   1      [     :         j  &   )   h      &   '   ^   �   �     �  �      �   8         j        �t�bhhK ��h��R�(KK,��h�C�      �   �      �     �   9     �  �            9      �      L      �     6   5      #   5   <   S      L            )   h   1  ^   �  o   "         �t�bhhK ��h��R�(KK��h�Cx7         D   5              )   h                 2   ^      �      )   h         �  o   "         �t�bhhK ��h��R�(KK��h�CP   1      [        #   5                  �  )   h   A   �        �t�bhhK ��h��R�(KK"��h�C�   M      1   e        )   e  ^               	  �  o   "      7   :         [     �        #   d  �           �t�bhhK ��h��R�(KK��h�CX   �   �  +  V   #               J  �   	   r     �  m  n   �  q         �t�bhhK ��h��R�(KK��h�CD	   +  e   +        K  +  V   �     �         A        �t�bhhK ��h��R�(KK��h�Cl�  +  V         U      �	     ?   x	     *   �   $   A  �         z  s   k  ?   %  R        �t�bhhK ��h��R�(KK)��h�C�   V   �   �      2   �   H     �      �  �   �   �     v  �   9   �
        V   �            4         �     2   �   9     
   	   0
        �t�bhhK ��h��R�(KK��h�C`*   O     3   �  �         J        U      �	     r  V   �  �   9                �t�bhhK ��h��R�(KK!��h�C�   V   Y  d  �        �          K  V   �     �         A        �      �  +   V      	  	   �   Z         �t�bhhK ��h��R�(KK��h�CH   V   �      �  :  
      h   $   �     �          ~        �t�bhhK ��h��R�(KK��h�Cd   3      �            �   V   �     X       %  v   O           {              �t�bhhK ��h��R�(KK��h�C\   1         U      x	          V   $   _        t     �	     [   �         �t�bhhK ��h��R�(KK3��h�C��   	   /   ;         k   V         �
                 �      	   $   �   %      �           _        7      $   -     �     	   �   e   4     $     �      R     �        �t�bhhK ��h��R�(KK&��h�C��   `   7  k   V   +         �  	   $   �         R     �   	   $      3   4   }   a      3         +     �  >      #     *        �t�bhhK ��h��R�(KK��h�CH   O         2  ;      $   _              �	  �   9         �t�bhhK ��h��R�(KK��h�ChY  	   d     �        4      K  V   �        �      �  +   V      	  	   �   Z         �t�bhhK ��h��R�(KK��h�CLV   <  1   <   [   S         	      (     5  +   C   s   a         �t�bhhK ��h��R�(KK��h�CPT     2  ;      $   ;  <            �        ;      ,            �t�bhhK ��h��R�(KK��h�CP�       ;         �        ;      p   �           ,            �t�bhhK ��h��R�(KK��h�C\�     �  ;      $   ;  <   �
     <     !   1  l   p         ?   t  �        �t�bhhK ��h��R�(KK��h�CL   �   �  �  �
     �  �   k         '   ;   u   k   =            �t�bhhK ��h��R�(KK9��h�C�      V            d   �        �
  L   ;            �   '   �      (               V   �  �        ;        '   �  =         *      1  h   �      �  �   I                     ;           �t�bhhK ��h��R�(KK/��h�C�   �  �                 �        V        	   �        "   d   D  "      	      )   �   H   f           �     �     �  �   X   '   h   �      "            �t�bhhK ��h��R�(KK��h�Ct   �      1  h      �   �         s
     P              �   �  ?            �          b         �t�bhhK ��h��R�(KK4��h�C�   9   f           V   :   
   $   �  h        �   	     �          7   h  p   �   �            U   �   �         .     y        w   �  �     �  F              �            �t�bhhK ��h��R�(KK,��h�C�   1   �  >            $   �   %         V      �         �  >   2   �   d  R           %   H     �  3     g         3     g   8     3   �	        �t�bhhK ��h��R�(KK(��h�C�      %     �   H     �  /     U      8     '   a      `   �      �  %   �         �  >     %   e   3   G   �      �         �        �t�bhhK ��h��R�(KK��h�CH*   V     A      �   	   �   T     [   �                   �t�bhhK ��h��R�(KK!��h�C�   �  >   2  F      �  0   %      �  ?   �     �      !      3  
   $   �   �   �  0   %      %   s     g        �t�bhhK ��h��R�(KK!��h�C�   T  1   �      	   $   �  E  �   %      G  %      v   	   2      �   C   6   �       �  O   0   %   K           �t�bhhK ��h��R�(KK��h�CX!      `  ]   �
  	   +   /   �            `   �  ;  0   %   K   �  >         �t�bhhK ��h��R�(KK"��h�C�   	            &     �   (   �              �   (      /        &   �  >   �   "   �        d      J  "         �t�bhhK ��h��R�(KK ��h�C�,   1   ?     H     �      �   W   D  H     ?     �  a         �   �   �      O   M      T   :              �t�bhhK ��h��R�(KK��h�CL�   o  T  Z      s   a      �  K              �              �t�bhhK ��h��R�(KK��h�C|!   *   �  >   �       �     �  �         '   �         -  %   t      �         �  %   T     ~        �t�bhhK ��h��R�(KK$��h�C�   Q    �        $   �   �     S      �                 
        }   �   %  �     F                     �        �t�bhhK ��h��R�(KK6��h�C�*   A   u   �     V        	   [   S      m   <   �            	   f   Z             �  	   0   %      (  K             *   V   $   4  0   %      �  K        h  `   %      �              �t�bhhK ��h��R�(KK ��h�C�!     �  b     S         V   �             �   �   H        e   �  �   9   �
     �	       	   e         �t�bhhK ��h��R�(KK/��h�C��  �      ?      �      �  �               T  F            |  �  �   I         f         .  �	     �  V   �  �      ~        T  �  �	                 �t�bhhK ��h��R�(KK+��h�C�   V   �   P   x     3   '           �  �     �  �      ,               �        ]	  1      1          	   �   F     3   �      X          �t�bhhK ��h��R�(KK'��h�C�   ]   �  �   	   F                            6                 v   V   K   �  �   4   �      O     V      C   ]   �      ~        �t�bhhK ��h��R�(KK��h�Cl�   �     �     #  ?   h           +     r               �
  f        K              �t�bhhK ��h��R�(KK ��h�C�   �      �     #              ;      +     r         9     �      
   $   2   |  �                   �t�bhhK ��h��R�(KK ��h�C�   �      �  ?   r     B   ,         9   
   $   c        c        �        	   ,   e      �	     �
        �t�bhhK ��h��R�(KK��h�CL�      S         u   	         {     ;            1  �         �t�bhhK ��h��R�(KK��h�CL`   p   f     �
     r                1     '   e  q         �t�bhhK ��h��R�(KK��h�C<!      ^  0   K   S         V         �  S         �t�bhhK ��h��R�(KK,��h�C�      V      T        o  }   S          �         S      3   a  g     �      w        �  (      �              �   �  �   �     �            �t�bhhK ��h��R�(KK,��h�C�T  c         M      �     �  s   a         �               D   �   k      m  D   �  h   H     �     D   �   f  H     �   9       �  <   S   H      �t�bhhK ��h��R�(KK��h�CtU  u   t  �  m        T     Q  �   T  F      )  �      [   S         f        �     ~        �t�bhhK ��h��R�(KK ��h�C�   T        V   P                 S   N  �  G  �   �   �  ~            �   N  &  �   n  �   �  9         �t�bhhK ��h��R�(KK��h�CX!   �       $   	      o       }      7   t  �  ,      �     T        �t�bhhK ��h��R�(KK��h�C4:   
   $   �  2  5         	   r  S         �t�bhhK ��h��R�(KK"��h�C�      V      5               �  �  �           �   A      !      1   )   e  @     7         -  �   �           �t�bhhK ��h��R�(KK��h�C4!      �      �     1                    �t�bhhK ��h��R�(KK'��h�C�   b      �      V      L        �         �   l  �     Z      "         �       F   +   "   2   
      d            T   "            �t�bhhK ��h��R�(KK��h�CD   m   �  t      V                        �            �t�bhhK ��h��R�(KKD��h�B  r        d      ]  �     �   �      E         �   �  �   j            �         �      j   �  �     E   @   �     o     �   �   �   �               @   �     �  �  [   6   �        1   �  n        x      
      a  (            �t�bhhK ��h��R�(KK$��h�C�V   c   �           #      X        !   �   (      �     @   q      7   '     #   �   X           d         �           �t�bhhK ��h��R�(KK��h�CL   �         o  �      S            n  �   ~      S           �t�bhhK ��h��R�(KK<��h�C�   5   �      �  K   ~        �        !   *   �           �     �      G     >     g           	                           #   �     �  1   )   q   �            @   �  �      ?                  �t�bhhK ��h��R�(KK.��h�C�*   1   V   ]  0   G   �      �   _   @   �  �    �      U     2      �     /   q      �  <   ~          	         8                 r      G   �        �t�bhhK ��h��R�(KKI��h�B$     V         5            ,   �      
         ]   �   �        #         
      �     �   :   @  #      !   `      D        :   X      �   H   �      D   5      M   )   q   �  %   K   (      D   �   ^      !      K   �   a               �               �t�bhhK ��h��R�(KK��h�Ch!   @   �     �     �      V      V   �   b   �      4  2   �  +                        �t�bhhK ��h��R�(KK��h�CH   V   m   �      �        �   
   �  $   j     @   �         �t�bhhK ��h��R�(KK!��h�C�      1     %   &      �   	   _            '   &  l   
   p              %      !                         �t�bhhK ��h��R�(KK!��h�C�   V   f            *         �   0      �   _   V      m   	   Z   �        �  r      �      s   �      V         �t�bhhK ��h��R�(KK-��h�C�   V                  �  (        B         )   e              B   �     2   �  +         �  (         E  	        M      �  �  �   ]            �t�bhhK ��h��R�(KK-��h�C�            V         r           M   O   D   �   U   T   :           _      �   3     "                   6           �     +  3              �t�bhhK ��h��R�(KK)��h�C�!   k   V   c            f        d           E  	     7      d      �   +         
   #   �         �     
         �                �t�bhhK ��h��R�(KK��h�CD   V   �   +         q  c  �   o  �         E  O        �t�bhhK ��h��R�(KK��h�C|   V   �  B   2   �  +         �       �     	   N              	   c           3   U     G        �t�bhhK ��h��R�(KK��h�C4      @   �  =     s   �  �               �t�bhhK ��h��R�(KK��h�CP      *   V   ^        $                        �  	   B         �t�bhhK ��h��R�(KK��h�Cd!   @   �     
   J   $   u  T           �     G     ?      �     �
     �        �t�bhhK ��h��R�(KK��h�C\D     V      �   o   �   �                     �  ,   	      @      �        �t�bhhK ��h��R�(KK��h�CT   V            �         �   ^   ,        �   �      6              �t�bhhK ��h��R�(KK"��h�C�   V         9   �   �  k     �  
   N     6   I         	   �        
   �   �  F   B            �   ^         �t�bhhK ��h��R�(KK��h�Ct   V      6                �	                       e   �     �             "           �t�bhhK ��h��R�(KK��h�CH                  7   �        �   y          V         �t�bhhK ��h��R�(KK8��h�C�V   �  \        D   ;     #   @           !   6  
         +      �    �  9              �               4           d   �   �     +               9  V           �  /   z        �t�bhhK ��h��R�(KK��h�CX   	   �     %   /   ;        �          2   ^   +         6   5         �t�bhhK ��h��R�(KK��h�Cl   V         /   ;              $   �             2   ^   +   @      D   �      �         �t�bhhK ��h��R�(KK.��h�C�!   @   �   f      (      	               r  C          n  V  �                2   ^   +      �      �         r     �   C     �         D   y        �t�bhhK ��h��R�(KK4��h�C�!   _      +   "      g     ;      	      �         9               �      �   �     4   G   �  =  �      7        	   �	             �        �   p  <   S      '   �         �t�bhhK ��h��R�(KK#��h�C�	        2   ^   +      �      	      N   D   ;               N   '   �               z  '      <   S      �  �         �t�bhhK ��h��R�(KK ��h�C�   �   1         "      D   ;      M      �   �     �     @      )   �      ^      8   	      �  &   "         �t�bhhK ��h��R�(KK ��h�C�M      �   x   "         �     *   	   }  "         <   S            "         �   @      )   �      (        �t�bhhK ��h��R�(KK&��h�C�         �   �     &      �     �   =      �     �  
         �   J         S      ,   �     �
     �        ,               �t�bhhK ��h��R�(KK:��h�C�   _            �        1         @   ^   2   �   �   d  �      �   ;  �   d  R     G     �     6  �   �   
   �         7      �   #               �        e            �   M      �   M        �t�bhhK ��h��R�(KK��h�Ch         e                             G  �	  a   
   #   �     C     �  �        �t�bhhK ��h��R�(KK��h�Cp   �     �              �   �   "  �     0         b               �         "   �         �t�bhhK ��h��R�(KK��h�CH�   �  V   4   6           �      '   ;        	            �t�bhhK ��h��R�(KK*��h�C�         -   5      #   �      -         u  -   �   �     4        7   	      �   �    ~     D   q         �      �         '   a            �t�bhhK ��h��R�(KK5��h�C�   +  1   �  !     -   ~                 -   5         &  0            �   8	           9   �     @   .     :   �  
   J     �   8	  t         ^   
         +   @   �            �t�bhhK ��h��R�(KK��h�CL   *   V   u   7           v   	   /   ;        k   <   S         �t�bhhK ��h��R�(KK��h�C8   	     4   6           e   �     �        �t�bhhK ��h��R�(KK��h�C|   �  K  �
        \  
   p   �  �   M  E   �        P   '     �     4        U     �     �         �t�bhhK ��h��R�(KK��h�Cl      `            	         Q      �         ?   @   ^         c  �   N   �     �        �t�bhhK ��h��R�(KK��h�C`&  �   Q   N         &  �   Q                  
         u  T                  �t�bhhK ��h��R�(KK��h�C@   V   �         �
  =   Q  l      �  "	     �        �t�bhhK ��h��R�(KK��h�C               r        �t�bhhK ��h��R�(KK��h�C<   l   p                           �  �         �t�bhhK ��h��R�(KK��h�CP   l   p                    �  �      `   p   ~        �        �t�bhhK ��h��R�(KK��h�CT      l   p         G                  `   p      l      �  &        �t�bhhK ��h��R�(KK��h�C|   ,               ,      �     !            $      �  >      �   �     O  �      t	        �        �t�bhhK ��h��R�(KK��h�C<P  l   p   f           2           �  &        �t�bhhK ��h��R�(KK,��h�C�   l   p   �      J         �   u     G   l      r  �               8                  r  �   �  �  o         T     o              '   �         �t�bhhK ��h��R�(KK
��h�C(!   z  �  l         �  �         �t�bhhK ��h��R�(KK��h�C �  l   p                  �t�bhhK ��h��R�(KK��h�C    l   p                  �t�bhhK ��h��R�(KK��h�CX      l   p                  $   Z  }   l      !      l   p   �  '        �t�bhhK ��h��R�(KK��h�C    l   p                  �t�bhhK ��h��R�(KK��h�C`   l   p                        �              �                 �        �t�bhhK ��h��R�(KK��h�C8   l   p   ~                       �        �t�be.