��vz      ]�(�numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i4�����R�(K�<�NNNJ����J����K t�b�C0   *      �     �  �     �           �t�bhhK ��h��R�(KK��h�C s      -   �              �t�bhhK ��h��R�(KK��h�C0@    �  .   �  �   z   �  >  I         �t�bhhK ��h��R�(KK	��h�C$�     �  6   �     %        �t�bhhK ��h��R�(KK��h�C�     �             �t�bhhK ��h��R�(KK��h�C<   H   2   7      P     �           
   �        �t�bhhK ��h��R�(KK��h�C\
      "   �   
   &   [            =         &   �                         �t�bhhK ��h��R�(KK��h�C      &   �       �t�bhhK ��h��R�(KK��h�C�  :  e     �t�bhhK ��h��R�(KK��h�C,(      <               <            �t�bhhK ��h��R�(KK��h�C[   X         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C[                    �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C   <              �t�bhhK ��h��R�(KK��h�C~            �t�bhhK ��h��R�(KK��h�C	        �t�bhhK ��h��R�(KK��h�C~       
     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�     C      �t�bhhK ��h��R�(KK��h�Cx$      �     $   U           @   �           �     
   �  Z   $   �  a      �     .   �   �         �t�bhhK ��h��R�(KK��h�C s   V  <  �              �t�bhhK ��h��R�(KK
��h�C(�     �  �  d  I               �t�bhhK ��h��R�(KK
��h�C(      7         *   Q   2         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cx�   s      $            �  	      t     )            E      s     �      �     �      �     �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK	��h�C$�   s      $                  �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK
��h�C(         B   �   Z   >            �t�bhhK ��h��R�(KK��h�C4      �      C   X      �  #     �         �t�bhhK ��h��R�(KK��h�C`&   �         �     L      �   	                     �   �  �  k     )         �t�bhhK ��h��R�(KK��h�C0p     D   i            9      !         �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8   *         �     '     �      n           �t�bhhK ��h��R�(KK��h�C8   <          *         �                �t�bhhK ��h��R�(KK��h�C4�   U   *      D   g           W   @        �t�bhhK ��h��R�(KK��h�CD   *      '   
     �     v   �      �                 �t�bhhK ��h��R�(KK��h�C@   �     B   -   @        v  >     �   P           �t�bhhK ��h��R�(KK��h�C,�     �   �   )      �   l  �        �t�bhhK ��h��R�(KK��h�CD   �     n  �      C      �  X      �  #     �        �t�bhhK ��h��R�(KK��h�CT      �     L      �   �      �  	   5  �  �  4           F
        �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C   X      �            �t�bhhK ��h��R�(KK��h�CA   
           �t�bhhK ��h��R�(KK��h�C[   X      �      �t�bhhK ��h��R�(KK��h�CL
         ?     I   �        @   f        M        q         �t�bhhK ��h��R�(KK��h�C<    x   /   
      4   "   '   �         �         �t�bhhK ��h��R�(KK��h�CD      -   �   
   W   �  	         F   �      Q  �         �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C     �     �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�Cz     �t�bhhK ��h��R�(KK��h�C   *                  �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C�  !        �t�bhhK ��h��R�(KK��h�C            �   �        �t�bhhK ��h��R�(KK��h�C8                     	            �        �t�bhhK ��h��R�(KK��h�CDD      9      .   t     }  v   B      �   �   Z   p        �t�bhhK ��h��R�(KK
��h�C(      7         9   Q   2         �t�bhhK ��h��R�(KK��h�C         z     �t�bhhK ��h��R�(KK��h�C0t  �   /  	   ^                       �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C*        �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�Cq     �t�bhhK ��h��R�(KK��h�CW   �     �t�bhhK ��h��R�(KK��h�C`   *   C     D  E           �      F   k   	   t          �      r  �         �t�bhhK ��h��R�(KK��h�C0p     �     �   �  �        �        �t�bhhK ��h��R�(KK	��h�C$               a  �         �t�bhhK ��h��R�(KK��h�C<   *         D           $      L   �   �        �t�bhhK ��h��R�(KK��h�C�     �        �t�bhhK ��h��R�(KK��h�C<   *   3     D           $      �   �   �         �t�bhhK ��h��R�(KK��h�C         W   �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�CG                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK
��h�C(�     $      *                 �t�bhhK ��h��R�(KK��h�CA   3        �t�bhhK ��h��R�(KK��h�C       $      ?           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK��h�C�     C      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CV           L      �t�bhhK ��h��R�(KK��h�Cz     �t�bhhK ��h��R�(KK��h�CW   �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK
��h�C(   *      �  �     �   �         �t�bhhK ��h��R�(KK��h�C   *      �   l        �t�bhhK ��h��R�(KK	��h�C$�   �     )                  �t�bhhK ��h��R�(KK��h�C8�  
   �  w  �   n    z   6   f     &        �t�bhhK ��h��R�(KK��h�CH
         F   D  O   �         �         i   
   l  �        �t�bhhK ��h��R�(KK��h�C4N      �   
   l  6              x        �t�bhhK ��h��R�(KK	��h�C$      D   g   �  M   �        �t�bhhK ��h��R�(KK��h�CP     �     *      D   g   �     v  $      9   	   !      8         �t�bhhK ��h��R�(KK��h�C,   6   c  �   �   J   `      *         �t�bhhK ��h��R�(KK	��h�C$      O      M   q   �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C`   
   d     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C                   �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C,   *   �       �        U        �t�bhhK ��h��R�(KK	��h�C$�   V     )                  �t�bhhK ��h��R�(KK��h�C,     �  B   a   M   *   Q   2         �t�bhhK ��h��R�(KK��h�C               �t�bhhK ��h��R�(KK��h�Cf     �             �t�bhhK ��h��R�(KK��h�CT   �   :        �         D   =         H         i                 �t�bhhK ��h��R�(KK��h�CP        H   2         �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C`                 �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK��h�C0   *      �     �  �     �           �t�bhhK ��h��R�(KK��h�C s      -   �              �t�bhhK ��h��R�(KK��h�C0@    �  .   �  �   z   �  >  I         �t�bhhK ��h��R�(KK	��h�C$�     �  6   �     %        �t�bhhK ��h��R�(KK��h�C�     �             �t�bhhK ��h��R�(KK��h�C<   H   2   7      P     �           
   �        �t�bhhK ��h��R�(KK��h�C\
      "   �   
   &   [            =         &   �                         �t�bhhK ��h��R�(KK��h�C      &   �       �t�bhhK ��h��R�(KK��h�C�  :  e     �t�bhhK ��h��R�(KK��h�C,(      <               <            �t�bhhK ��h��R�(KK��h�C[   X         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C[                    �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C   <              �t�bhhK ��h��R�(KK��h�C~            �t�bhhK ��h��R�(KK��h�C	        �t�bhhK ��h��R�(KK��h�C~       
     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�     C      �t�bhhK ��h��R�(KK��h�Cx$      �     $   U           @   �           �     
   �  Z   $   �  a      �     .   �   �         �t�bhhK ��h��R�(KK��h�C s   V  <  �              �t�bhhK ��h��R�(KK
��h�C(�     �  �  d  I               �t�bhhK ��h��R�(KK
��h�C(      7         *   Q   2         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cx�   s      $            �  	      t     )            E      s     �      �     �      �     �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK	��h�C$�   s      $                  �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK
��h�C(         B   �   Z   >            �t�bhhK ��h��R�(KK��h�C4      �      C   X      �  #     �         �t�bhhK ��h��R�(KK��h�C`&   �         �     L      �   	                     �   �  �  k     )         �t�bhhK ��h��R�(KK��h�C0p     D   i            9      !         �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8   *         �     '     �      n           �t�bhhK ��h��R�(KK��h�C8   <          *         �                �t�bhhK ��h��R�(KK��h�C4�   U   *      D   g           W   @        �t�bhhK ��h��R�(KK��h�CD   *      '   
     �     v   �      �                 �t�bhhK ��h��R�(KK��h�C@   �     B   -   @        v  >     �   P           �t�bhhK ��h��R�(KK��h�C,�     �   �   )      �   l  �        �t�bhhK ��h��R�(KK��h�CD   �     n  �      C      �  X      �  #     �        �t�bhhK ��h��R�(KK��h�CT      �     L      �   �      �  	   5  �  �  4           F
        �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C   X      �            �t�bhhK ��h��R�(KK��h�CA   
           �t�bhhK ��h��R�(KK��h�C[   X      �      �t�bhhK ��h��R�(KK��h�CL
         ?     I   �        @   f        M        q         �t�bhhK ��h��R�(KK��h�C<    x   /   
      4   "   '   �         �         �t�bhhK ��h��R�(KK��h�CD      -   �   
   W   �  	         F   �      Q  �         �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C     �     �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�Cz     �t�bhhK ��h��R�(KK��h�C   *                  �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C�  !        �t�bhhK ��h��R�(KK��h�C            �   �        �t�bhhK ��h��R�(KK��h�C8                     	            �        �t�bhhK ��h��R�(KK��h�CDD      9      .   t     }  v   B      �   �   Z   p        �t�bhhK ��h��R�(KK
��h�C(      7         9   Q   2         �t�bhhK ��h��R�(KK��h�C         z     �t�bhhK ��h��R�(KK��h�C0t  �   /  	   ^                       �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C*        �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�Cq     �t�bhhK ��h��R�(KK��h�CW   �     �t�bhhK ��h��R�(KK��h�C`   *   C     D  E           �      F   k   	   t          �      r  �         �t�bhhK ��h��R�(KK��h�C0p     �     �   �  �        �        �t�bhhK ��h��R�(KK	��h�C$               a  �         �t�bhhK ��h��R�(KK��h�C<   *         D           $      L   �   �        �t�bhhK ��h��R�(KK��h�C�     �        �t�bhhK ��h��R�(KK��h�C<   *   3     D           $      �   �   �         �t�bhhK ��h��R�(KK��h�C         W   �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�CG                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK
��h�C(�     $      *                 �t�bhhK ��h��R�(KK��h�CA   3        �t�bhhK ��h��R�(KK��h�C       $      ?           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK��h�C�     C      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CV           L      �t�bhhK ��h��R�(KK��h�Cz     �t�bhhK ��h��R�(KK��h�CW   �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK
��h�C(   *      �  �     �   �         �t�bhhK ��h��R�(KK��h�C   *      �   l        �t�bhhK ��h��R�(KK	��h�C$�   �     )                  �t�bhhK ��h��R�(KK��h�C8�  
   �  w  �   n    z   6   f     &        �t�bhhK ��h��R�(KK��h�CH
         F   D  O   �         �         i   
   l  �        �t�bhhK ��h��R�(KK��h�C4N      �   
   l  6              x        �t�bhhK ��h��R�(KK	��h�C$      D   g   �  M   �        �t�bhhK ��h��R�(KK��h�CP     �     *      D   g   �     v  $      9   	   !      8         �t�bhhK ��h��R�(KK��h�C,   6   c  �   �   J   `      *         �t�bhhK ��h��R�(KK	��h�C$      O      M   q   �        �t�bhhK ��h��R�(KK��h�C         1     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C`   
   d           �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C                   �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C,   *   �       �        U        �t�bhhK ��h��R�(KK	��h�C$�   V     )                  �t�bhhK ��h��R�(KK��h�C,     �  B   a   M   *   Q   2         �t�bhhK ��h��R�(KK��h�C               �t�bhhK ��h��R�(KK��h�Cf     �             �t�bhhK ��h��R�(KK��h�CT   �   :        �         D   =         H         i                 �t�bhhK ��h��R�(KK��h�CP        H   2         �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C`                 �t�bhhK ��h��R�(KK��h�C[   X      �t�bhhK ��h��R�(KK��h�C0   *      �     �  �     �           �t�bhhK ��h��R�(KK��h�C s      -   �              �t�bhhK ��h��R�(KK��h�C0@    �  .   �  �   z   �  >  I         �t�bhhK ��h��R�(KK	��h�C$�     �  6   �     %        �t�bhhK ��h��R�(KK��h�C�     �             �t�bhhK ��h��R�(KK��h�C<   H   2   7      P     �           
   �        �t�bhhK ��h��R�(KK��h�C\
      "   �   
   &   [            =         &   �                         �t�bhhK ��h��R�(KK��h�C      &   �       �t�bhhK ��h��R�(KK��h�C�  :  e     �t�bhhK ��h��R�(KK��h�C,(      <               <            �t�bhhK ��h��R�(KK��h�C[   X         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C[                    �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C   <              �t�bhhK ��h��R�(KK��h�C~            �t�bhhK ��h��R�(KK��h�C	        �t�bhhK ��h��R�(KK��h�C~       
     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�     C      �t�bhhK ��h��R�(KK��h�Cx$      �     $   U           @   �           �     
   �  Z   $   �  a      �     .   �   �         �t�bhhK ��h��R�(KK��h�C s   V  <  �              �t�bhhK ��h��R�(KK
��h�C(�     �  �  d  I               �t�bhhK ��h��R�(KK
��h�C(      7         *   Q   2         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�Cx�   s      $            �  	      t     )            E      s     �      �     �      �     �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK	��h�C$�   s      $                  �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK
��h�C(         B   �   Z   >            �t�bhhK ��h��R�(KK��h�C4      �      C   X      �  #     �         �t�bhhK ��h��R�(KK��h�C`&   �         �     L      �   	                     �   �  �  k     )         �t�bhhK ��h��R�(KK��h�C0p     D   i            9      !         �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�C%            �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8   *         �     '     �      n           �t�bhhK ��h��R�(KK��h�C8   <          *         �                �t�bhhK ��h��R�(KK��h�C4�   U   *      D   g           W   @        �t�bhhK ��h��R�(KK��h�CD   *      '   
     �     v   �      �                 �t�bhhK ��h��R�(KK��h�C@   �     B   -   @        v  >     �   P           �t�bhhK ��h��R�(KK��h�C,�     �   �   )      �   l  �        �t�bhhK ��h��R�(KK��h�CD   �     n  �      C      �  X      �  #     �        �t�bhhK ��h��R�(KK��h�CT      �     L      �   �      �  	   5  �  �  4           F
        �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C   X      �            �t�bhhK ��h��R�(KK��h�CA   
           �t�bhhK ��h��R�(KK��h�C[   X      �      �t�bhhK ��h��R�(KK��h�CL
         ?     I   �        @   f        M        q         �t�bhhK ��h��R�(KK��h�C<    x   /   
      4   "   '   �         �         �t�bhhK ��h��R�(KK��h�CD      -   �   
   W   �  	         F   �      Q  �         �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C     �     �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�Cz     �t�bhhK ��h��R�(KK��h�C   *                  �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C�  !        �t�bhhK ��h��R�(KK��h�C            �   �        �t�bhhK ��h��R�(KK��h�C8                     	            �        �t�bhhK ��h��R�(KK��h�CDD      9      .   t     }  v   B      �   �   Z   p        �t�bhhK ��h��R�(KK
��h�C(      7         9   Q   2         �t�bhhK ��h��R�(KK��h�C         }     �t�bhhK ��h��R�(KK��h�C0t  �   /  	   ^                       �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C*        �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�Cq     �t�bhhK ��h��R�(KK��h�CW   �     �t�bhhK ��h��R�(KK��h�C`   *   C     D  E           �      F   k   	   t          �      r  �         �t�bhhK ��h��R�(KK��h�C0p     �     �   �  �        �        �t�bhhK ��h��R�(KK	��h�C$               a  �         �t�bhhK ��h��R�(KK��h�C<   *         D           $      L   �   �        �t�bhhK ��h��R�(KK��h�C�     �        �t�bhhK ��h��R�(KK��h�C<   *   3     D           $      �   �   �         �t�bhhK ��h��R�(KK��h�C         R     �     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�CG                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK
��h�C(�     $      *                 �t�bhhK ��h��R�(KK��h�CA   3        �t�bhhK ��h��R�(KK��h�C       $      ?           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C  �      �t�bhhK ��h��R�(KK��h�C�         �     �t�bhhK ��h��R�(KK��h�Cj          �t�bhhK ��h��R�(KK��h�C7     �t�bhhK ��h��R�(KK��h�Ck     &     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C<   *      �         O  .
  B           1         �t�bhhK ��h��R�(KK��h�C4.      �  {      E     �      Y  k
        �t�bhhK ��h��R�(KK��h�C8.   8  a          }               >            �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C`d      �   ;     .     s      @      �   	   5        �  .
  B     H   �         �t�bhhK ��h��R�(KK��h�C0      g   �   �      *   M      �        �t�bhhK ��h��R�(KK��h�Cv     !     �t�bhhK ��h��R�(KK��h�Cv     !           �t�bhhK ��h��R�(KK��h�C�      *           �t�bhhK ��h��R�(KK��h�C�      *           �t�bhhK ��h��R�(KK��h�C<
                 @      �           *         �t�bhhK ��h��R�(KK��h�C@�             X  x  y           %              �t�bhhK ��h��R�(KK��h�Cy        �t�bhhK ��h��R�(KK��h�C �      z                 �t�bhhK ��h��R�(KK��h�C �      z                 �t�bhhK ��h��R�(KK��h�CH   �      �t�bhhK ��h��R�(KK��h�C@H   �      O     B  �     B         �      w        �t�bhhK ��h��R�(KK��h�CX.      �  Z      �   
   H   �     x     �       :   M  O      �         �t�bhhK ��h��R�(KK��h�C             �  �        �t�bhhK ��h��R�(KK��h�C8H   �         D    �     D    �           �t�bhhK ��h��R�(KK��h�CT
      �   i   
      �   	   �        x     �      D      2         �t�bhhK ��h��R�(KK��h�C4      -        �     D              �t�bhhK ��h��R�(KK
��h�C(      D   @   �     �           �t�bhhK ��h��R�(KK��h�CD  �      @      �         r   M       �     �        �t�bhhK ��h��R�(KK��h�CP       �  i   
      �   d   �   	   �      �  {      w  '   I         �t�bhhK ��h��R�(KK��h�C(      <            �t�bhhK ��h��R�(KK��h�C `      I        n        �t�bhhK ��h��R�(KK��h�C<g  .   �      g  J   `   
      $     g  �         �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�CA   �          �t�bhhK ��h��R�(KK��h�C `   
   �      +           �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�CH   !                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C8   "     Z         {     *      *  v        �t�bhhK ��h��R�(KK��h�C4   
   �     �   7         j   �           �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C\
      �   
         	   5      '            �   
         *      9            �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C=  "         *         �t�bhhK ��h��R�(KK	��h�C$      7            2         �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C  �      �t�bhhK ��h��R�(KK��h�C4   *      Z   >      v   B      �          �t�bhhK ��h��R�(KK��h�C           �         �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK
��h�C(                  E      �     �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�C`
   J   �   "   �     F      �     �     �     �     �  �  �  :   �  �        �t�bhhK ��h��R�(KK
��h�C(=   r     .  N   �  "   �        �t�bhhK ��h��R�(KK��h�Cl      �      �t�bhhK ��h��R�(KK��h�Cd
        J   �  G  l   p  /      �  /      l   	         =   q   �     �           �t�bhhK ��h��R�(KK��h�C0�  �      �  �      /        $         �t�bhhK ��h��R�(KK��h�C�     q      �t�bhhK ��h��R�(KK��h�C�  �  �     �t�bhhK ��h��R�(KK��h�C(   �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK	��h�C$         y      �     /     �t�bhhK ��h��R�(KK��h�C0      �   �        �t�bhhK ��h��R�(KK��h�C(         �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK
��h�C(+      �     �                 �t�bhhK ��h��R�(KK��h�CP
              "   ,   �  	         =   �   	  
  !  _   (        �t�bhhK ��h��R�(KK��h�C"        �        �t�bhhK ��h��R�(KK��h�C:   _   (     �t�bhhK ��h��R�(KK��h�C(      <      C     �t�bhhK ��h��R�(KK��h�C�   	  
        �t�bhhK ��h��R�(KK��h�C :   _   #                 �t�bhhK ��h��R�(KK��h�Cj          �t�bhhK ��h��R�(KK��h�CX       	      F   q     �   	   "   {      D     :   |  }  �   +         �t�bhhK ��h��R�(KK��h�CXY      "   �  S     *      @          *      	      F         �        �t�bhhK ��h��R�(KK��h�C,�  ;   x          D  a      �        �t�bhhK ��h��R�(KK��h�CXq     �      4   �         �  W  	      �     '              Y        �t�bhhK ��h��R�(KK��h�C         j          �t�bhhK ��h��R�(KK��h�C@
      "   �   :        �   	   =         *            �t�bhhK ��h��R�(KK��h�C*   Q         �t�bhhK ��h��R�(KK��h�C|	        <            �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C      �                 �t�bhhK ��h��R�(KK��h�CD
      "   �   :        �   	   =   *   Q   c      S        �t�bhhK ��h��R�(KK��h�C*   Q   c      S     �t�bhhK ��h��R�(KK��h�C(      <            �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C      "                 �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C   
     �           �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C    
   �      _           �t�bhhK ��h��R�(KK��h�C7     �t�bhhK ��h��R�(KK��h�C4
          	   =   *   Q   �              �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C �                        �t�bhhK ��h��R�(KK��h�C@
           	         -   =   0      �      *         �t�bhhK ��h��R�(KK��h�C0      �      �t�bhhK ��h��R�(KK��h�Cs  �      �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C(      <      D     �t�bhhK ��h��R�(KK��h�CA            �t�bhhK ��h��R�(KK��h�C 0                       �t�bhhK ��h��R�(KK��h�C         7     �t�bhhK ��h��R�(KK��h�Ck     &     �t�be.