underhållsbidrag (8/8)
länge (27/27)
handikapporganisationer (1/1)
verka (2/2)
kom (18/18)
Nuortennettifinska (1/1)
breddgraderna (1/1)
nätbankskoderfinska (1/1)
kejsarsnitt (3/3)
medborgarskapet (1/1)
redaktioner (1/1)
parförhållanden (3/3)
delat (1/1)
djur (1/1)
trivas (1/1)
fett (1/1)
firas (11/11)
HSL (2/2)
socialverk (2/2)
serviceställena (1/1)
garantipension (2/2)
skriftlig (7/7)
tema (1/1)
Hedersrelaterat (1/1)
Eira (1/1)
efterskott (4/4)
lagakraftvunnet (1/1)
ansökningstider (2/2)
rötterna (1/1)
kön (22/22)
digitalbox (1/1)
redogörelsen (1/1)
styrkor (1/1)
Begravningbyråers (1/1)
tandklinikerna (1/1)
gren (1/1)
trappuppgången (1/1)
uppsikt (3/3)
Insurance (1/1)
byråer (3/3)
skryter (1/1)
tidningar (9/9)
äter (4/4)
byggnader (2/2)
förväntar (5/5)
polikliniker (2/2)
bekantat (1/1)
ungdomsgårdarna (4/4)
nära (13/13)
sparas (2/2)
dekorerat (1/1)
Väestöliitto (6/6)
handikappservicen (2/2)
uppstartsföretagare (11/11)
etc (1/1)
presidentens (1/1)
datoranvändningen (1/1)
skick (7/7)
infödda (1/1)
daghemfinska (1/1)
personliga (3/3)
folkpensionens (1/1)
Spa (1/1)
praktiska (7/7)
tagalog (1/1)
examensnivåerna (1/1)
följeslagare (1/1)
kerho (1/1)
vigseltillfället (1/1)
räknats (1/1)
framför (1/1)
säkerhetstjänster (1/1)
musikgrupper (1/1)
työpaikat (2/2)
arbetefinska (1/1)
nattetid (1/1)
söderifrån (1/1)
vanligtvis (47/47)
vinster (1/1)
arbetsintygfinska (1/1)
allmänheten (2/2)
vetenskapsbibliotek (1/1)
finnas (10/10)
är (1322/1322)
ansökningstiderna (2/2)
planen (1/1)
förebyggande (6/6)
bekänna (1/1)
startpenning (5/5)
välsignas (1/1)
tillfällen (1/1)
åkrarna (1/1)
turist (2/2)
finansieringsandelar (1/1)
uppgjort (1/1)
underhålla (1/1)
företagskulturen (2/2)
föräldrarnafinska (1/1)
uppstår (5/5)
förbundet (2/3) Förbundet (1)
justitieministeriets (2/2)
verksamhet (40/40)
Brottsofferjourens (2/2)
noll (1/1)
barnfamiljerfinska (2/2)
operation (2/2)
kommunernafinska (2/2)
Vanttauskoski (1/1)
freelancer (1/1)
preparaten (1/1)
världen (2/2)
uppdateringen (1/1)
tillstånden (1/1)
tvungen (8/8)
egenskaper (1/1)
hallitus (1/1)
tryggt (5/5)
förbrukning (3/3)
frivilliga (4/4)
dessutom (25/25)
regionkontorfinska (1/1)
finansierar (1/1)
identitetsnummer (1/1)
förfaller (2/2)
innehas (2/2)
legalisering (2/2)
vilka (37/37)
fortbildning (5/5)
ett (963/965) Ett (2)
kartong (1/1)
studielinjer (1/1)
bokhandlar (1/1)
ansökning (5/5)
kiosker (4/4)
Utbildningsstyrelsen (3/3)
mitt (9/9)
inreseförbud (2/2)
kommersiellt (1/1)
barnens (7/7)
viga (1/1)
metspö (3/3)
giftermål (1/1)
fågelungar (2/2)
verkets (1/1)
fulla (1/1)
driver (3/3)
säljer (9/9)
ammatti- (3/3)
kvinnorna (3/3)
arvolaki (1/1)
närståendevårdare (1/1)
säljaren (7/7)
specialyrkesläroanstalter (1/1)
kränker (1/1)
självstyre (2/2)
allmäneuropeisk (1/1)
nationellt (1/1)
flyga (1/1)
bostadsägaren (2/2)
yrkesinstitutet (1/1)
Genève- (2/2)
sannolikt (2/2)
länkarna (2/2)
avlidit (1/1)
utbildats (1/1)
bistå (2/2)
bostadsrättsbostaden (1/1)
republikens (1/1)
makar (2/2)
lagarna (5/5)
arvsskattfinska (1/1)
koulu (2/2)
straffa (1/1)
säkerställer (1/1)
hen (28/28)
yrkesutbildningfinska (4/4)
insamlat (2/2)
betraktas (5/5)
bibliotekskunderna (1/1)
akut (22/22)
livmoderns (1/1)
grammatikengelska (1/1)
bankonto (1/1)
Sodankylä (1/1)
medeltemperaturen (1/1)
ingripa (3/3)
skatteavdrag (1/1)
varhaiskasvatushakemus (1/1)
avled (1/1)
nättjänsterna (2/2)
alakoulu (1/1)
utkomstskydd (9/11) Utkomstskydd (2)
uppskattar (4/4)
kedja (1/1)
ljusa (1/1)
stugan (1/1)
samlaget (1/1)
centret (5/5)
faderskapspenningdagar (4/4)
säkerhets- (1/1)
åka (5/5)
social- (26/26)
lämnat (3/3)
Familjeledighet (2/4) familjeledighet (2)
levnadskostnaderna (1/1)
handlingarna (3/3)
heminkvartering (1/1)
kreditupplysningsregistret (2/2)
närbibliotek (1/1)
tidsbokningen (5/5)
videoklipp (3/3)
servicevägledning (1/1)
bedöms (7/7)
nås (2/2)
sträckte (1/1)
utbetalning (4/4)
organisera (1/1)
Soldatskär (1/1)
skyddshemmet (5/5)
förvärvsarbeta (3/3)
betalats (3/3)
handlar (2/2)
fritid (4/5) Fritid (1)
lantdag (1/1)
Haartmanska (4/4)
verksamhetsprogram (1/1)
företedde (1/1)
kranen (1/1)
Oodi (2/2)
valdagen (8/8)
tempus (1/1)
magistraten (87/88) Magistraten (1)
företags (1/1)
eija.kyllonen (1/1)
juli (7/7)
hälsa (63/69) Hälsa (6)
utförande (1/1)
arbetsvillkoret (2/2)
myndig (5/5)
bidra (2/2)
mamma- (1/1)
festivalerfinska (1/1)
anordnar (1/1)
stödboende (3/3)
företagshälsovården (7/8) Företagshälsovården (1)
turvakoti (4/6) Turvakoti (2)
hänvisa (1/1)
förbjuda (1/1)
-stiftelser (1/1)
yrkesutbildning (35/36) Yrkesutbildning (1)
invandrarmän (3/3)
fått (44/44)
nationalpark (2/2)
universitetssjukhus (2/2)
omänsklig (1/1)
samtliga (11/11)
arbetskulturen (5/5)
samfällighets (3/3)
handikappservice (2/2)
vintrarna (1/1)
slutit (1/1)
långvarig (3/3)
åringar (5/5)
undersökningar (4/4)
bibliotekstjänstfinska (1/1)
intressebevakare (1/1)
plastkasse (2/2)
produktionsmedel (2/2)
prioriteten (1/1)
genom (47/47)
tvingas (5/5)
ändamål (1/1)
röst (3/3)
Omatila (4/4)
lånet (7/7)
väderleksrapporterna (1/1)
lågstadiet (2/2)
Rovaniemen (2/2)
midsommareldar (1/1)
mallarfinska (1/1)
belastad (1/1)
emellan (1/1)
avgift (2/2)
där (110/110)
bostadsförmedlingar (1/1)
utreder (10/10)
upplagan (1/1)
arbets- (58/59) Arbets- (1)
utvecklat (1/1)
säljs (6/6)
drivs (5/5)
reservationsavgifter (1/1)
ekonomi (4/4)
tapaturmavakuutus (1/1)
terapin (2/2)
upphört (6/6)
repertoar (1/1)
töms (1/1)
rättvist (3/3)
avdrag (5/5)
visumets (1/1)
församlingar (10/10)
kurator (1/1)
grad (1/1)
europeiska (11/18) Europeiska (7)
begär (2/2)
tillhandahåller (19/19)
sak (5/5)
oavslutad (1/1)
fakturera (2/2)
integritetsskydd (1/1)
Pyhäjoki (1/1)
förlossningssjukhuset (2/2)
rutterna (1/1)
leksaker (2/2)
könssjukdom (3/3)
inkomster (34/34)
yngsta (2/2)
serbiska (1/1)
självständiga (3/3)
magisterprogram (4/4)
insikt (1/1)
rester (1/1)
framskrida (1/1)
landets (6/6)
EU:s (2/2)
jämställdhetsombudsmannen (3/3)
cookies (1/1)
konkurrenter (1/1)
bostadsrättsbostadfinska (1/1)
videoklippet (12/12)
husets (8/8)
islam (1/1)
marker (1/1)
insjöar (1/1)
asylprocessen (1/1)
yläkoulu (1/1)
kostnader (9/9)
Avfallshantering (3/4) avfallshantering (1)
bedrivs (1/1)
markområden (1/1)
skolhälsovårdenfinska (1/1)
nyttiga (2/2)
servicepunkt (1/1)
ingås (5/5)
internetsidor (1/1)
blanketten (18/18)
ni (42/42)
ryssarna (1/1)
biljetter (2/2)
tidigare (21/21)
giltiga (2/2)
insjuknandet (4/4)
hälsostationerna (10/10)
synagoga (1/1)
siktar (1/1)
inbringar (2/2)
centralernafinska (1/1)
gravkontor (1/1)
drogbruk (1/1)
elva (3/3)
utkomstskyddet (4/4)
perheasioiden (2/2)
faderns (4/4)
norra (2/2)
Abfinska (1/1)
innebära (1/1)
minderåriga (7/7)
en (1442/1442)
sovittelu (2/2)
liten (11/11)
medelhög (1/1)
girering (1/1)
demonstrationer (1/1)
magistratfinska (1/1)
Asianajajaliitto (1/1)
lägga (5/5)
vård (57/57)
karttjänstfinska (1/1)
översättare (4/4)
lekparker (3/3)
ekonomibranschen (2/2)
två (97/97)
Väestörekisterikeskus (1/1)
disponenten (3/3)
förflyttningstillstånd (1/1)
fre (22/22)
midsommaren (1/1)
utkomststödfinska (1/1)
bostadsrätten (2/2)
vårdande (1/1)
pensionsärenden (1/1)
bort (4/4)
daghemsdagen (1/1)
yrkeshögskolanfinska (2/2)
sammanhängande (1/1)
aktörer (1/1)
oppilaitos (1/1)
stadissa.fi (2/2)
familjeförhållande (1/1)
kunskapscentret (1/1)
religion (31/31)
belägen (1/1)
tillställning (1/1)
skillnad (1/1)
dagtid (3/3)
ansökningar (4/4)
palveluasuminen (1/1)
Business (5/5)
bereda (1/1)
persiska (25/25)
skolhälsovården (2/2)
trupper (1/1)
inkomstbeskattningfinska (1/1)
bo (55/55)
Schengenvisumfinska (1/1)
bistår (2/2)
skattepengar (1/1)
sitt (53/53)
källan (1/1)
läkarremiss (2/2)
hyrt (1/1)
avvisas (1/1)
ålderspensionsålder (1/1)
ägo (1/1)
representera (1/1)
skåp (1/1)
prepaid (2/2)
landsomfattande (1/1)
Fulbright (2/2)
binder (2/2)
sjöstad (1/1)
naturstigar (1/1)
utmärkta (1/1)
webbläsarinställningar (1/1)
längd (3/3)
målarfärg (1/1)
tolk (40/40)
Alkoholister (2/3) alkoholister (1)
spel (4/4)
flaggdagarna (1/1)
tillbringa (1/1)
Ristin (2/2)
delas (15/15)
trygghet (13/13)
mall (1/1)
kielikahvila (1/1)
spelande (3/3)
uppehållskortet (3/3)
överföringen (1/1)
museidagen (1/1)
tolkförbund (2/2)
Omena (4/4)
Museiverkets (2/2)
bastulaven (1/1)
turneringar (1/1)
Schengenländerna (1/1)
behöva (6/6)
svenskspråkigt (4/4)
Resultatenheten (1/1)
industrin (1/1)
överbefälhavare (1/1)
Jourhjälpen (1/1)
ulkomaalaisten (1/1)
dari (2/2)
växel (1/1)
uppfylls (4/4)
härsken (1/1)
socialt (1/1)
äktenskapet (29/29)
pedagogiska (3/3)
-lokaler (1/1)
miljon (1/1)
densamma (1/1)
II (1/1)
besiktigas (1/1)
fjärde (13/13)
kulturer (6/6)
informationen (6/6)
stiftelsen (2/2)
Schengen (1/1)
familjefrågorfinska (2/2)
vuokrasopimus (1/1)
bank (4/5) Bank (1)
registrerats (3/3)
omhändertas (1/1)
över (82/82)
näringsbyrå (14/14)
fötts (3/3)
brottsmål (1/1)
pdf (25/26) PDF (1)
central (2/2)
återkallas (6/6)
Internetuppkoppling (1/1)
slutbetyget (1/1)
beskattningen (24/24)
anslutet (2/2)
Nordea (1/1)
förmedlingsarvodet (3/3)
försäkringsintyg (1/1)
Simundervisnings- (1/1)
allmänbildande (3/3)
FöPL (1/1)
lääkäri (2/2)
böjs (2/2)
Kannus (1/1)
avlider (4/4)
garanterar (1/1)
hälsomyndighet (1/1)
pappaledig (1/1)
längs (1/1)
medborgarinstitut (8/8)
befolkningsregistret (5/5)
konventioner (1/1)
tidigast (2/2)
fyll (4/4)
tekniska (1/1)
människorna (3/3)
sjukförsäkrad (2/2)
flickor (5/5)
utan (101/101)
näringsbyråns (9/9)
högtidligt (1/1)
branschen (2/2)
halt (2/2)
statsministern (2/2)
beslut (47/47)
riskabelt (1/1)
byarna (1/1)
taxa (1/1)
utvecklingsstadium (1/1)
preventionen (1/1)
avancemang (2/2)
skadad (1/1)
utnyttjande (1/1)
vägande (5/5)
byggas (1/1)
brottmålet (1/1)
serviceboendefinska (1/1)
diskuteras (1/1)
teaterstad (1/1)
utifrån (10/10)
anmälas (5/5)
yrkeshögskola (18/18)
tänkande (1/1)
Konvaljvägen (1/1)
verkar (2/2)
avgiftsfria (8/8)
låna (10/10)
anlänt (2/2)
trafik- (1/1)
lektioner (2/2)
specialtillstånd (1/1)
hyresbostäderengelska (1/1)
preliminär (1/1)
länders (5/5)
inhemsk (1/1)
Versofinska (1/1)
vigseltiden (1/1)
km (1/1)
startsida (1/1)
skiljasfinska (1/1)
skogsindustrin (1/1)
brutit (2/2)
såväl (5/5)
Centria (1/1)
befinner (5/5)
samlas (3/3)
samtidigt (25/25)
Kronoby (1/1)
arbetspensionssystemet (1/1)
körkortfinska (1/1)
Norden (1/1)
beslutsfattarna (1/1)
förhandlare (1/1)
hurdana (6/6)
marknaden (1/1)
tjeckiska (1/1)
vårdåtgärder (1/1)
undersöka (1/1)
sommar- (1/1)
ansökte (2/2)
Australien (1/1)
per (60/60)
mentor (2/2)
Optia (1/1)
religioner (3/4) Religioner (1)
lisensiaatti (1/1)
hälsovårdstjänster (23/26) Hälsovårdstjänster (3)
storlek (16/16)
middag (1/1)
konstaterar (1/1)
raskauden (1/1)
återvinning (6/6)
premier (1/1)
sådant (16/16)
Skatteförvaltningens (9/12) skatteförvaltningens (3)
sosiaali- (4/6) Sosiaali- (2)
slutföra (1/1)
resurscenter (1/1)
reparation (1/1)
kirkko (2/2)
tillfrågad (1/1)
pappersblanketter (1/1)
motions- (1/1)
efterlevandes (1/1)
Ullava (3/3)
åldern (11/11)
vederbörligt (1/1)
avgörs (1/1)
roll (2/2)
boendeträffpunkter (1/1)
kartläggningar (1/1)
ängre (1/1)
skärgårdenfinska (1/1)
säker (5/5)
företagsformen (3/3)
Oulun (1/1)
kronologisk (2/2)
medicinskt (1/1)
työntekijä (1/1)
noggrann (2/2)
utkomststöd (18/18)
stanna (10/10)
förvaltningsdomstolen (5/5)
självständighetsdagen (1/1)
kosthålls- (2/2)
rundvandringarna (1/1)
grundskolebaserad (4/4)
eläke (1/1)
datorn (1/1)
kontot (1/1)
Celia (1/1)
garantipensionens (1/1)
utarbetats (1/1)
familjecentret (4/4)
enskilde (1/1)
biografer (3/3)
webbtjänsten (7/7)
resekostnaderna (2/2)
hon (47/47)
eleven (2/2)
varifrån (1/1)
gälla (2/2)
brand (9/9)
perheneuvonta (1/1)
färdtjänsten (1/1)
låg (1/1)
steg (5/5)
lite (11/11)
elarbeten (1/1)
närstående (20/20)
arbetsinkomster (2/2)
ansöks (4/4)
spalt (1/1)
registreras (20/20)
förvaltningen (2/2)
fackets (1/1)
situation (31/31)
utbildningskoncern (1/1)
skulder (10/10)
bibliotekarien (2/2)
sammanfattning (3/3)
skickas (8/8)
anställningsoptioner (1/1)
största (16/16)
delen (10/10)
begår (4/4)
olycksfall (5/5)
konfessionslösa (2/2)
flest (2/2)
åriga (10/10)
ortodoxa (13/13)
asylprocessens (1/1)
högskoleexamen (18/18)
gymnasie- (1/1)
itsehoitolääke (1/1)
meddelar (4/4)
d.v.s. (14/14)
bostadsaktiebolaget (6/6)
begravningfinska (1/1)
telefonrådgivning (3/3)
länderfinska (1/1)
öppna (55/55)
avsett (10/10)
busstidtabellerna (1/1)
fakulteten (1/1)
socialarbetaren (2/2)
bioprogram (1/1)
flyttgodsfinska (1/1)
orterna (1/1)
närliggande (2/2)
problem (83/90) Problem (7)
bibliotekskort (7/7)
rådgivningen (23/23)
studierfinska (2/2)
ungdomsgård (2/2)
skoldagarna (1/1)
företagsformer (2/3) Företagsformer (1)
tjänste- (1/1)
metalli (1/1)
sagotimmar (1/1)
oljemängden (1/1)
ensamstående (3/3)
anställningsförhållande (1/1)
användande (1/1)
Köpcentret (1/1)
kvällarna (1/1)
drogmissbruk (1/1)
kansli (7/7)
inriktningar (1/1)
Migrationsverkets (27/27)
bestämda (1/1)
tittar (1/1)
Rysslands (2/2)
råkar (7/7)
framgå (3/3)
summa (4/4)
bekräftas (1/1)
vaccineras (1/1)
mottagit (1/1)
minipiller (1/1)
stärka (1/1)
gör (30/30)
kallt (3/3)
specialiserade (1/1)
turism (4/4)
bostadsrådgivning (1/1)
centralerna (1/1)
tidskrifter (3/3)
VR:s (2/2)
omsorg (2/2)
studiemiljö (2/2)
ändrade (1/1)
sökandens (2/2)
somliga (1/1)
webbläsare (1/1)
romerna (1/1)
genast (9/9)
din (511/511)
mottagningscenter (1/1)
inlärningssvårigheter (1/1)
försörjer (1/1)
utflykter (6/6)
startandet (1/1)
insulin (1/1)
ansvar (8/8)
löneanspråk (1/1)
skjuta (1/1)
matkulturer (1/1)
bör (18/18)
Kylämaja (1/1)
hälsorådgivningen (2/2)
uppdragsavtal (2/2)
tips (3/3)
piller (2/2)
arbetsliv (1/1)
möjliga (1/1)
pensionärsrabatten (1/1)
utgångstid (1/1)
änkling (2/2)
samboförhållandet (6/6)
sysslor (1/1)
RIKU (1/1)
januari (12/12)
utgöra (4/4)
uppehållstillståndskortet (1/1)
assistent (1/1)
fördjupa (1/1)
uppehållstillståndsärenden (1/1)
startpeng (5/5)
planerar (10/10)
preparat (1/1)
erbjuder (79/79)
högskolorna (7/7)
gränserna (2/2)
poliisi (1/1)
arbetslöshet (2/2)
faktum (1/1)
höra (5/5)
café (1/1)
Herman (1/1)
pysyvä (1/1)
ungdomsledare (1/1)
fadernfinska (1/1)
försenad (2/2)
specialdagvård (1/1)
simhallen (1/1)
gruppmöten (1/1)
fackevenemang (1/1)
yrkesbevis (1/1)
utexamineras (1/1)
högskolan (4/4)
kollektivtrafiken (4/4)
bestämmer (4/4)
lyfta (3/3)
studietid (1/1)
doulaverksamheten (1/1)
verklig (2/2)
kreditgivning (1/1)
parentes (1/1)
hamnverksamheten (1/1)
räntestödetfinska (1/1)
påbyggnadsutbildning (4/4)
läsas (2/2)
hemresan (2/2)
rekommendera (2/2)
telefonnumren (1/1)
revisionsbyrå (1/1)
ASE (7/7)
visumcentral (1/1)
förtjänade (1/1)
stipendier (4/4)
och (2619/2619)
studentmössor (1/1)
betalda (1/1)
dokument (4/4)
tillväxtföretagare (2/2)
bostadslånet (3/3)
försäljning (1/1)
arbetssäkerheten (2/2)
besökarna (1/1)
utöver (5/5)
brottsoffret (1/1)
telefonjouren (1/1)
kursutbudet (1/1)
kundtjänsten (7/7)
nödvändig (3/3)
Pro (3/3)
saknas (2/2)
servicenivån (1/1)
användningsdatumet (1/1)
hälsovårdsministeriet (3/3)
tala (14/14)
missbrukat (1/1)
rehabiliteringsplan (2/2)
naturhistoriska (1/1)
arvo (1/1)
konsertsalar (1/1)
mån.-tors. (1/1)
utbildningfinska (2/2)
sen (1/1)
arabisktalande (1/1)
Barnsjukhuset (2/3) barnsjukhuset (1)
följa (19/19)
lämningar (1/1)
samtycker (2/2)
riksdagenfinska (1/1)
föreslog (1/1)
ålderdom (1/1)
svenskan (2/2)
Barnskydd (1/1)
symtomen (1/1)
vardagsmotion (1/1)
förrätta (1/1)
självständig (2/2)
frilansarefinska (1/1)
vardags- (1/1)
uppehälle (5/5)
skolbarn (2/2)
skaffa (26/26)
företagarutbildningar (1/1)
bostadsansökan (3/3)
Korso (3/3)
lekverksamhet (1/1)
bussbiljetter (1/1)
yrket (1/1)
långtidssjuka (2/2)
internationalisering (1/1)
anställdafinska (1/1)
fri (1/1)
bedömning (6/6)
rf:s (3/3)
integritetsskyddet (1/1)
gjort (5/5)
firandet (1/1)
vigslar (2/2)
företett (1/1)
informellt (1/1)
vart (10/10)
privatläkare (4/4)
vuxengymnasier (2/2)
kostnadsfria (11/11)
arbetsoförmögen (2/2)
fart (1/1)
biologi (1/1)
försätts (1/1)
surfplatta (1/1)
EMMAfinska (1/1)
Ilmonet.fi (1/1)
ge (23/23)
valtion (1/1)
Eiran (1/1)
kartlägga (2/2)
trafikförsäkring (1/1)
lör (1/1)
fortbildar (1/1)
existensminimum (2/2)
yliopistollinen (1/1)
Bredvikens (1/1)
familjeplaneringfinska (2/2)
anses (10/10)
invandrarbyrå (2/2)
begäras (2/2)
inbördeskrig (1/1)
riktnummer (1/1)
arbetsintyg (12/14) Arbetsintyg (2)
komma (53/53)
tvätt- (1/1)
servicesedlar (1/1)
folkmängd (1/1)
bokföringsskyldighet (1/1)
utvecklingsstörda (3/3)
socialstationen (1/1)
straffas (1/1)
inresereglerna (1/1)
drogproblemfinska (1/1)
läder- (1/1)
bolag (6/6)
socialskyddsavtal (2/2)
ert (1/1)
folkpensionen (1/1)
föräldrarna (51/51)
felen (1/1)
institutfinska (1/1)
kommuntilläggfinska (1/1)
gruppfamiljedagvården (1/1)
näring (1/1)
sammankallas (1/1)
skattenumret (3/3)
ljusaste (1/1)
boendetfinska (1/1)
ledande (2/2)
receptbelagda (1/1)
högteknologisk (1/1)
informationsservice (1/1)
parförhållandet (14/14)
assistans (1/1)
barnskötare (3/3)
förorsakat (1/1)
besöka (35/35)
mödra- (8/8)
mån (16/16)
telefonservicefinska (1/1)
invandrarföreningar (3/3)
strävar (3/3)
Kompetenscentret (1/1)
gardet (1/1)
farliga (2/2)
förutsatt (1/1)
skapade (1/1)
arbetslöshetsförmån (7/7)
indoeuropeiska (1/1)
kopiera (2/2)
hjälpa (26/26)
skriva (16/16)
räntan (2/3) Räntan (1)
hyresdepositionen (3/3)
elpriserfinska (1/1)
löneperioden (1/1)
korta (4/4)
anställa (3/3)
distansgymnasiet (1/1)
FPA.I (1/1)
menar (1/1)
omedelbar (5/5)
arbetsmarknadsstödet (1/1)
bodelning (1/1)
självständighet (2/2)
betalat (10/10)
regel (7/7)
vikens (1/1)
längden (1/1)
företag (101/101)
storlekar (1/1)
verifierats (1/1)
permanent (17/17)
utbetald (1/1)
fattas (10/10)
statsborgen (1/1)
hänvisas (1/1)
tidsbokningssystem (1/1)
pass (23/23)
kanaler (5/5)
urologisk (1/1)
arbetslöshetsförsäkringen (2/2)
ursprung (12/12)
jakttillstånd (1/1)
bostadslån (7/7)
kontanter (5/5)
deltagarna (1/1)
funderar (5/5)
baserade (1/1)
era (2/2)
fritt (14/14)
Steinerskola (2/2)
blanketter (1/1)
responssystemfinska (1/1)
intressebevakning (1/1)
sökanden (3/3)
oroliga (1/1)
häva (2/2)
flygplatsen (1/1)
trots (6/6)
anspråkslös (1/1)
väntat (1/1)
byggherren (1/1)
förvärvar (1/1)
sköterskan (1/1)
miljöer (1/1)
inverkar (6/6)
sista (6/6)
Ryssland (9/9)
Olkkarifinska (1/1)
sökmotorer (1/1)
nytt (26/26)
uppenbart (1/1)
korrigera (1/1)
Institutet (2/3) institutet (1)
ry:s (2/2)
arbetskamraterna (1/1)
dubbade (1/1)
lunchpaus (1/1)
dag (27/27)
bekräfta (1/1)
idrottscentret (1/1)
flyktingar (14/14)
barns (19/23) Barns (4)
fisketillstånd (3/3)
personförsäkring (1/1)
tecknat (1/1)
bondgård (1/1)
sjukdomsfall (1/1)
tryggheten (61/61)
Norge (7/7)
motionsdosen (1/1)
ingen (22/22)
invandrat (2/2)
hedersrelaterade (2/2)
släktning (1/1)
öppnar (11/11)
internet (40/61) Internet (21)
bodelningsman (2/2)
samtalar (3/3)
sjunga (2/2)
passfoto (2/2)
Domus (1/1)
nöjd (1/1)
avlönat (1/1)
förbjudet (2/2)
kulturen (10/10)
utföra (9/9)
vin (1/1)
upphovsrätts- (1/1)
bank- (1/1)
hemifrån (2/2)
engelskspråkigt (1/1)
församlingen (1/1)
knappsatsen (1/1)
skuldrådgivningen (1/1)
InfoFinland (21/21)
industristad (1/1)
föreningarfinska (1/1)
damm (1/1)
Pejas (2/2)
samkommunens (1/1)
lokalförvaltningfinska (1/1)
skorna (1/1)
utgång (1/1)
A1.3 (1/1)
tills (16/16)
karensen (1/1)
exakt (2/2)
titta (5/5)
religionen (2/2)
äe (1/1)
systerdotter (1/1)
feber (1/1)
lönekvittona (1/1)
kl. (1/1)
sätta (1/1)
hyresbostäderfinska (5/5)
medling (6/6)
andelslag (6/6)
pilkning (1/1)
avvägs (1/1)
testamente (5/5)
förslossningsdatumet (1/1)
fastlagen (1/1)
Salutorget (1/1)
olycka (10/10)
värderingar (1/1)
flyktingorganisation (2/2)
Kehitysvammaliittos (1/1)
informering (1/1)
bildas (4/4)
lönen (16/16)
hammashoidon (3/3)
parförhållandets (1/1)
medborgare (138/139) Medborgare (1)
syfte (2/2)
vaccination (1/1)
västerut (1/1)
myndighetsärenden (1/1)
MinSkatt (3/3)
integritet (3/3)
Lahtis (1/1)
sökmotor (6/6)
parken (1/1)
förlossningsavdelningen (1/1)
berättar (9/9)
gå (36/36)
dagar (35/35)
anlita (14/14)
instrument (2/2)
hemkommun (104/114) Hemkommun (10)
anmäl (2/2)
anmälningsdagen (2/2)
hälsovårdsstiftelses (1/1)
idrottsmöjligheter (2/2)
butiken (1/1)
missbruksproblemfinska (2/2)
stiftelser (3/3)
Esbos (1/1)
bedömningar (1/1)
guidade (3/3)
bilskola (1/1)
helgerna (2/2)
samerna (1/1)
sjukförsäkring (8/8)
tyska (38/38)
blankett (15/15)
jordbruk (1/1)
lukiopohjainen (1/1)
Tavastehus (1/1)
webbplats (174/174)
filmvisningarfinska (1/1)
rättshjälpen (1/1)
jourmottagning (1/1)
uppskattning (2/2)
klimatet (1/2) Klimatet (1)
bemötts (1/1)
hyressed (1/1)
civilvigsel (1/1)
teatrarnas (2/2)
Virtanen (2/2)
finansiärerna (1/1)
arbetarinstitutens (1/1)
definierar (1/1)
reparationsarbeten (1/1)
överskridits (1/1)
direktör (1/1)
Hautaustoimistojen (1/1)
be (44/44)
misstänkt (1/1)
sörja (4/4)
staden (32/32)
nationalmuseum (1/1)
extra (4/4)
spisen (4/4)
aktier (2/2)
kurs (4/4)
socialtjänsterna (2/2)
pensionsåldern (1/1)
utsänd (1/1)
helsingforsare (1/1)
skolbarns (4/4)
demensfinska (1/1)
teckenspråk (3/3)
förrättas (14/14)
munsjukdomar (1/1)
talet (15/15)
semester (4/4)
Arctica (3/3)
livssituation (7/7)
större (13/13)
månatliga (1/1)
häradsskrivare (1/1)
sakkunniga (1/1)
arbetskontrakt (1/1)
fiskebyn (1/1)
underhållsbidraget (4/4)
eläkekassa (1/1)
men (71/71)
lägre (9/9)
leder (8/8)
RAOS (1/1)
intervjuerna (1/1)
numret (9/9)
prioriteras (2/2)
kriget (4/4)
utvecklingsidéer (1/1)
video (2/2)
postfinska (1/1)
pauserna (1/1)
HelsingforsHels (1/1)
märker (1/1)
besöksförbud (3/3)
kontaktspråk (1/1)
hygienen (1/1)
uhrien (1/1)
utbildningskoncernfinska (1/1)
fotografi (1/1)
insamlingsställen (1/1)
konflikterna (2/2)
regiontaxi (1/1)
medan (5/5)
kulturförening (1/1)
känns (1/1)
militärunderstöd (1/1)
adopterar (1/1)
lånord (1/1)
rättigheterfinska (1/1)
artigt (2/2)
källskatt (1/1)
vattenkran (1/1)
nätbankskoderna (1/1)
nationell (1/1)
kursavgiften (2/2)
studiekraven (1/1)
tätskikt (1/1)
sektorn (10/10)
ersättning (16/16)
rumänska (12/12)
vattenmätare (1/1)
barntillsynsmannen (1/1)
erbjuds (13/13)
åt (22/22)
personalen (5/5)
risker (2/2)
oroar (1/1)
förskoleundervisningfinska (3/3)
To (4/4)
förövaren (1/1)
caféer (1/1)
högst (37/37)
Ihmiskaupan (1/1)
lekparkerna (1/1)
parkeringsbiljetten (1/1)
bildkonstskolor (1/1)
teckna (9/9)
dubbelnamn (1/1)
nomineras (2/2)
RFV (1/1)
talas (8/8)
hyresvärd (2/2)
Vionoja (1/1)
Lastensuojelulaki (1/1)
vigselceremonin (1/1)
tälta (1/1)
höga (1/1)
misstänker (11/11)
förarexamen (1/1)
utbyten (1/1)
barnatillsynsmannen (1/1)
kränkande (1/1)
logi (1/1)
sjukvårdskostnader (2/2)
populäraste (1/1)
administrativa (2/2)
koulunkäyntiavustaja (1/1)
toleransen (1/1)
telefontid (1/1)
betalningsstörningfinska (1/1)
jämte (1/1)
vårdens (1/1)
biografens (1/1)
upplevt (1/1)
kostnaderna (15/15)
undantag (4/5) Undantag (1)
ingått (6/6)
läsa (16/16)
förskoleplats (4/4)
tolksbehovet (1/1)
samboskap (1/1)
telefontjänst (11/11)
krismottagningen (1/1)
intresse (4/4)
apparater (2/2)
företagarguider (1/1)
utförandet (5/5)
pappersblankett (5/5)
precis (2/2)
drogfritt (1/1)
förhandsröstningstiden (1/1)
autonoma (1/1)
slotten (2/2)
tandkliniken (3/3)
varar (20/20)
ungdomspsykiatriska (1/1)
rådgivningsbyrån (21/21)
arbetsavtal (8/8)
surfplattan (1/1)
appen (2/2)
förhållandena (1/1)
bouppteckningen (3/3)
klä (4/4)
karneval (1/1)
kontrolleras (3/3)
minoriteter (3/3)
slutarbete (2/2)
anhöriga (10/10)
myhelsinki.fi (1/1)
inslag.Om (1/1)
miljöministeriet (1/1)
kopplas (2/2)
delvis (10/10)
förebygga (1/1)
motorfordon (3/3)
informationfinska (1/1)
inkluderar (1/1)
hemvårdsstödet (3/3)
utgår (3/3)
lönenivån (1/1)
varmaste (1/1)
HIV (2/2)
julafton (2/2)
började (6/6)
användningen (6/6)
ryskspråkiga (1/1)
inkomsterna (6/6)
sorteringen (1/1)
försäljningen (4/4)
värnplikt (1/1)
rörelsehindradefinska (1/1)
moderskapsunderstöd (6/6)
Kokkola (2/2)
Korset (6/6)
sjunger (1/1)
delta (35/35)
sjukledighetsdagen (1/1)
skapandet (1/1)
Rovaniemifinska (2/2)
betalades (2/2)
jordbruks- (1/1)
ingrepp (1/1)
apoteken (1/1)
känner (12/12)
finskspråkig (3/3)
2:a (1/1)
idkar (1/1)
hälsostationsläkare (1/1)
långvarigt (1/1)
daghemsföreståndarna (2/2)
medeltida (1/1)
försvara (2/2)
Gloet (2/2)
Yrkenas (1/1)
kortti (2/2)
beskattningsärenden (1/1)
ängarna (1/1)
kollektivavtal (4/4)
trygg (5/5)
sopbehållare (1/1)
tillfällig (9/9)
anslöts (2/2)
förvaltning (1/1)
inredningsarkitekt (1/1)
hyreskontrakt (2/2)
läkemedelfinska (1/1)
kunnallisvaalit (1/1)
fönstret (1/1)
uppfyller (5/5)
affärsidé (1/1)
leverans- (1/1)
uppdragsgivare (1/1)
skriftligt (27/27)
förlossningsdatumet (3/3)
textning (1/1)
dra (3/3)
progressivt (1/1)
återbetalas (1/1)
Luetaan (1/1)
Akademi (1/1)
insjuknade (1/1)
förändringsarbeten (2/2)
beskattningsbara (3/3)
upprepade (1/1)
ärenden (58/58)
yta (1/1)
Företagarna (1/1)
överens (43/43)
medborgaren (1/1)
ämnena (1/1)
bostadssökande (1/1)
tog (3/3)
Banvägen (1/1)
biograf (2/2)
ehkäisyneuvola (1/1)
räcker (11/11)
bolagsvederlag (1/1)
skötseln (6/6)
Förenta (1/1)
kl (73/73)
familjemedlems (1/1)
samhällslivet (1/1)
familjepensionen (1/1)
inför (11/11)
särbehandlas (2/2)
industrialisering (1/1)
Apostille (1/1)
behovsprövat (2/2)
lämna (39/39)
fortsätta (8/8)
människogrupp (1/1)
Kaustarviken (1/1)
EK (2/3) Ek (1)
seurakuntien (1/1)
ifyllda (3/3)
förstå (2/2)
bosättningsort (1/1)
övervakar (10/10)
stilla (1/1)
databas (1/1)
situationerna (1/1)
Lapin (1/1)
dagliga (12/12)
värdefull (1/1)
livligare (1/1)
utbytesprogrammetengelska (1/1)
transportera (1/1)
badrumsrenovering (1/1)
registreringsintyg (2/2)
äger (11/11)
hjälper (63/63)
Tallinn (2/2)
skriver (11/11)
tingsrätten (9/9)
startade (1/1)
STTK (1/1)
inkassokostnader (1/1)
luterilainen (1/1)
bedömningsskalan (1/1)
ansökningsförfarandena (1/1)
föräldraledigheten (7/7)
föremål (2/2)
skolgången (2/2)
rasismi (1/1)
besöker (10/10)
viseringsskyldiga (1/1)
preventivrådgivning (1/1)
auktoriserad (1/1)
opintotuki (2/2)
miljön (3/3)
humanitärt (1/1)
människor (37/37)
insamlingsställe (1/1)
godkännas (1/1)
klart (1/1)
hushållfinska (1/1)
bostadslösa (5/5)
erkänns (1/1)
plötsliga (1/1)
listan (2/2)
enspråkiga (2/2)
sent (4/4)
framgångsrikt (1/1)
välityspalkkio (1/1)
sysselsättningsplan (4/4)
radhus (3/3)
oleskeluoikeuden (1/1)
betala (88/88)
livet (11/12) Livet (1)
underhyresgäst (3/3)
stödfunktioner (1/1)
lånetiden (1/1)
Tankkari (1/1)
Myrbackahuset (1/1)
referensramen (1/1)
lämplighetsprov (1/1)
skogsbruksområden (1/1)
bostäderfinska (2/2)
lärokurs (5/5)
sosiaalineuvonta (1/1)
föreningen (12/14) Föreningen (2)
inleds (8/8)
yrkeshögskolestudier (1/1)
ungafinska (8/8)
inkorporerades (1/1)
turism- (2/2)
lärare (4/4)
matka.fi (1/1)
far (9/9)
sexuell (5/5)
ökar (1/1)
matfinska (1/1)
glasögon (1/1)
var (48/56) Var (8)
barnlösheten (1/1)
delaktig (1/1)
ungdomsgården (2/3) Ungdomsgården (1)
hävs (1/1)
enkelt (2/2)
upprättar (3/3)
grupper (11/11)
linkkiFörsamlingen (1/1)
Dödsfall (1/1)
Opintopolku.fi (3/3)
betänketiden (5/5)
skattedeklarationen (6/6)
tonåringar (1/1)
länk (3/3)
lättläst (1/1)
utrymmen (1/1)
tjänsteleverantör (1/1)
Familjeledigheter (1/1)
nya (40/40)
Handikappforums (1/1)
unionenfinska (1/1)
minimilöner (4/4)
sökfunktionen (1/1)
hyresvärdar (5/5)
rutten (1/1)
studieplaner (1/1)
befann (1/1)
hyresgästen (4/4)
läroverket (1/1)
lö (1/1)
receptet (1/1)
hoppas (1/1)
annars (5/5)
ger (82/83) GER (1)
påsk (1/1)
asuntosäätiö (2/2)
ställs (5/5)
fortare (1/1)
grund (122/122)
grupplivförsäkring (1/1)
hit (1/1)
vräka (1/1)
aning (1/1)
arbetskraftsutbildningen (2/2)
varvid (1/1)
osuuskunta (1/1)
högtidlig (1/1)
bostadsrättsavtalet (1/1)
majoriteten (1/1)
Vvo (1/2) VVO (1)
uppförande (1/1)
antingen (35/35)
livscykel (1/1)
bosättningsland (1/1)
försöker (6/6)
musikhus (1/1)
hämtas (1/1)
sedan (11/11)
asylsökande (22/22)
ligger (22/22)
tingsrättfinska (2/2)
bostad (102/102)
huvudsak (3/3)
hemhjälp (1/1)
förväg (22/22)
Ristrand (1/1)
handikappat (8/8)
barnrådgivningens (1/1)
intjänade (3/3)
kielioppi (1/1)
perintövero (1/1)
Esbo (100/100)
kamratförening (1/1)
pappa (1/1)
samboende (1/1)
rättsskyddsförsäkring (1/1)
vigselförrättningen (1/1)
diabetes (2/2)
hänsyn (5/5)
försäljningsmetoder (1/1)
privata (45/45)
mångkulturella (6/6)
stängda (2/2)
månaders (5/5)
boendemöjligheter (1/1)
cycling (1/1)
skaffat (1/1)
stulits (1/1)
anhörigas (1/1)
nekande (1/1)
motionsslingorna (1/1)
byggnaderna (1/1)
webbplatserna (1/1)
fastställa (1/1)
tidningarna (1/1)
studiestödetengelska (1/1)
kommanditbolag (4/4)
till (1547/1553) Till (6)
tidsbokningfinska (1/1)
musik (18/18)
vidtar (1/1)
Alexandersgatan (1/1)
integrationsplanfinska (1/1)
Centralorganisation (1/1)
tidiga (3/3)
starta (17/17)
työeläkelaitokset (1/1)
tillverkas (2/2)
fick (12/12)
baserat (4/4)
magistratet (1/1)
lämnar (12/12)
hemmetfinska (1/1)
kurser (36/36)
köra (6/6)
apotekens (1/1)
skilda (1/1)
hörseln (1/1)
offentliga (56/56)
stämman (1/1)
vuxenutbildning (8/8)
dagvårdstjänster (2/2)
familjeverksamhet (1/1)
yrke (16/16)
problematiska (5/6) Problematiska (1)
flyttar (86/86)
vad (22/24) Vad (2)
varje (35/35)
produktionen (1/1)
medborgarorganisation (1/1)
h (1/1)
FIRMAXI (1/1)
statsöverhuvud (1/1)
brotten (1/1)
salar (1/1)
prövningfinska (2/2)
toalettstolen (1/1)
ibland (11/11)
C2 (1/1)
jämställdhet (12/14) Jämställdhet (2)
brandsläckaren (1/1)
Karleby (56/56)
Trafiksäkerhetsverkets (1/1)
styrgrupp (1/1)
dragits (1/1)
koulupsykologit (1/1)
arbetarskyddsföreskrifterna (2/2)
kärnkraftverket (3/3)
lunchsedlar (1/1)
mervärdesskatt (3/3)
ovanliga (1/1)
barn (315/319) Barn (4)
vattendrag (3/3)
myndigheterfinska (1/1)
studentkort (1/1)
DVD (1/1)
upphovsmannen (1/1)
hem (34/34)
mottagningen (5/5)
kommunvalfinska (1/1)
handeln (4/4)
avläggas (5/5)
skrivit (1/1)
språkcaféerna (2/2)
ökade (1/1)
relationsrådgivningstjänsterfinska (1/1)
Uunofinska (1/1)
idrottsanläggningarna (1/1)
bil (12/12)
användas (6/6)
tukiverkko (1/1)
muslimska (1/1)
penningbelopp (1/1)
lätt (5/5)
paluun (1/1)
vattenavgiften (3/3)
givet (1/1)
ositus (1/1)
kielitutkinto (3/3)
försäkringar (9/9)
skattebyråns (1/1)
självrisk (1/1)
fyrverkerier (1/1)
avancerad (1/1)
Muurola (1/1)
grannländer (2/2)
jobbsajterfinska (1/1)
Karlebynejden (1/1)
slutliga (3/3)
hitar (2/2)
tasa (2/3) Tasa (1)
hävas (2/2)
stärker (1/1)
kontaktspråket (1/1)
vuotiaan (1/1)
landsbygden (3/3)
misstänks (2/2)
förverkligas (3/3)
hälsovården (18/18)
uträttar (3/3)
företagande (12/12)
familjeförmåner (2/2)
orsak (7/7)
utvisad (1/1)
närarbetets (1/1)
besiktningsstationer (2/2)
invandrarkvinnor (10/10)
medborgarskapsanmälan (4/4)
sön (2/2)
äktenskapfinska (2/2)
museum (3/3)
deltar (6/6)
samarbetsområdet (1/1)
litet (6/6)
pakolainen (1/1)
allmänna (18/18)
ämnar (2/2)
samhörighet (1/1)
levereras (1/1)
Västerkulla (1/1)
resurser (2/2)
invandrareleverna (1/1)
Ruokavirasto (1/1)
euro (23/23)
byrån (54/54)
standardblanketter (1/1)
grenarna (1/1)
säsongsarbete (2/2)
folkpension (6/6)
spårvagnarna (1/1)
ut (113/113)
mobbad (1/1)
arbetslöshetskassan (6/6)
högklassig (1/1)
publicerades (1/1)
relationerna (3/3)
nordlig (1/1)
belagt (1/1)
Ammatilliseen (1/1)
mörkare (1/1)
som (1265/1266) Som (1)
vidaredistribuera (1/1)
settlementföreningen (1/1)
Rex (2/2)
rusmedelsberoende (1/1)
affärsmodell (1/1)
umgängetfinska (1/1)
hamnade (1/1)
början (16/16)
Vandakanalen (1/1)
nordiska (13/13)
halvt (1/1)
bosniska (2/2)
grannen (1/1)
beakta (7/7)
hjälptelefonen (2/2)
yrkesstudier (1/1)
stödperson (4/4)
kansalaisen (1/1)
sjukvårdsdistrikt (3/3)
pensionskassor (2/2)
seniorrådgivningen (4/5) Seniorrådgivningen (1)
at (3/3)
några (24/24)
hand (60/60)
kulturcenter (1/1)
vårdnadshavarna (2/2)
rättshjälpsbyrån (4/4)
studerandefinska (5/5)
tillståndet (17/17)
HNS (3/3)
löfte (1/1)
utarbetandet (1/1)
kvinnans (2/2)
Kalkkers (1/1)
auttamisjärjestelmä (1/1)
kallade (3/3)
går (43/43)
registrerar (7/7)
psykoterapeut (1/1)
skolelevers (1/1)
sådan (9/9)
ord (4/4)
funktionalitet (1/1)
engångskaraktär (1/1)
anor (1/1)
kunskapscenter (1/1)
behandlas (28/28)
friluftsliv (4/4)
skolkuratorn (2/2)
lapsilisä (1/1)
genomgått (1/1)
familjeförmånerna (1/1)
digital- (1/1)
säkerheten (3/3)
utrikespolitik (1/1)
aldrig (2/2)
förskolanfinska (1/1)
krisjourenfinska (2/2)
husbolaget (2/2)
Ajovarmas (2/2)
Lichtenstein (1/1)
arbetsinkomsten (1/1)
ber (1/1)
höghus (10/10)
byggplats (1/1)
riksväg (1/1)
just (4/4)
denna (22/23) Denna (1)
patientförening (1/1)
skala (1/1)
hemvårdsstöd (13/13)
statsstöd (1/1)
använda (79/79)
sälj (1/1)
volym (1/1)
universitetscenter (1/1)
hel.fi (2/2)
USA (4/4)
skolämnen (1/1)
Inre (4/4)
avlägga (56/56)
konto (13/13)
elektroniskt (11/11)
böckerna (1/1)
skydd (12/12)
Österbotten (2/2)
YTHS (1/1)
ungdom (1/1)
tillsvidareanställning (1/1)
föreningsmedlemmar (1/1)
fullsatta (1/1)
förekommer (2/2)
sämre (3/3)
treårigt (2/2)
biografkedjan (1/1)
ändringsarbeten (2/2)
material (13/13)
tidsbokning (11/11)
anställningsavtalets (1/1)
förening (9/9)
därifrån (1/1)
muntligt (2/2)
säkert (3/3)
bidragen (1/1)
lärokursen (2/2)
motionshobbyer (1/1)
Inkomstregistret (1/1)
vet (6/6)
startande (1/1)
skyldigheter (23/23)
kallelse (1/1)
bevisar (2/2)
uppsägningstid (2/2)
eleverna (5/5)
tolkningsspråket (1/1)
skyddshus (10/10)
nätverk (9/9)
september (3/3)
ordnas (81/81)
Anon (1/1)
vuxen (5/5)
pimpla (2/2)
barnet (160/160)
översatt (2/2)
arbetslöshetsersättning (10/10)
jaga (1/1)
privatvårdsstöd (2/2)
familjerådgivningfinska (1/1)
livförsäkring (1/1)
testamentsgåva (1/1)
nycklarna (1/1)
vidimeras (1/1)
expertråd (1/1)
Mielenterveysseura (3/3)
social (12/12)
bästa (11/11)
änka (2/2)
kontakta (116/116)
nättjänst (1/1)
köptjänst (1/1)
fyllt (29/29)
inga (9/9)
friluftsmuseum (1/1)
ogiltigt (1/1)
skolgång (4/4)
syrjintä (1/1)
mobiltelefontillverkaren (1/1)
arbetarskydd (2/3) Arbetarskydd (1)
god (11/12) God (1)
infopankki (1/1)
bostadsform (1/1)
käpp (1/1)
redogörs (1/1)
domstolen (4/4)
myndigheter (35/35)
enskilda (6/6)
slidan (1/1)
använts (2/2)
klädregler (1/1)
tolktjänster (5/5)
Estnäs (1/1)
inkvartering (2/2)
työsuojelun (1/1)
medborgarskapsansökan (2/2)
utformas (1/1)
vinnare (2/2)
gymnasium (13/14) Gymnasium (1)
socialmyndigheters (1/1)
motionsevenemang (1/1)
integrationsåtgärderna (1/1)
händer (2/2)
bankärendenfinska (1/1)
ministrarna (1/1)
åtalas (1/1)
regiontrafiken (1/1)
förorter (1/1)
täydennyskoulutus (1/1)
strax (1/1)
allmäneuropeiskt (1/1)
bostadsbidraget (3/3)
eget (62/62)
datumet (2/2)
lånat (1/1)
hyresgästenfinska (1/1)
musikinstitutet (1/1)
antagning (1/1)
sällskapar (1/1)
regelbundna (3/3)
visumfritt (2/2)
nödvändigt (4/4)
bilagorna (4/4)
arbetspensionsutdragfinska (1/1)
huvudsakligen (2/2)
grädde (1/1)
grundutbildning (2/2)
hoidon (1/1)
länderna (18/18)
pojkvän (1/1)
upphovsmannens (1/1)
affärer (1/1)
kvinnan (5/5)
intagen (1/1)
bokföringen (6/6)
Liikenteen (1/1)
förlorat (1/1)
fortsättningskriget (1/1)
otrogenhet (1/1)
Indien (1/1)
tvåspråkiga (4/4)
förföljd (2/2)
elevverksamhet (1/1)
förhöjd (1/1)
parets (1/1)
väder (1/1)
progressiv (4/4)
upprätthåll (1/1)
asylsökandefinska (2/2)
lönsamheten (1/1)
ohälsa (1/1)
utbetalningen (2/2)
arbetsmarknadsstöd (4/4)
slott (4/4)
kompetens (3/3)
röster (2/2)
affärsmannen (1/1)
Miehen (6/6)
yrken (11/11)
oktober (2/2)
mannens (1/1)
Punaisen (2/2)
trädgårdsskötsel (1/1)
handläggning (1/1)
Kiinteistöyhtiö (1/1)
hemma (39/39)
utgående (8/8)
borealis (1/1)
konfidentiella (2/2)
församlingssammansutning (1/1)
webblanketten (1/1)
dött (2/2)
föräldrar (37/37)
hälsorisk (1/1)
förbereder (3/3)
tillfoga (2/2)
kommandiittiyhtiö (1/1)
grenförbunden (1/1)
behöver (266/270) Behöver (4)
utvecklas (2/2)
uppstod (1/1)
lähdevero (1/1)
mera (5/5)
metron (2/2)
yrkesbeteckning (1/1)
regnar (1/1)
bemötande (3/3)
förändring (1/1)
acceptansen (1/1)
beaktande (2/2)
vistas (35/35)
gynekolog (4/4)
vakuus (1/1)
maximitiden (1/1)
dammsugaren (1/1)
slutexamen (1/1)
vuxenutbildningsinstitut (4/4)
studiematerial (1/1)
invånarlokalen (1/1)
grekiska (2/2)
barnpassning (1/1)
utfärdat (1/1)
medicinsk (13/13)
öppning (1/1)
specialfall (1/1)
inom (99/99)
lastensuojelu (1/1)
tilläggsstudier (1/1)
tillfälligt (21/22) Tillfälligt (1)
marknadsföring (1/1)
minnesproblemen (1/1)
ansökningsblanketter (2/2)
förhand (19/19)
sjukvårdskort (1/1)
bereder (2/2)
lämpliga (2/2)
TE (73/74) te (1)
bestyren (1/1)
jämlikt (4/4)
innehållet (4/7) Innehållet (3)
alkoholism (1/1)
beskattningsrätt (1/1)
ansikte (2/2)
faderskapspenning (3/3)
billigast (1/1)
byrå (17/17)
vilken (39/39)
arbetarinstitutet (1/1)
pensionering (1/1)
kotoutumissuunnitelma (1/1)
närskolan (2/2)
portfölj (1/1)
Karlebynejdens (2/2)
baltiska (1/1)
tillräckligt (25/25)
skolpsykologerna (1/1)
språkkunskaper (27/28) Språkkunskaper (1)
väntar (6/6)
IB (1/1)
förtrogen (1/1)
valomgången (3/3)
utlänningars (1/1)
förklarade (1/1)
livsåskådningskunskap (2/2)
mentala (12/12)
välbefinnandeområden (1/1)
gav (2/2)
Sport (5/7) sport (2)
tidsperioder (1/1)
Hörselförbundetfinska (1/1)
intressebevakningsorganisationer (1/1)
servicebolag (1/1)
lyckades (2/2)
rekisterihallitus (1/1)
månader (71/71)
arbetarskyddsfrågor (1/1)
MERCURIA (1/1)
härkomst (4/4)
osasairauspäiväraha (1/1)
karriären (1/1)
upphörde (1/1)
neuvontapalvelu (1/1)
kista (1/1)
terveysasema (13/13)
Easyfinnishfinska (1/1)
integrationsplanen (9/9)
ammattiopisto (4/4)
plågor (1/1)
högerextrema (1/1)
webbankkoder (4/4)
avdragsgill (2/2)
återförening (1/1)
Kemi (1/2) kemi (1)
invandrare (86/86)
närståendevård (6/6)
kommunalval (9/9)
akutpreventivmedel (1/1)
kristna (3/3)
Danske (1/1)
effektiva (1/1)
bestraffas (1/1)
inträffat (2/2)
hälsovårdenfinska (1/1)
riskfaktorer (1/1)
förlossningsavdelning (1/1)
överinspektören (1/1)
initiala (2/2)
ur (8/8)
lähityön (1/1)
Patentti- (1/1)
pågår (16/16)
yrkeskvalifikationer (1/1)
översättningstjänsterfinska (1/1)
regeringen (2/2)
kollegor (3/3)
personal (2/2)
ylioppilaskokeet (1/1)
CV (13/13)
tvättstuga (2/2)
fira (1/1)
tåg (3/3)
eller (1301/1301)
neuvola (4/4)
jobbar (1/1)
århundradet (1/1)
arbetarskyddsinspektioner (1/1)
förbindelse (2/2)
utställningarfinska (1/1)
hälsotillstånd (7/7)
skrivfärdigheter (1/1)
gravplats (1/1)
ogift (3/3)
Karlebys (2/2)
asiointipiste (1/1)
strategier (1/1)
bebott (3/3)
utlandsprefix (1/1)
förhindra (1/1)
konkret (1/1)
studerar (21/21)
motionstjänsternafinska (1/1)
tfn (16/17) Tfn (1)
etälukio (1/1)
språkexaminafinska (4/4)
FIRST (1/1)
servicestyrcentral (1/1)
det (475/476) Det (1)
investerare (1/1)
brann (1/1)
bidragens (1/1)
studiepenning (2/2)
förenings (1/1)
kemikaler (1/1)
invandrarförening (1/1)
springa (1/1)
utrustningen (2/2)
dans (6/6)
stunder (1/1)
rättsbiträde (3/3)
tidsbundet (7/7)
havsvik (1/1)
Foreigners (2/2)
elevernas (3/3)
utreda (5/5)
stiger (4/4)
välfärds- (1/1)
faderskapserkännande (1/1)
gym (3/3)
sjukhuset (17/17)
säkerhet (11/11)
registrerades (2/2)
banker (3/3)
eduskunta (2/2)
ungdomsväsendet (1/1)
arbetsavtalfinska (1/1)
Nivavaara (1/1)
centraler (1/1)
varit (22/22)
bussbolag (1/1)
integrationsprocessen (1/1)
grundas (3/3)
Soites (4/4)
Europaparlamentsval (4/4)
inget (21/21)
försäkringen (4/4)
Wilma (6/6)
svårigheter (3/3)
mottagningar (2/2)
ekonomiplaneringen (1/1)
finansieringsvederlag (1/1)
villkor (18/18)
bekostar (1/1)
depression (2/2)
krigsskadeståndet (1/1)
saker (27/27)
turvapaikkapuhuttelu (1/1)
tvärvetenskapliga (1/1)
jämkning (1/1)
information (337/342) Information (5)
kräva (10/10)
ställena (1/1)
ungefär (16/16)
identifieras (1/1)
jobba (2/2)
ons. (1/1)
vårens (1/1)
samjour (1/1)
kemikalier (2/2)
beräkning (1/1)
svenskafinska (2/2)
begåtts (2/2)
överenskommelse (3/3)
själva (12/12)
inkomstrelaterad (9/9)
ägare (6/6)
nuvarande (7/7)
bostadsrättsbostad (10/11) Bostadsrättsbostad (1)
Turku (1/1)
avses (16/16)
Advokatförbund (1/2) advokatförbund (1)
Kors (9/11) kors (2)
beskattning (6/10) Beskattning (4)
minimikraven (1/1)
på (1686/1687) På (1)
terrängen (1/1)
barnrådgivning (1/1)
80:e (1/1)
prov (6/6)
fiska (2/2)
fordonfinska (1/1)
lånas (1/1)
synskadades (1/1)
fyller (17/17)
taket (1/1)
vårdnaden (8/8)
grunden (5/5)
positiva (1/1)
tycker (1/1)
vidimera (1/1)
fastställts (5/5)
påbörjas (2/2)
undervisningstjänster (2/2)
besökare (1/1)
dagpenning (13/13)
spelberoende (3/3)
accepterade (1/1)
betalningsanmärkning (2/2)
tänker (2/2)
bor (84/84)
ställning (9/9)
riktad (1/1)
rättigheter (40/41) Rättigheter (1)
yrkesvägledning (1/1)
bostadsaktie (2/2)
upphör (18/18)
efternamn (48/48)
välmående (3/3)
trafik (3/3)
maahanmuuttajapalvelut (1/1)
brott (48/50) Brott (2)
ungdomarnas (2/2)
Noux (1/1)
avtog (1/1)
kvarskatten (1/1)
krig (4/4)
dess (18/18)
fullgjort (1/1)
frånskild (1/1)
släkting (6/6)
kollaps (1/1)
hälsocentralläkarens (1/1)
egnahemshus (5/5)
umgås (1/1)
vattenledningar (2/2)
hyr (8/8)
gonorré (1/1)
född (1/1)
bredvid (1/1)
psykologi (1/1)
klagar (1/1)
förstörs (2/2)
integrera (2/2)
infektion (1/1)
myndighets (1/1)
Helsingforsbor (1/1)
fött (3/3)
talen (2/2)
år (260/260)
påbrå (1/1)
väg (2/2)
könssjukdomarfinska (1/1)
engelska (783/783)
oppisopimus (1/1)
korrigerande (1/1)
jourmottagningarna (1/1)
klinikka (3/3)
linkkiFörbundet (1/1)
företagstjänsterna (1/1)
ännu (10/10)
dagstidningar (2/2)
utfärdad (1/1)
onyktert (1/1)
hobbyer (4/4)
yrkessjukdom (1/1)
ordentlig (2/2)
biograferna (1/1)
kärren (1/1)
vänta (8/8)
välbefinnandet (1/1)
reser (5/5)
begränsningarna (4/4)
utfärdats (10/10)
orsaken (6/6)
grader (3/3)
tis (2/2)
antecknar (1/1)
uppehållsrätten (18/18)
återhämtar (3/3)
hemlandet (2/2)
samarbeta (1/1)
tillsammans (56/56)
företagarhandböcker (1/1)
inkomst (12/12)
gränsöverskridande (1/1)
dela (5/5)
organisationer (15/15)
relativt (4/4)
utveckla (12/12)
meningar (1/1)
tidsbeställningen (2/2)
bostadsbyrå (1/1)
förmedling (1/1)
socialskyddet (3/3)
bostadslösafinska (2/2)
mark (3/3)
gångtrafiken (1/1)
finskspråkiga (14/14)
Uudenmaan (1/1)
återvändandefinska (1/1)
lokal (1/1)
finansieras (1/1)
behärska (1/1)
språkversionerna (2/2)
arbetarskyddet (2/2)
förlovningen (1/1)
hjärtat (1/1)
parktanterna (1/1)
historia (6/6)
bedriver (5/5)
kostnad (1/1)
skarvsladd (1/1)
kvalifikationer (4/4)
Vionojas (1/1)
bibliotek (16/17) Bibliotek (1)
arbetsamhet (1/1)
städning (1/1)
sexualitetfinska (1/1)
stred (2/2)
åren (6/6)
Kvinnokliniken (1/1)
områden (17/17)
peruskoulutukseen (1/1)
säkerheter (1/1)
upptagna (1/1)
ombud (1/1)
Nupoli (4/4)
familjemedlem (28/30) Familjemedlem (2)
anställningar (4/4)
ansökan (145/147) Ansökan (2)
operera (1/1)
förhållanden (2/2)
vigseln (9/9)
straffbart (2/2)
mobbning (1/1)
lekpark (2/2)
stadsdelfinska (3/3)
organisationen (1/1)
rättelserna (2/2)
hälsovårdstjänsterfinska (1/1)
ansökningstiden (3/3)
vägar (1/1)
skatter (9/9)
studenthälsovårdarna (1/1)
skenäktenskap (1/1)
parkerna (1/1)
modern (20/20)
Utvecklingsstörning (1/2) utvecklingsstörning (1)
lönebesked (1/1)
kontor (4/4)
uppförandet (1/1)
lagringsavgifter (1/1)
kortfattade (1/1)
r.f. (4/4)
folkhögskolorfinska (1/1)
ingå (10/10)
inkorporerade (1/1)
båtlivfinska (1/1)
bolagsordningen (1/1)
förbereds (1/1)
person (64/64)
småbarnspedagogik (11/11)
omedelbart (3/3)
omfattning (5/5)
äldrefinska (1/1)
färdas (4/4)
korttidsrehabilitering (1/1)
studentexpeditionen (1/1)
skräp (1/1)
stadslotsen (1/1)
panelen (2/2)
sitter (3/3)
anmält (4/4)
utländska (17/20) Utländska (3)
sjöfästning (1/1)
Suomenkielisen (1/1)
fostras (2/2)
pensionsinkomster (1/1)
ej (1/1)
semesterna (1/1)
kustregionerna (1/1)
bindande (6/6)
anknyter (4/4)
nio (5/5)
fruktan (1/1)
fysioterapeut (1/1)
ca (4/4)
utsidan (1/1)
besiktningskontor (1/1)
rusmedelsmottagning (1/1)
kulturarvet (1/1)
tjänst (11/11)
ugnen (1/1)
varma (4/4)
morbror (1/1)
papperslöshetfinska (1/1)
närståendevåld (1/1)
syns (4/4)
överklagas (1/1)
Romppu (1/1)
översättas (3/3)
fuktproblem (1/1)
myndighetens (2/2)
högskolor (12/13) Högskolor (1)
tingsrättenfinska (1/1)
ytmaterial (1/1)
följd (5/5)
hemvist (2/2)
gammalt (6/6)
Liechtenstein (12/12)
möjlighet (23/23)
visumärenden (1/1)
julen (2/2)
gymnasiestudierfinska (1/1)
gottgörelse (1/1)
utgången (4/4)
karens (1/1)
Runeberg (1/1)
hallen (1/1)
kostnadsersättningfinska (1/1)
begått (4/4)
finansieringen (4/4)
fås (14/14)
packas (2/2)
utbildningsväsendet (2/2)
beräkna (3/3)
främmande (9/9)
föregående (1/1)
urspråken (1/1)
uppträder (2/2)
germanska (1/1)
Marthaförbundetfinska (1/1)
Startup (1/1)
heltidsarbete (2/2)
kursstart (1/1)
egendom (28/28)
styrker (2/2)
sju (8/8)
stödpersoner (1/1)
stegen (1/1)
areal (3/3)
intresserad (8/8)
målsättningen (1/1)
perhe (1/1)
rådgivningsställe (1/1)
tatarer (1/1)
kundtjänstfinska (1/1)
invånarantalet (1/1)
vinterskor (1/1)
elev (2/2)
överallt (1/1)
skilsmässoansökan (6/6)
länkar (5/5)
handelsstad (2/2)
arbetarinstitut (11/11)
vandrarhem (1/1)
tjänstemännen (2/2)
uppsöka (1/1)
grunda (31/31)
medlemsländer (1/1)
nätbankkoder (1/1)
felaktiga (3/3)
rökfria (1/1)
underhållsstöd (4/4)
omfattar (24/24)
maksuhäiriömerkintä (1/1)
fördröjas (1/1)
utbildningen (53/53)
stödjer (5/5)
yrkesutbildade (1/1)
ungerska (8/8)
idrottsväsendet (1/1)
kultur (13/13)
stället (2/2)
döva (1/1)
kassan (5/5)
gymnasiestudierna (2/2)
miljoner (1/1)
understöd (10/10)
servicehus (5/5)
mötesplatsen (1/1)
socialhandledningfinska (1/1)
tillsvidare (6/6)
bostadsförmedlaren (4/4)
egenföretagare (1/1)
Mona (4/4)
andra (185/185)
borgare (1/1)
hinder (15/15)
flyttservice (1/1)
europeiskt (2/2)
lyder (1/1)
filmfestival (1/1)
omskärelse (6/6)
bakgrund (5/5)
studerandeengelska (1/1)
tidningsannonser (2/2)
anslagstavlor (1/1)
dubbelexamen (1/1)
Akatemia (3/3)
människa (2/2)
dygn (3/3)
institutets (7/7)
haltijakohtainen (1/1)
cykling (4/4)
bland (38/38)
konstnären (1/1)
undgår (1/1)
avgiftningsvård (1/1)
överenskomna (2/2)
utomstående (3/3)
ske (2/2)
dröjsmål (1/1)
Rovalan (7/7)
skild (1/1)
hyresgarantin (2/2)
P (3/5) p (2)
cykelkarta (1/1)
BY (2/2)
föräldradagpenningar (3/3)
appar (2/2)
narkotika (1/1)
daggymnasiet (1/1)
fester (3/3)
Akava (1/2) AKAVA (1)
arbetstagarens (5/5)
asylansökanfinska (1/1)
avser (6/6)
hälsofrämjande (1/1)
Marthaförbundet (1/1)
födelseattest (6/6)
avbryts (3/3)
osäker (2/2)
företagarefinska (6/6)
start (1/1)
par- (1/1)
behörig (1/1)
servicenumret (1/1)
besvären (4/4)
lösgjorde (1/1)
ordningsreglerna (7/7)
dig (368/368)
varierar (18/18)
företagshälsovårdenfinska (1/1)
laddat (1/1)
ungdomar (27/27)
nedsättande (2/2)
lokaltidningarna (1/1)
gymnasiestudier (6/6)
anställningsvillkoren (2/2)
familjehusen (1/1)
picknick (1/1)
införde (2/2)
familjeförening (2/2)
utsätta (1/1)
slutligen (1/1)
studentbostadsstiftelser (1/1)
välfärd (6/6)
Startpunkter (1/1)
ersatts (1/1)
gäller (40/40)
så (63/63)
lämnade (4/4)
integrationsspråk (1/1)
cykel- (1/1)
olaglig (1/1)
höjs (1/1)
självständighetens (1/1)
van (1/1)
arbetsmotivation (1/1)
Rooska (1/1)
tillväga (1/1)
individer (1/1)
uppsägningen (1/1)
egendomsfördelning (1/1)
mödrahem (2/2)
värdesätts (4/4)
bevåg (1/1)
fisket (1/1)
upp (67/67)
ockuperade (1/1)
bedömningsgrunder (1/1)
hälsovårdsstationen (1/1)
näringsbyråer (2/2)
Barnkliniken (3/3)
kvinnorfinska (1/1)
originalexemplaren (5/5)
festföremålet (1/1)
byråerna (1/1)
vuxnafinska (3/3)
färdmedel (1/1)
orsaka (5/5)
koncentrerad (1/1)
resa (7/7)
Livsmedelsverket (1/1)
pappersansökan (1/1)
tidsbokningstjänst (1/1)
Asunnot (6/12) asunnot (6)
finländarna (19/19)
sjukdagpenningfinska (2/2)
jobbet (3/3)
betyder (24/24)
kierrätyspiste (1/1)
lisä (1/1)
utöva (8/8)
främja (9/9)
upphovsrätt (6/6)
hobbygrupper (1/1)
rötter (1/1)
vårdsystemet (1/1)
grunddagpenningen (1/1)
YouTube (2/2)
privatvårdsstödet (1/1)
K.H.Renlunds (3/3)
industriprodukter (1/1)
handelstrafik (1/1)
begravningen (3/3)
socialväsen (2/2)
anmälningsblanketten (2/2)
löften (1/1)
museiområden (1/1)
ramen (1/1)
översättningarna (1/1)
FRK (1/1)
likabehandling (12/12)
Tulli (1/1)
legaliserad (2/2)
kierratys.info (2/2)
se (16/16)
börja (16/16)
skattebyrå (3/3)
videkvistar (1/1)
offentlig (8/8)
industri (2/2)
barndagvård (8/8)
föreskrivas (1/1)
servicen (1/1)
vardera (2/2)
transport (1/1)
följer (12/12)
psykoterapeutti (1/1)
sjukvårdstjänster (5/5)
någon (71/71)
befolkningen (3/3)
samhälleliga (1/1)
verkställande (1/1)
befriats (2/2)
avfallet (5/5)
vokabulär (2/2)
följs (11/11)
grundlag (2/2)
förskottsinnehållning (2/2)
rimliga (1/1)
föreningsmötet (1/1)
lekens (1/1)
flygplatser (1/1)
översättning (1/1)
gymnasiebaserad (2/2)
elbolaget (1/1)
affärsverksamhetsplan (9/9)
kulturproducenter (1/1)
intervjuar (1/1)
hennes (9/9)
arbetskollektivavtal (1/1)
arbetets (2/2)
tillväxt (4/4)
pappfabrik (1/1)
disk- (1/1)
lån (23/23)
slussar (1/1)
identitetskort (7/7)
skadegörelse (1/1)
antalet (5/5)
sådana (14/14)
preventivmedel (12/12)
lyfter (1/1)
uttrycka (2/2)
ändringar (6/6)
kauniainen.fi (1/1)
Reittiopas (2/2)
matburkar (1/1)
almanacksbyrå (2/2)
sjukdom (20/20)
hamnar (2/2)
Hyresboende (1/1)
Opetushallitus (5/7) opetushallitus (2)
graviditetstest (2/2)
Navigatorn (5/5)
dagpenningenfinska (1/1)
lastensairaala (1/1)
bestäms (6/6)
Silkinportin (1/1)
bristfälliga (1/1)
blivit (30/30)
anhörigvård (1/1)
fre. (1/1)
kosthållsbranschen (1/1)
språkstudier (1/1)
App (1/1)
persons (3/3)
tjänsteleverantörers (1/1)
moderns (7/7)
medborgares (7/7)
tilläggsundervisning (2/2)
högskolornas (3/3)
sjukhusvård (2/2)
värms (1/1)
sökfält (1/1)
webbtjänstfinska (1/1)
Grankullafinska (1/1)
pensionärer (4/4)
Tyskland (1/1)
matlagning (3/3)
skuld (1/1)
Nyföretagarcentral (1/1)
organ (1/1)
självrisktiden (2/2)
presidentvalfinska (1/1)
tredjelandsmedborgare (1/1)
anmäler (14/14)
slags (17/17)
arbetslösfinska (1/1)
samkönade (2/2)
översättar- (3/3)
kypsyysnäyte (1/1)
Mt (2/2)
tävlingsdeltagaren (1/1)
kalla (2/2)
privatpersoners (1/1)
resekortet (2/2)
flerårigt (1/1)
avsätts (1/1)
työehtosopimukset (1/1)
arbetsdagen (2/2)
familjerådgivningscentralen (1/1)
vardagkvällar (1/1)
smarta (1/1)
kommunfullmäktige (5/5)
snön (1/1)
avstängda (1/1)
högsta (8/8)
sökordet (1/1)
andraspråk (3/3)
psykoterapifinska (1/1)
barnpassningshjälpen (1/1)
skal (1/1)
barnets (93/94) Barnets (1)
erforderliga (1/1)
parterapi (1/1)
kontinuerlig (1/1)
projektet (1/1)
registrera (36/36)
kontrollerar (1/1)
takt (2/2)
garantipensionen (2/2)
småbarn (1/1)
Befolkningsregistercentralen (1/1)
nödsituation (11/11)
seder (5/5)
rättsväsendet (1/1)
kaupunginvaltuusto (1/1)
pääkaupunkiseudun (1/1)
ägodelarna (1/1)
brandvarnare (6/6)
registreringsblanketten (1/1)
skattskyldiga (1/1)
idrott (3/3)
maka (31/31)
ersättningarfinska (1/1)
bolagsmän (1/1)
grannmedlingfinska (1/1)
frivilligt (8/8)
utrikes (1/1)
uskonnonvapaus (1/1)
befogade (1/1)
ägda (1/1)
remiss (12/12)
graviditeten (16/16)
senast (25/25)
Helsingforsregionen (5/5)
när (196/202) När (6)
minnestest (1/1)
Komihåglista (2/4) komihåglista (2)
tillfrågas (1/1)
lyftandet (1/1)
rättshjälpfinska (1/1)
politik (1/1)
bilen (6/6)
bolagsman (2/2)
också (308/308)
kesäteatterifinska (1/1)
köpeanbudet (2/2)
lönesystemet (1/1)
oman (1/1)
ventilation (1/1)
känslofyllda (1/1)
rehabiliteringfinska (5/5)
avliden (1/1)
servicerådgivningen (1/1)
sammanlagda (2/2)
aborten (1/1)
Estland (1/1)
värme (1/1)
stiftas (1/1)
symtom (1/1)
begravas (3/3)
Yle (1/1)
mannen (5/5)
misstänka (1/1)
trygga (8/8)
svårare (4/4)
avgifter (5/5)
avtalad (2/2)
godkänts (3/3)
uppbära (1/1)
överlåter (2/2)
gränssnittetfinska (1/1)
Företagsrådgivning (2/4) företagsrådgivning (2)
genomgå (2/2)
riksdag (1/1)
republik (2/2)
kyrkliga (5/5)
oklarheter (3/3)
höghusfinska (1/1)
må (1/1)
syn (2/2)
verksamhetsformerna (1/1)
centralsjukhus (3/3)
linkkiBybiblioteken (1/1)
keskus (1/1)
Åboregionen (1/1)
siviilisäätytodistus (1/1)
ungdomars (1/1)
A1 (5/5)
upptäcka (1/1)
utövar (7/7)
kommer (62/62)
Migrationsverket (28/31) migrationsverket (3)
kondylom (1/1)
HRT:s (2/2)
sjukfall (3/3)
väestötietojärjestelmä (1/1)
anställningsskyddet (1/1)
temperaturen (2/2)
lätta (1/1)
löner (2/2)
öppettider (8/8)
videon (1/1)
därom (1/1)
färdig (1/1)
makes (5/5)
församlingfinska (1/1)
föräldrarnas (10/10)
pappersrecept (1/1)
inkomstgränsen (1/1)
befolkningsdatasystem (4/4)
patients (1/1)
personligt (6/6)
populärare (1/1)
börjar (34/34)
säkerhetsanvisningar (1/1)
verkställer (1/1)
nationalitet (9/9)
anställdas (5/5)
högskolestudier (8/8)
fortsatte (1/1)
företagarkurser (1/1)
Alkoholistit (1/1)
bostadfinska (3/3)
yhdistys (1/1)
järnaffärer (1/1)
Begravningsbyråers (1/1)
arbetarskyddsmyndigheter (1/1)
psykiatrisk (2/2)
respons (6/6)
emigranter (2/2)
jobbsökningenfinska (1/1)
lönesättning (1/1)
FöretagsEsbo (1/1)
riksdagens (1/1)
påskdagen (1/1)
mellanmål (1/1)
syskon (4/4)
färdighetsnivå (2/2)
pompa (1/1)
kaavinta (1/1)
rådgivningsbyråernas (2/2)
ämbetsverk (1/1)
kroatiska (4/4)
statsrådet (2/2)
www.teosto.fi (1/1)
distansundervisning (1/1)
kvotflyktingar (8/8)
ammattiliitto (1/1)
ekonominfinska (1/1)
krigsskadestånd (1/1)
toimisto.fi (1/1)
sjukpenning (1/1)
hissa (1/1)
regionförvaltningsverken (1/1)
resmålet (1/1)
äldsta (2/2)
kontakttolkar (1/1)
eftersom (19/19)
forskningen (1/1)
katastrofer (1/1)
uppgift (8/8)
ämnen (10/10)
informationstjänst (1/1)
önskar (5/5)
berättigad (2/2)
motionsalternativfinska (1/1)
Opiskelija (4/4)
chatten (2/2)
faderskapet (12/12)
beteendefinska (3/3)
avsluta (1/1)
lista (7/9) Lista (2)
Spafinska (2/2)
sjukhusen (1/1)
ingång (3/3)
Esbotillägget (1/1)
närmaste (20/20)
Nokia (1/1)
bostadsrättsavgift (1/1)
medeltalet (1/1)
skogar (1/1)
rutter (5/5)
linkkiFinnkino (1/1)
åtgärdande (1/1)
grundade (2/2)
scenkonst (1/1)
tandläkaren (3/3)
sopsortering (1/1)
instruktioner (1/1)
invånarantal (1/1)
stadiluotsi (1/1)
hörselundersökning (1/1)
kulturhistoria (2/2)
heltidsarbetande (1/1)
hälscentralsavgifter (1/1)
studiebetyg (1/1)
miljö (5/5)
isdubbar (1/1)
osittainen (1/1)
hammashoitola (2/2)
tutkinta (1/1)
julskinka (1/1)
uppehållstillståndetfinska (1/1)
norska (9/9)
lika (15/15)
arbetstagare (32/33) Arbetstagare (1)
bisyssla (2/2)
vakinaista (2/2)
familjehem (2/2)
Schengenområdet (6/6)
förälderns (3/3)
smärtjouren (1/1)
handlingen (2/2)
hemmet (36/36)
nationella (2/2)
upplösande (1/1)
samkommunen (3/3)
undervisningfinska (2/2)
lokaltrafikens (1/1)
koncentrationssvårigheter (1/1)
känslor (1/1)
resepti (1/1)
fortsätter (2/2)
tjänstemän (1/1)
upplöses (1/1)
skett (1/1)
sätter (2/2)
Psykologiförbund (1/1)
tidskriften (1/1)
guiden (2/2)
läkemedelsförpackningen (1/1)
kursen (4/4)
kuntoutustuki (1/1)
spis (1/1)
välkomna (3/3)
spisfläkten (1/1)
idkandet (1/1)
stad (47/47)
arbetskraft (2/2)
gymnasiet (21/21)
diskriminerande (2/2)
folkhögskolanfinska (1/1)
värdesätter (3/3)
bestraffning (2/2)
arbetstiderna (1/1)
gårdsområdet (1/1)
bolagsmannen (1/1)
estniska (51/51)
arbetskraftsmyndigheten (1/1)
låneräknare (1/1)
påverkan (5/5)
namnskylt (1/1)
beredningen (1/1)
mening (1/1)
Tysklands (1/1)
skilt (3/3)
yhtiö (1/1)
undrar (1/1)
hantverk (3/3)
semesterersättning (2/2)
elatustuki (1/1)
förskottsskatt (1/1)
enklast (1/1)
hyrs (9/9)
välbefinnande (1/1)
läckaget (1/1)
överklagan (1/1)
InfoFinlands (289/289)
fristående (9/9)
alternativ (8/8)
läroboken (1/1)
vi (11/15) Vi (4)
hembygdsmuseer (1/1)
språkkurser (3/3)
fortsättningen (1/1)
skatteräknare (1/1)
besvärlig (1/1)
beställer (7/7)
tolkningstjänsten (1/1)
enligt (53/53)
uppsägningsvillkor (3/3)
för- (1/1)
Nuorisoasiainkeskus (1/1)
kropps (1/1)
handikapp (18/18)
perustamisilmoitus (1/1)
tågbiljetter (1/1)
träffarna (1/1)
stödåtgärderfinska (1/1)
hårt (1/1)
suomi.fi (2/3) Suomi.fi (1)
desto (1/1)
besökt (3/3)
peruskoulupohjainen (1/1)
droganvändning (1/1)
skivor (1/1)
dras (4/4)
provar (1/1)
själv (93/93)
Studenternas (1/1)
utländsk (15/16) Utländsk (1)
delaktighet (1/1)
gravida (8/8)
besluten (1/1)
droger (5/5)
viitekehys (1/1)
kvalitet (2/2)
Oy (9/9)
matematik (1/1)
telefon (38/38)
normalt (4/4)
högersinnade (1/1)
dagvårdsproducenten (1/1)
skrift (1/1)
hälsotjänsterna (3/4) Hälsotjänsterna (1)
patientens (2/2)
utvecklingsstördafinska (1/1)
västliga (1/1)
språketfinska (6/6)
hörselskadade (5/5)
beslutsorganet (1/1)
rehabiliteringar (1/1)
djuren (1/1)
satsat (1/1)
gäst (2/2)
avslutas (1/1)
forna (1/1)
elev- (1/1)
konstruktionen (1/1)
tillväxten (1/1)
tjära (3/3)
makan (8/8)
klubbarfinska (1/1)
hälsostationernas (2/2)
omsorgsfullt (2/2)
paus (1/1)
uppges (3/3)
missbruksfrågor (1/1)
flyktingfinska (1/1)
grundlagen (2/2)
fots (2/2)
semestern (2/2)
NA (1/1)
läroavtalscenter (3/3)
Yritys (2/2)
mitten (3/3)
begravningsplats (8/8)
reservera (4/4)
flyttning (1/1)
hälsoundersökning (1/1)
uppgifterna (12/12)
erkände (1/1)
centralt (1/1)
stängt (6/6)
välartat (1/1)
utomlands (61/61)
föräldraledig (3/3)
skidåkning (2/2)
biljettkontoren (1/1)
satt (2/2)
skolhälsovårdaren (4/4)
presidenten (3/3)
utbilda (5/5)
stödundervisningen (1/1)
motsätter (2/2)
ITE (1/1)
upplever (7/7)
psykoterapi (4/4)
tågen (1/1)
synnerhet (1/1)
underskrifterna (1/1)
-kuntayhtymä (1/1)
teckenspråketfinska (1/1)
sorani (3/3)
ensam (15/15)
ägaren (1/1)
specialfinansieringsbolag (1/1)
Clubs (1/1)
konsumentens (3/3)
smärtan (1/1)
tjänsterna (31/31)
konditionen (2/2)
studierna (26/26)
musikhobby (1/1)
lähetetty (1/1)
konstruktioner (2/2)
tillverkning (1/1)
sakkunskap (1/1)
avslag (2/2)
Unionin (1/1)
sanning (1/1)
startas (1/1)
hjälpt (1/1)
myndighetshandlingen (1/1)
drogs (1/1)
taitavan (1/1)
läkemedlen (1/1)
ansökningsbilagorna (6/6)
bostadsaktier (1/1)
innevarande (1/1)
kyrkoherdeämbetet (1/1)
fars (1/1)
plastförpackningarna (1/1)
plan (1/1)
vars (20/20)
kö (1/1)
upphävande (1/1)
ärlighet (3/3)
fram (13/13)
löntagar- (1/1)
äitiysavustus (2/2)
rekreationsområde (1/1)
helgons (3/3)
sistnämnda (1/1)
historiska (4/4)
framförd (1/1)
sjukdomar (8/8)
varat (5/5)
försvårar (1/1)
årligen (1/1)
ändring (1/1)
servicehandledning (1/1)
anvisa (1/1)
säätiö (1/1)
beviljar (4/4)
arbetspensionsutdraget (1/1)
ledigheterna (1/1)
postadressen (1/1)
Förbundfinska (1/1)
kombineras (1/1)
mängd (5/5)
flerfaldiga (1/1)
pappersformat (1/1)
konstuniversitet (2/2)
Sammallahdenmäki (1/1)
medlemskortetfinska (1/1)
praktiskt (1/1)
lokala (8/8)
handelskammare (2/2)
kulturgrupper (1/1)
vintersporterna (1/1)
mån. (1/1)
ägarskapet (1/1)
Lapplands (21/21)
samtalskostnad (1/1)
människohandel (12/12)
måltidstjänster (1/1)
sommaruniversitetet (2/2)
biljettjänstens (1/1)
patientjournalen (1/1)
väderförhållanden (1/1)
museums (1/1)
grammatikfinska (1/1)
räknar (1/1)
relaterade (1/1)
utsatta (2/2)
avdragen (1/1)
hälsoproblem (1/1)
medarbetare (1/1)
olja (1/1)
kommunikationskanal (1/1)
bostadsrättskontraktet (1/1)
läkarutlåtande (2/2)
sinsemellan (1/1)
skattepliktiga (1/1)
utbildningar (7/7)
veckoslut (15/15)
magistraternafinska (1/1)
Perho (1/1)
avloppet (1/1)
japanska (6/6)
tulkkaus (1/1)
huvudsyssla (3/3)
originalspråk (1/1)
hur (93/94) Hur (1)
skadas (1/1)
magistratens (7/7)
API (1/1)
moder (1/1)
Folkdans (1/1)
Ceremonier (1/1)
ämne (3/3)
avlyssnas (1/1)
ändrat (1/1)
stiftelsens (2/2)
fyllda (1/1)
upphängningsbygel (1/1)
allmänt (6/6)
kommunikationen (1/1)
kontaktuppgifterna (15/15)
Residuum (2/2)
informerar (5/5)
SERI (2/2)
läkarstation (14/14)
Ohjaamo (1/1)
bäst (9/9)
suppleanter (1/1)
Fennovoimas (1/1)
etniskt (7/7)
inbyggd (1/1)
blir (59/59)
personbeteckningar (1/1)
öppningsoperation (3/3)
applikationsbutiken (1/1)
rösten (1/1)
skolkuratorerna (2/2)
undervisningen (26/26)
hjälpsystemet (1/1)
jourmottagningen (17/17)
oikeus (1/1)
stödengelska (1/1)
pensionsförsäkring (3/3)
godkänt (4/4)
bouppteckningfinska (1/1)
organen (1/1)
yrkeshögskoleexamina (1/1)
hyresgaranti (1/1)
omhändertagande (1/1)
vaccinationer (4/4)
sjukförsäkringen (13/13)
skulden (2/2)
konkurs (3/3)
studentskrivningarna (1/1)
utbildningsplats (2/2)
bassjälvrisk (1/1)
förskoleenheter (1/1)
civil (2/2)
löneutbetalningen (4/4)
förpackningsmaterial (1/1)
A (25/26) a (1)
hobbyklubbar (1/1)
driva (5/5)
sälja (6/6)
ordningsnummerfinska (1/1)
medlem (20/20)
beskriver (5/5)
förmåga (2/2)
åstadkomma (1/1)
skräpa (1/1)
lokaltrafiken (1/1)
specialiserat (2/2)
kraft (13/13)
30l (1/1)
licentiat- (1/1)
vårdbidrag (1/1)
förtrogna (1/1)
garanti (2/2)
bildkonst (8/8)
jourtidsbeställning (1/1)
Karlebystöd (1/1)
kontinuerliga (3/3)
kran (1/1)
händelsen (1/1)
pimpelfiske (1/1)
förlossning (8/8)
Health (1/1)
renkött (1/1)
prövningsbaserat (1/1)
beaktas (14/14)
huvudbiblioteket (1/1)
ugriska (1/1)
vuxengymnasiums (1/1)
avboka (2/2)
förbereda (2/2)
anskaffningspris (1/1)
Tukiliittos (1/1)
tietopankki (1/1)
försörjningen (4/4)
medverkat (4/4)
både (24/24)
dygnet (25/25)
tolkförbunds (1/1)
civilstånd (1/1)
Chydenius (2/2)
förhandlar (1/1)
parkeringsautomat (1/1)
specialundervisning (5/5)
yrkesval (1/1)
enlighet (7/7)
hälsostationsläkaren (1/1)
arbetar (40/40)
nackdel (1/1)
studietakt (1/1)
seniorer (6/6)
vinterkriget (1/1)
alternativt (2/2)
återresa (2/2)
asylansökan (15/15)
ambulans (1/1)
låga (4/4)
höger (1/1)
butiker (2/2)
hälsovårdsverket (1/1)
grannarna (1/1)
strejk (1/1)
lägger (2/2)
biblioteksnätverket (1/1)
studievägledarna (2/2)
patientombudsmannen (2/2)
psykiska (6/6)
nödvändigtvis (10/10)
invånarparker (1/2) Invånarparker (1)
musikundervisning (1/1)
lönsam (3/3)
papperspåse (1/1)
turistersvenska (1/1)
Internetanslutningar (1/1)
skatteprocenten (2/2)
kommunaval (1/1)
å (3/3)
augusti (6/6)
Centralförbundet (1/1)
resorna (1/1)
Ylikylä (1/1)
naturcenter (1/1)
vuxenstuderande (4/4)
misslyckades (1/1)
handling (4/4)
webbenkäter (1/1)
högt (4/4)
skydda (3/3)
Kervo (2/2)
idkas (2/2)
fukt (2/2)
tillgångar (4/4)
bruksvederlaget (2/2)
arbetsuppgiften (4/4)
varderas (1/1)
sorgfinska (1/1)
brottsmisstänkta (3/3)
yrkena (1/1)
populära (4/4)
basis (11/11)
kotihoito (1/1)
osakliga (1/1)
arbetstagaren (16/16)
kansalaisuusilmoitus (2/2)
hemtjänster (1/1)
läst (4/4)
läroanstalterna (2/2)
huvudhälsostationen (1/1)
lånekostnaderna (1/1)
medeltiden (1/1)
läkarhjälp (1/1)
kortkurser (1/1)
tolken (13/13)
fortsättningsvis (1/1)
medicinska (2/2)
statliga (9/9)
dagvården (13/13)
medborgarinstitutets (4/4)
arbetet (49/49)
avgiften (4/4)
Korsets (1/1)
boendeform (1/1)
bruk (3/3)
läser (8/8)
transporttjänst (1/1)
bådas (2/2)
trästadshelheter (1/1)
helsinki.fi (1/1)
heder (1/1)
Sportkort (1/1)
eftermiddagsverksamhet (3/3)
arbetspensionsanstalt (1/1)
vare (5/5)
läggs (1/1)
socialservice (1/1)
specialtjänster (1/1)
abort (8/9) Abort (1)
grundundervisning (2/2)
talar (6/6)
antas (3/3)
doula (1/1)
högskola (7/7)
Espoon (7/7)
helger (6/6)
räkna (2/2)
utmattade (1/1)
sjukhuskostnaderna (1/1)
diskrimineringfinska (1/1)
västeuropéer (1/1)
göra (73/73)
grundande (3/3)
turvallisuusvirasto (1/1)
fritiden (1/1)
husdjur (1/1)
förekomma (2/2)
Osviitta (1/1)
visning (1/1)
skolarbete (1/1)
Kitfinska (1/1)
IHH (1/1)
ylletröja (1/1)
babyns (1/1)
linor (1/1)
hälsocentralsjouren (1/1)
diskriminerings- (2/2)
työväenopisto (4/4)
Mielenterveys (1/1)
tjänsteställen (1/1)
ingåtts (5/5)
styrelsemedlem (1/1)
modersmålsundervisning (1/1)
båtliv (1/1)
vården (11/11)
tävlingens (3/3)
vattentrafiken (1/1)
konstundervisningfinska (1/1)
begå (2/2)
dina (112/113) Dina (1)
måltidsstödet (1/1)
sjunde (1/1)
tigga (1/1)
Finlandfinska (28/28)
utanför (17/17)
stödtjänsterna (2/2)
lantdagsmannen (1/1)
vindruta (1/1)
missbruk (2/2)
utfärdades (1/1)
tyger (1/1)
boendetjänster (2/2)
pensionsanstalt (3/3)
lands (5/5)
resan (2/2)
arbetslösafinska (3/3)
Lappland (6/6)
förvärvats (1/1)
administration (1/1)
eftermiddagen (2/2)
yrkeskunskaper (2/2)
beräknas (10/10)
teaterföreställningar (2/2)
förutsätta (1/1)
tolktjänst (2/2)
bruttoinkomster (1/1)
socialskyddsförmånerna (1/1)
honom (3/3)
erhöll (1/1)
polisanmäla (1/1)
konsumenter (1/1)
fordon (1/1)
hyresboendefinska (1/1)
utevistelse (1/1)
steril (2/2)
starttiraha (1/1)
arbetarskyddschef (1/1)
viktig (15/15)
hör (26/26)
asunto (2/2)
redaktionen (1/1)
tillhandahålla (2/2)
rödbetssallad (1/1)
republiken (1/1)
brandvarnaren (2/2)
banken (11/11)
bosättningsbaserade (1/1)
rättegången (2/2)
huvudstad (3/3)
läroanstalternas (2/2)
Garantistiftelsen (1/1)
sjukvårdstjänsterna (4/4)
karttjänsten (2/2)
holländska (10/10)
tand- (1/1)
arbetsplatserfinska (1/1)
familjeplaneringsrådgivningarna (1/1)
röstningsställe (1/1)
överklagar (1/1)
tillgängligheten (1/1)
sommarlov (1/1)
hammashoito (1/1)
pensionärerfinska (1/1)
hemspråksundervisning (5/5)
äidinkielen (1/1)
farföräldrarna (1/1)
linkkiLapplands (1/1)
medlemmar (15/15)
hälsocentralen (2/2)
dessa (56/56)
jobb (55/55)
pensionen (2/2)
upprättandet (3/3)
lågstadiets (1/1)
rollen (1/1)
oartigt (3/3)
medlemskommunernas (1/1)
krävande (5/5)
Hanhikivi (1/1)
dyrare (11/11)
skyldighet (7/7)
klinikerna (1/1)
kännedom (1/1)
italienska (15/15)
uppståndelse (1/1)
hittat (3/3)
fisk (1/1)
tal (1/1)
ljust (1/1)
föregår (1/1)
FPA.Som (1/1)
anrika (1/1)
internetionellt (1/1)
stadiet (6/6)
betalas (44/44)
likaberättigandefinska (1/1)
taxitjänster (1/1)
bekanta (6/6)
främjande (2/2)
tidsbestämt (8/8)
dansa (3/3)
vakuutus (2/2)
invandrarens (1/1)
tandläkarkontroll (2/2)
handelsmän (1/1)
fullt (1/1)
Aalto (2/2)
kända (1/1)
behålla (1/1)
tillförlitligt (2/2)
studerandena (1/1)
paddling (1/1)
herraväldet (1/1)
hobbystudier (2/2)
specialdiakoner (1/1)
Kunta (5/5)
resedokument (3/3)
hälsocentraler (1/1)
servicesställen (1/1)
nyheter (2/2)
Iso (5/5)
indriver (1/1)
Maahanmuuttovirasto (9/9)
rehabiliterande (2/2)
påverkar (14/14)
träffa (8/8)
gymnasieskolorna (2/2)
registrerat (12/12)
ll (1/1)
trafikfinska (1/1)
återflyttarefinska (1/1)
tvingats (1/1)
karriärmentorskap (1/1)
kremeras (1/1)
åtminstone (13/13)
föräldrapenning (3/3)
socialnämnden (1/1)
oss (1/1)
läkarrecept (3/3)
handelsregisterutdraget (1/1)
upprätthålls (5/5)
löpning (1/1)
bulgariska (6/6)
menas (1/1)
synskadade (4/4)
myndighetstjänst (1/1)
latauspiste (1/1)
giltighetstiden (2/2)
grundats (2/2)
Määräaikainen (1/1)
moderskapsförpackning (1/1)
servicebostäder (1/1)
finsk- (1/1)
familjerfinska (3/3)
batteriinsamlingslådor (1/1)
rösta (16/16)
Backas (1/1)
viktigt (30/30)
ventilationssystem (1/1)
intresserade (6/6)
månad (24/24)
fastställt (1/1)
sättet (4/4)
hanteras (2/2)
makten (4/4)
källa (1/1)
anknutna (1/1)
läsår (4/4)
fastlagsbullar (1/1)
informations- (2/2)
lyftanordningar (1/1)
CD- (1/1)
gruppen (5/5)
ständigt (1/1)
yleinen (3/3)
internationellt (8/8)
familjemedlemmar (21/21)
läsårsavgiften (2/2)
discipliner (1/1)
paperi (1/1)
textfält (1/1)
påverkafinska (3/3)
fackman (1/1)
skulle (9/9)
ombeds (1/1)
betydande (1/1)
något (71/71)
läroplanen (1/1)
reparationer (5/5)
producerar (1/1)
asylsamtal (1/1)
förra (1/1)
rad (1/1)
avstå (1/1)
invånarhusen (1/1)
besöken (1/1)
kassakvittot (1/1)
offentligt (7/7)
Perheiden (2/2)
Andelsbanken (1/1)
släckningsfilt (2/2)
hända (2/2)
ersätter (12/12)
aktiebolag (4/4)
missbruks- (1/1)
-trivsel (1/1)
CC (1/1)
ettdera (1/1)
lasi (1/1)
kontaktuppgifterfinska (7/7)
funktionsförmågan (2/2)
uppgöra (1/1)
begära (14/14)
folkhögskolafinska (1/1)
Havukoski (1/1)
offer (24/24)
judarna (1/1)
hårdare (1/1)
valkretsar (1/1)
flygeln (1/1)
delges (1/1)
lagarfinska (1/1)
sekajäte (1/1)
behovet (6/6)
landsvägsförbindelsermed (1/1)
arbetsolycksfall (1/1)
akuta (5/5)
Ungdomspolikliniken (1/1)
sidor (18/18)
utsökningfinska (1/1)
fungerar (5/5)
källskattekort (1/1)
lokaltrafik (1/1)
anser (3/3)
B (7/7)
förskrivningsrätt (1/1)
könummer (4/4)
äldre- (1/1)
kulturkontor (1/1)
Furumo (3/3)
flertal (1/1)
råkat (4/4)
språkkaféerna (1/1)
vardagsum (1/1)
männen (1/1)
reglerat (4/4)
observera (3/3)
tjänsten (64/64)
ljus (2/2)
skriven (1/1)
hjälpen (8/8)
förlossningen (18/18)
betalningen (1/1)
Mejlansvägen (1/1)
representerar (6/6)
handikapptjänster (2/2)
spelar (1/1)
skattmyndigheten (1/1)
grundare (2/2)
överförda (1/1)
läkaren (20/20)
källorna (1/1)
granskningar (1/1)
tolkar (2/2)
universitetskurser (1/1)
medverka (1/1)
skuldrådgivare (1/1)
Österbottens (17/17)
kunnig (1/1)
strid (1/1)
kör (1/1)
omskurits (2/2)
full (4/4)
ungdomarna (2/2)
fortlöpande (2/2)
gärna (3/3)
innehållits (1/1)
flyg (3/3)
vårdar (16/16)
handredskapsavgiften (1/1)
asuminen.fifinska (2/2)
Varia (3/3)
innefattar (1/1)
Ingående (2/3) ingående (1)
personen (9/9)
beskickningar (10/10)
uppsökande (3/3)
garantier (1/1)
regionutvecklingen (1/1)
påfrestande (2/2)
Utbildningsstyrelsens (13/17) utbildningsstyrelsens (4)
fördelningen (3/3)
tidigt (6/6)
skrivas (3/3)
smälter (1/1)
modersmål (35/35)
olyckor (2/2)
språkkunskapskraven (1/1)
principerna (1/1)
patienter (1/1)
Nuorten (3/3)
ladda (7/7)
byråerfinska (1/1)
övningar (1/1)
Vandatillägget (1/1)
buddhism (1/1)
kamratstöd (2/2)
letade (1/1)
lagrar (1/1)
A1.1 (1/1)
separata (4/4)
intyget (11/11)
Schengenland (1/1)
ålder (13/13)
asiointi (1/1)
ska (417/417)
publikationer (1/1)
välhållen (1/1)
rusmedelsberoendefinska (2/2)
hautausavustus (1/1)
försök (1/1)
språkinlärning (1/1)
högskolexamen (1/1)
daghem (34/34)
lönespecifikationen (2/2)
utom (4/4)
arbetslöshetsförmånfinska (1/1)
finansiera (1/1)
språken (5/5)
varmt (2/2)
tas (23/23)
uppväxt (4/4)
friluftsleder (1/1)
maken (10/10)
barnskyddsmyndigheten (2/2)
tvingande (2/2)
socken (1/1)
cykla (4/4)
förmedlare (1/1)
caféerna (1/1)
fiske (3/3)
biljettpriser (2/2)
undersöker (3/3)
Lochteå (1/1)
tors (5/5)
legaliserade (1/1)
könen (2/2)
telefoner (1/1)
granska (1/1)
telegram (1/1)
börjat (3/3)
handikappadefinska (3/3)
småstad (1/1)
klasserna (1/1)
högteknologiska (1/1)
riskerna (1/1)
G (1/1)
gäster (1/1)
deltid (5/5)
boendefrågor (1/1)
genomtänkta (1/1)
gymnasieböckerna (3/3)
brottsanmälan (7/7)
pensionstagarefinska (1/1)
tillåter (3/3)
hoitotakuu (1/1)
avbokat (1/1)
utföras (3/3)
arbetsuppgifterna (2/2)
utövat (2/2)
ulosotto (1/1)
fackföreningsverksamhet (1/1)
undersökningen (3/3)
peruskielitaito (1/1)
Rinteenkulmafinska (1/1)
pauser (2/2)
Registreringsanmälan (1/2) registreringsanmälan (1)
uppdrag (3/3)
utevistelser (2/2)
kvällen (4/4)
representant (2/2)
vartannat (3/3)
työtulo (1/1)
arbetslöshetspenning (1/1)
disponibla (3/3)
efter (88/88)
renoveringskostnaden (1/1)
företagsläkare (1/1)
missbrukstjänster (1/1)
huruvida (7/7)
liv (15/15)
stadigvarande (45/45)
finskakunskaper (1/1)
koulumatkatuki (1/1)
fiskelov (1/1)
kraftiga (1/1)
månatligen (2/2)
kopplat (1/1)
kursernas (1/1)
Tavataan (1/1)
försvunna (1/1)
konst (11/12) Konst (1)
klinikens (5/5)
Baltikum (1/1)
Al (1/1)
behörighet (4/4)
utlänningar (19/19)
Jesusbarnet (1/1)
musicera (1/1)
föräldrapenningperioden (3/3)
upplevs (1/1)
arbetsgivare (63/63)
kaffe (1/1)
godta (1/1)
ansvarsområden (1/1)
innerstad (1/1)
sommaren (10/10)
lähestymiskielto (1/1)
jourtid (1/1)
metodstudier (2/2)
polisstationernafinska (1/1)
klubben (2/2)
stadens (53/53)
konserter (1/1)
firma (1/1)
arbete (78/82) Arbete (4)
funktionsförmåga (1/1)
kärnkompetens (2/2)
verk (1/1)
arbetsuppgifter (8/8)
arbetsavtalslagen (2/2)
förbudet (1/1)
flygresor (1/1)
nuorisoasunnot (2/2)
äktenskapsförord (4/5) Äktenskapsförord (1)
sorts (2/2)
ungdomspolitiken (1/1)
betjänar (29/29)
bemött (1/1)
leda (1/1)
apteekki (1/1)
annanstans (10/10)
natur (1/1)
planer (1/1)
postpositioner (1/1)
aktuella (6/6)
anställningsavtal (1/1)
föräldramöten (2/2)
avtalet (21/21)
trafiken (2/3) Trafiken (1)
april (4/4)
Sporttia (1/1)
jämföra (4/4)
visering (1/1)
rekreationsdagar (1/1)
preventivmedelsrådgivningens (1/1)
ägarbostäder (1/1)
Studentkårers (1/1)
avsedda (27/27)
familjeåterförening (6/6)
toisena (1/1)
kortet (8/8)
dörrar (1/1)
band (1/1)
verifiera (1/1)
utrikespolitiken (1/1)
ansvarar (12/12)
görs (37/37)
medier (3/4) Medier (1)
diplomingenjörsexamen (1/1)
medlemskap (2/2)
betalningsanmärkningar (2/2)
temperaturerna (1/1)
grundskolanengelska (1/1)
hamnat (2/2)
skatt (21/21)
skicka (27/27)
Anonyymit (1/1)
volontärarbete (1/1)
grenar (3/3)
invandrarfamiljer (1/1)
vårdledig (3/3)
sjukvården (11/11)
osakeyhtiö (1/1)
godtar (1/1)
läroavtal (3/3)
allmän (8/9) Allmän (1)
Kopparbergsvägen (1/1)
grundläggande (43/45) Grundläggande (2)
uppstartsföretag (2/2)
facket (1/1)
oberoende (5/5)
ramper (1/1)
samband (10/10)
metallindustrin (1/1)
Arbisfinska (1/1)
inbrottstjuvar (1/1)
obetald (1/1)
semesterdagar (1/1)
anledningarna (1/1)
perustoimeentulotuki (1/1)
räkningar (2/2)
Inkomstregistrets (1/1)
universitetets (2/2)
fientlig (1/1)
eKirjasto (1/1)
anmärkning (2/2)
barnatillsyningsmannen (10/10)
sevärdheter (1/1)
Flickornas (2/2)
synnerligen (1/1)
elevens (8/8)
Uleåborgs (1/1)
kortfattad (1/1)
identitet (14/14)
företagets (8/8)
landskapsmuseumfinska (1/1)
berättigar (2/2)
hurudan (2/2)
idrottsplaner (2/2)
studenthem (1/1)
vaccinationsprogrammet (1/1)
placerar (2/2)
tänka (2/2)
ägodelar (2/2)
lagligt (5/5)
hög (7/7)
litar (1/1)
besvaras (2/2)
efterfrågan (1/1)
Patent- (2/3) patent- (1)
intressant (2/2)
förbjuden (2/2)
brottsofferfinska (2/2)
tryggare (1/1)
vårdkostnadsförsäkring (1/1)
grannskapet (1/1)
is (1/1)
stadgar (1/1)
krävs (32/32)
ämnet (6/6)
mathjälp (1/1)
mor (11/11)
hälsovårdsbranschen (1/1)
servicepunkterna (1/1)
socialjouren (2/2)
motiverade (1/1)
läs (2/2)
dödsorsaken (2/2)
Infopankki.fi (1/1)
om (1845/1851) Om (6)
tjänstens (2/2)
brinna (3/3)
elapparater (1/1)
utfärda (6/6)
hundratals (1/1)
kräver (21/21)
yrkeshögskolor (9/12) Yrkeshögskolor (3)
hemvården (2/2)
kartläggningfinska (1/1)
rådgivningstjänst (5/5)
identifiera (2/2)
krismottagning (2/2)
oåterkalleligt (1/1)
mentalvårdstjänsterna (1/1)
samtalsstöd (1/1)
minimibelopp (1/1)
pääomatulo (1/1)
fylla (19/19)
syssla (2/2)
trähus (1/1)
elektronisk (5/5)
endast (44/44)
personuppgifter (5/5)
rajoitetusti (1/1)
tydliga (1/1)
avgifterna (1/1)
näringar (1/1)
hälsostation (37/37)
inlärning (4/4)
förknippade (2/2)
sairauspäiväraha (2/2)
-Förbundet (1/1)
näyttötutkinto (4/4)
minoritetsspråk (1/1)
tillnyktrings- (1/1)
diskrimineringsombudsmannens (2/2)
www.tuotos.fi (1/1)
krigen (2/2)
sopsäck (1/1)
etnisk (2/2)
återfå (1/1)
julgran (1/1)
Kafnetin (1/1)
inomhus (1/1)
vårdkostnaderna (1/1)
näringslivstjänsterna (1/1)
lokaler (7/7)
guld (1/1)
farfinska (1/1)
jaktfinska (1/1)
mat (18/18)
vandring (2/2)
samhällsvetenskaper (2/2)
perustuslaki (1/1)
arbetsgivarens (4/6) Arbetsgivarens (2)
sekretessplikt (2/2)
utländskt (2/2)
land (140/140)
kollektivavtalen (3/3)
Finavia (1/1)
Apostilleavtaletengelska (1/1)
lilla (1/1)
hyran (14/14)
stambyte (1/1)
Ateneum (1/1)
palvelu (1/1)
arbetspraktik (3/3)
underhåll (5/5)
möjligtvis (1/1)
skilsmässafinska (2/2)
står (11/11)
Mannerheims (2/2)
fastän (5/5)
farförälder (2/2)
veckovisa (1/1)
opetus (2/2)
utkomst (6/6)
vetenskaps- (3/3)
hemfrid (1/1)
Regionförvaltningsverket (2/2)
skor (1/1)
vitsord (5/5)
ting (3/3)
normal (2/2)
uttalas (1/1)
intressen (7/7)
diskuterar (2/2)
ansluta (10/10)
musikskolor (1/1)
utlandsresa (1/1)
kalkyleras (1/1)
spela (4/4)
göras (29/29)
vårdenheter (1/1)
familjepension (5/5)
myndigheten (18/18)
olägenhet (1/1)
grundval (1/1)
landskapsplanerare (1/1)
tolka (1/1)
tillträde (2/2)
fördelas (1/1)
oikeusaputoimisto (4/4)
endera (4/4)
föreningarna (1/1)
bönestund (1/1)
påbyggnadsnivå (1/1)
moderskaps- (1/1)
kt (5/5)
luggas (1/1)
registreringen (6/6)
vän (7/7)
nätetfinska (1/1)
dagpenningens (1/1)
stödtjänsterfinska (1/1)
medborgarskapfinska (3/3)
jobbförmedlingssidor (2/2)
födelse (10/10)
marken (1/1)
närtågen (1/1)
vårda (1/1)
partier (1/1)
lägg (2/2)
hälsan (13/13)
korkein (1/1)
försörjning (12/12)
terminsavgift (1/1)
borta (1/1)
resten (3/3)
urval (1/1)
genomsnitt (4/4)
befunnit (1/1)
tomt (1/1)
Eija (2/2)
båda (20/20)
tillåtna (2/2)
bikulturellt (1/1)
Vantaalla.info (1/1)
ungdomen (1/1)
liksom (2/2)
bidrag (11/11)
förlora (7/7)
frivillig (5/5)
spelproblem (4/4)
saken (9/9)
barnmorska (1/1)
verksamheter (1/1)
hobby (7/7)
erkänts (3/3)
konstämnen (3/3)
pedagogik (5/5)
hjälpbehovet (2/2)
familjecenter (1/1)
hinner (3/3)
betalt (2/2)
separeras (1/1)
hyrorna (1/1)
treårig (1/1)
oväntat (2/2)
födelsedagar (1/1)
armé (1/1)
röstar (2/2)
idka (4/4)
pappor (1/1)
grundskolor (4/4)
avsnitt (5/5)
publicus (2/2)
behandling (9/9)
Suomen (12/13) suomen (1)
tunnustaminen (1/1)
skriftliga (5/5)
l (3/3)
baseras (1/1)
läroplikten (2/2)
bromsas (1/1)
Kärlek (1/1)
lyhytkurssi (1/1)
inresa (1/1)
underuthyrning (1/1)
ennakonpidätys (2/2)
hengenvaara (1/1)
norr (1/1)
utbildningsstöd (1/1)
palvelutalo (1/1)
återkallar (2/2)
ABC (2/2)
läkarundersökning (4/4)
individuella (1/1)
väcker (3/3)
mycket (66/66)
kliniken (7/8) Kliniken (1)
förpackningar (3/3)
lindras (1/1)
ikäihmisten (1/1)
annonserar (1/1)
työvoimakoulutus (1/1)
delägarbostadfinska (2/2)
handledningstjänster (1/1)
ålderspension (5/5)
skaffas (1/1)
kurserna (16/16)
bryter (4/4)
affärsverksamhetsplanen (5/5)
privatsektorn (1/1)
innehavarkort (1/1)
gatan (1/1)
detta (95/95)
högutbildade (1/1)
toimeentulotuki (1/1)
tillräcklig (10/10)
Twitter (1/1)
isen (7/7)
personlig (8/8)
publiceras (1/1)
arbetslivsfärdigheter (2/2)
fritidsverksamhet (1/1)
invandrares (2/2)
kommunsidor (1/1)
hälsorelaterade (1/1)
dags (1/1)
tjänat (1/1)
kaupunki (1/1)
partnern (2/2)
anhörigfinska (1/1)
utlänning (2/2)
näringsbyråeran (1/1)
fritidsaktiviteterna (1/1)
HIVfinska (1/1)
systemet (1/1)
samtal (4/4)
älvarna (1/1)
resesättet (1/1)
fara (6/6)
giftorätt (1/1)
vara (146/146)
poliklinik (1/1)
YEL (1/1)
Helsingforsregionen.fi (1/2) HelsingforsRegionen.fi (1)
sidoapotek (1/1)
billigare (2/2)
övernatta (5/5)
ämnesområden (1/1)
besök (8/8)
tidtabellerna (1/1)
teknik (2/2)
brinnande (1/1)
yrittäjien (1/1)
allra (2/2)
bostadsrättsavgiften (4/4)
3D (1/1)
hittar (202/202)
äventyras (1/1)
insjuknar (10/10)
Lapset (1/1)
fadern (10/10)
svagheterna (1/1)
mödrarådgivning (1/1)
förtida (3/3)
vokabulär- (1/1)
Schweiz (31/31)
gåvor (1/1)
med (667/667)
flyttsakerna (1/1)
föreslå (2/2)
känna (6/6)
tillsyn (1/1)
arbetstillstånd (1/1)
hushållspapper (2/2)
fördela (2/2)
pojkes (1/1)
regnbågsfamiljerfinska (1/1)
koder (1/1)
seger (1/1)
studiestöd (8/8)
skapar (1/1)
ofött (1/1)
absolut (1/1)
pitkä (1/1)
sakkunnig (2/2)
hemspråksundervisningfinska (1/1)
invaliditet (1/1)
vaccinerar (1/1)
EES (35/35)
månaden (6/6)
tis. (1/1)
arbetssökning (1/1)
biträdande (1/1)
landet (32/32)
förlängas (3/3)
beordra (1/1)
anpassa (1/1)
grupp (9/9)
Korkalovaara (1/1)
ränta (1/1)
genomförandet (1/1)
koordinatoren (1/1)
hens (1/1)
Flerspråkiga (2/2)
terapibesök (1/1)
följande (48/48)
universitetet (19/19)
veronpalautus (2/2)
minuter (1/1)
ganska (1/1)
delar (11/11)
följ (1/1)
barnrådgivningen (8/8)
tillståndsärenden (4/4)
övertidsarbete (1/1)
kontrollera (19/19)
kistor (1/1)
obligatoriskt (3/3)
föräldrapenningperiodens (1/1)
tingsrätts (2/2)
diskmaskinen (2/2)
stödnät (1/1)
fackförbund (14/16) Fackförbund (2)
oavsett (7/7)
köpare (2/2)
avgiftsbelagt (4/4)
narkos (1/1)
konsthusen (1/1)
borgensmän (1/1)
insamlingskärl (2/2)
omständigheter (4/4)
bosatta (16/16)
tjänster (128/133) Tjänster (5)
dröjsmålsränta (1/1)
studieregisterutdrag (1/1)
arbetspensionsanstalten (3/3)
värmeaggregat (1/1)
lekparkernas (1/1)
perhehoito (1/1)
värmeelement (1/1)
tvingade (1/1)
Petäjävesi (1/1)
440kt (1/1)
kartläggningen (14/14)
arbetsgivaren (49/49)
nyttar (1/1)
försäkringspremierna (4/4)
denne (3/3)
sända (1/1)
universitetsutbildningar (1/1)
aptit (1/1)
intersexuella (1/1)
ansökningsprocessen (1/1)
Anders (1/1)
avvisa (2/2)
jämkas (1/1)
varorna (1/1)
söder (1/1)
upprättade (1/1)
sommartid (1/1)
förmiddagar (1/1)
uppfattas (1/1)
fingeravtryck (1/1)
hälsostationens (1/1)
grundundervisningenfinska (1/1)
genetiska (1/1)
ingår (23/23)
hyra (21/21)
arbetslöshetsförmåner (1/1)
EU- (6/6)
nybörjareengelska (1/1)
preventivmetoder (1/1)
pensionerad (1/1)
personer (96/96)
sår (1/1)
formulerad (1/1)
framställning (1/1)
Oikarainen (1/1)
sammanlagt (2/2)
stressyndromfinska (1/1)
hjälp (183/183)
passar (7/7)
flicka (1/1)
finansierat (1/1)
anställningstiden (1/1)
arbetssökande (25/25)
siffror (1/1)
plötsligt (4/4)
brottsoffer (1/1)
medelst (2/2)
cyklister (1/1)
Vailla (1/1)
vid (450/450)
gjorda (1/1)
klarar (11/11)
r.f (1/1)
räntorna (1/1)
avslår (2/2)
mentalvårdstjänsternafinska (1/1)
fastställas (3/3)
flit (1/1)
vårdnadshavares (1/1)
plastföremål (1/1)
permanenta (2/2)
gångfinska (1/1)
samfund (17/17)
svensk (1/1)
Gammelstadsforsen (1/1)
handelsläroanstalten (1/1)
förete (1/1)
bostaden (62/62)
avfallsåtervinningfinska (1/1)
ons (3/3)
värnpliktiga (1/1)
nationalspråk (2/2)
kemiska (1/1)
del (65/65)
Kvarkens (1/1)
privatskolor (1/1)
socialarbete (6/6)
drog- (1/1)
skogsbruksingenjör (1/1)
franskan (1/1)
undervisningstillstånd (1/1)
minns (4/4)
fallit (3/3)
exakta (3/3)
kväll (1/1)
traumatiska (1/1)
barnskyddslagen (1/1)
Konsumentrådgivningen (1/2) konsumentrådgivningen (1)
möjligheterna (3/3)
Luksia (1/1)
sjukdomsattack (1/1)
obegränsad (2/2)
exempel (355/355)
skogen (2/2)
elever (9/9)
papperslösa (6/6)
utför (4/4)
ser (8/8)
byggdes (1/1)
hyresgäster (3/3)
förändras (1/1)
introduktion (1/1)
kultur- (2/2)
påtryckningar (1/1)
verksamhetsplanen (1/1)
sökandena (1/1)
utveckling (15/18) Utveckling (3)
ändra (6/6)
valuta (4/4)
tiotals (1/1)
syften (1/1)
kejsaren (1/1)
bostadslösas (1/1)
affären (1/1)
belopp (23/23)
tilläggsdagar (1/1)
besvara (1/1)
maskinmästare (1/1)
agera (1/1)
språk (85/85)
stadinasunnot.fi (1/1)
födelsedatum (3/3)
Avia (1/1)
urologiska (1/1)
Vandas (2/2)
tobak (1/1)
böcker (16/16)
bankernas (1/1)
Stenängens (1/1)
Vardagslivet (1/1)
responssystemet (1/1)
diplomi (1/1)
Dövas (3/3)
husbolagets (2/2)
utfärdas (1/1)
reseplaneraren (3/5) Reseplaneraren (2)
kuntoutuspsykoterapia (1/1)
FPA:s (55/57) Fpa:s (2)
avgiftsbelagd (12/12)
igång (2/2)
barnbidrag (8/9) Barnbidrag (1)
guidar (1/1)
naturen (11/11)
privatskola (2/2)
Vuokra (1/1)
skolelever (1/1)
tingsrättens (5/5)
medlemmarna (3/3)
arbetskraftsutbildningfinska (1/1)
bröstsmärtor (1/1)
Kehitysvammaisten (1/1)
fest (3/3)
Barnskyddsförbund (4/5) barnskyddsförbund (1)
etableringsanmälan (2/2)
badstränder (1/1)
fiskeområden (1/1)
färdigt (2/2)
European (1/1)
varan (1/1)
införskaffat (1/1)
hemsidorfinska (1/1)
föbund (1/1)
tiderna (1/1)
tryggat (2/2)
Äkta (1/2) äkta (1)
kontoutdrag (1/1)
understiger (1/1)
telefonnummer (8/8)
begränsar (2/2)
barnskyddslagenfinska (1/1)
juristhjälp (1/1)
företagsrådgivningen (4/4)
munhälsans (1/1)
tillståndsärende (1/1)
tandläkare (8/8)
automatik (1/1)
länder (36/36)
händerna (1/1)
Island (7/7)
spelproblemfinska (1/1)
tredje (6/6)
domstolsbeslut (4/4)
gällande (6/6)
kullfallna (1/1)
företagarnas (6/6)
anmäla (40/40)
polisstationen (6/6)
kommunikationsteknik (1/1)
anarki (2/2)
läkarmottagningen (3/3)
skattas (1/1)
ordningen (1/1)
diskriminera (3/3)
förberedande (39/41) Förberedande (2)
flesta (29/29)
svenskspråkig (8/8)
kaksoistutkinto (1/1)
dagvårdfinska (3/3)
olika (179/179)
fruktar (2/2)
ordföranden (3/3)
omskärelsen (2/2)
anmälningsblankett (1/1)
uppsägningstiden (7/7)
invandrarkunder (1/1)
nödvändiga (5/5)
aikuiskoulutuskeskus (1/1)
Björkby (2/2)
praktikant (1/1)
verksamhetsstället (1/1)
invandrafamiljer (1/1)
högtid (1/1)
höja (4/4)
sammanställts (1/1)
väljas (4/4)
registerstyrelsens (1/1)
familjerådgivning (5/5)
veta (4/4)
välgrundad (3/3)
äventyra (1/1)
immateriella (1/1)
återgå (3/3)
äktenskapsförordet (2/2)
skolåldern (21/21)
uppgifter (37/39) Uppgifter (2)
betalningskrav (1/1)
rådgivningstjänsterna (3/3)
sydkusten (1/1)
skald (1/1)
personbeteckning (31/31)
påsken (1/1)
födelsedatumet (1/1)
dagvårdsplats (8/8)
jag (54/54)
granskas (1/1)
stads (61/61)
sexuellt (7/7)
svalt (2/2)
påföljder (1/1)
skatten (2/2)
vattenkranarna (1/1)
maistraatti (16/16)
socialskyddsförmåner (1/1)
affärsverksamhet (3/3)
rutt (4/4)
frihet (1/1)
sed (2/2)
förlänga (3/3)
albanska (7/7)
goda (10/10)
fullföljer (1/1)
hygienpass (1/1)
alkohol (6/6)
orsakat (4/4)
länken (3/3)
Sinettä (1/1)
kulturhistorisk (1/1)
blind (1/1)
utbud (1/1)
barnen (25/25)
arbetsmarknadsstödets (1/1)
senioruniversitetet (2/2)
vårdnadshavaren (1/1)
vanliga (12/12)
tillämpas (6/6)
enfas (2/2)
terveysministeriö (2/2)
Alberga (1/1)
smittsamma (2/2)
yttranderätt (1/1)
skör (1/1)
närheten (4/4)
studentexamenfinska (1/1)
stadenfinska (3/3)
verotoimisto (3/3)
förtroendeman (4/4)
återflyttning (1/1)
teatrar (4/4)
betonat (1/1)
papper (5/5)
Nettineuvola (1/1)
skötare (5/5)
isländska (1/1)
mödrahemsverksamheten (1/1)
sätt (44/44)
nattcaféet (1/1)
pågå (1/1)
fysiska (4/4)
Vantaa (1/1)
tvingades (1/1)
rådgivningsbyråns (1/1)
motarbeta (3/3)
hindersprövningen (6/6)
uppväxtmiljö (1/1)
skatterelaterade (1/1)
stadshus (2/2)
firar (1/1)
tohtori (1/1)
nödcentraloperatörens (1/1)
utvisning (1/1)
kostnadsfritt (5/5)
berör (5/5)
polska (13/13)
dator (5/5)
närskola (3/3)
moderskapspenningperioden (1/1)
Nuorisosäätiö (2/2)
juridik (2/2)
porten (1/1)
hobbymöjligheterna (1/1)
förknippas (1/1)
sysselsättnings- (1/1)
tvisten (1/1)
arbetserfarenheten (1/1)
doseras (1/1)
utlandetfinska (1/1)
orsaker (8/8)
moderskapspenning (9/9)
Vandafinska (1/1)
bolsjevikregeringen (1/1)
upprätthåller (4/4)
nödnumretfinska (1/1)
skyldig (10/10)
handläggningsavgiften (1/1)
primärhälsovård (2/2)
östra (2/3) Östra (1)
modersmålsprovet (2/2)
hav (1/1)
antecknats (3/3)
personers (3/3)
vederlagets (1/1)
lånesumman (1/1)
alltså (25/25)
arbetstid (10/10)
Nimettömät (1/1)
lovade (1/1)
lön (46/46)
agerar (1/1)
inkräktar (1/1)
åldersspannet (1/1)
kriisipäivystys (3/3)
åldringspension (1/1)
examensnivån (1/1)
betalningsplan (2/2)
grundat (2/2)
pensionfinska (1/1)
gentemot (2/2)
lämnats (3/3)
mer (418/418)
Axxell (2/2)
brådskande (27/27)
bostadsbehov (4/4)
omkring (1/1)
andel (6/6)
näringfinska (1/1)
rådgivare (1/1)
make (27/27)
socialtjänst (1/1)
moderskapsledig (3/3)
försiktig (1/1)
framstegsvänligt (1/1)
reklammedel (1/1)
byar (1/1)
utlänningarfinska (3/3)
månadsskift (1/1)
fordonsskatten (1/1)
äktenskapengelska (1/1)
Suomessa (2/2)
regeringarna (1/1)
serviceställen (2/2)
vårdledigheten (2/2)
hemförsäkring (5/5)
lastenvalvoja (3/3)
hantera (2/2)
illegalt (1/1)
smarttelefonen (1/1)
ställe (9/9)
färdigheter (22/22)
graviditetsintyg (1/1)
stödbostad (3/3)
fel (12/12)
vidimerad (1/1)
närvarar (1/1)
nytta (5/5)
interna (1/1)
musiker (1/1)
bostadens (9/9)
ja (19/19)
Omnia (3/3)
kort (21/22) Kort (1)
utbildningstiden (2/2)
Hilma (1/1)
utgör (2/2)
utbildningsväsendetfinska (1/1)
utbildningsanordnare (1/1)
bankerna (1/1)
berusad (1/1)
vårdnadshavarens (1/1)
arbetsplatserna (7/7)
parrådgivning (1/1)
gammal (13/13)
definieras (4/4)
Chile (1/1)
praktiken (5/5)
in (81/85) In (4)
tjänstekollektivavtal (1/1)
arbetsmiljö (1/1)
nödfall (8/8)
tillståndsansökan (4/4)
itsenäisen (1/1)
klara (16/16)
nettolönen (1/1)
invånarnas (1/1)
avslå (1/1)
harkinnanvarainen (1/1)
royaltyn (1/1)
tillgängliga (3/3)
verket (9/9)
passa (1/1)
annans (2/2)
räkning (3/3)
minska (1/1)
riksdagsledamöter (1/1)
utredningen (3/3)
pyssel (1/1)
begravningsplatser (4/4)
undernivåer (1/1)
enda (1/1)
diskussioner (2/2)
beslutar (13/13)
innan (75/75)
familjeterapi (1/1)
kylskåpet (2/2)
hitta (28/28)
demokratin (1/1)
umgängesrätt (6/6)
helgjour (1/1)
dagen (15/15)
sälfångst (1/1)
kliniker (2/2)
socialarbetarefinska (1/1)
taxin (1/1)
stödja (2/2)
vilket (44/44)
midsommartraditionerna (1/1)
B1 (2/2)
lönar (17/17)
sö (1/1)
vinterlov (1/1)
kartläggs (1/1)
kallelsen (1/1)
grunder (9/9)
penningunderstödfinska (1/1)
föråldrade (1/1)
viktigaste (9/9)
apotek (4/4)
formella (1/1)
makas (4/4)
Kejsardömet (1/1)
barnskyddsmyndigheterna (2/2)
tvinga (8/8)
skiftarbetstillägg (1/1)
mobil (1/1)
PISA (1/1)
psykiatriskötare (1/1)
läkarens (2/2)
anknytning (2/2)
föreningens (3/3)
yrkesutövning (2/2)
tämligen (1/1)
styrka (9/9)
studiefärdigheter (1/1)
högstadiet (4/4)
simpass (1/1)
varningsmärke (1/1)
kommande (1/1)
bankkonto (14/14)
skattebyrån (13/13)
ordningsnumret (1/1)
Rösa (1/1)
urvalsbaserade (1/1)
snitt (1/1)
skapa (7/7)
integrationsutbildning (5/5)
camping (1/1)
Seure (1/1)
beskrivs (2/2)
sjukvård (8/8)
hanke (1/1)
grundandet (1/1)
övertidstillägg (1/1)
världsarv (2/2)
flyttrörelsen (1/1)
varannan (1/1)
Kafnettis (1/1)
religionsutövande (1/1)
frivilligarbete (5/6) Frivilligarbete (1)
undertecknade (1/1)
krissituationer (8/8)
hälsovårdens (1/1)
nuortenkeskus (2/2)
A2.2 (1/1)
slag (2/2)
högljudd (1/1)
skyddshem (15/18) Skyddshem (3)
barndomen (1/1)
samhällsvetenskapliga (3/3)
amorteras (1/1)
internationell (2/3) Internationell (1)
betjäna (1/1)
november (4/4)
kommunalt (3/3)
familjedagvård (2/2)
instans (3/3)
påvisa (3/3)
ekonomi- (3/3)
engelskspråkiga (3/3)
överstiga (2/2)
vanhempainvapaa (1/1)
träning (1/1)
tullens (1/2) Tullens (1)
kostnadsfri (12/12)
måla (1/1)
deltidsarbeta (1/1)
förmånligaste (1/1)
flyttat (9/9)
sida (270/270)
dömer (1/1)
förnya (4/4)
föräldralediga (1/1)
vägg (1/1)
återvänder (3/3)
daghemmen (3/3)
fattar (15/15)
evenemangskalendrarna (3/3)
möjlig (2/2)
förvänta (1/1)
polisanmälan (1/1)
finländska (60/64) Finländska (4)
spårvagnar (1/1)
ansvara (1/1)
varsel (1/1)
bostadslös (3/3)
arbetslösa (25/25)
Clinic:s (1/1)
färger (1/1)
invånarna (10/10)
relationer (1/1)
stämning (1/1)
verksamhetssätt (1/1)
territorium (2/2)
kuntoutuspäätös (1/1)
beviljandet (1/1)
rusmedel (2/2)
tisdagar (3/3)
förtroende (1/1)
jour (1/1)
tulkki (1/1)
hemlig (1/1)
upptäckt (1/1)
centrum (9/9)
databank (1/1)
skatteåterbäring (4/4)
bönder (1/1)
center (5/5)
seniorineuvonta (2/2)
undertecknas (1/1)
skaffar (6/6)
verkliga (2/2)
lokalförvaltning (3/3)
motionsrutter (1/1)
bekostat (1/1)
arbetslöshetsdagpenning (2/2)
danskonst (1/1)
eläkevakuutus (2/2)
snabba (1/1)
tuki (5/5)
län (3/3)
CV:t (2/2)
avgångsbetyget (1/1)
skyddsåldersgränsen (1/1)
jobbsökningen (11/11)
handikappbidrag (5/5)
Uusi (1/1)
studiepenningen (1/1)
historiafinska (1/1)
avlagda (1/1)
fågelbon (2/2)
prövotiden (2/2)
förteckning (5/5)
baserar (1/1)
förs (3/3)
beloppet (5/5)
fastighetsförmedlare (1/1)
skötandet (2/2)
inlärnings- (1/1)
läkemedel (25/29) Läkemedel (4)
missbruksproblem (6/7) Missbruksproblem (1)
moderskapsledigheten (5/5)
tolkcentral (3/3)
tvåspråkigt (2/2)
mångsidig (2/2)
vaginalt (2/2)
tiotusentals (2/2)
finskspråkigt (2/2)
museot.fi (1/1)
Kotoutumiskeskus (1/1)
kunna (38/38)
kejsare (1/1)
apotekets (3/3)
Helsinkis (1/1)
halsduk (1/1)
felfri (1/1)
arrangerar (1/1)
religionssamfund (4/4)
huvudansvaret (1/1)
sydkust (1/1)
ID (5/5)
uppehållstiden (1/1)
examensinriktad (1/1)
beviljades (3/3)
jokamiehen (1/1)
studentkårens (1/1)
varainsiirtovero (1/1)
Takuusäätiös (1/1)
Nylands (10/10)
betald (1/1)
tvättmaskinen (1/1)
hyresgäst (1/1)
registrering (20/29) Registrering (9)
bebiskläder (1/1)
följas (1/1)
via (103/103)
småbarnspedagogisk (1/1)
klarlägga (1/1)
ifrån (5/5)
kranvatten (1/1)
tvärtom (1/1)
stadsbiblioteken (1/1)
mognadsprov (2/2)
franska (60/60)
F (1/1)
V (2/2)
haft (7/7)
utlåtandet (3/3)
sommarteatern (1/1)
kylskåpets (1/1)
affärsförhandlingar (1/1)
väster (2/2)
lådor (1/1)
dörrklocka (1/1)
års (16/16)
slidmynningen (1/1)
pålitligt (3/3)
gymnasieutbildningen (1/1)
folkhögskolan (3/3)
perioder (5/5)
kollektivtrafikförbindelser (4/4)
ordning (2/2)
skäl (14/14)
gjorts (1/1)
viss (20/20)
fem (24/24)
rekreation (1/1)
gratis (22/22)
andelar (1/1)
vem (15/15)
läcker (1/1)
osaomistusasunto (2/2)
ansiotulovähennys (1/1)
utbytesstudenter (1/1)
rädsla (1/1)
vårdnadshavare (23/23)
radhuslägenheter (1/1)
studieplatsen (1/1)
försäkringspremier (1/1)
mödrarådgivningen (8/8)
akutvården (1/1)
stor (10/10)
kallad (2/2)
familjeplanering (5/5)
kärnkraftverksprojekt (1/1)
Schengenländer (1/1)
måltiden (1/1)
lämplighet (1/1)
ifrågavarande (4/4)
torra (2/2)
motiverat (1/1)
arbetslöshetskassor (1/1)
österut (1/1)
marknadsundersökning (1/1)
barndom (1/1)
bostadsort (2/2)
bibliotekarienfinska (1/1)
konkurrerar (2/2)
stämmor (1/1)
vetenskap (1/1)
hushållsapparater (1/1)
motionsplatserna (1/1)
reaali (1/1)
ned (6/6)
omfattande (6/6)
nybörjare (1/1)
uppfylla (3/3)
hälsostationen (38/38)
korrigerar (1/1)
igenom (5/5)
arbetsgivarna (4/4)
51:a (2/2)
el (3/3)
beslutas (5/5)
människovärde (1/1)
Verla (1/1)
ortodox (4/4)
fungera (2/2)
specialvårdspenning (1/1)
läroinrättning (2/2)
vila (1/1)
föreskriver (1/1)
Rovaniemi (42/42)
framgår (3/3)
stressyndrom (1/1)
handläggarna (1/1)
cykel (1/1)
gårdar (1/1)
inkomstrelaterade (5/5)
arbetslöshetsstöd (1/1)
utrikesministeriet (2/2)
ägs (9/9)
erfarenheter (3/3)
cirkuskonst (2/2)
arabiska (59/59)
småbarnspedagogiken (12/12)
uppehållsrätt (28/28)
Sato (2/2)
Finland (1008/1008)
flyttfirmorna (1/1)
långfredagen (1/1)
doktorsexamen (4/4)
friluftsområden (1/1)
Pensionsskyddscentralen (6/6)
vuxenutbildningscentra (1/1)
alltför (3/3)
servicebostadsgrupp (1/1)
joustava (1/1)
linjekartor (1/1)
tillfälliga (3/3)
beror (42/42)
vårdkostnader (1/1)
födas (1/1)
säsongsarbetsvisum (1/1)
skador (3/3)
nuorisoasema (1/1)
invandrarbakgrund (5/5)
kommunernas (4/4)
uppvisa (1/1)
öppnas (1/1)
läroämnen (4/4)
näringslivet (1/1)
-eller (1/1)
ordböckerfinska (2/2)
tillståndskort (1/1)
prevention (5/5)
stannar (5/5)
E101 (2/2)
räkningen (5/5)
busstation (1/1)
hälsovård (3/3)
filmer (8/8)
hälsostationer (10/10)
arkivet (1/1)
trafikerar (1/1)
finskt (30/34) Finskt (4)
dock (54/54)
stadgas (3/3)
arkitektur (2/2)
laitos (2/2)
avlidnes (2/2)
avslutade (2/2)
reseförsäkring (1/1)
landsbygd (1/1)
NewCo (5/5)
behåller (2/2)
Konsumentförbunds (1/1)
pendlar (1/1)
studiepenningens (1/1)
förman (1/1)
Villa (1/1)
varierande (1/1)
bemanningsbolag (1/1)
Nationalgalleriet (1/1)
självrisken (2/2)
praktik (4/4)
diskrimineringen (1/1)
valkretsen (1/1)
arbetspensionsutdragen (1/1)
godtagbar (3/3)
Asokoditfinska (2/2)
tysta (4/4)
utbytesstudent (2/2)
yrkesprov (1/1)
HRT (3/3)
köper (13/13)
företagsformerfinska (1/1)
språkanvändares (2/2)
penningspelproblemfinska (1/1)
utbildningslinjer (1/1)
överenskommelsen (3/3)
inredning (1/1)
skattepliktig (2/2)
utbudet (3/3)
leker (1/1)
mikrovågsugnen (1/1)
tillåtelse (1/1)
snart (1/1)
käyttövastike (1/1)
uppehållstillståndfinska (6/6)
mammor (1/1)
kortvarig (4/4)
sexåringar (2/2)
bildar (1/1)
köpt (3/3)
parten (3/3)
inrättas (1/1)
mobilcertifikat (3/3)
ansökningstid (1/1)
samtalspriset (1/1)
elektrisk (2/2)
bestämd (4/4)
rasistiskt (5/5)
anlitar (1/1)
folkpensionerna (1/1)
intygen (1/1)
arbetarskyddsfullmäktige (2/2)
idrottshobbyer (1/1)
stater (2/2)
överlåtits (1/1)
klubbar (6/6)
ner (4/4)
bortgång (1/1)
anställningsvillkor (1/1)
modersmålsundervisningen (1/1)
handelsregistret (2/2)
någonting (2/2)
före (52/52)
tvillingar (1/1)
tider (10/10)
trossamfund (5/5)
prick (1/1)
ungdomsgrupper (1/1)
kuntoutussuunnitelma (1/1)
hotar (9/9)
remixa (1/1)
språket (50/50)
verksamheten (14/14)
umgängesrättfinska (2/2)
avoimet (2/2)
Project (1/1)
undersökningarna (5/5)
visas (5/5)
vårdfinska (1/1)
stödspråkfinska (1/1)
RAMK (2/2)
invandrarbyrån (4/4)
konstmuseum (2/2)
FRK:s (1/1)
tågtidtabellerna (1/1)
målet (4/4)
Vuxeninstitut (1/1)
lukio (4/4)
data- (1/1)
Gustav (3/3)
TTS (1/1)
rörande (3/3)
eventuellt (11/11)
Seremoniat (1/1)
arbetslivetfinska (1/1)
bussar (4/4)
möter (1/1)
officiell (4/4)
Poikien (1/1)
vigselfinska (2/2)
inspiration (1/1)
sättas (1/1)
förskolan (4/4)
biljettpriserna (2/2)
avfallshanteringen (1/1)
texttelefon (1/1)
femte (2/2)
sukupuolitautien (1/1)
festmat (1/1)
ändamålet (1/1)
hälso- (20/20)
bilda (1/1)
fisketillståndfinska (1/1)
näringsbyråerfinska (1/1)
sortering (1/1)
svår (5/5)
dit (6/6)
mousserande (1/1)
målsättningar (1/1)
skilsmässan (5/5)
arbetsgivarförbundet (1/1)
ringa (58/58)
vise (1/1)
kunskaper (27/27)
dagars (1/1)
ungdomsfullmäktige (1/1)
slovakiska (1/1)
ångest (1/1)
mellanrum (4/4)
planering (2/2)
blivande (3/3)
föras (2/2)
rehabiliteringscenter (1/1)
viseringspliktigt (1/1)
lärandet (1/1)
ledda (2/2)
skadligt (1/1)
temadagar (1/1)
studiemöjligheter (5/5)
avtalas (1/1)
förlorar (3/3)
vårdinrättning (2/2)
nutidskonst (1/1)
nivå (7/7)
Helsinki (11/11)
nedsatt (1/1)
apoteket (8/8)
nationalmuseumfinska (1/1)
borgerliga (1/1)
boenderegistret (2/2)
studiestödetfinska (1/1)
växlande (1/1)
yttrandefrihet (1/1)
påtryckning (1/1)
dem (64/64)
Näringsliv (3/3)
rädd (3/3)
familjebandfinska (2/2)
innehåll (5/5)
äktenskap (52/54) Äktenskap (2)
åldrarna (2/2)
jourmottagningfinska (1/1)
allaktivitetscentret (1/1)
bärbar (1/1)
muovi (1/1)
kvällar (6/6)
dagvårdsenhet (1/1)
beslutsfattandet (6/6)
handpenning (1/1)
rätt (226/226)
regionen (3/3)
järnvägsstation (1/1)
handskar (1/1)
miljö- (1/1)
romanifinska (1/1)
oppisopimuskoulutus (1/1)
centralsjukhuset (1/1)
flyktingläger (2/2)
uppleva (1/1)
aktiva (5/5)
D (1/1)
beräknade (6/6)
vapaarahoitteinen (1/1)
hjälpmedel (18/18)
högklassiga (1/1)
sjukvårdsersättningar (1/1)
undersökning (8/8)
mångkulturellt (2/2)
talets (1/1)
utsända (1/1)
avgöras (1/1)
avvika (3/3)
nu (1/1)
bilskatten (1/1)
hyresvärden (18/18)
släkten (1/1)
uppehållstillstånden (1/1)
delegation (1/1)
besvärsanvisning (1/1)
inriktning (1/1)
saknar (6/6)
kyrkor (1/1)
linkkiLaNuti (1/1)
arbetstider (5/5)
gymnasiernas (1/1)
telefonservice (2/2)
EVK (1/1)
belönas (1/1)
uppfyllas (1/1)
webbapotek (1/1)
betraktar (1/1)
yrkeshögskoleexamenfinska (1/1)
lapsikaappaus (1/1)
linkkiMiljöministeriet (1/1)
www.kopiosto.fi (1/1)
upphörande (2/2)
samverkan (1/1)
godkännande (1/1)
hushållets (1/1)
typ (4/4)
språkkurserna (1/1)
Sveriges (2/2)
återkallats (2/2)
mielenterveysseuran (1/1)
skrivna (1/1)
funderingar (1/1)
sjuksköterska (2/2)
demonstration (1/1)
farlig (1/1)
utfärdar (2/2)
sköter (23/23)
hot (12/12)
konflikter (5/5)
säsongtopp (1/1)
nyligen (5/5)
olycksfallsstation (2/2)
gränser (2/2)
sysslorna (3/3)
kandiderar (1/1)
skötaren (2/2)
grundlagenfinska (1/1)
uppstartsföretagarefinska (1/1)
avgångsbetyg (5/5)
föds (18/18)
slutat (1/1)
avträdelseanmälan (1/1)
fönstren (2/2)
besöket (3/3)
Yrittäjän (1/1)
ehkäisyneuvonta (1/1)
sederengelska (1/1)
varor (5/5)
kombinerat (5/5)
bifogas (1/1)
Förbund (5/5)
tolv (6/6)
sökningen (1/1)
lagman (1/1)
överhuvudtaget (1/1)
sällskapande (3/3)
VALMA (13/13)
Infobank (1/1)
asylansökningsblankett (1/1)
status (1/1)
råd (89/89)
hyresbostadfinska (1/1)
Monika (3/3)
museer (10/10)
ärva (2/2)
kapital (2/2)
bastuugn (2/2)
ländernafinska (1/1)
placera (2/2)
hindersprövning (5/5)
studerat (3/3)
möjliggör (1/1)
tingsdomare (1/1)
når (1/1)
viken (3/3)
materialet (4/4)
delarna (2/2)
nämna (1/1)
hotfull (1/1)
beskickningarna (1/1)
bara (13/13)
psykoterapin (1/1)
fatta (5/5)
därmed (2/2)
skidåkningfinska (1/1)
mäklararvode (1/1)
sköts (4/4)
förmåner (28/28)
innehåller (14/14)
godkänner (4/4)
teckenspråkstolk (1/1)
fax (3/3)
annonsen (2/2)
gymnasieutbildningfinska (1/1)
förvärvsinkomstavdrag (1/1)
utrikesministeriets (4/4)
tillsätter (1/1)
tingsrätt (3/3)
användarpanel (2/2)
pojken (2/2)
sairausvakuutus (4/4)
läkarcentral (1/1)
inskrivet (1/1)
sjukdomstid (2/2)
kollektiv (1/1)
orolig (2/2)
har (1057/1057)
uppehålla (1/1)
handikapprådgivningen (2/2)
samfunden (1/1)
kravet (3/3)
främst (5/5)
ansvariga (5/5)
överlåtelse (1/1)
tillfrisknande (1/1)
finlandssvenska (2/2)
tillfälle (1/1)
rådgivningspunkt (1/1)
födseln (4/4)
föreskrivs (2/2)
filosofi (1/1)
försenade (2/2)
angett (1/1)
efternamnen (1/1)
legaliseras (4/4)
nioårig (1/1)
huvudsakliga (1/1)
arbetsplatser (13/13)
former (4/4)
statligt (1/1)
arbetslöshetskassa (9/10) Arbetslöshetskassa (1)
företagstjänster (1/1)
barnskyddet (4/4)
trauma (1/1)
vardagssysslor (2/2)
årfinska (2/2)
växande (1/1)
lös (1/1)
osakligt (3/3)
kvarskatt (3/3)
kastrullock (1/1)
thai (10/10)
förplikta (1/1)
slutsyn (1/1)
Nordplus (1/1)
namnen (3/3)
platsansökan (1/1)
naken (1/1)
rättshjälpsbyrå (10/10)
Koivuhaan (1/1)
kundrådgivningen (1/1)
mellanskillnaden (1/1)
musikverksamhet (1/1)
perheneuvola (6/6)
makars (1/1)
älvar (1/1)
taasengelska (1/1)
villasamhället (1/1)
Sverige (16/16)
följebrev (1/1)
Europaparlamentsvalet (1/1)
socialtjänster (4/4)
valkrets (1/1)
ställningen (1/1)
alls (1/1)
stapelrättigheter (1/1)
skäliga (4/4)
smittats (1/1)
insjöarna (1/1)
rikt (1/1)
familjeband (25/25)
starkt (2/2)
kontakter (2/2)
skattenummer (5/5)
verkosto (1/1)
nödinkvartering (2/2)
kaffesump (1/1)
underhålls (1/1)
husfinska (2/2)
skiljer (5/5)
samtalshjälp (4/4)
smidig (1/1)
familj (22/22)
ägarbostäderfinska (2/2)
lottar (1/1)
Pensionsskyddscentralens (1/1)
tidsbunden (2/2)
pensioner (2/2)
simma (1/1)
psykoterapeutens (1/1)
framskrider (3/3)
lånegaranti (1/1)
samtals- (1/1)
detsamma (1/1)
hemvård (6/6)
papperspåsar (1/1)
inhämta (4/4)
täckande (1/1)
insatt (2/2)
framhäver (1/1)
tåg- (1/1)
intelligenta (1/1)
konfidentiellt (3/3)
kompletterar (2/2)
publicera (1/1)
nivån (5/5)
Avara (2/2)
ansiotulo (1/1)
kosta (1/1)
upprätthållande (1/1)
myndiga (2/2)
matkakortin (1/1)
juridisk (7/7)
valts (1/1)
placeras (1/1)
klassificerats (1/1)
cykelleder (1/1)
resehandling (2/2)
säkring (1/1)
förmyndarskap (2/2)
stöttar (1/1)
faderskapsärendet (1/1)
förmånlig (2/2)
ungas (26/26)
skuldlinjen (1/1)
hette (1/1)
mentalvårdsenheten (1/1)
vårdledighet (4/4)
Esbobor (1/1)
flygstationen (1/1)
musikinstitut (3/3)
koppling (1/1)
besvarar (2/2)
samboförhållande (14/16) Samboförhållande (2)
bostadsbidrag (20/25) Bostadsbidrag (5)
söka (138/138)
gåva (1/1)
kompletterande (2/2)
isännöitsijä (1/1)
revisionsbyråer (1/1)
integrations- (2/2)
umgänget (4/4)
banklån (4/4)
Hollihaan (1/1)
Rinteenkulma (1/1)
chefer (1/1)
skolor (18/18)
erillinen (1/1)
verben (1/1)
ekonomisk (1/1)
sistone (1/1)
psykiskt (1/1)
åsikt (8/8)
Hakunilan (1/1)
arbetslivet (20/20)
aktörerna (1/1)
ihåg (25/25)
specialundervisningen (1/1)
peruspäiväraha (1/1)
ange (8/8)
Västra (8/11) västra (3)
låta (7/7)
perioden (2/2)
förföljelse (2/2)
förmodligen (1/1)
specialvårdpenning (2/2)
Rovala (2/2)
väsentlig (3/3)
balansera (1/1)
finskakurser (3/3)
handikappade (35/36) Handikappade (1)
centralmuseetfinska (1/1)
barnklubbar (3/3)
startpaket (1/1)
barnfostran (1/1)
medlemsfamiljerna (1/1)
umgängesarrangemanget (1/1)
utbildnings (1/1)
gymnasiumfinska (1/1)
fackliga (1/1)
företaget (18/18)
kuljetuspalvelu (1/1)
hyresbostad (33/35) Hyresbostad (2)
jourtelefon (1/1)
förvärvsarbete (2/2)
migration (1/1)
statens (9/9)
invandrartjänster (1/1)
religiöst (9/9)
servicenummer (1/1)
förvärvsinkomster (1/1)
mediciner (2/2)
stöds (1/1)
akademiskt (1/1)
samlar (1/1)
önskemål (6/6)
motionfinska (1/1)
uppstå (1/1)
islamska (1/1)
chattenfinska (1/1)
personaltjänsteföretag (1/1)
företagsservicecentralerna (1/1)
registerstryrelsen (1/1)
döden (1/1)
måltider (4/4)
Verso (1/1)
papprullar (1/1)
åtföljs (2/2)
England (1/1)
flexibel (7/7)
respekteras (1/1)
tvåspråkig (1/1)
infödd (4/4)
cykelvägar (2/2)
Tölö (2/2)
etablerades (2/2)
beroende (10/10)
verohallinto (1/1)
tullanmälan (1/1)
krav (4/4)
tandvårdens (2/2)
rättshjälp (5/5)
graviditetsprevention (2/2)
avfallshanteringfinska (1/1)
älv (1/1)
föddes (1/1)
avsnitten (1/1)
spara (2/2)
ryskaryska (1/1)
hemhjälpfinska (1/1)
helhetsbetonat (1/1)
religionstillhörigheten (1/1)
val (13/16) Val (3)
snittbetyg (1/1)
problematiskt (1/1)
frånvaro (1/1)
Medelhavet (1/1)
mental- (2/2)
leta (7/7)
sammanhang (2/2)
Bottniska (2/2)
sjukvårdskortet (6/6)
partiella (3/3)
föräldrarfinska (1/1)
gift (12/12)
barnomsorgen (1/1)
grannmedlingscentret (1/1)
språkkursernas (1/1)
orättvist (1/1)
program (8/8)
erhålla (3/3)
tillhandahålls (9/9)
sjukvårdskortetfinska (2/2)
fostran (18/21) Fostran (3)
anstaltsvårdenfinska (1/1)
prövotid (1/1)
stadsrättigheter (1/1)
klarspråk (1/1)
College (1/1)
beviljande (1/1)
priser (5/5)
arbetsinkomst (2/2)
info (8/8)
boendeservice (2/2)
serviceplanen (1/1)
stadsmuseum (1/1)
stipendiesystem (2/2)
Kuluttajansuojalaki (1/1)
kvinnlig (2/2)
vammaistuki (2/2)
adresserna (1/1)
växer (2/2)
Silkesportens (1/1)
metrostationer (1/1)
kouluterveydenhoitaja (1/1)
flyktingbakgrund (1/1)
förlossningsdatum (1/1)
hyresförhållandet (2/2)
skyddshusfinska (2/2)
toimintaohjelma (1/1)
finansieringsalternativ (3/3)
kansalaisopisto (2/2)
framföra (2/2)
samtycke (4/4)
genomförs (2/2)
kölapp (1/1)
diabetesfinska (1/1)
vistelsen (4/4)
sjöar (1/1)
linjen (1/1)
klient (1/1)
församling (7/7)
hemvårdens (5/5)
kuntoutus (2/2)
specialkompetens (1/1)
snabel (1/1)
skattefria (1/1)
näringstjänsterfinska (2/2)
öppettiderfinska (2/2)
Kristinestad (1/1)
reparera (1/1)
stödformer (1/1)
morgon (2/2)
prövning (11/13) Prövning (2)
folkhögskola (2/2)
funktionell (1/1)
tilläggsinformation (1/1)
föreslår (3/3)
rabatter (1/1)
fackförbundsverksamhetfinska (2/2)
veckan (4/4)
skattar (1/1)
rehabiliteringen (5/5)
stöder (8/8)
blev (17/17)
vilkas (1/1)
hemfriden (1/1)
ibruktagande (1/1)
heltidsstuderande (1/1)
meritförteckning (5/5)
släktens (1/1)
vädra (1/1)
biblioteken (6/6)
vitsorden (1/1)
läget (1/1)
mot (36/36)
forskarefinska (1/1)
passfinska (1/1)
Företagsfinlands (2/3) FöretagsFinlands (1)
www.gramex.fi (1/1)
vuxengymnasierna (1/1)
händelser (5/5)
antagningen (1/1)
mottagningscentral (4/4)
advokater (1/1)
centrala (8/8)
brottsmålsvittnen (1/1)
sambon (4/4)
tobaksprodukter (1/1)
bokföring (1/1)
kulturell (1/1)
oktoberrevolutionen (1/1)
boendefinska (1/1)
tideräkningen (1/1)
sidan (36/36)
arbetsintervju (1/1)
Bio (1/1)
arbetsintyget (2/2)
proffs (2/2)
partner (12/12)
hans (10/10)
styrkorna (1/1)
funktionsnedsättning (7/7)
skadats (4/4)
het (1/1)
nyfödda (1/1)
integrationsplaner (1/1)
hembesök (2/2)
sömnskola (1/1)
församlingssammanslutnings (2/2)
sjukdagpenningen (3/3)
freden (1/1)
Jesu (3/3)
resenärerfinska (1/1)
besluta (10/10)
ortodoksinen (1/1)
oljud (3/3)
fritidsaktiviteter (3/3)
intyg (26/26)
UNHCR (4/4)
taget (3/3)
rådgivning (54/54)
barnförhöjning (1/1)
hålla (4/4)
alle (1/1)
servicecentret (1/1)
yrkesskolorna (1/1)
teknisk (1/1)
teaterfinska (1/1)
Finlands (67/67)
Håkansböle (6/6)
emellertid (9/9)
bastuugnen (3/3)
utbildade (4/4)
äitiyspakkaus (1/1)
likadant (1/1)
kansainvälinen (1/1)
bifaller (1/1)
industrialiserades (1/1)
dödsfallet (1/1)
cirka (31/31)
föreläsningsserier (1/1)
centralförbund (1/2) Centralförbund (1)
relationsrådgivning (2/2)
befolkningsdataregistret (1/1)
polisstation (1/1)
Infobanken (5/5)
bidraget (2/2)
bekantskaper (1/1)
bygga (6/6)
Åbo (7/7)
speciell (2/2)
bekräftar (5/5)
produkter (5/5)
uppvärmningen (1/1)
stödtjänster (6/6)
konstaktiviteter (1/1)
parkeringsbiljett (1/1)
filmens (1/1)
inhemska (3/3)
uppskatta (4/4)
avlidne (4/4)
kopior (2/2)
Medborgarrådgivning (1/1)
verifieras (1/1)
långa (6/6)
andelslaget (1/1)
skedet (1/1)
svar (1/1)
bostadsvisning (2/2)
födelsen (1/1)
färdtjänst (7/7)
montera (1/1)
bevittnat (1/1)
EMMA (1/1)
utbetalad (2/2)
angelägenheter (5/5)
bostadsrättsavgifter (1/1)
vardagar (17/17)
avtal (30/30)
igen (2/2)
webbtjänst (9/9)
identitetsbevis (8/8)
nättjänsten (2/2)
tandhälsan (1/1)
verkstäder (1/1)
varmare (1/1)
kunden (6/6)
päivystys (3/3)
socialväsendet (1/1)
handikappservicefinska (4/4)
hindi (1/1)
Europaparlamentsvalfinska (1/1)
bibliotekfinska (1/1)
hautaustoimisto (2/2)
barnlöshetspolikliniken (1/1)
vårdenhet (2/2)
underleveransarbete (1/1)
salu (3/3)
familjepensionsskydd (1/1)
regioner (1/1)
bostäder (38/38)
politiskt (1/1)
närvara (1/1)
åtagit (1/1)
existerande (1/1)
telefontjänsten (6/6)
bostadsrättsavtal (1/1)
ungdomsbostäder (5/5)
Närpes (1/1)
samtalet (5/5)
tjänsteman (1/1)
livsmedel (2/2)
system (3/3)
yrkesläroanstalter (6/6)
underhåller (1/1)
avgör (3/3)
lagen (26/26)
opetuksen (1/1)
hurdan (2/2)
farföräldrar (2/2)
hoppat (1/1)
kostar (12/12)
stadssund (1/1)
helst (23/23)
ovanför (2/2)
problemet (1/1)
betjänas (1/1)
värden (1/1)
efterhand (5/5)
bilskatt (1/1)
ställt (2/2)
kandidat- (1/1)
upphävs (2/2)
karaoke (1/1)
vederlag (2/2)
rådgivningstelefon (1/1)
fuktisolering (1/1)
lampa (1/1)
CVfinska (2/2)
hela (27/27)
aluekoordinaattori (2/2)
insinööri (1/1)
vuxensocialarbetetfinska (1/1)
kartläggning (17/17)
territoriet (3/3)
behov (38/38)
jämlika (1/1)
efternamnfinska (1/1)
registret (1/1)
markägarna (1/1)
text (1/1)
utbildningens (1/1)
offentliggöra (1/1)
rådgivningsbyrå (2/2)
torteras (1/1)
Villenpirtti (1/1)
bl.a. (7/7)
isär (3/3)
bioavfall (2/2)
huset (4/4)
hälsafinska (2/2)
avtalsperioden (1/1)
Flyktingrådgivningen (3/3)
Galoppbrinken (1/1)
tulosyksikkö (1/1)
innehållen (1/1)
toimisto (4/4)
skattedeklaration (1/1)
vilja (1/1)
lettiska (1/1)
skidspår (2/2)
Karl (1/1)
tidsbegränsade (1/1)
torgsidan (1/1)
asunnotfinska (1/1)
socialservicecenter (1/1)
textade (1/1)
Vinge (2/2)
bostadsförmedlingen (1/1)
innebär (20/20)
familjeträning (1/1)
bolagsavtal (1/1)
upprättat (3/3)
SOA (1/1)
giltig (2/2)
sidorna (9/9)
asumisoikeusmaksu (1/1)
abortti (1/1)
allvarliga (1/1)
kundtjänst (1/1)
nyttig (8/8)
matkakortti (2/2)
Metropolia (1/1)
olycksfallsförsäkring (3/3)
elapparat (2/2)
Setlementti (7/7)
tretton (1/1)
läsåret (2/2)
webben (2/2)
beskickning (16/16)
kvinnor (34/34)
anhörigafinska (1/1)
läggas (1/1)
industrialiseringen (2/2)
Pakolaisneuvonta (2/2)
förmånen (1/1)
fakturor (1/1)
servicestället (10/10)
rekommendabelt (1/1)
Nylandfinska (1/1)
4:e (2/2)
bekymmer (1/1)
genomför (1/1)
öppenvården (1/1)
upplysningar (2/2)
lättföretagande (1/1)
lägenheter (1/1)
köa (1/1)
regelbundet (5/5)
säsongsarbetstillstånd (1/1)
förvärvsrelaterad (1/1)
administrerar (1/1)
makarfinska (1/1)
mopedkort (1/1)
arbetsgivarförbunden (1/1)
omständighet (1/1)
tillståndsansökningarfinska (1/1)
uppföljning (1/1)
Jorv (10/10)
räddningsverk (1/1)
fanns (3/3)
hemlika (1/1)
bekymrar (1/1)
regionförvaltningsverk (1/1)
uppehållstillståndet (14/14)
rummet (1/1)
yhdenvertaisuus- (1/1)
bröllopsdagen (1/1)
Företagsfinland (1/1)
Helsingin (5/5)
teckenspråket (1/1)
stå (1/1)
intressebevakningsorganisationfinska (1/1)
rundvandringar (2/2)
ammattitutkinto (1/1)
danska (2/2)
förnamn (1/1)
spänning (2/2)
yrkeshögskolan (9/10) Yrkeshögskolan (1)
utmärkt (1/1)
arbetarinstitutets (1/1)
undantagsfall (4/4)
företagare (51/54) Företagare (3)
fast (10/10)
Mellersta (11/13) mellersta (2)
inhyste (1/1)
drag (1/1)
medlare (2/2)
konstskola (1/1)
pepparkakor (1/1)
psykologhjälp (1/1)
finansieringsbolag (1/1)
annonser (4/4)
sjukledigheten (3/3)
leva (6/6)
ryska (146/146)
guldåldern (1/1)
Linja (7/10) linja (3)
Sveaborgsfärjorna (2/2)
Sovjetunionen (8/8)
giltigt (12/12)
förlängning (2/2)
kyrkan (21/21)
särskild (6/6)
värkjouren (1/1)
förlossningssjukhus (1/1)
snöar (1/1)
Finlex (2/2)
bikulturella (1/1)
telefonnumret (2/2)
löneutbetalningfinska (1/1)
garantin (1/1)
vuxenutbildningsstöd (1/1)
biblioteketfinska (2/2)
läkarstationfinska (1/1)
Internetfinska (8/10) internetfinska (2)
disponent (2/2)
exceptionellt (2/2)
medborgarskap (70/70)
kväv (1/1)
midsommar (1/1)
högre (26/26)
koncernen (1/1)
förläggning (1/1)
lagstadgad (2/2)
medlemmars (2/2)
mellannivån (1/1)
politisk (2/2)
ges (42/42)
nyttigt (2/2)
brottfinska (1/1)
humanistiska (4/6) Humanistiska (2)
konst- (1/1)
webbutik (1/1)
museet (3/3)
bostadsaktiebolag (5/5)
mental (8/9) Mental (1)
kartor (1/1)
anpassningsbara (1/1)
äts (1/1)
förvärvat (2/2)
hemort (17/17)
terminen (1/1)
www.infopankki.fi (1/1)
undervisningsväsendet (1/1)
tävlingsarrangören (1/1)
egentliga (4/4)
klinikstiftelsens (2/2)
hyresbostaden (2/2)
jourtelefonen (2/2)
speciellt (9/9)
stödmottagarens (1/1)
undervisningssektorn (1/1)
Trapesa (2/2)
punktlighet (3/3)
motionsspår (1/1)
AUS (1/1)
arbetslöshetskassafinska (1/1)
stunderna (1/1)
språkkaféer (1/1)
originalhandlingen (1/1)
adoptera (1/1)
Musikantitfinska (1/1)
dagvård (10/11) Dagvård (1)
Helsingfors (169/169)
avlopp (2/2)
lämplig (14/14)
gifter (4/4)
Bostadslöshet (1/1)
Ab (2/2)
växter (1/1)
gynekologiska (2/2)
snabbare (3/3)
hälsosam (1/1)
pris (6/6)
högskolekoncern (1/1)
Religionerna (1/1)
arbetsavtalet (15/15)
universitets (3/3)
uppfattning (1/1)
planerad (1/1)
elinkeinotoimisto (4/4)
samman (2/2)
Lumon (2/2)
kvadratmeter (2/2)
våldet (1/1)
Kela (11/11)
kunnat (2/2)
delbeslut (3/3)
Myyrinki (1/1)
arvsskatt (1/1)
hyrsvärden (1/1)
anledning (5/5)
post (32/32)
områdeskoordinatorerna (1/1)
vandra (1/1)
krama (1/1)
arrangerades (1/1)
överenskommen (1/1)
Renlunds (1/1)
köparen (2/2)
hälsovårdarens (3/3)
förebyggandet (1/1)
meddelats (1/1)
arbetsgivarförbund (1/1)
viseringsfria (1/1)
undervisar (4/4)
närståendevårdfinska (6/6)
flyktingens (1/1)
samarbetar (1/1)
konkreta (1/1)
delägarbostad (2/3) Delägarbostad (1)
pensionens (1/1)
potilasasiamies (2/2)
återhämta (2/2)
förtroendemannen (4/4)
förflutit (1/1)
Oy:s (6/6)
faktor (1/1)
kortvarigt (1/1)
förskoleundervisning (14/15) Förskoleundervisning (1)
inledningsvis (1/1)
erfarenhetstillägg (1/1)
gemensamma (37/37)
vetenskaplig (1/1)
legitimerad (1/1)
slutar (9/9)
utbildningarfinska (2/2)
jurist (14/14)
lunch (3/3)
stöd (81/92) Stöd (11)
skol- (1/1)
flyktingstatus (16/16)
evankelis (1/1)
misstag (1/1)
ljudböcker (2/2)
fallet (2/2)
slås (1/1)
förskolebarn (2/2)
individuellt (3/3)
familjeskäl (4/4)
flaggan (2/2)
nätverka (1/1)
likvärdiga (2/2)
avgiftsbelagda (9/9)
häxor (1/1)
boningsort (1/1)
wc (1/1)
friluftsmuseumfinska (1/1)
form (11/11)
övervaka (1/1)
variera (4/4)
semesterresor (1/1)
avlidna (4/4)
ersättas (1/1)
skolhälsovårdarna (1/1)
barnkapning (1/1)
krisen (1/1)
måndagar (3/3)
aktiveringsmodellen (1/1)
Wien (2/2)
adoption (3/3)
yrkesinstitut (8/8)
påverkas (7/7)
tolkningen (8/8)
Huvudstadens (3/3)
anges (11/11)
biIdkonstskola (1/1)
frågor (51/51)
äldre (14/19) Äldre (5)
uppvisande (1/1)
språkexamen (10/10)
istiden (1/1)
exempelvis (15/15)
föreningsmöten (1/1)
använd (2/2)
utvecklingsstörd (3/3)
sökas (4/4)
lördagar (1/1)
enskild (4/4)
återförenas (1/1)
ordna (23/23)
bli (27/29) Bli (2)
medborgarna (2/2)
antagen (4/4)
företagaren (5/5)
rusmedelsbruk (1/1)
måsta (1/1)
diskrimineras (6/6)
plastprodukter (2/2)
telefontjänster (1/1)
verksamma (5/5)
återvinningsstationer (1/1)
intagning (1/1)
billigaste (1/1)
julstjärnor (1/1)
Pääkaupungin (2/2)
unga (72/72)
kontakt (51/51)
ungdomsstation (1/1)
avsätta (1/1)
stödpersonen (1/1)
stiftar (1/1)
nödsituationer (8/8)
valt (1/1)
sociala (74/74)
pension (16/17) Pension (1)
snö (1/1)
motionsslingor (3/3)
täcker (3/3)
inkomstgräns (1/1)
abikurssi (1/1)
hörde (2/2)
Smith (2/2)
krisarbetare (1/1)
plastförpackningar (1/1)
ansökt (4/4)
utser (3/3)
förpackningen (1/1)
institut (6/6)
den (588/602) Den (14)
psykiater (1/1)
Suomenlinna (1/1)
dagsgymnasierna (1/1)
sysselsättningen (1/1)
familjemedlemmen (1/1)
korttidsvård (1/1)
värdegrunden (1/1)
behandlar (4/4)
ambassaden (1/1)
ändå (25/25)
upprätta (6/6)
förbjuder (5/5)
YH (2/2)
adressen (10/10)
yrityksen (1/1)
examen (68/68)
livssituationen (1/1)
utrikesflygen (1/1)
omfatta (5/5)
vore (2/2)
budskap (1/1)
barnlöshetsklinik (1/1)
åtta (3/3)
hurdant (4/4)
öarna (2/2)
förverkligandet (1/1)
årervinns (1/1)
föräldraledighet (2/2)
tävlingen (4/4)
våningen (4/4)
bevisa (6/6)
stödåtgärder (1/1)
förlorade (2/2)
träna (1/1)
godkänns (3/3)
mångsidigt (1/1)
järnvägsstationer (1/1)
anmälan (25/25)
finsk (51/51)
motionsmöjligheter (2/2)
resor (2/2)
kielenkäyttäjän (2/2)
himmelsfärdsdag (1/1)
blommor (2/2)
telefonabonnemang (1/1)
varav (6/6)
väst- (2/2)
dagvårdens (2/2)
grunderfinska (1/1)
skollov (1/1)
Oma (1/1)
chef (8/8)
gången (2/2)
sommaruniversitetetfinska (1/1)
bestämmanderätt (1/1)
beslutsmakt (1/1)
paret (2/2)
sin (75/75)
våldsamt (3/3)
kulturcentret (1/1)
ju (1/1)
uppringd (2/2)
Sveaborgs (1/1)
här (32/32)
maistraatti.fi (2/2)
tukipiste (2/2)
inloggning (1/1)
studieresor (1/1)
oavlönad (3/3)
automatiskt (7/7)
examensnivå (1/1)
utbildningssystemet (1/1)
parterna (7/7)
fornlämningsområde (1/1)
inskolning (3/3)
fungerande (1/1)
mottagning (4/4)
utlåtande (9/9)
loven (1/1)
motionslokaler (1/1)
skatterna (1/1)
kvällstid (4/4)
PUK (1/1)
specialsmåbarnspedagogiken (1/1)
undersida (1/1)
oppisopimustoimisto (1/1)
tull (1/1)
allmänhet (10/10)
förvaltningsrätten (1/1)
översättningen (4/4)
informationsförmedlare (1/1)
digital (1/1)
omgivningen (1/1)
kapitalinkomsten (1/1)
konsumenträttigheterfinska (1/1)
avgiftsfri (10/10)
rörelsenedsättning (2/2)
handlingar (11/11)
beskickningen (14/14)
faktureringstjänst (1/1)
texter (1/1)
universitets- (1/1)
Kylämajafinska (1/1)
platsen (1/1)
detalj (1/1)
pensionsanstalten (1/1)
utbildningsprogrammet (1/1)
brottsanmälanfinska (1/1)
kulturevenemang (1/1)
tillgång (5/5)
användning (2/2)
beviljas (36/36)
oavlönat (1/1)
regler (5/5)
högskolexamenfinska (1/1)
ända (3/3)
bensinstationer (2/2)
slottfinska (1/1)
jourens (1/1)
barnfinska (7/7)
juridiskt (2/2)
återflyttare (2/2)
näringsbyråerna (4/4)
rehabiliteringsbeslut (1/1)
tidtabellerfinska (1/1)
backe (1/1)
dåligt (1/1)
emot (13/13)
kommunalskatt (1/1)
nog (1/1)
ansökningen (7/7)
affärsidén (2/2)
frispråkighet (1/1)
samlingar (3/3)
Laurea (2/2)
områdena (1/1)
rådgivningsbyråerna (3/3)
tandklinik (4/4)
harmoniska (1/1)
Europaskolan (1/1)
underhållsbehov (3/3)
resedokumentfinska (1/1)
Isyysraha (1/1)
operationen (5/5)
Brottsofferjouren (4/5) brottsofferjouren (1)
pensionsskyddet (2/2)
kalendern (1/1)
kämpade (1/1)
Kyllönen (2/2)
tillstånd (57/57)
yrkenfinska (1/1)
självrisktid (2/2)
anhålla (1/1)
utesluta (1/1)
skriftligen (2/2)
finskafinska (2/2)
fastighetsägare (1/1)
näringstjänsten (1/1)
skadan (2/2)
isolering (1/1)
fler (10/10)
skyddfinska (4/4)
transformera (1/1)
yrkesläroanstalterfinska (1/1)
svenskspråkiga (10/10)
någondera (3/3)
människohandelns (2/2)
Elfvik (1/1)
Myyrinkis (1/1)
lära (21/21)
klockslaget (1/1)
avslutar (1/1)
telefonen (2/2)
poliklinikka (3/3)
klass (5/5)
timmarna (1/1)
stödcentret (3/3)
moderna (1/1)
tryckta (1/1)
föräldradagpenningens (1/1)
tillhandahållas (1/1)
invalidpension (4/4)
skaka (1/1)
vån (14/14)
rubrik (1/1)
uppehållskort (5/5)
komplettera (2/2)
åligger (2/2)
förändringar (2/2)
anställningsrådgivningen (1/1)
förgiftningfinska (1/1)
Esbofinska (3/3)
bilagor (6/6)
brandlarm (1/1)
sång (1/1)
inskärper (1/1)
ordnar (66/66)
organiserade (1/1)
ersättningen (1/1)
dispens (2/2)
Vantaan (10/10)
välfungerande (1/1)
medför (1/1)
Olofsborg (1/1)
uppföljningen (1/1)
mamman (1/1)
flexibla (1/1)
invid (1/1)
perukirja (1/1)
försämrar (1/1)
hektar (1/1)
arbetafinska (2/2)
anledningar (1/1)
skolbarnfinska (3/3)
bokar (11/11)
markägaren (1/1)
dyrt (1/1)
läge (1/1)
fordrar (1/1)
smidigt (1/1)
barnlöshet (1/1)
yhdenvertaisuusvaltuutettu (1/1)
storfurstendömets (1/1)
betänketid (2/2)
advokat (1/1)
magistrat (4/4)
medlemsländerna (1/1)
näringsministeriet (8/8)
växte (1/1)
motionärer (1/1)
alla (120/120)
familjeåterföreningen (1/1)
reseersättning (1/1)
patienten (4/4)
kommunallagen (1/1)
kommunsidorna (1/1)
ungdomsledarna (1/1)
arbetstagarna (3/3)
Helsingforsregionens (10/10)
advokatförbundfinska (1/1)
ställas (3/3)
arbetsförhållanden (3/3)
Soite (5/5)
integrationsutbildningen (2/2)
utgifter (5/5)
LUVA (3/3)
statsgaranti (2/2)
meriterna (1/1)
invånare (45/45)
papparollen (1/1)
byggen (1/1)
biljettpriset (1/1)
Kyrkbacken (1/1)
personerlinkkiEsbo (1/1)
tullmyndigheterna (1/1)
krävas (1/1)
tidsgränser (1/1)
Maahanmuuttajanuorten (1/1)
våren (14/14)
borgarna (1/1)
fakulteterna (1/1)
äänioikeusrekisteri (1/1)
förskott (1/1)
ytterligare (9/9)
nybörjarkurser (1/1)
vuxensocialarbetet (1/1)
grundskolorna (1/1)
behovsprövad (3/3)
sökmotorns (2/2)
polisen (18/19) Polisen (1)
förtagaren (1/1)
svars (1/1)
työsuojelupiiri (1/1)
gårdsbyggnader (1/1)
Rovanapa (2/2)
bättre (5/5)
arbetspension (6/6)
löneintyg (4/4)
officiellt (11/15) Officiellt (4)
bankgiroblankett (1/1)
grannkommunen (1/1)
svartsjuka (1/1)
eventuell (2/2)
samfundfinska (2/2)
studiestödfinska (1/1)
arbetslöshetskassorfinska (1/1)
genomgår (1/1)
bortfaller (1/1)
naturskyddsområde (2/2)
ingreppet (1/1)
dubbelrum (1/1)
intressebevakningsorganisation (3/3)
sluta (6/6)
ställen (3/3)
lagstiftningen (6/6)
avbryta (2/2)
badrum (1/1)
psykolog (3/3)
misstanken (1/1)
lider (2/2)
storprojekt (1/1)
min (5/7) Min (2)
sjukförsäkringsersättningen (1/1)
levnadskostnader (2/2)
haku (1/1)
examenstillfällen (1/1)
produkt (1/1)
spanska (37/37)
hälsovårdare (19/19)
egenskaperna (1/1)
ylempi (1/1)
vigselhandlingarna (1/1)
bok (1/1)
rehabiliteringsinrättning (1/1)
upphöra (2/2)
söks (4/4)
posttraumatiskt (2/2)
tionde (5/5)
intill (3/3)
seglare (1/1)
upprättas (5/5)
sairaala (2/2)
skilja (3/3)
baserad (2/2)
partnerskap (2/2)
påminnelse- (1/1)
finansiering (12/12)
utsätts (1/1)
erityisammattioppilaitos (1/1)
frysen (1/1)
jobbsökningfinska (1/1)
filmfestivaler (2/2)
universitetsstudier (3/3)
arbetslöshetsförmånerfinska (1/1)
lokaltidningen (3/3)
bilteknik (1/1)
förgiftats (1/1)
äktenskapsintyg (4/4)
hemlands (4/4)
kulturföreningar (2/2)
seniorrådgivning (1/1)
löntagare (1/1)
erityisäitiysraha (1/1)
förmedlingsarvode (1/1)
studieprogrammet (1/1)
skrapning (2/2)
dagvårdsstart (1/1)
medlas (1/1)
hemvårdsavgiften (1/1)
jympa (1/1)
beredd (1/1)
sagts (1/1)
religiös (5/5)
utnyttja (13/13)
yrkesutbildningar (1/1)
musikskolorna (1/1)
natt (1/1)
ståt (1/1)
parternas (1/1)
särskilt (15/15)
garantipensionerna (1/1)
TyEL (1/1)
åtalsprövning (1/1)
sommaruniversitetfinska (2/2)
elavtal (4/4)
vårdpenning (10/10)
gifte (1/1)
mekanisk (1/1)
minderårig (2/2)
flyktingkvoten (1/1)
skoltiden (1/1)
månaderna (5/5)
österifrån (1/1)
vägra (7/7)
bristen (2/2)
vuxengymnasium (12/13) Vuxengymnasium (1)
tullanmäla (1/1)
missbrukarproblem (2/2)
Sveaborg (2/2)
arbetspensionsanstalter (1/1)
handikapptjänsternafinska (1/1)
anställningsintervju (1/1)
anordnad (2/2)
utvecklades (2/2)
handläggningsavgift (1/1)
magisterexamen (3/3)
stranden (1/1)
yrkeskunskap (1/1)
brottmål (3/3)
minnas (2/2)
serviceboendet (2/2)
Kelviå (5/5)
uppriktighet (1/1)
ärendena (1/1)
enas (2/2)
kontaktar (3/3)
farligt (4/4)
studiebyrå (1/1)
begäran (6/6)
ungdomsarbetare (1/1)
portugisiska (18/18)
stödcentretfinska (1/1)
säger (12/12)
skilsmässa (50/54) Skilsmässa (4)
traditionsarbetefinska (1/1)
Päihdelinkki (2/2)
redskapet (1/1)
bodelningen (4/4)
verksamhetscenter (2/2)
samiska (8/8)
centraliserade (3/3)
Vasagatan (1/1)
ens (3/3)
HelMet (3/4) Helmet (1)
barnskyddfinska (1/1)
rådgivningsbyråer (6/6)
riksdagen (2/2)
presidentval (4/4)
midnattssolens (1/1)
vapaaehtoisen (1/1)
högskoleutbildning (5/5)
antibiotika (1/1)
roliga (1/1)
invandrarkvinnorfinska (1/1)
blödande (1/1)
kommunikationssvårigheter (1/1)
toiminimi (2/2)
lämnas (13/13)
anställda (45/45)
omavastuuaika (2/2)
betalar (71/71)
polisens (8/9) Polisens (1)
budget (1/1)
flyktingarna (2/2)
boendekostnaderna (6/6)
varandras (1/1)
förmögnare (1/1)
avfall (10/10)
tystnadsplikt (2/2)
rådgivnings- (2/2)
grunddagpenning (8/8)
städer (22/26) Städer (4)
nämnda (3/3)
ambassad (1/1)
narkomaner (2/2)
expert (1/1)
föda (3/3)
sker (14/14)
anställningsintervjun (1/1)
uppmärksammar (1/1)
flygplats (7/7)
bortföranden (1/1)
dokumentmallar (1/1)
lapsettomuusklinikka (1/1)
dagpenningen (4/4)
sommaruniversitetets (1/1)
flyttade (6/6)
specialist (6/6)
programmeringsgränssnitt (1/1)
service (2/3) Service (1)
rekisteröintitodistus (2/2)
studentbostad (2/2)
film (4/4)
museikvarterens (1/1)
övningsskola (1/1)
lekar (1/1)
notaries (1/1)
lågkonjunkturen (1/1)
sevärt (1/1)
näringsidkare (5/5)
ärvs (1/1)
palveluohjaaja (1/1)
måltidservice (1/1)
mångformigt (1/1)
beredskap (1/1)
kommit (12/12)
espoo.fi (1/1)
opetustoimi (1/1)
familjedagvårdare (7/7)
intervjuer (1/1)
vrida (1/1)
familjsvenska (1/1)
tio (3/3)
livsfara (2/2)
handikappad (4/4)
framtidens (1/1)
päivystysajanvaraus (1/1)
invånarverksamheten (1/1)
hemland (20/20)
språkversioner (1/1)
biometriska (1/1)
kommun (19/19)
exemplar (1/1)
regelbunden (2/2)
invandrarungdomar (1/1)
försäljningsmetoderna (1/1)
utfärder (2/2)
boendekostnader (5/5)
livsmiljö (1/1)
förhandsröstningsställe (1/1)
gruppera (1/1)
föräldern (23/23)
depressionen (1/1)
kommunikationsfärdigheter (1/1)
tidtabeller (2/2)
språk- (3/3)
bastun (4/4)
sexuella (6/6)
tolkning (3/3)
slogs (1/1)
organisationerna (1/1)
inkomstrelaterat (1/1)
försäkring (7/7)
rehabiliteringspenning (2/2)
fastställer (2/2)
yttra (1/1)
skolläkaren (3/3)
kontorstjänster (1/1)
Petikkos (1/1)
snöskottande (1/1)
nätter (1/1)
kung (4/4)
avstånd (1/1)
kulturstad (1/1)
förmynderskap (2/2)
vanligen (46/46)
vak (1/1)
begränsad (4/4)
hemstad (2/2)
läkare (35/35)
hälsocentral (1/1)
förstår (1/1)
enheter (2/2)
idrottsplatser (5/5)
stöd- (2/3) Stöd- (1)
utrustning (3/3)
linkkiRovaniemi (3/3)
matsäck (1/1)
vardagen (7/7)
lönerna (3/3)
instanser (2/2)
webbplatsen (19/19)
viktigare (1/1)
yrkesläroanstalt (8/8)
tim. (1/1)
tvåspråkighet (1/1)
utmätning (3/3)
förhandsmeddelande (1/1)
förskoleundervisningenfinska (3/3)
Ambassader (2/2)
intresseorganisationfinska (1/1)
pratar (4/4)
framtid (2/2)
hösten (9/9)
huvudstadsregionen (12/12)
dagvårdsplatsfinska (2/2)
barnrådgivningsbyråns (1/1)
nationer (1/1)
jobbsökning (4/4)
herpes (1/1)
handleder (8/8)
e (29/30) E (1)
webbsida (2/2)
hemkommunen (3/3)
barnatillsyningsmännen (1/1)
bevilja (1/1)
ammatillinen (3/3)
Fjällrävsstigen (1/1)
invandrararbete (1/1)
Struves (1/1)
initiativtagande (1/1)
försörja (3/3)
kring (9/9)
synskada (1/1)
Nöteborgsfreden (1/1)
sparat (1/1)
boendetid (1/1)
lutherska (19/19)
idrottsanläggningar (1/1)
antecknas (4/4)
ungdomsarbete (3/3)
oavbrutet (1/1)
paddlare (1/1)
arbetstagarnas (5/5)
läkar- (1/1)
bestå (6/6)
affärsresa (1/1)
ansluter (4/4)
riksdagsledamot (1/1)
kontaktinformation (1/1)
fyllning (1/1)
skyddsbehov (1/1)
Myrkytystietokeskus (1/1)
bestämma (10/10)
responslänk (1/1)
&quot; (14/14)
Ludvig (1/1)
opintolinja (1/1)
utbildar (2/2)
nyföretagarcentralerna (1/1)
tandvårdsjouren (1/1)
grundtryggheten (1/1)
larm (1/1)
kämpades (1/1)
arbetarinstituten (2/2)
anvisningar (19/19)
strängare (1/1)
vänner (6/7) Vänner (1)
svårt (17/17)
lovat (2/2)
kommunalvalet (2/2)
anhörig (9/9)
hyresgästerna (1/1)
slidmynning (1/1)
läkemedelskostnaderna (1/1)
uppehållstillstånd (269/274) Uppehållstillstånd (5)
laga (3/3)
Sporttikortti (1/1)
köket (1/1)
arbeten (1/1)
invandrarbarn (4/4)
arbetarskyddsmyndigheternafinska (1/1)
civiltjänstgörare (2/2)
tandvårdsjourenfinska (1/1)
vidare (10/10)
vuxenläroanstalter (2/2)
åtgärder (4/4)
studieplats (29/29)
uppgiften (3/3)
medborgarinstituten (1/1)
självständigt (14/14)
Kaustby (2/2)
musiikkiopisto (1/1)
övriga (28/28)
negativt (4/5) Negativt (1)
branschspecifika (1/1)
kansanopisto (2/2)
sjukhus (31/31)
utgångsläge (1/1)
adresser (3/3)
illegala (1/1)
betalningssvårigheter (1/1)
förstasida (1/1)
integrationsplan (14/14)
bibehålla (2/2)
arbetarskyddsdistriktet (1/1)
fredagar (2/2)
familjeförhållanden (4/4)
försvar (1/1)
såsom (23/23)
tecknar (2/2)
invandrararbetefinska (1/1)
kvar (10/10)
Myyringin (1/1)
väst (2/2)
trygghetfinska (1/1)
C1 (1/1)
ateriatuki (1/1)
utbildningenfinska (1/1)
intervju (1/1)
läroanstalter (17/17)
idrotts- (1/1)
solen (3/3)
tjänstestyrningen (1/1)
Yhdenvertaisuuslaki (1/2) yhdenvertaisuuslaki (1)
köp (5/5)
tvätta (2/2)
responsen (1/1)
byråfinska (1/1)
psykiatrian (1/1)
bevara (2/2)
arbetsförmåga (1/1)
babyresa (1/1)
skyddshuset (1/1)
hälsostations (1/1)
telefonsamtal (1/1)
tel (2/2)
skolresor (1/1)
möjligheter (11/11)
februari (5/5)
pojkar (4/4)
ekonomiskt (4/5) Ekonomiskt (1)
lek (2/2)
hyvinvoinnin (1/1)
PB (1/1)
studentexamen (7/7)
längre (23/23)
återflyttningfinska (1/1)
yrkeskunnighet (7/7)
initiativ (1/1)
delägare (1/1)
äitiysneuvola (2/2)
stort (8/8)
pålitlig (3/3)
livskompetensen (1/1)
anslutningsledning (1/1)
bekantar (1/1)
S2 (4/4)
vatten (4/4)
okomplicerat (1/1)
samborna (3/3)
hemkommunfinska (1/1)
ersätta (8/8)
underlätta (2/2)
beaktar (2/2)
folkomröstningar (1/1)
knöt (1/1)
orten (4/4)
kontonummerfinska (1/1)
sjukförsäkringskort (1/1)
våld (57/61) Våld (4)
familjeärenden (2/2)
tull- (1/1)
webbplatsfinska (4/4)
yrkeshögskoleexamen (10/10)
resmål (1/1)
namnlag (1/1)
påverka (25/25)
vittnen (4/4)
existerar (3/3)
undervisning (43/43)
asyl (20/20)
Räckhals (1/1)
företagsekonomi (1/1)
äitiysraha (2/2)
förmögen (1/1)
tid (148/148)
sittunderlag (1/1)
fortsatta (9/9)
grundskolans (12/12)
skolpsykologen (2/2)
vårdanstalter (1/1)
arbetstagarefinska (1/1)
priset (2/2)
bassjälvrisken (1/1)
minderårigt (4/4)
offret (1/1)
kollektivbostäder (1/1)
hälsopunkterfinska (1/1)
fall (62/62)
noggrant (2/2)
språkkunniga (1/1)
seudun (3/3)
tjänstestället (11/11)
närvarande (3/3)
journumret (2/2)
uthyrning (1/1)
eld (2/2)
Sovjetunionens (1/1)
kroppsaga (2/2)
flyttades (2/2)
IT (1/1)
bekräftande (1/1)
nordliga (3/3)
talo (2/2)
problemavfall (1/1)
döda (2/2)
tack (4/4)
kinesiska (36/36)
stödet (12/12)
plats (26/26)
programmeringsgränssnittfinska (1/1)
byråns (13/13)
fåglar (1/1)
försvunnit (1/1)
förvärvsinkomst (2/2)
arbetslivsguide (1/1)
försäljningsställen (1/1)
receptfinska (1/1)
ditt (254/254)
varandra (16/16)
fastställs (15/15)
deras (36/36)
utkommer (3/3)
lääkinnällinen (1/1)
framhävs (2/2)
atmosfär (1/1)
studerandehälsovården (2/2)
psykologen (2/2)
arbetsverksamhet (2/2)
frånluftsventilerna (1/1)
lämpar (2/2)
Saarnio (2/3) saarnio (1)
skede (5/5)
köpingen (1/1)
prata (12/12)
övertygelse (5/5)
hälsovårdaren (9/9)
samlat (1/1)
päivälukio (1/1)
helhet (3/3)
biblioteket (17/17)
omfattas (43/43)
identifiering (2/2)
erhållit (2/2)
Lumo (1/1)
FPA (94/108) Fpa (14)
vårdutgifterna (1/1)
skolväsendet (1/1)
evenemang (9/9)
onsdag (1/1)
anställer (1/1)
studentkårer (2/2)
rekommendationer (1/1)
pensionerna (3/3)
obekvämt (1/1)
graviditetsmånaden (5/5)
brandsläckare (1/1)
Nordisk (3/4) nordisk (1)
läkarstationer (4/4)
förmånligare (9/9)
bostäderna (4/4)
förhållandet (1/1)
består (8/8)
tutkiminen (2/2)
märkningen (1/1)
kunderna (10/10)
uppfostrande (1/1)
kommunal (6/6)
egendomen (16/16)
dagverksamhet (4/4)
veckor (12/12)
hyreslägenheten (1/1)
vaccinationerna (2/2)
botas (1/1)
klädskåp (1/1)
symptom (2/2)
Svartskär (1/1)
klassen (4/4)
arbetsgivares (1/1)
handelsflotta (1/1)
diskrimineringsfall (1/1)
undervisnings- (1/1)
subventionerade (1/1)
avausleikkaus (2/2)
egnahemshuset (1/1)
yrkesutbildningenfinska (1/1)
invandrarenheten (2/2)
antal (4/4)
situationen (14/14)
växelvis (1/1)
skolkuratorer (1/1)
Helsingforsfinska (9/9)
hyresetta (1/1)
handelscentra (1/1)
märkts (1/1)
biojäte (1/1)
socialskydd (1/1)
motioner (1/1)
inkludera (1/1)
möbler (4/4)
västländerna (1/1)
vakuutusyhtiö (1/1)
stat (4/4)
oljevärme (1/1)
universitetetfinska (1/1)
väljs (12/12)
gränssnittet (1/1)
Finnishcourses.fi (2/4) finnishcourses.fi (2)
examensdel (2/2)
jobbsökningscoachning (1/1)
institution (1/1)
samling (1/1)
typer (4/4)
hälsotjänster (3/3)
restauranger (1/1)
avancerade (1/1)
installera (1/1)
ihop (1/1)
synskadadefinska (1/1)
avlägsnande (1/1)
startar (5/5)
lånekort (1/1)
Kilo (2/2)
mödravården (2/2)
understöds (1/1)
egenfinansieringsandel (1/1)
respektive (2/2)
teoretiskt (1/1)
behärskar (2/2)
rusmedels- (1/1)
förlängd (1/1)
Spektr (1/1)
anvisning (1/1)
sigfinska (1/1)
förskottsuppbördsregister (1/1)
nummer (6/6)
studieprogram (2/2)
tillverkningen (1/1)
rättshjälpsbyråer (1/1)
pedagogiskt (1/1)
beslutsfattande (3/3)
flytta (16/21) Flytta (5)
gynekologisk (1/1)
anslutna (1/1)
föra (12/12)
lediga (12/12)
hämta (6/6)
ris (1/1)
sjukdomen (1/1)
väl (8/8)
utvecklar (2/2)
fastställande (2/2)
barnatillsyningsmännenfinska (2/2)
webbundervisning (1/1)
ritualer (1/1)
efternamnet (2/2)
ungdomstjänster (6/6)
Europa (3/3)
skidor (2/2)
huvudjärnvägsstation (1/1)
statsförvaltningens (5/5)
företagshälsovård (8/9) Företagshälsovård (1)
återvinns (1/1)
bedömningen (1/1)
gården (1/1)
möjligt (41/41)
först (50/50)
köpte (1/1)
pensionssystem (1/1)
pengar (10/10)
kondomer (1/1)
startpengen (1/1)
nattjour (3/3)
arbetarskyddsmyndigheterna (3/3)
grupperna (1/1)
funktionshinder (1/1)
arbetssökandefinska (2/2)
huvudstadsregionens (3/3)
nätverket (1/1)
alkuomavastuu (1/1)
handpenningen (1/1)
skattemedel (1/1)
snabbköp (1/1)
kunskap (2/2)
järnvägsstationerna (1/1)
stadsbor (1/1)
smärtlindring (1/1)
ungdomstjänsterfinska (1/1)
länsbaserade (1/1)
kortare (5/5)
hälsorådgivningens (1/1)
studiemetoder (1/1)
avsikt (2/2)
SHVS (1/1)
gymnasieutbildning (6/6)
råder (2/2)
vattenskada (5/5)
miljötjänster (1/1)
nivåer (7/7)
stängd (1/1)
inträde (3/3)
Dublinprocessen (1/1)
privat (46/46)
tillståndstjänstenfinska (1/1)
söndagen (1/1)
entreprenörskap (5/5)
Konstskolanfinska (1/1)
ersättningsgill (1/1)
Itä (1/1)
tillgången (2/2)
ovanlig (1/1)
punktskriftsböcker (1/1)
köparens (1/1)
studietiden (1/1)
visa (12/12)
ha (119/119)
skolan (43/43)
rör (40/40)
motivera (1/1)
Renlund (1/1)
indelat (4/4)
medborgarinstitutet (1/1)
patientavgift (1/1)
medicinerna (1/1)
försäkrad (3/3)
uppmuntras (1/1)
yrkesinriktad (31/31)
minnesbilderna (1/1)
visst (6/6)
begagnade (1/1)
väljer (10/10)
röstning (2/2)
grannmedling (1/1)
jämställda (3/3)
talous- (1/1)
sommargymnasium (1/1)
kollektivtrafikens (5/5)
ersättningar (1/1)
LinkedIn (1/1)
graviditetenfinska (1/1)
invandringsfrågor (1/1)
privatpersoner (8/8)
TV:n (1/1)
jobbansökan (5/5)
ympärileikkaus (3/3)
lastenneuvola (5/5)
färdigheterna (1/1)
vägnar (1/1)
moderskapsledighet (2/2)
yliopisto (4/4)
biblioteks (1/1)
inledande (27/27)
förhöjningsdelen (1/1)
Tyttöjen (1/1)
arbetslivets (1/1)
vittna (1/1)
visumansökningsblankett (1/1)
hembygdsmuseerna (1/1)
mamma (1/1)
restaurangbranschen (1/1)
semesterresa (1/1)
kulturministeriet (4/4)
rasism (4/4)
hjälptelefon (3/3)
kvotflykting (4/4)
visumansökan (1/1)
rådgivningarna (2/2)
krisområden (1/1)
reda (22/22)
sjöfartsbranschen (1/1)
följeslagartjänstfinska (2/2)
tjänstemannafinska (1/1)
Pulkamontiefinska (1/1)
inlärningen (1/1)
Infobankens (3/3)
rosoll (1/1)
folk (2/2)
Livräddningsförbund (1/1)
partiellt (2/2)
matställen (1/1)
flyktingarfinska (3/3)
motsvarar (11/11)
boendet (9/9)
energiavfall (2/2)
transvestiter (1/1)
användaren (2/2)
dagvårdsplatsen (1/1)
i (2699/2701) I (2)
grannar (1/1)
meddelandet (2/2)
familjefrågor (4/4)
människohandelfinska (1/1)
sysselsättningstjänster (1/1)
betalningar (3/3)
behandlingsmetoder (1/1)
Uskonnot (2/2)
tre (83/83)
arbetssätt (1/1)
språkexamina (5/5)
trafikförbindelser (1/1)
identiska (3/3)
förvärvsarbetar (2/2)
arbetarna (2/2)
undervisas (3/3)
rokotus (1/1)
religiösa (10/10)
serbokroatiska (1/1)
namn (21/21)
-motion (1/1)
beskattningenfinska (2/2)
hyötyliikunta (1/1)
åtal (1/1)
överföras (1/1)
allmänläkare (3/3)
frågorfinska (1/1)
sukupuolitauti (1/1)
långt (4/4)
skada (8/8)
NTM (3/3)
kriser (1/1)
föreningar (13/14) Föreningar (1)
identitetshandling (6/6)
Päivystysapu (1/1)
utexaminerats (1/1)
familjemedlemmarnas (2/2)
enkel- (1/1)
församlingens (1/1)
licentiatexamen (1/1)
oikeusturvavakuutus (1/1)
Kansa (1/1)
företagsledning (1/1)
utsatt (23/23)
lov (1/1)
arbetslandet (1/1)
Kanada (1/1)
ärendehantering (2/2)
InfoFinland.fi (2/2)
Olkkari (1/1)
bröstcancer (2/2)
hyresavtal (16/18) Hyresavtal (2)
vattenavgift (1/1)
branscher (10/10)
försäkringsbolag (11/11)
vårdnad (16/16)
storfurstendöme (1/1)
Konttisen (1/1)
koulu- (1/1)
aktivt (4/4)
översätta (1/1)
överklaga (7/7)
högskolors (1/1)
vederbörliga (2/2)
graviditet (10/10)
foto (1/1)
nordligaste (2/2)
medborgarefinska (11/11)
neutral (1/1)
berättelse (1/1)
broschyrer (2/2)
Israel (1/1)
gånger (13/13)
ordningsnummer (1/1)
meneefinska (1/1)
licensen (2/2)
samjouren (1/1)
smal (1/1)
konstarter (3/3)
överväger (7/7)
borde (2/2)
profil (2/2)
Clinic (7/7)
examenfinska (1/1)
förmån (2/2)
efteråt (1/1)
kvotflyktingarna (1/1)
arvonlisävero (1/1)
drivas (1/1)
säljas (1/1)
företagfinska (2/2)
Sininauha (1/1)
Ounasälv (1/1)
villkoren (15/15)
eventuella (7/7)
undervisningenfinska (2/2)
Creative (1/1)
sjukvårdfinska (1/1)
AA (2/2)
barnskyddets (2/2)
sträcker (1/1)
ungdomscentralen (1/1)
utöka (2/2)
upptäcks (2/2)
anställning (21/21)
samlats (1/1)
serviceboende (12/12)
ammattikorkeakoulututkinto (1/1)
beroendeproblem (1/1)
Arbetseffektivitetsföreningen (2/2)
ordnade (1/1)
familjerådgivningen (18/18)
yrkeshögskolafinska (3/3)
bekostas (1/1)
työttömyyskorvaus (2/2)
identiteten (2/2)
bearbetningar (1/1)
anslutningsblankett (1/1)
överskrids (1/1)
genomsnittliga (1/1)
grammatikövningar (1/1)
gravid (7/7)
alternativen (1/1)
födelseattester (3/3)
Metropolias (1/1)
Kuntien (1/1)
busslinjer (2/2)
hindrar (1/1)
döms (1/1)
Tammerfors (2/2)
dolda (1/1)
mest (3/3)
bostadssökandet (1/1)
universiteten (3/3)
byta (8/8)
nia (2/2)
elledningar (2/2)
dyrast (1/1)
stöda (4/4)
friska (1/1)
väldigt (4/4)
ålders- (1/1)
idrottstjänster (5/5)
Adolf (1/1)
MB (10/10)
kraven (2/2)
traditionell (2/2)
hoitoraha (2/2)
läroplikt (3/3)
stadshuset (2/2)
ena (16/16)
fredag (8/8)
helhetsbetonade (1/1)
familjens (21/21)
flyttas (1/1)
registrerad (3/3)
aktiviteter (10/10)
fastighetsskötseln (3/3)
brev (5/5)
medium (1/1)
möte (5/5)
användarråd (1/1)
köpebrevet (1/1)
studieområden (4/4)
hota (1/1)
kredituppgifterna (1/1)
åsikter (3/3)
Sello (1/1)
meddelandekortet (1/1)
nummerserie (1/1)
många (143/143)
hemförsäkringen (4/4)
bostadsköpet (1/1)
kyrkanfinska (1/1)
mataffären (1/1)
kristendomen (1/1)
giftorätten (1/1)
barnuppfostran (1/1)
flytten (7/7)
Handelsbanken (1/1)
fordonsföreskrifter (1/1)
anvisar (2/2)
personligen (11/11)
jämställdheten (1/1)
skridskobanor (1/1)
detaljerna (1/1)
dagstidning (1/1)
plastleksaker (1/1)
förutsätter (5/5)
studielinjerna (1/1)
makans (1/1)
programmet (1/1)
rekrytering (1/1)
heltid (8/8)
batterierna (1/1)
posta (3/3)
specialbibliotek (1/1)
utreds (4/4)
avgår (2/2)
uppge (5/5)
slutfört (1/1)
kesäyliopisto (1/1)
föreningsverksamhet (2/2)
tjänsteprocesserna (1/1)
kontrollen (1/1)
du (2752/2757) Du (5)
skyldigheterfinska (1/1)
gardena (1/1)
världskriget (2/2)
besegrat (1/1)
myndighet (11/11)
könsstympning (2/2)
hälsovårdscentraler (1/1)
festlokal (1/1)
medlemsavgift (2/2)
färre (1/1)
integreras (1/1)
veroilmoitus (1/1)
Danmark (1/1)
ute (3/3)
projekt (3/3)
individualism (1/1)
internettjänsten (1/1)
tillhörande (1/1)
finns (411/411)
läkarpriserfinska (1/1)
handarbete (4/4)
tillhörighet (3/3)
avoin (7/7)
ungdomsarbetet (3/3)
partiregistret (1/1)
läsning (2/2)
gymnasiekurser (1/1)
traditioner (1/1)
stridig (1/1)
terveydenhoitaja (2/2)
bostadssidor (1/1)
specifikationsdel (2/2)
skolans (10/10)
biljetten (1/1)
könsidentitet (3/3)
Suomipassi (1/1)
Finnish (2/2)
arbetarskyddfinska (2/2)
tandkliniker (4/4)
besvärstillstånd (2/2)
Kiasmafinska (1/1)
tagit (2/2)
abonnemang (4/4)
gamla (8/9) Gamla (1)
Schengenvisum (1/1)
avkoppling (1/1)
grundinformation (1/1)
föräldraskapet (4/4)
dessafinska (1/1)
diakoniarbetaren (1/1)
utlandet (13/13)
bedömer (16/16)
förhandla (2/2)
SIMHE (4/4)
sakerna (1/1)
fullgjorts (2/2)
vigselintyg (1/1)
bostadslånfinska (1/1)
beslutat (2/2)
Strandväg (1/1)
läsämnena (1/1)
brottet (1/1)
päiväkoti (2/2)
inkomsten (2/2)
styrelse (2/2)
förseningsavgift (1/1)
förskola (2/2)
samhället (14/14)
festivalen (1/1)
säga (23/23)
betalning (1/1)
Stadin (4/4)
mål (3/3)
utskrivna (1/1)
förtroendeuppdrag (1/1)
virkatodistus (1/1)
familjedagvården (2/2)
oleskelulupa (1/1)
tidsbeställning (7/7)
bero (1/1)
köpas (6/6)
bedrivit (1/1)
tidsfrist (2/2)
familjehus (1/1)
lekparksverksamhetfinska (1/1)
snabbt (11/11)
studeranden (7/7)
tuberkulosfinska (2/2)
samarbete (4/4)
liikenne (1/1)
jämlikhet (4/6) Jämlikhet (2)
diskrimineringsombudsmannen (2/3) Diskrimineringsombudsmannen (1)
ärendet (11/11)
får (399/399)
rekommenderas (2/2)
elbolag (1/1)
samma (72/72)
kunnanvaltuusto (1/1)
käräjäoikeus (3/3)
inleddes (2/2)
informera (1/1)
ledamöter (5/5)
genus (1/1)
skolresestödetfinska (1/1)
organisationsverksamhet (1/1)
ersättningsgilla (1/1)
bygger (1/1)
inflyttningen (2/2)
Naiset (1/1)
vända (7/7)
Kluuvi (1/1)
elvärme (1/1)
vita (4/4)
samhällsmedlem (1/1)
R (1/1)
föder (4/4)
förutsättning (1/1)
arbetspensionsutdrag (1/1)
renoveringen (1/1)
onsdagar (4/4)
nämnden (1/1)
skrämma (1/1)
legalisera (1/1)
skatteförvaltningenfinska (1/1)
vårdare (1/1)
rakt (3/3)
sosiaaliohjaaja (1/1)
ytan (1/1)
register (1/1)
vintern (7/7)
hålls (8/8)
betydelse (1/1)
träffar (1/1)
högskolestuderandefinska (1/1)
faderlöst (2/2)
andelslagets (3/3)
återhämtningen (3/3)
utvecklingsstörningar (1/1)
asuntoa (2/2)
tilläggsutbildning (3/3)
ansökningarna (2/2)
organisationens (2/2)
finansierade (3/3)
viktiga (7/9) Viktiga (2)
Haag (1/1)
gårdsområden (1/1)
Hagalunds (1/1)
faderskap (4/4)
skattefritt (1/1)
meta (1/1)
Quebec (1/1)
nödläge (1/1)
klienten (2/2)
navigator (1/1)
bilplatser (1/1)
morgonen (7/7)
punkt (1/1)
arbetsförsök (1/1)
håller (11/11)
gränsen (1/1)
veronumero (2/2)
utbildning (87/92) Utbildning (5)
abonnemanget (1/1)
domstol (2/2)
framställningen (2/2)
studieresultat (1/1)
tjänsteställe (11/11)
returnera (1/1)
Grani (2/2)
kund (12/12)
problemsituationer (1/1)
jobbannonsen (3/3)
självfinska (2/2)
känt (1/1)
Översättningar (1/1)
matkulturenengelska (1/1)
finländskt (5/5)
insjuknat (1/1)
läroanstalten (11/11)
slut (4/4)
bostadsområde (4/4)
ntresserad (1/1)
tolkcentraler (2/2)
loss (1/1)
byggs (1/1)
tjänstekollektivavtalet (1/1)
specialgymnasier (1/1)
problemfinska (2/2)
familjemedlemmarna (2/2)
utbildningsprogrammen (2/2)
asevelvollisuus (1/1)
kommuns (3/3)
studier (80/81) Studier (1)
demokratiska (1/1)
någonstans (3/3)
stadsbibliotek (7/7)
slutade (1/1)
integration (13/18) Integration (5)
brottsoffrets (1/1)
hygienföreskrifter (1/1)
tidpunkt (2/2)
föräldraskap (2/2)
av (1120/1120)
fryser (1/1)
företagarpensionsförsäkringenfinska (1/1)
arbetssäkerhets- (1/1)
organisationers (2/2)
somaliska (46/46)
konventionerna (2/2)
tillvalsämnen (1/1)
kyrka (5/5)
hoitoapupalvelu (1/1)
betraktats (1/1)
tidsbeställningfinska (1/1)
aikuislukio (4/4)
Helsingforstilläggetfinska (1/1)
uträtta (3/3)
återvändande (1/1)
släktingar (9/9)
naturkunskap (1/1)
UNHCR:s (3/3)
museerna (4/4)
hemsidor (2/2)
bekant (2/2)
faderskapsledigheten (3/3)
studentbostadsstiftelse (6/6)
heller (14/14)
sähköinen (1/1)
turvakaukalo (1/1)
lokaltidningar (2/2)
idrottssällskap (2/2)
korrekta (3/3)
familjen (49/49)
drabbats (1/1)
umgänge (2/2)
återvinningsstation (1/1)
on (2/2)
mor- (4/4)
Folkmusik (1/1)
ordningsregler (2/2)
respektera (1/1)
käsiraha (1/1)
oftast (22/22)
kompetensområden (1/1)
rörelser (1/1)
mångfald (2/2)
anonymt (2/2)
MoniNet (4/4)
livlig (1/1)
fullmäktiges (2/2)
skattepengarna (1/1)
byggd (1/1)
tandvården (6/6)
gick (2/2)
International (2/2)
Klockarmalmens (1/1)
samråd (2/2)
cirkus (1/1)
högskolenivå (1/1)
flera (61/61)
områdets (2/2)
näringsidkande (1/1)
annat (135/135)
Card (1/1)
teaterfestivaler (1/1)
vanligaste (8/8)
höstens (1/1)
beskattningsbeslutet (4/4)
blåser (1/1)
bytet (1/1)
rättvisa (1/1)
nationernas (2/2)
Valvira (3/3)
handledning (21/21)
rättighet (2/2)
begränsat (1/1)
säkerställa (5/5)
semesterpenning (1/1)
läroavtalscenterfinska (1/1)
psykisk (3/5) Psykisk (2)
beträffande (2/2)
ovan (4/4)
nätbankskoder (4/4)
samtalsklubbar (1/1)
bra (54/54)
staterna (1/1)
yrkesexamen (11/11)
värd (1/1)
funktionellt (1/1)
Apteekkariliitto (1/1)
erbjuda (3/3)
varuhus (1/1)
rasistiska (2/2)
avtalat (4/4)
befolkning (2/2)
församlingarna (4/4)
släktband (1/1)
lagt (1/1)
lägenhetshotell (2/2)
bakgaller (1/1)
särskilda (5/5)
dagvårdplats (1/1)
ljudet (1/1)
Mariegatan (1/1)
inte (661/661)
Arbetslöshetsförsäkring (5/9) arbetslöshetsförsäkring (4)
naturvetenskapliga (2/2)
intrång (1/1)
begravningsplatsfinska (1/1)
Unescos (1/1)
avbokar (1/1)
församlings (3/3)
arbeta (80/82) Arbeta (2)
oväsen (1/1)
Advokatförbunds (1/1)
föräldrars (2/2)
lager (1/1)
begravning (4/4)
kommersiella (2/2)
rättsliga (1/1)
boenderådgivare (1/1)
diskriminering (37/39) Diskriminering (2)
period (5/5)
statlig (1/1)
tjänsterfinska (9/9)
ärekränkning (1/1)
voimavarakeskus (1/1)
chefredaktör (2/2)
hotell (1/1)
bekräftade (1/1)
politiska (6/6)
köpeanbud (1/1)
åldrar (5/5)
Fpas (1/1)
populär (1/1)
landskommunen (1/1)
datum (2/2)
undertrycka (1/1)
utbildningsprogram (8/8)
Matkahuoltos (4/4)
obligatoriska (4/4)
dömas (5/5)
automat (1/1)
tukiasuminen (1/1)
bevis (4/4)
arbetsmarknaden (1/1)
tvätten (1/1)
årskurser (1/1)
inhämtat (1/1)
räknas (10/10)
finska (348/355) Finska (7)
hyresavtalet (16/16)
läs- (1/1)
rådgivningens (1/1)
förmögenhet (3/3)
sluttexterna (1/1)
babyn (3/3)
körning (1/1)
personerfinska (1/1)
skyddar (1/1)
konventionsstaterna (1/1)
studiemiljön (1/1)
intressanta (1/1)
köksskåpen (1/1)
t.ex. (18/18)
bilplats (1/1)
jobbsökande (2/2)
fostrets (2/2)
skadar (1/1)
uppsägning (4/4)
badar (4/4)
vattenkonsumtionen (1/1)
WC:n (1/1)
webbsidor (8/8)
åker (5/5)
beskrivningar (1/1)
gymnasieskolor (2/2)
slutet (14/14)
hyresbostäder (32/32)
organisation (4/4)
slussa (1/1)
ry. (1/1)
tillgodoräknas (2/2)
grannkommuner (1/1)
sjöss (3/3)
hotfullt (1/1)
bibehålls (1/1)
km2 (5/5)
biogas (1/1)
arktiska (3/3)
obligatorisk (2/2)
borgen (6/6)
bindestreck (1/1)
arbetslöshetstförmån (1/1)
kommunicerar (1/1)
inkassobyrån (1/1)
resväg (1/1)
kommunsida (1/1)
civilvigslar (1/1)
hundra (1/1)
växelverkan (2/2)
bildkonstskola (1/1)
Laureas (1/1)
hobbymöjligheter (2/2)
presenteras (3/3)
sökte (1/1)
förmiddagen (1/1)
sommarsolståndet (1/1)
ensikoti (1/1)
broschyren (1/1)
bildats (2/2)
Tammerforsregionen (1/1)
utträda (1/1)
kalendermånad (2/2)
näringsbyrån (40/40)
kulturcentral (1/1)
studera (89/89)
MoniNets (4/4)
jouren (6/6)
minimivillkor (1/1)
anstalt (2/2)
studieområde (1/1)
barnförhöjningen (1/1)
original (6/6)
området (18/18)
grundskola (1/1)
semestrar (3/3)
mångfacetterad (1/1)
sjukdagpenning (11/11)
underskridas (1/1)
rektorn (1/1)
sommarkollon (1/1)
handledd (2/2)
rådgivningstjänsten (1/1)
mödrar (1/1)
integrationfinska (1/1)
kära (1/1)
kymppiluokka (2/2)
arbetstiden (4/4)
Kampen (2/2)
bokas (1/1)
Takuusäätiö (3/3)
arbetslöshetsförmånen (2/2)
skeden (2/2)
vårdartiklar (1/1)
Valviras (1/1)
någons (1/1)
vietnamesiska (7/7)
burmesiska (1/1)
Isyyden (1/1)
återkallande (1/1)
betjänad (1/1)
frukter (1/1)
klär (1/1)
esteiden (3/3)
bollplaner (1/1)
stödundervisning (3/3)
miljöcentralerna (1/1)
underteckna (4/4)
frånvarande (2/2)
motionera (1/1)
dialekterfinska (1/1)
tillståndsenhet (1/1)
samhällelig (1/1)
slottets (1/1)
annons (1/1)
svag (1/1)
uttryck (2/2)
avtalats (2/2)
mörkt (1/1)
veckoslutet (2/2)
henne (4/4)
lärt (3/3)
kan (1874/1875) Kan (1)
registerstyrelsen (5/5)
flaskor (1/1)
samorganisation (1/1)
från (235/235)
Suomi (1/2) suomi (1)
missbruksvård (1/1)
himmelsfärd (1/1)
akutmottagningen (1/1)
esiopetus (3/3)
tungt (1/1)
arrangören (1/1)
godkänd (3/3)
avvecklas (1/1)
friare (1/1)
efterlevande (2/2)
Halloween (1/1)
restaurang (3/3)
Clinicin (1/1)
postfack (1/1)
Advisor (1/1)
gymnasieskolans (1/1)
verkställa (1/1)
alkoholdrycker (2/2)
parkeringsautomater (1/1)
orsakar (4/4)
halvsyskon (1/1)
skötsel (2/2)
skolresa (1/1)
tulkkikeskus (1/1)
filmvisningar (1/1)
fysiskt (1/1)
ansöker (72/72)
senare (11/11)
undervisningsgrupper (1/1)
strykjärnet (1/1)
uppgår (1/1)
främjar (5/5)
underhållsskyldigafinska (1/1)
dagvårdsavgifter (2/2)
studieort (1/1)
vanligt (9/9)
heltidsstudier (4/4)
träffpunkten (1/1)
preventivmedels- (1/1)
rederiverksamheten (1/1)
hyreshusbolaget (1/1)
dyra (6/6)
kust (1/1)
monteringsarbetsplats (1/1)
fostret (1/1)
present (1/1)
måltidstjänst (1/1)
sosiaalivirasto (1/1)
december (6/6)
priserna (5/5)
icke (5/6) Icke (1)
läroanstaltens (2/2)
repetera (1/1)
VAV (2/2)
studentkår (1/1)
befrämjande (1/1)
kvälls- (2/2)
lärande (4/4)
arvolautakunta (1/1)
julens (1/1)
flickorfinska (2/2)
Nelonen (1/1)
studentrabatter (1/1)
kläder (6/6)
allt (17/17)
första (40/40)
arbetsoförmögenhet (2/2)
nedan (1/1)
aikuiskoulutustuki (1/1)
tv (5/6) TV (1)
investerat (1/1)
gruppfamiljedaghem (4/4)
vägguttaget (1/1)
Kokkolan (1/1)
hel (1/1)
kommuntillägg (4/4)
öka (2/2)
läsesal (1/1)
U2 (1/1)
valet (3/3)
flytt (8/8)
flyttningsdagen (1/1)
skola (18/18)
packa (1/1)
barnrådgivningsbyrån (1/1)
djurskötarexamen (1/1)
elbolags (1/1)
ledig (1/1)
Vandainfo (1/1)
kontakttolkcentral (1/1)
mobiltelefonens (1/1)
äta (1/1)
hemvårdsstödets (1/1)
mottagningscentret (1/1)
ljud (1/1)
distansstudier (1/1)
församlingars (1/1)
kulturhus (1/1)
Kieppi (2/2)
finskundervisning (2/2)
världsarven (1/1)
livsåskådning (1/1)
bilaga (1/1)
ställa (6/6)
sjukt (6/6)
rörlighet (3/3)
Facebook (1/1)
fiskeavfall (1/1)
storstäderna (1/1)
familjeträningen (1/1)
tandläkarkontroller (1/1)
kommunala (18/18)
invånarinitiativ (1/1)
Juristförbunds (2/2)
ofrånkomliga (1/1)
turistbyrån (1/1)
redaktör (1/1)
dricks (1/1)
krishjälp (1/1)
besitter (1/1)
hyresstöd (2/2)
hemsjukvården (1/1)
läggning (6/6)
underhållsförmåga (2/2)
beskattningsbeslutfinska (1/1)
representeras (1/1)
part (5/5)
andras (3/3)
egenvårdsläkemedel (1/1)
bistånd (1/1)
namnändring (3/3)
työterveyshuolto (1/1)
södra (5/5)
er (8/8)
vardagliga (4/4)
hjälpsystem (1/1)
gemensamt (11/11)
region (2/2)
allemansrätten (2/2)
bilhandlare (1/1)
privatsfär (1/1)
hyresvärder (1/1)
finlandssvenskarna (1/1)
fortsatt (13/15) Fortsatt (2)
affärspartner (1/1)
skolorna (5/5)
terapi (2/2)
utarbeta (3/3)
läroavtalsutbildning (5/5)
besöksförbudfinska (1/1)
Migrationsverketfinska (1/1)
sosiaalitoimisto (3/3)
juni (9/9)
grundar (6/6)
ålderspensionen (3/3)
drar (1/1)
huvuddukar (1/1)
vattenkannor (1/1)
skoldagen (3/3)
utredning (15/15)
MIELI (2/2)
samhällsgrupp (2/2)
Karlebystödet (1/1)
barnlöst (1/1)
mataffärer (1/1)
skiljas (3/3)
måndag (9/9)
slå (3/3)
körkort (11/11)
utbetalas (9/9)
frysens (1/1)
handikappet (1/1)
Stensvik (1/1)
fattats (4/4)
allvarligt (4/4)
kriisipalvelu (1/1)
hobbyverksamhet (5/5)
bokad (1/1)
vandringfinska (1/1)
upplevelser (1/1)
A2 (2/2)
tillverka (1/1)
kommunfinska (1/1)
meddelande (4/4)
yrkesexamenfinska (1/1)
bokbussarna (1/1)
mobilabonnemang (1/1)
äktenskapshinder (6/6)
kierrätys.info (1/1)
kreditgivningfinska (1/1)
självständighetsdagens (1/1)
starka (2/2)
konsumtionsskatt (1/1)
skedda (1/1)
flyttsak (2/2)
uppgett (1/1)
undgås (1/1)
mylla (1/1)
lähikoulu (1/1)
ungdomsväsende (1/1)
tag (1/1)
kotihoidon (2/2)
lösa (2/2)
styr (1/1)
bärande (1/1)
kurdiska (24/24)
livshotande (2/2)
letar (5/5)
tandborstar (2/2)
klinikkaan (1/1)
lyckas (1/1)
vårdplats (3/3)
hyresvärdens (2/2)
redan (30/30)
kristen (1/1)
språktest (1/1)
varhaiskasvatuspäällikkö (1/1)
vistelse (9/9)
bastu (6/6)
handikapptolkar (1/1)
avbrott (9/9)
tatarerna (1/1)
arbetsplats (27/27)
skattemyndigheten (3/3)
Europafinska (1/1)
språkkunskapskrav (1/1)
barnpassningsservicen (1/1)
koulukuraattorit (1/1)
arbetsför (1/1)
mödrarådgivningar (1/1)
måltid (2/2)
öva (2/2)
tidsbegränsat (2/2)
öppet (38/39) Öppet (1)
ringer (13/13)
gravt (1/1)
hemvårdsstödfinska (2/2)
kvotflyktingarfinska (1/1)
miljöområdet (2/2)
museets (1/1)
gravkvarter (1/1)
sjukhusavgifter (1/1)
mån.-fre. (4/4)
förlikning (2/2)
fastighet (4/4)
kotikunta (6/6)
idrottsområdet (4/4)
ansökningssättet (1/1)
diskriminerat (2/2)
uppkommer (1/1)
rådfråga (2/2)
bostadsförsäljningsannonser (2/2)
nedtecknas (2/2)
verovelvollisen (1/1)
kvotflyktingens (1/1)
skyddshemfinska (3/3)
kyrkans (3/4) Kyrkans (1)
giltighetstid (1/1)
hårdaste (1/1)
landskapsbibliotek (3/3)
reliefbilder (1/1)
hudfärg (3/3)
studieförmåga (1/1)
Liitto (4/4)
nödsamtal (1/1)
festivaler (1/1)
inleda (3/3)
yrkes- (2/2)
asukastila (1/1)
samfällighet (3/3)
arvodet (1/1)
övervåningen (1/1)
stadsdirektören (1/1)
religionssamfunds (2/2)
bokat (4/4)
rabatt (5/5)
gjorde (1/1)
milda (1/1)
övergår (1/1)
ammattikorkeakoulu (4/4)
Caisa (1/1)
sysselsättningsstöd (2/2)
skolanfinska (2/2)
förblir (3/3)
sjukskötarens (2/2)
rätten (11/11)
naturhuset (1/1)
medel (17/17)
allmännyttiga (1/1)
trappan (1/1)
sök (1/1)
testamentti (2/2)
bilder (3/3)
klienter (8/8)
ylioppilastutkinto (1/1)
vänskap (1/1)
böter (4/4)
batteri (2/2)
sorg (1/1)
hallinto (1/1)
Giftinformationscentralen (1/1)
kreditkort (3/3)
tandvård (19/19)
föräldrapenningsperioden (1/1)
Böle (4/4)
likvidation (1/1)
specialyrkesexamen (3/3)
lampor (2/2)
luthersk (1/1)
riksdagsval (2/2)
reglerar (1/1)
tusen (2/2)
for (2/2)
Trafi (1/1)
notarius (1/1)
rullator (1/1)
verksamhetsställe (6/6)
fyra (26/26)
punkten (1/1)
vikt (1/1)
skärgård (1/1)
skilts (1/1)
trafikverkets (1/1)
namnet (2/2)
bekänner (2/2)
näromgivning (2/2)
Erasmus (2/2)
självständighetsdag (1/1)
sönder (1/1)
brottsligt (1/1)
människors (5/5)
ville (2/2)
sjukskötare (6/6)
försvarandet (1/1)
frånvaron (1/1)
livmoderhalscancer (2/2)
ofta (44/44)
psykiatriska (1/1)
sex (22/22)
kontaktperson (1/1)
mössa (1/1)
tryggar (8/8)
möten (6/6)
finansiärer (2/2)
religionsfrihet (2/2)
Schengenstat (1/1)
kallas (12/12)
ingriper (1/1)
arbetsplatsintroduktion (1/1)
arbetsplatssajtfinska (1/1)
ägarbostad (17/20) Ägarbostad (3)
Mundus (1/1)
ta (117/117)
förutsättningar (3/3)
prövas (2/2)
R3 (2/2)
redogörelse (5/5)
Väestöliittos (2/2)
erövrats (1/1)
intagna (1/1)
experterna (1/1)
därför (5/5)
familjer (25/28) Familjer (3)
jourhavande (2/2)
tidpunkten (5/5)
socialbyrå (2/2)
larmar (1/1)
medlemsland (1/1)
måltidsstöd (1/1)
tillåtet (6/6)
handlägger (1/1)
elden (1/1)
flyktinghjälp (3/3)
recept (15/15)
jobbfinska (1/1)
därefter (12/12)
bostadsrättsbostäder (4/4)
svarat (1/1)
avläggs (1/1)
prat (2/2)
tiden (25/25)
hobbyutbud (1/1)
används (7/7)
studielån (4/4)
uppgå (2/2)
kvarter (1/1)
rösträtt (13/13)
än (106/106)
utvisningfinska (1/1)
universitetens (1/1)
rösträttsregistret (6/6)
familjelivet (1/1)
pappersformulär (1/1)
företagsverksamhet (15/15)
företagsrådgivningscentra (1/1)
diskriminerad (1/1)
försäkringsbolaget (1/1)
Europaparlamentet (4/4)
handläggningen (2/2)
nödnumret (32/32)
löptid (1/1)
underhållsbehovet (1/1)
tätorterna (1/1)
ort (5/5)
kopia (4/4)
studiepoäng (2/2)
medgivande (3/3)
bekräftats (2/2)
hus (7/7)
flyttsaker (4/4)
uppmuntrar (2/2)
förpliktelser (1/1)
bilens (1/1)
kilometer (2/2)
skyddskårerna (1/1)
förutsättningarna (3/3)
tvätt (1/1)
kyrklig (2/2)
träsliperi (1/1)
driftställe (1/1)
bedrevs (1/1)
sköta (21/21)
män (25/25)
utredningar (5/5)
tacka (2/2)
utarbetas (5/5)
medborgarorganisationer (1/1)
skolornas (2/2)
ansökningsblanketten (3/3)
öppnad (1/1)
kunnandet (2/2)
akademiska (1/1)
stadsfullmäktige (7/7)
autovero (1/1)
legaliserat (2/2)
medicineringen (1/1)
torka (1/1)
Konsumentförbund (1/1)
valmistava (1/1)
anger (3/3)
kaffepaus (2/2)
vuxna (33/33)
hälsovårdsministeriets (3/3)
delgivits (1/1)
sorggrupper (1/1)
övrig (2/2)
arbetar- (1/1)
uppgifterfinska (1/1)
anställd (15/15)
specialboende (1/1)
biografen (1/1)
bevisas (4/4)
öster (2/2)
rehabiliteringsbehovet (1/1)
gymnasierna (2/2)
delägarbostäder (4/4)
trapphuset (2/2)
ordnades (1/1)
kommunerna (18/18)
lönespecifikation (1/1)
tortyr (1/1)
tyngdpunkt (1/1)
kontorenfinska (1/1)
underlättar (6/6)
varken (1/1)
verksamhetfinska (3/3)
utses (3/3)
årstider (2/2)
inriktade (3/3)
vuxenutbildningen (1/1)
konsulat (3/3)
ombord (1/1)
postadress (1/1)
missnöjd (1/1)
rehabilitering (42/43) Rehabilitering (1)
utrymme (1/1)
bekosta (3/3)
arrangeras (4/4)
säsongsarbetefinska (1/1)
rådgivningstjänster (4/4)
skattekort (20/20)
att (1223/1233) Att (10)
deltidsarbete (1/1)
kulturtjänster (2/2)
sopsorterar (1/1)
dåliga (1/1)
kapitalinkomst (1/1)
tyst (3/3)
riket (1/1)
buss (1/1)
Global (7/7)
yhteispäivystys (1/1)
ansvaret (9/9)
yngre (5/5)
året (19/19)
kb (4/5) kB (1)
hemmaarbete (1/1)
köpta (1/1)
skatteprocent (6/6)
kuntoutuslaitos (1/1)
hemsjukvård (1/1)
knapp (1/1)
avsnittet (1/1)
kristelefon (3/3)
företagsverksamheten (9/9)
svenska (890/890)
upphovsrättsavgifter (1/1)
företagarutbildning (4/4)
missgynnas (1/1)
entrédörren (2/2)
gått (10/10)
sairaalan (1/1)
audiovisuella (1/1)
missbrukarefinska (2/2)
amatörteatrar (2/2)
verksamhetsspråk (1/1)
frågorna (1/1)
närmotion (1/1)
idrottsföreningar (1/1)
beter (2/2)
dagarna (1/1)
utförs (4/4)
huvudhälsostation (1/1)
noga (13/13)
mindre (24/24)
tandvårdstjänster (1/1)
arbetsprov (2/2)
utgift (1/1)
vähennykset (1/1)
samt (81/81)
ändras (4/4)
campingområdenfinska (1/1)
bett (2/2)
hobbyredskap (1/1)
vill (149/149)
förhållande (1/1)
likaså (2/2)
resekorten (1/1)
ovanligt (1/1)
konfidentiell (1/1)
pedagoger (2/2)
VR (1/1)
ansvarig (4/4)
lekparksträffar (1/1)
mars (6/6)
underlättas (1/1)
behandlats (1/1)
parts (1/1)
närundervisning (1/1)
Grankulla (40/40)
Vanda (115/115)
peruskoulu (3/3)
aktiv (2/2)
parter (1/1)
företer (1/1)
ledamöterna (1/1)
särställning (1/1)
velkaneuvonta (1/1)
ungdomsverksamheten (1/1)
betalningsdagar (1/1)
lär (16/16)
beträda (2/2)
dvs. (3/3)
förutom (2/2)
invånaren (1/1)
kundens (2/2)
KOSEKs (1/1)
städa (1/1)
åldringshem (1/1)
utbildnings- (1/1)
B2 (1/1)
servicetorget (1/1)
överklagande (1/1)
penningunderstöd (2/2)
lönetillägg (1/1)
uppdatera (2/2)
medverkar (2/2)
försörjningsförutsättningen (2/2)
underhållsskyldiga (1/1)
Veroprosentti (1/1)
beviljats (11/11)
ovannämnda (1/1)
bokfinska (1/1)
arbetssökanden (1/1)
filmerfinska (1/1)
motsvarighet (2/2)
hälsorådgivningfinska (2/2)
mödrahemmet (2/2)
arbetsförmögen (1/1)
finansrådgivningen (1/1)
MTV3 (1/1)
katolska (2/2)
A1.2 (1/1)
hemkommuns (3/3)
avslagits (1/1)
toimipiste (1/1)
stora (15/16) Stora (1)
symboler (1/1)
färdighetsnivåerna (1/1)
flaggar (1/1)
fråga (68/68)
ombyggnadsarbeten (1/1)
senaste (9/9)
utvidgar (1/1)
mandatperioder (1/1)
tillkalla (1/1)
kollektivavtalet (14/14)
konkurrera (1/1)
format (4/4)
fullständigt (1/1)
inlärningsgrupp (1/1)
ansökningsblankett (9/9)
läkemedelsbutikerna (1/1)
företagshälsovårdens (1/1)
motsvarande (5/5)
nöjaktiga (3/3)
kvinna (3/3)
möblerade (1/1)
Naapuruussovittelun (1/1)
fördel (2/2)
seniorerfinska (1/1)
polikliniken (8/8)
borgerlig (2/2)
bedriva (1/1)
exporterade (2/2)
trafikeras (1/1)
turvatalo (3/3)
integrationsrelaterade (4/4)
runt (29/29)
nordiskt (7/7)
socialhandledarna (1/1)
beskattningsbeslut (1/1)
all (1/1)
årskurserna (12/12)
ansökanfinska (2/2)
aktiivimalli (1/1)
underrättelse (2/2)
servicecenter (1/1)
könumret (1/1)
ordkonst (1/1)
hälsomotionsgrupper (1/1)
kontaktade (1/1)
anspråkslöshet (1/1)
VAU (1/1)
kännas (1/1)
direkt (55/55)
www.infofinland.fi (1/1)
påsen (2/2)
utbetalat (1/1)
vissa (88/88)
forststyrelsens (1/1)
ökat (3/3)
förödmjukande (1/1)
helt (5/5)
läkartid (4/4)
stadsdirektörer (1/1)
överenskommits (3/3)
krisjour (3/3)
hätänumero (2/2)
prepositioner (1/1)
glasförpackningar (1/1)
modersmålet (6/6)
EHIC (1/1)
belägna (3/3)
handikappråd (1/1)
kunnande (16/16)
installeras (1/1)
makthavaren (1/1)
utlänningarengelska (1/1)
helgdagar (4/4)
höst (1/1)
yrkesskola (1/1)
ny (12/12)
annorlunda (2/2)
flerfaldigt (5/5)
yrkeshögskolorna (2/2)
trafikreglerna (2/2)
nej (1/1)
tjänstetid (2/2)
grupps (1/1)
enhet (7/7)
registrerade (6/6)
norrsken (3/3)
resmålen (1/1)
skönhetsvård (1/1)
bolaget (1/1)
klarläggs (1/1)
erityishoitoraha (1/1)
examina (8/8)
ras (2/2)
servicepunkter (1/1)
klicka (1/1)
gymnasieelever (1/1)
avgiftsfritt (3/3)
Kivenkolo (5/5)
inleder (6/6)
rf (11/11)
inslag (1/1)
under (232/232)
beredning (2/2)
behandlingen (7/7)
medlingen (1/1)
stjälande (1/1)
sommaruniversitet (2/2)
påverkat (1/1)
socialbyrån (15/15)
Mina (4/4)
serveras (3/3)
par (17/17)
boka (57/57)
Östersjön (1/1)
läger (3/3)
skogsmuseumfinska (1/1)
jäte (1/1)
uppförs (1/1)
opiskeluterveydenhoitajat (1/1)
luftfartsyrken (1/1)
utbytesstudier (1/1)
blombukett (1/1)
gett (2/2)
situationer (32/32)
bosatt (19/19)
dennes (4/4)
minst (61/61)
karta (1/1)
sosiaalipäivystys (1/1)
arbetslagstiftningen (2/2)
begravningsbyråer (2/2)
civilståndsintyg (1/1)
enkla (1/1)
ämbetsbevis (2/2)
familjevåldfinska (2/2)
inletts (1/1)
innanför (1/1)
tempel (1/1)
köping (1/1)
brett (1/1)
yrkesbenämning (1/1)
grunderna (2/2)
lever (4/4)
webbplatsens (1/1)
serviceproducent (1/1)
servicepunkten (3/3)
sund (1/1)
kommunens (18/18)
reseplanerare (1/1)
oumbärliga (1/1)
Sanomat (1/1)
kansliet (1/1)
hemkommunens (1/1)
officiella (5/5)
skrivs (4/4)
makarnas (6/6)
valmansförening (1/1)
Kasabergsområdet (1/1)
forskning (5/5)
Vasa (6/6)
presenter (2/2)
levt (1/1)
tillbaka (6/6)
verksamhetsställen (9/9)
bygget (1/1)
snabb (1/1)
fördelning (2/2)
rörelsehandikappad (1/1)
ingenjör (1/1)
autonomt (1/1)
upphovsrättsliga (1/1)
bemärkelsedagar (1/1)
avgörande (3/3)
skuldrådgivning (3/3)
kartanfinska (1/1)
flyttanmälan (3/3)
samarbetsmöjligheter (1/1)
sjukskrivning (1/1)
mångfaldigades (1/1)
gardinerna (1/1)
SOS (1/1)
brister (3/3)
fallen (1/1)
tvingar (1/1)
vänskapsförening (1/1)
massörexamen (1/1)
beskattas (2/2)
förråd (1/1)
äktenskapslagen (1/1)
fiskeredskap (1/1)
swahili (2/2)
avlägger (10/10)
elektriska (2/2)
problemen (1/1)
24h (3/3)
erkännande (12/14) Erkännande (2)
meddelas (8/8)
telefonledes (4/4)
typen (1/1)
bibliotekets (3/3)
vardag (2/2)
använder (17/17)
utgörs (3/3)
nödcentralen (2/2)
bestämmelser (2/2)
kontinuerligt (8/8)
avioliiton (2/2)
reserverad (1/1)
terapeut (1/1)
sjuk (20/20)
införd (1/1)
webbplatser (13/13)
visum (20/20)
landfinska (1/1)
asumisoikeussopimus (1/1)
kortvariga (2/2)
kommunicera (1/1)
motionsform (1/1)
uteblir (1/1)
jakt (2/2)
nämn (1/1)
läskunnighet (1/1)
avslås (1/1)
ungdomslokalerna (1/1)
ry (16/16)
alternativa (1/1)
annan (65/65)
närserviceprincipen (2/2)
fortfarande (9/9)
hälften (1/1)
varumärkesrätt (1/1)
OYS (1/1)
familjebostäder (1/1)
godtagbara (1/1)
energibesparingslampor (1/1)
könsminoriteters (1/1)
lagenliga (1/1)
upptäckande (1/1)
vädret (2/2)
bioprogrammet (1/1)
tillgänglig (2/2)
följaktligen (1/1)
församlingenfinska (1/1)
procent (26/26)
aurora (1/1)
gravområde (2/2)
terminsavgifter (1/1)
gripa (1/1)
försäkringarna (1/1)
Jakobstad (2/2)
söker (41/41)
Rovalas (1/1)
invandrarefinska (20/20)
nationalparker (1/1)
möjligheten (3/3)
fyrverkerierna (1/1)
Celsiusgrader (3/3)
förarutbildning (1/1)
obegränsat (1/1)
Skatteförvaltningen (4/5) skatteförvaltningen (1)
hemsida (1/1)
ställer (2/2)
skolors (1/1)
konstindustri (2/2)
Kaapatut (1/1)
kommanditbolaget (1/1)
ledare (1/1)
sökt (3/3)
kuvataidekoulu (1/1)
julsånger (1/1)
undertecknar (4/4)
universitetfinska (6/6)
idrottsklubbar (6/6)
handelsplats (1/1)
låter (1/1)
erfarenhet (2/2)
äktenskapslagenfinska (1/1)
underhållet (1/1)
rahoitusvastike (1/1)
estetiska (1/1)
liknande (2/2)
ledigheten (1/1)
övertid (2/2)
minimilönerna (1/1)
fort (8/8)
minskar (3/3)
babyskydd (1/1)
grundskolan (33/33)
återvända (5/5)
upptäcker (8/8)
regeringenfinska (1/1)
arbetspensionsförsäkringarna (1/1)
toimintakeskus (1/1)
skuldrådgivningfinska (1/1)
socialarbetare (10/10)
rehabiliteringsstöd (1/1)
1500kt (1/1)
gård (1/1)
dagligen (1/1)
rädda (1/1)
luopumisilmoitus (1/1)
sorteras (1/1)
innehar (2/2)
område (28/28)
narkomaanit (1/1)
samarbetet (2/2)
rätta (4/4)
han (44/44)
magisterstudierna (1/1)
sammanslutning (1/1)
belysta (1/1)
ägande (1/1)
välja (16/16)
internetanslutning (1/2) Internetanslutning (1)
sökande (6/6)
ungdomsgårdar (5/5)
startpenningen (1/1)
vigsel (11/11)
parkeringsavgiften (1/1)
ansöka (206/206)
mångsidiga (3/3)
tar (52/52)
familjerådgivningsbyråerna (1/1)
underhållsskyldighet (2/2)
kallare (1/1)
Studieinfo.fi (9/9)
trivsamt (1/1)
författningar (1/1)
ring (10/12) Ring (2)
gemensam (8/8)
medelstora (1/1)
skattekortet (6/6)
orter (20/20)
skattefriheten (1/1)
frågar (2/2)
vägledning (5/5)
reglerna (4/4)
områdeskoordinatorn (1/1)
ungdomsstationen (3/3)
flykting (8/9) Flykting (1)
specialdiet (1/1)
punktligt (1/1)
servicerådgivare (1/1)
assistentens (1/1)
ung (7/7)
bygg- (1/1)
meddelanden (1/1)
könsminoriteterfinska (1/1)
försvarsmakt (1/1)
snöa (1/1)
Myrbacka (2/2)
skuldfria (1/1)
underlivet (1/1)
arbetsplatsen (25/25)
ledd (5/5)
fortsättare (1/1)
preventivrådgivningen (1/1)
utvisas (2/2)
universitetsutbildningfinska (1/1)
serviceställe (5/5)
seurakunnan (1/1)
staten (8/8)
unionens (2/2)
identifierats (1/1)
työ- (3/4) Työ- (1)
sopkärlen (1/1)
förskoleundervisningen (13/13)
verkligen (3/3)
yttre (1/1)
vårdtillägg (1/1)
frukta (1/1)
Terveyden (1/1)
bär (4/4)
växa (2/2)
arbetslös (34/34)
Sandudd (1/1)
likvärdigt (4/4)
Veikko (1/1)
vaarallinen (1/1)
sysselsättning (5/5)
Työväen (2/2)
turkiska (15/15)
finländsk (18/18)
låneräntan (1/1)
grund- (1/1)
ungdomsbostadsföreningen (1/1)
träd (3/3)
moderskapspenningperiodens (1/1)
syn- (1/1)
mellan (40/40)
tidtabellen (1/1)
jurister (4/4)
förkortat (1/1)
researrangemangen (1/1)
hyresdeposition (2/2)
viktigast (1/1)
representerade (4/4)
faktorer (2/2)
civiltjänstgöring (1/1)
lönearbete (3/3)
tung (1/1)
utdrag (3/3)
bild (2/2)
realiseringen (1/1)
svåra (2/2)
torsdagar (2/2)
koululaisten (1/1)
batterier (1/1)
cykeln (1/1)
vanlig (3/3)
Nuorisoasuntoliitto (1/1)
självständigheten (1/1)
koulukuraattori (1/1)
språkcaféer (2/2)
turistbyrå (1/1)
mentorprogram (1/1)
erbjudande (1/1)
beställa (14/14)
tvunget (1/1)
ELY (1/1)
övernattar (1/1)
yöpäivystys (2/2)
sina (57/57)
betalningspåminnelse (1/1)
Välkommen (1/1)
aikuisopisto (6/7) Aikuisopisto (1)
skyldiga (4/4)
egen (83/83)
timmar (14/14)
fritidsintressen (3/3)
Nödcentralsverkets (1/1)
telefonabonnemangfinska (1/1)
parkera (1/1)
publicerats (3/3)
servicehandledaren (1/1)
löneinkomster (2/2)
rimligt (2/2)
lösas (3/3)
styrs (2/2)
bruksföremål (1/1)
planeras (1/1)
upprepa (1/1)
integrering (1/1)
hyresbeloppet (1/1)
tror (2/2)
lättare (6/6)
småbarnsfostran (4/4)
anställningens (3/3)
värmesystem (1/1)
öst (2/2)
kommunen (34/34)
språkfinska (2/2)
Informationscentralen (2/2)
platser (5/5)
arbetsoförmåga (1/1)
tjänstebehörighet (2/2)
kommunikation (4/4)
varieteter (1/1)
ekonomin (1/1)
sortera (1/1)
ögonkontakt (2/2)
jobbsajter (2/2)
invandrarmänfinska (1/1)
tillhör (11/11)
huvudpolisstation (1/1)
debiteras (1/1)
webbaserade (1/1)
stadgarna (1/1)
praxis (1/1)
fenomen (1/1)
kielenä (1/1)
sig (184/184)
helgdag (1/1)
Finlandengelska (6/6)
försöka (1/1)
sökandes (1/1)
stickkontakt (1/1)
webbankkoderna (1/1)
makens (4/5) Makens (1)
pensionstagare (3/3)
redovisning (2/2)
rehabiliteringstjänster (1/1)
intyga (1/1)
rekryteringen (1/1)
kunde (2/2)
studentteaters (1/1)
separat (23/23)
då (82/82)
överlåtelseskatt (3/3)
täckjacka (1/1)
förlängs (3/3)
universitet (43/48) Universitet (5)
servicerådgivning (1/1)
erövrade (2/2)
sålt (1/1)
yrkeshögskolekurser (1/1)
familjeledigheten (2/2)
förändrades (1/1)
arv (2/2)
död (2/2)
duger (3/3)
hyrestiden (3/3)
förhistoria (1/1)
parkgympa (1/1)
återkalla (1/1)
sjukhusjouren (1/1)
tron (2/2)
högsommarens (1/1)
työkyvyttömyyseläke (1/1)
dateras (1/1)
-årigt (1/1)
lääkärintodistus (1/1)
insjukna (1/1)
motion (26/27) Motion (1)
faderskapsledighet (3/3)
unionen (6/6)
Novgorod (2/2)
näst (1/1)
rullstol (1/1)
studerande (52/54) Studerande (2)
mossa (1/1)
Karlebyfinska (5/5)
Tullrådgivningen (1/1)
företagsekonomiska (1/1)
undervisningstimmar (1/1)
somrarna (1/1)
Kipinä (2/2)
stavelsen (1/1)
undersökas (1/1)
stipendium (4/4)
evangelisk (17/17)
uttryckligen (1/1)
yrkesutbildningen (1/1)
markägarens (1/1)
förfaringssätten (1/1)
pyntas (1/1)
hyresvärdarnas (1/1)
hälsovårdssamkommun (7/7)
visar (2/2)
Monde (1/1)
Rovaniemiområdet (1/1)
kaikille (1/1)
hörselnfinska (1/1)
förts (1/1)
lokalerna (1/1)
arvingarna (1/1)
hemförlossning (1/1)
kraftig (1/1)
gifta (23/23)
myndigheterna (16/16)
tisdag (1/1)
flytväst (1/1)
förbinder (1/1)
läkarintyg (5/5)
godtas (1/1)
Firmaxifinska (1/1)
faktiska (1/1)
egna (44/44)
personbolag (1/1)
fackförbundet (5/5)
ombes (1/1)
folkhögskolor (3/3)
Rosatom (1/1)
krisjouren (11/11)
åldringar (4/4)
posten (2/2)
demokrati (1/1)
avsedd (39/39)
sammanträden (3/3)
stadgade (1/1)
diskutera (7/7)
gott (7/7)
tryggad (3/3)
allvarlig (1/1)
integrationsstöd (1/1)
avtala (1/1)
praktiknära (2/2)
priserfinska (1/1)
notering (1/1)
mentalvårdstjänster (2/2)
lyssna (2/2)
aktuell (4/4)
kieli (1/1)
planera (2/2)
byggbranschen (1/1)
påverkanfinska (1/1)
positivt (4/4)
ungdomsevenemang (1/1)
Internetberoende (1/1)
bytas (1/1)
Duo (1/1)
svarar (6/6)
sambo (17/17)
erityisammattitutkinto (1/1)
ingendera (1/1)
ägt (1/1)
arbetat (10/10)
klockan (10/10)
storleken (4/4)
tolktjänsterna (4/4)
tandkirurgi (1/1)
ansökningsproceduren (1/1)
speciella (1/1)
examensstuderande (2/2)
familjfinska (1/1)
inträdesprov (2/2)
bifoga (7/7)
työttömyyskassa (1/1)
angående (3/3)
halvvägs (1/1)
gymnasier (6/6)
upplösning (2/2)
idag (2/2)
färdtjänster (1/1)
städerna (7/7)
bott (22/22)
utomlandsfinska (2/2)
institutioner (2/2)
arbetsplatsens (4/4)
tillgångarna (1/1)
utlämnad (1/1)
textinnehåll (1/1)
hänt (1/1)
anslutning (8/8)
hemskickad (1/1)
enheten (4/4)
sägs (1/1)
Hyvin (1/1)
förmedlar (2/2)
hotad (1/1)
Sanduddsgatan (1/1)
metall (1/1)
hälstocentralen (1/1)
högljutt (3/3)
centraliserat (1/1)
bakgrundsmusik (2/2)
regent (1/1)
meddela (18/18)
störa (1/1)
työttömyysturvan (1/1)
för (1620/1622) För (2)
-svenska (1/1)
mödrarådgivningstjänsterna (1/1)
kost (2/2)
alltid (66/66)
fortbildningfinska (1/1)
närmare (13/13)
trottoaren (1/1)
originalspråket (1/1)
Mårtensdal (1/1)
förvaltas (1/1)
pensionspremierna (1/1)
ärende (3/3)
pensionssystemen (1/1)
webbtjänster (2/2)
regionkontor (1/1)
kris (2/2)
daghemmet (7/7)
frivilligarbeta (1/1)
Finnkinos (1/1)
Asuntosäätiös (1/1)
Menyn (1/2) menyn (1)
barnfamiljer (7/7)
Apostilleintyg (1/1)
förbättra (12/12)
formen (1/1)
jobbsajt (1/1)
stadigt (1/1)
betalningstiden (3/3)
könssjukdomar (8/8)
rubriken (8/8)
juristens (1/1)
arbetslagstiftningenfinska (1/1)
valmentava (1/1)
hälsomotionskalendern (1/1)
närarbetefinska (1/1)
bransch (9/9)
idrottsgrenar (3/3)
medborgarnas (2/2)
företagarens (3/4) Företagarens (1)
nätterna (3/3)
behövs (28/28)
resekort (9/9)
människovärdet (1/1)
täcka (5/5)
E303 (1/1)
ärver (2/2)
man (251/251)
köpet (4/4)
medlemskommuner (1/1)
nätet (13/13)
straffpåföljd (1/1)
responsiv (1/1)
de (328/335) De (7)
samarbetsavtal (2/2)
kulturella (1/1)
fysik (1/1)
pojkens (1/1)
teoretiska (1/1)
FPAfinska (1/1)
femton (1/1)
skyldigheterna (2/2)
gång (14/14)
chefen (1/1)
plast (1/1)
begränsa (1/1)
amatörer (1/1)
skuldrådgivarefinska (1/1)
begravningsbidrag (1/1)
Tukinainen (1/1)
läraren (3/3)
anställningen (9/9)
lagstadgade (1/1)
föräldradagpenning (5/5)
bostadsaktiebolagets (2/2)
yksityisen (1/1)
åldersgränser (1/1)
centralen (2/2)
underskrift (2/2)
nuorisopsykiatrian (1/1)
reglerade (4/4)
kök (1/1)
Apotekareförbundets (1/1)
trafikknutpunkt (1/1)
röra (20/20)
munhälsovårdfinska (1/1)
folks (1/1)
hälsovårdscentralen (7/7)
inlärningsresultaten (1/1)
professionella (1/1)
bereds (1/1)
tandhälsovårdenfinska (1/1)
ansvarsområde (1/1)
helheter (1/1)
utvecklingsplan (2/2)
vuxengymnasiet (5/5)
användarna (4/4)
Varias (1/1)
antagits (2/2)
beskriva (1/1)
värde (1/1)
familjerådgivningscentral (3/4) Familjerådgivningscentral (1)
redaktion (2/2)
verokortti (3/3)
lägsta (1/1)
Enter (26/26)
tryggaste (2/2)
rättegång (1/1)
glaset (1/1)
Monikas (1/1)
tilltalar (1/1)
huvudstaden (2/2)
mångkulturell (3/3)
maximibelopp (1/1)
president (4/4)
psykoterapitjänst (1/1)
utlänningsbyrån (3/3)
förberedelserna (2/2)
promenader (1/1)
förslag (3/3)
förvaltningsmyndigheter (1/1)
roligt (1/1)
måste (206/206)
få (338/338)
kondition (1/1)
Yrittäjät (1/1)
kompletteras (2/2)
bedöma (3/3)
högskolestuderande (1/1)
livmodern (1/1)
-flickor (1/1)
avgjorts (1/1)
flyttningen (3/3)
normala (1/1)
krissituation (5/5)
personefterforskningen (1/1)
fasta (3/3)
närmast (5/5)
åring (1/1)
vårt (2/2)
A2.1 (1/1)
buffert (1/1)
blödningar (3/3)
inträdesprovet (2/2)
maj (1/1)
hälft (1/1)
tillräckliga (25/25)
döma (1/1)
komposteras (1/1)
lugga (1/1)
kontrakt (1/1)
Vionojafinska (1/1)
kiinteistövero (1/1)
sjuk- (1/1)
universitetsexamen (2/2)
hotat (2/2)
våldssituationer (1/1)
bruksvederlag (3/3)
hälsovårdstjänsterna (21/21)
affärsverksamheten (2/2)
vårdas (8/8)
familjepensionfinska (1/1)
rättigheterna (2/2)
jämnt (5/5)
berätta (5/5)
undervisningsspråket (7/7)
mig (3/3)
vistats (6/6)
individuell (1/1)
familjebidrag (1/1)
personbeteckningen (7/7)
enhetlig (1/1)
grundexamen (7/7)
erövrades (1/1)
Fernissan (1/1)
förnyas (1/1)
bolagets (1/1)
parförhållande (24/24)
trakasserar (1/1)
beslutet (13/13)
våldsam (3/3)
rekryteringsevenemang (1/1)
avlagt (38/38)
Dickursby (4/4)
vågar (2/2)
diskmaskin (1/1)
påvisas (1/1)
VSB (1/1)
betjäning (3/3)
tandvårdstjänsterna (1/1)
evenemangskalenderfinska (1/1)
Tullen (1/1)
utställningar (7/7)
hörsel (2/2)
HOAS (8/8)
hobbyverksamheter (2/2)
Finnvera (3/3)
ansökningens (1/1)
stationen (1/1)
förfallodagen (2/2)
olydiga (1/1)
kielitaito (2/2)
studiekamrater (1/1)
stämma (3/3)
glömde (1/1)
oikeudet (1/1)
samfundet (1/1)
rum (4/4)
kommissionen (1/1)
skiftesvård (1/1)
webbsidan (1/1)
kristelefonfinska (1/1)
tillslutas (1/1)
Pojkarnas (1/1)
idrottshallar (2/2)
judiska (1/1)
fängelsestraff (3/3)
kommunstyrelsen (1/1)
flyktingen (1/1)
tillrådligt (1/1)
EU (117/117)
kommunerer (1/1)
även (347/347)
grundlagfinska (1/1)
läkemedlet (3/3)
tusentals (2/2)
arbetslösheten (4/4)
arbetskraftsutbildning (18/19) Arbetskraftsutbildning (1)
Nyland (8/8)
Jönsasvägen (1/1)
förskottsuppbördsregistret (2/2)
nivåerna (2/2)
vattenånga (1/1)
adress (27/27)
webbsidorna (1/1)
alkukartoitus (2/2)
Peijaksen (2/2)
årskurs (5/5)
kompetensbaserat (2/2)
samtala (2/2)
Loktorget (2/2)
hos (167/167)
avsevärt (3/3)
ingick (1/1)
litauiska (1/1)
kotivakuutus (1/1)
våning (4/4)
yhdessä (1/1)
lokal- (1/1)
koulutus (3/3)
lagar (13/13)
betyg (4/4)
duar (3/3)
Röda (10/15) röda (5)
runtom (3/3)
makarna (18/18)
förtjänat (1/1)
torsdag (2/2)
pengarna (1/1)
arbetserfarenhet (10/10)
kandidat (4/4)
brännskador (1/1)
partiell (9/9)
jämställdhetsnämnden (4/4)
visumcentralen (1/1)
simhallar (4/4)
internationella (19/21) Internationella (2)
trakasserier (2/2)
familjeförhållandena (1/1)
bosättning (2/2)
kyrkoherden (1/1)
engelskspråkig (6/6)
fundera (8/8)
familjerna (1/1)
experter (3/3)
hälsoåvård (1/1)
handarbeten (3/3)
obetalda (2/2)
utrikeshandel (1/1)
teater (8/8)
vecka (7/7)
löper (4/4)
vite (1/1)
juridiska (6/6)
dagvårdenfinska (1/1)
applikationer (1/1)
fyllde (1/1)
förmånliga (3/3)
påse (1/1)
såvida (1/1)
Martinus (1/1)
Flyktingrådgivningens (1/1)
ledighet (4/4)
situationerfinska (1/1)
kriscentret (1/2) Kriscentret (1)
löpt (2/2)
inverka (1/1)
befogad (1/1)
befolkningsdatasystemet (14/14)
ansökningspraxis (1/1)
städernas (1/1)
varför (4/4)
bokbussar (1/1)
klasser (5/5)
handikappidrott (1/1)
hörselskada (3/3)
tätorter (2/2)
Sparbanken (1/1)
små (15/15)
grundskoleinstitutionen (1/1)
studielivet (1/1)
språketengelska (1/1)
Torggatan (1/1)
handel (1/1)
filmarkiv (1/1)
bygg (1/1)
ses (1/1)
förälder (36/36)
riksomfattande (4/4)
alkoholisterfinska (1/1)
byggherrar (1/1)
flytthjälp (1/1)
finskakurs (1/1)
linje (2/2)
elektroniska (5/5)
joggingbanor (1/1)
ArPL (1/1)
hjälpmedlen (2/2)
nästan (12/12)
svara (1/1)
sambor (5/5)
Commons (1/1)
Kehitysvammahuollon (1/1)
stödhandtag (1/1)
informationsmöten (3/3)
hälsovårdsenhet (1/1)
omständigheterna (1/1)
storindustrin (1/1)
resekostnader (1/1)
specialutbildning (1/1)
lång (17/17)
volontärarbetefinska (1/1)
förvalta (2/2)
öppen (13/13)
boende (44/48) Boende (4)
ekonomiska (22/24) Ekonomiska (2)
smärtor (3/3)
religionsundervisningen (2/2)
anordnas (5/5)
yhdenvertaisuus (1/1)
personbeskattning (1/1)
kontaktuppgifter (6/6)
dör (6/6)
syskonrabatt (1/1)
framsteg (1/1)
dagvårdsplatserfinska (1/1)
överenskommit (1/1)
hade (7/7)
nettopalkka (1/1)
dagvårdsplatser (1/1)
skickar (12/12)
företagsform (2/2)
alkohol- (3/3)
kandidater (1/1)
ålderfinska (1/1)
hormonella (2/2)
integrationen (4/4)
lag (37/37)
producera (3/3)
tydlig (1/1)
vice (1/1)
pappret (1/1)
invaliditetspension (6/6)
förbundets (2/2)
begränsas (2/2)
separation (1/1)
Vanhemman (2/2)
håll (10/10)
kunder (5/5)
Chydeniusfinska (1/1)
tabletdator (1/1)
Nuppi (3/3)
vitas (1/1)
juristen (1/1)
fyllas (1/1)
fotot (1/1)
House (2/2)
terapeuten (1/1)
natten (2/2)
utvecklingen (5/5)
skolgångsbiträde (1/1)
församlingarfinska (1/1)
gränsövergång (2/2)
hushållsmaskin (1/1)
årstiderna (2/2)
granne (6/6)
empirestil (1/1)
mete (1/1)
kommuner (20/20)
enbart (3/3)
läroavtalsbyrån (1/1)
vändagen (2/2)
Raumo (1/1)
Seniorinfo (1/1)
hushåll (7/7)
ungdomarfinska (2/2)
förmånligast (1/1)
familjeplaneringsrådgivningen (1/1)
kompletteringsutbildning (1/1)
yrkesinriktade (6/6)
ruokakunta (1/1)
köpa (32/33) Köpa (1)
finländare (11/11)
övrigt (2/2)
tillståndsenheter (1/1)
avtalade (2/2)
läroanstalt (12/12)
yrkeshögskolorfinska (4/4)
Yhden (2/2)
sägas (2/2)
förvärvsarbetande (1/1)
kortfinska (1/1)
etniska (3/3)
läkarintyget (1/1)
ehkäisy (1/1)
räknare (1/1)
avger (1/1)
