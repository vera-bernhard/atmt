��      ]�(�numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i4�����R�(K�<�NNNJ����J����K t�b�C<      �      �  :   M     (      x   "   �        �t�bhhK ��h��R�(KK��h�CD1        A   �     K  ?      
   &           F         �t�bhhK ��h��R�(KK��h�C4      J   a      �  &                    �t�bhhK ��h��R�(KK��h�C8   �         L  �      �   ]   )   d   �         �t�bhhK ��h��R�(KK��h�C8�     N  �     8   E  y      �               �t�bhhK ��h��R�(KK��h�C4#   !      x   (      :   %        �        �t�bhhK ��h��R�(KK��h�CT   b      �   G   �        J   �   <     �         .                  �t�bhhK ��h��R�(KK��h�CP   (   -   x               �     [      8   �      �     o         �t�bhhK ��h��R�(KK��h�CL      5   �   9   �   �  &      U     �   
   �  *     �        �t�bhhK ��h��R�(KK��h�C4   .   �           �  �  =     @         �t�bhhK ��h��R�(KK��h�C�  �   �  �
        �t�bhhK ��h��R�(KK��h�C0�  �
     �  �     
      :   O        �t�bhhK ��h��R�(KK��h�C�
     �t�bhhK ��h��R�(KK��h�CD      =         =  M  *         
  8   �  :   O        �t�bhhK ��h��R�(KK	��h�C$      )   F  >  
   &        �t�bhhK ��h��R�(KK��h�C<      '     �  
   ?           
   A   }         �t�bhhK ��h��R�(KK��h�C`	  (  �     p            �             �     $   �     @     $  	        �t�bhhK ��h��R�(KK&��h�C�      )   \  N  "         �        
         O  �  j   �  �       �      �           �   �     �  �      �              �t�bhhK ��h��R�(KK��h�CdA        �
  �
                   �         �
     �              �  F        �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C    >   
  L   "   �        �t�bhhK ��h��R�(KK��h�CX�
     �
                 �   �  �   "   @      X      e                �t�bhhK ��h��R�(KK��h�C�     X      �t�bhhK ��h��R�(KK��h�CD      ~      P     �     �
  @   '      "   Q  �        �t�bhhK ��h��R�(KK��h�C4M     
   R  y         �   �              �t�bhhK ��h��R�(KK��h�C<�      �  �     �
     �     0   <   "   �
        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CD      2        �  �   �   "   �       '  O  7         �t�bhhK ��h��R�(KK��h�C P  5   �   3  :   +          �t�bhhK ��h��R�(KK��h�C0      &   �   �            G  ]  �     �t�bhhK ��h��R�(KK��h�C              �t�bhhK ��h��R�(KK
��h�C(�  �       B       �        �t�bhhK ��h��R�(KK��h�C   �  �  �         �t�bhhK ��h��R�(KK��h�C/   "   �      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C4   �  �  $     �     l   9     7         �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK	��h�C$H   �     (  S  -   �        �t�bhhK ��h��R�(KK	��h�C$)     �   *   Q     �        �t�bhhK ��h��R�(KK��h�C0   X   �   )   H      V   C    m        �t�bhhK ��h��R�(KK��h�CD        �          �t�bhhK ��h��R�(KK��h�CP  j      	         �t�bhhK ��h��R�(KK��h�C�   E  	         �t�bhhK ��h��R�(KK	��h�C$T        �                 �t�bhhK ��h��R�(KK��h�C4U  4     A   F     *     �
  +   n         �t�bhhK ��h��R�(KK��h�C<"   �              (      <      �     G        �t�bhhK ��h��R�(KK��h�C\$     �     +         5      V        �      �   :            O           �t�bhhK ��h��R�(KK��h�C�   �     �      �     �t�bhhK ��h��R�(KK��h�C�  �  	      	         �t�bhhK ��h��R�(KK	��h�C$�     L  �      �  �         �t�bhhK ��h��R�(KK��h�CH      O         Y      Q      Q     Q      x              �t�bhhK ��h��R�(KK��h�C`      0   R  <   "      �
  )   
               )               G     )        �t�bhhK ��h��R�(KK��h�C W     �
  	      	         �t�bhhK ��h��R�(KK��h�C\
   �     �     F   '      H     %        *  �      *         �   �         �t�bhhK ��h��R�(KK��h�C@)     /      �   L   G   �     0      �     �        �t�bhhK ��h��R�(KK��h�CI           �t�bhhK ��h��R�(KK��h�C8#   !      �     �  ?      
   3   6            �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK%��h�C�X  �        �  a  �      �     �  
   Z                    
   �        M   �      �
              �  >     �         �t�bhhK ��h��R�(KK��h�CT"           /      �   z   �     "     �
     /      ^  z           �t�bhhK ��h��R�(KK	��h�C$+  �   �  �
  �      �         �t�bhhK ��h��R�(KK��h�C�  Y  �      Z       �t�bhhK ��h��R�(KK��h�C          H   o            �t�bhhK ��h��R�(KK��h�C�  �
  [     �t�bhhK ��h��R�(KK��h�C0#   !         (      
   3   6   �        �t�bhhK ��h��R�(KK��h�C      �  �        �t�bhhK ��h��R�(KK��h�Cb     �      �        �t�bhhK ��h��R�(KK��h�C       �                  �t�bhhK ��h��R�(KK��h�Cd      ~      ,     �
  &      �   -   �   �     �    �                          �t�bhhK ��h��R�(KK
��h�C(      &   \     �  
   c        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C8d  S  \   �  ]     �      �  �  �           �t�bhhK ��h��R�(KK��h�C�  	         �t�bhhK ��h��R�(KK��h�C<�  (   %      R  H        �                    �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C0   '      .   
   e     5     y        �t�bhhK ��h��R�(KK��h�C{         S   4      �t�bhhK ��h��R�(KK��h�C~   +           �t�bhhK ��h��R�(KK	��h�C$      f     �      �  f     �t�bhhK ��h��R�(KK��h�C@  &   N   ^         /      �     J     &        �t�bhhK ��h��R�(KK��h�C0�  �     T  
   �     �     @         �t�bhhK ��h��R�(KK��h�C\�   f     g  (  �   )   _     /      �      �                   �
        �t�bhhK ��h��R�(KK��h�CL   �    
   \   H   �        �     \   H   _  %      �        �t�bhhK ��h��R�(KK
��h�C(-   K     ;      �     �        �t�bhhK ��h��R�(KK��h�C0�     �        �
  M     �   �
        �t�bhhK ��h��R�(KK��h�C0      -   �   '     6  
   �            �t�bhhK ��h��R�(KK��h�C   &   N      �      �t�bhhK ��h��R�(KK��h�CH      5   !      �           �   �         �               �t�bhhK ��h��R�(KK��h�C@   
   �   �   -  �   :              �  q   �        �t�bhhK ��h��R�(KK	��h�C$�     z      ,         �      �t�bhhK ��h��R�(KK��h�C<         �      �     �
     �     �  
   �     �t�bhhK ��h��R�(KK��h�C`     �     �         �t�bhhK ��h��R�(KK��h�C,     �t�bhhK ��h��R�(KK��h�C@U   t   
   $   �     �
     U       S     +         �t�bhhK ��h��R�(KK��h�CDV     �     .    �     >   �  *                     �t�bhhK ��h��R�(KK��h�C �   [      �     �          �t�bhhK ��h��R�(KK
��h�C(   �  �      �        �        �t�bhhK ��h��R�(KK��h�C<      z     a     L  z  {  a       b        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK	��h�C$�  h  H   R      �           �t�bhhK ��h��R�(KK��h�CD�   7  (   2      
  �  �   s  :   ?  �  Q     �        �t�bhhK ��h��R�(KK��h�C8"   m   G   �      -  �   �  /  i              �t�bhhK ��h��R�(KK��h�CT   (   <      �  
   �      (        �  �          |      �         �t�bhhK ��h��R�(KK��h�C 2     �
  	      	         �t�bhhK ��h��R�(KK��h�CTj     �  �        �  M  �   �      �
       �   �  }      �
        �t�bhhK ��h��R�(KK��h�CH      w   �       �   �             &  *      �        �t�bhhK ��h��R�(KK��h�C4N  c   I  
   �  F      �                �t�bhhK ��h��R�(KK��h�C`        �     �t�bhhK ��h��R�(KK��h�C0�     �     =         �  G   P        �t�bhhK ��h��R�(KK��h�CO              �t�bhhK ��h��R�(KK��h�Cx   �  9     �  g  �   �  (      !      \         �     �     c  
      k  �     �
  �
           �t�bhhK ��h��R�(KK��h�C �   "   T     �      �     �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK#��h�C�   5   �           8   �                    �      �  P  
   c                 �   �     �
     �             �t�bhhK ��h��R�(KK	��h�C$1   #       *      �  /         �t�bhhK ��h��R�(KK��h�C          �              �t�bhhK ��h��R�(KK��h�CD            �  G      �        =      [   G   H        �t�bhhK ��h��R�(KK��h�CP   %   0  �     2   z  W        �     1        %   �  �        �t�bhhK ��h��R�(KK��h�C �      f   �             �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C!      �        �t�bhhK ��h��R�(KK��h�C         .   �        �t�bhhK ��h��R�(KK��h�C  E      �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C@   (   #   !      X     k   
   3   6   2              �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C/      8     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C �  )                   �t�bhhK ��h��R�(KK��h�CT�  �     N   �      �  �  �     J  
   C   �  -   �                �t�bhhK ��h��R�(KK��h�C     �     �     �t�bhhK ��h��R�(KK��h�C   �     `   �     �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK	��h�C$
     �  %     Q          �t�bhhK ��h��R�(KK��h�C`      R  �
       �   R         �  9   �  �        :            �  �        �t�bhhK ��h��R�(KK��h�CL   X   '   -   H   A   F     L  %   .           �     �        �t�bhhK ��h��R�(KK��h�CP2                �   �         .      S     �        �        �t�bhhK ��h��R�(KK��h�C@�                   �   �        �              �t�bhhK ��h��R�(KK��h�C          W        @      �t�bhhK ��h��R�(KK��h�C%      ~               �t�bhhK ��h��R�(KK��h�C`   l               l      A           �
     0   <      d     %   �          �t�bhhK ��h��R�(KK��h�CD�  �     q   .    V   2      e  C   h   H   B   3        �t�bhhK ��h��R�(KK��h�C  	      	   K      �t�bhhK ��h��R�(KK��h�C4K       �       �      �     9        �t�bhhK ��h��R�(KK
��h�C(!      	        	      	         �t�bhhK ��h��R�(KK��h�C �
        	      	         �t�bhhK ��h��R�(KK��h�C`4                �   �         0   �  �  -                        .         �t�bhhK ��h��R�(KK��h�Clf  
     �  	      	      	   K   	   �   	   �   	     	   I  	   �  	   U  	   �  	   �      �t�bhhK ��h��R�(KK��h�C0      �  �
     �   >        �         �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6            �t�bhhK ��h��R�(KK��h�C0
   �   F   '   !           �  �         �t�bhhK ��h��R�(KK
��h�C(�      /         	      	         �t�bhhK ��h��R�(KK��h�C!            �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C<        {      �     )  +      |      �         �t�bhhK ��h��R�(KK��h�CP   (   �  3  "   @        T     8   �     �  �                 �t�bhhK ��h��R�(KK��h�C�
     �t�bhhK ��h��R�(KK��h�CLY  h     �     h        O     g              �  U        �t�bhhK ��h��R�(KK��h�C�      �   0   <   r      �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�CL         9   9  7      5   �     M   �      �  "   $           �t�bhhK ��h��R�(KK��h�C8   (   �     *      �  +        G   t         �t�bhhK ��h��R�(KK��h�C�
     	      	         �t�bhhK ��h��R�(KK$��h�C�            �  4      �     �               Z        0      k            �
           $        �   �               �t�bhhK ��h��R�(KK��h�C8      �  h     
   �  (   %   )   �           �t�bhhK ��h��R�(KK	��h�C$   [  :     ?  �
  �        �t�bhhK ��h��R�(KK��h�CT   �
     J    /   &   %   �   5     �  |  
   �        "   �         �t�bhhK ��h��R�(KK	��h�C$H   �        �   �           �t�bhhK ��h��R�(KK ��h�C�            i  
   4  P  �   +      �  �     C      6     P               \  L   y      ]  �         �t�bhhK ��h��R�(KK	��h�C$   �      L                 �t�bhhK ��h��R�(KK��h�C@   �   �
  '   �        V         i  �             �t�bhhK ��h��R�(KK��h�C,   f   �    )   �   �      �
        �t�bhhK ��h��R�(KK��h�Cl:   ?  �  Q     �  (      M      +            j  �     �   �
     �  A  �   k  �
        �t�bhhK ��h��R�(KK��h�C<      �        �   j   �     �   9     7         �t�bhhK ��h��R�(KK��h�C    	      	         �t�bhhK ��h��R�(KK��h�C@  �  c                          f   A   �
        �t�bhhK ��h��R�(KK��h�CH           &  *      �        �       �   �  w         �t�bhhK ��h��R�(KK��h�C0�  �  �     �  �        �           �t�bhhK ��h��R�(KK��h�C�     �  r      �t�bhhK ��h��R�(KK��h�CD      �  5   <               �  &      �   j  /        �t�bhhK ��h��R�(KK
��h�C(�   q   7     �     `  �
        �t�bhhK ��h��R�(KK��h�C,      �      P     �   
           �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C@"   �   �   2        G   %  K  D      �   l          �t�bhhK ��h��R�(KK��h�C �           V     u      �t�bhhK ��h��R�(KK��h�CD�  a     �   W  �     �   f   W  >      w   =            �t�bhhK ��h��R�(KK��h�CX            N  �                             5      �  �  �        �t�bhhK ��h��R�(KK
��h�C(      �           J  E         �t�bhhK ��h��R�(KK��h�C!          �t�bhhK ��h��R�(KK��h�CX      0   �      8   �  �  �  �
     �     "     V     �      �         �t�bhhK ��h��R�(KK!��h�C�   �   �     0   4   -      �      �      �         t        6        l           y   �  �   W              �t�bhhK ��h��R�(KK��h�Cp      M     �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�Cb     �t�bhhK ��h��R�(KK��h�CL   �    �     7   �
     �     g      �     �     �        �t�bhhK ��h��R�(KK��h�C8#   !      �                               �t�bhhK ��h��R�(KK��h�C1   #       �         �t�bhhK ��h��R�(KK��h�C@1   #         }     o   
   3   6   7  }     o         �t�bhhK ��h��R�(KK	��h�C$�
           C   
   �        �t�bhhK ��h��R�(KK
��h�C(   m  )  �   *   Q     �        �t�bhhK ��h��R�(KK��h�C4      �  �     �      �                 �t�bhhK ��h��R�(KK��h�C  X     �t�bhhK ��h��R�(KK��h�C<�         e  +   
   �     �      v      �         �t�bhhK ��h��R�(KK��h�C �         �  �           �t�bhhK ��h��R�(KK��h�C<      -   �   8        �   o      �      n        �t�bhhK ��h��R�(KK��h�CY            �t�bhhK ��h��R�(KK��h�C4      �
  8  �
     Z       �  �        �t�bhhK ��h��R�(KK��h�CT*      �           �              )        n        ,           �t�bhhK ��h��R�(KK��h�Co     �t�bhhK ��h��R�(KK��h�C,1   #   
   3   6   �        �         �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C0�  �  �   �  �       [     �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�Cp^   \        a   �      d   ]     0   !      d   �     ^        �   p     �                  �t�bhhK ��h��R�(KK��h�C0      n      \  L   y                  �t�bhhK ��h��R�(KK	��h�C$�      )   v         0        �t�bhhK ��h��R�(KK��h�C0D   (   �  o  �   "   �     �   �          �t�bhhK ��h��R�(KK��h�CT   ]   �   &      =         �   ~     �  $        t      �           �t�bhhK ��h��R�(KK��h�C8#   !      �  ?      
   3   6   �             �t�bhhK ��h��R�(KK	��h�C$           �
              �t�bhhK ��h��R�(KK��h�C|   L     `     �  �       7   m  �
  7      �
          `     �       9  7      �  �  �        �t�bhhK ��h��R�(KK
��h�C(B    #             +         �t�bhhK ��h��R�(KK��h�C\   <      �           P        �     ,      @      X      e              �t�bhhK ��h��R�(KK��h�C8   ]   �   >      �           �
     H        �t�bhhK ��h��R�(KK��h�CT   S   G         
           $  �  '   �     *           �
        �t�bhhK ��h��R�(KK��h�C�  O      �t�bhhK ��h��R�(KK��h�CHq           %  +         S      q              @         �t�bhhK ��h��R�(KK��h�C 1   #       �     _        �t�bhhK ��h��R�(KK
��h�C(   �  k    
   ,               �t�bhhK ��h��R�(KK��h�C<p     �  �   �  �  �      �  "   �   �   �        �t�bhhK ��h��R�(KK��h�C    @   '   �             �t�bhhK ��h��R�(KK��h�C,   "   �   n        	      	         �t�bhhK ��h��R�(KK��h�C@
   &     �      �  �  +        c   �     �
        �t�bhhK ��h��R�(KK��h�C,      �      �  �  �  �   �
        �t�bhhK ��h��R�(KK��h�CL`  �  :              d   �  ^     �     D   �  N  7         �t�bhhK ��h��R�(KK��h�CP   ?   1     #   !      E      4      �  
   �     q  q   _        �t�bhhK ��h��R�(KK��h�C<                  �     9   '     $   E         �t�bhhK ��h��R�(KK��h�CP   .   r  C      �   O     �     �     u     :  �              �t�bhhK ��h��R�(KK	��h�C$(  s  (   J     I           �t�bhhK ��h��R�(KK��h�CT
   3   6   )  ?   �   �   r   '   !      \         �     �               �t�bhhK ��h��R�(KK��h�C,�         0   [      �              �t�bhhK ��h��R�(KK��h�C,1   #   
   3   6   �     �  m         �t�bhhK ��h��R�(KK��h�CXR  M        �     ]     �   �                 ,            �        �t�bhhK ��h��R�(KK
��h�C(               a  j   �
        �t�bhhK ��h��R�(KK��h�CD#   !      �  �  ?      
   3   6   �          �        �t�bhhK ��h��R�(KK��h�C�         �     u      �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   6   �  "   �         �t�bhhK ��h��R�(KK��h�CL�   �
     �   �              !  �      "     �      #        �t�bhhK ��h��R�(KK��h�CT         2                      +      ;  +         o  <        �t�bhhK ��h��R�(KK��h�C8         �         P   +  ^   =  b  *        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C 1   #       `     t        �t�bhhK ��h��R�(KK��h�C<u  �
     $         %  &  �        '  (        �t�bhhK ��h��R�(KK��h�C,   (   T   )     �        v        �t�bhhK ��h��R�(KK
��h�C(      *  +  +         ,        �t�bhhK ��h��R�(KK��h�Ct�        �             %   w  �      �  �         �  �   �  C  !  >     8        -        �t�bhhK ��h��R�(KK��h�C<�
     x       c  	   U  	   �   	   �  	         �t�bhhK ��h��R�(KK��h�C+     �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CL
   3   6   �
     �
        '   !      �        �              �t�bhhK ��h��R�(KK��h�C<
   �        e  �
  �
  �   �      ?             �t�bhhK ��h��R�(KK��h�C0�     �     d  <            .        �t�bhhK ��h��R�(KK	��h�C$%      �     �  �           �t�bhhK ��h��R�(KK
��h�C(   �  �   �          �           �t�bhhK ��h��R�(KK��h�C/  	         �t�bhhK ��h��R�(KK��h�Ce     �     �t�bhhK ��h��R�(KK��h�C4*           '   �  H   �     8   S        �t�bhhK ��h��R�(KK��h�CT      �      �  C         �   +     "  g            �              �t�bhhK ��h��R�(KK
��h�C(
   �  6   '   !         ,        �t�bhhK ��h��R�(KK��h�CD   @         �  �  G   k              W              �t�bhhK ��h��R�(KK��h�C0]   P     %         ;      �   �        �t�bhhK ��h��R�(KK��h�Cb   #   "   $            �t�bhhK ��h��R�(KK
��h�C(      -      :  g   0  p        �t�bhhK ��h��R�(KK��h�C4'   !      \         �     �               �t�bhhK ��h��R�(KK��h�C a        	      	         �t�bhhK ��h��R�(KK��h�C4   $   k      X         �   Q  �   �        �t�bhhK ��h��R�(KK��h�C      y  �   �      �     �t�bhhK ��h��R�(KK��h�C4      ,  "   T     :     $   �  �        �t�bhhK ��h��R�(KK
��h�C(I     :   `   3  �      �         �t�bhhK ��h��R�(KK��h�C0�   _        f  �   
   A  �  z        �t�bhhK ��h��R�(KK��h�C g  �  �
        �         �t�bhhK ��h��R�(KK��h�C0�  �     �                 ^        �t�bhhK ��h��R�(KK��h�C</            S   X  i   ,            0   0        �t�bhhK ��h��R�(KK
��h�C(X   �   p  9   W  7     �        �t�bhhK ��h��R�(KK��h�C        �t�bhhK ��h��R�(KK��h�C �     �  	      	         �t�bhhK ��h��R�(KK��h�C�   -     �t�bhhK ��h��R�(KK��h�C1  	      	         �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C
   ,   �
  2   �        �t�bhhK ��h��R�(KK��h�C<      �        {  �        �   2     "        �t�bhhK ��h��R�(KK��h�C<H        h     u            3  C   
            �t�bhhK ��h��R�(KK��h�CP      ~         +  &      �   �     �  �   $   .  n      L         �t�bhhK ��h��R�(KK��h�CD   /            |  �      q          �     �        �t�bhhK ��h��R�(KK��h�C1   #       i        �t�bhhK ��h��R�(KK
��h�C(      �      �
  @  N  �         �t�bhhK ��h��R�(KK	��h�C$�   �   �  A  :        �     �t�bhhK ��h��R�(KK��h�Cl   2   J     :  �     �   �  B     >   2   �   �  C   �   7      A  :   �   �     �         �t�bhhK ��h��R�(KK
��h�C(�   >   4  c   
   _      �         �t�bhhK ��h��R�(KK��h�C!         	         �t�bhhK ��h��R�(KK��h�CX%   �          j     �        k     R                    /         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CD4  �     \   �  �      �   +      �      -  d   �        �t�bhhK ��h��R�(KK��h�C5  	      	         �t�bhhK ��h��R�(KK#��h�C�         �   G      t  &      =      n     �     Y      O   
   _      �     �   �        
   �     �     �        �t�bhhK ��h��R�(KK��h�C�
     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CL
   t   C  2            "     F     k      l        +         �t�bhhK ��h��R�(KK��h�Ch      ;      �   �      �  R            
  0  4      �        +  4      m           �t�bhhK ��h��R�(KK	��h�C$      }           �        �t�bhhK ��h��R�(KK��h�C`   r     �  +     �  �     �  L         2         �       �
     e        �t�bhhK ��h��R�(KK��h�CL
        �
  6  n     �     �
  �     �     ?      !         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C4D      )   2     �  �      �     �        �t�bhhK ��h��R�(KK��h�C@m     Y      �     )      
   �   �     +  4         �t�bhhK ��h��R�(KK��h�C   5   �   �         �t�bhhK ��h��R�(KK��h�Ch~     �
     M  	      	      	   K   	   �   	   �   	     	   I  	   �  	   U  	   �      �t�bhhK ��h��R�(KK��h�C             �t�bhhK ��h��R�(KK��h�C!         	         �t�bhhK ��h��R�(KK��h�C T      �  R     +         �t�bhhK ��h��R�(KK��h�C�      �     /      �t�bhhK ��h��R�(KK��h�C1        7  �  r      �t�bhhK ��h��R�(KK
��h�C(   v     
     �   $   o        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C1   #       p     �     �t�bhhK ��h��R�(KK��h�C4   '   -      V   8     �     �   &        �t�bhhK ��h��R�(KK
��h�C(   	      	      	   K   	   U     �t�bhhK ��h��R�(KK��h�C�  q        �t�bhhK ��h��R�(KK��h�C`   �     �
        8     �
     9  V      {  $   �     $   :     �  �        �t�bhhK ��h��R�(KK��h�C;        �t�bhhK ��h��R�(KK��h�C0
      ]  T  '   !      .     �         �t�bhhK ��h��R�(KK	��h�C$      �     �  r  	         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�CDb  �
     b      s  �
     �   2      2  �               �t�bhhK ��h��R�(KK��h�C M      +   3     4         �t�bhhK ��h��R�(KK��h�C,   {  �          �     �        �t�bhhK ��h��R�(KK��h�C8      -   �  +              <  =           �t�bhhK ��h��R�(KK
��h�C(W   �   t     �  �              �t�bhhK ��h��R�(KK��h�Cd�      
   4  	      	      	   K   	   �   	   I  	   �  	   U  	   /  	   s  	   �     �t�bhhK ��h��R�(KK��h�C    �        8   �        �t�bhhK ��h��R�(KK��h�C4/      -   6        �        >           �t�bhhK ��h��R�(KK��h�C4�  �   +   x      5        `             �t�bhhK ��h��R�(KK��h�C`*      �         D  l        �   f        �      �   ;      0   �     �        �t�bhhK ��h��R�(KK��h�C      2         �        �t�bhhK ��h��R�(KK��h�C u     �  �  �   E        �t�bhhK ��h��R�(KK��h�C,   2   �  Y  ?     2   0   �        �t�bhhK ��h��R�(KK��h�C          	      	         �t�bhhK ��h��R�(KK��h�C8�      =      [      v    ^   �               �t�bhhK ��h��R�(KK��h�C06  �        F     G     C  /         �t�bhhK ��h��R�(KK��h�CT%   �   .  w  @     
   �        2      �   t     �   �      O        �t�bhhK ��h��R�(KK��h�CH      D  =         �  4      m  >      a      �  �         �t�bhhK ��h��R�(KK��h�C      �            �t�bhhK ��h��R�(KK	��h�C$      A  ?                �t�bhhK ��h��R�(KK��h�CH      c     `   m      /     B  i     %   ^  "   �        �t�bhhK ��h��R�(KK��h�CH      J         )     �   �   S        �     5           �t�bhhK ��h��R�(KK��h�C4     �      5   �      �         C        �t�bhhK ��h��R�(KK��h�C�   -     �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�CT
        2   �   0  p  
   z  �   7      �  �  p  
   z  s   7         �t�bhhK ��h��R�(KK��h�CL@   �   �        /      �  M     {     e     �  g           �t�bhhK ��h��R�(KK��h�CZ   D     �t�bhhK ��h��R�(KK��h�C,�  1        4   �   �      �         �t�bhhK ��h��R�(KK��h�C0]   �     E     F                    �t�bhhK ��h��R�(KK��h�CD   (   H              R  H     4   
   �   �   _         �t�bhhK ��h��R�(KK��h�C4      6  +      �  �        d  G        �t�bhhK ��h��R�(KK��h�Cx     �t�bhhK ��h��R�(KK��h�C�  H     �     �t�bhhK ��h��R�(KK��h�C q               I        �t�bhhK ��h��R�(KK��h�C�   !      �  	         �t�bhhK ��h��R�(KK��h�C0      �     0      k                   �t�bhhK ��h��R�(KK	��h�C$�   �  �  �  �               �t�bhhK ��h��R�(KK��h�C,     1        '   
   �  F         �t�bhhK ��h��R�(KK��h�CD
     (      [      "   >  x      �         0   <         �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C�   J     �t�bhhK ��h��R�(KK��h�C1   #       �        �t�bhhK ��h��R�(KK��h�C8�     K  �     C   �      �     �  �        �t�bhhK ��h��R�(KK��h�Cp�  L  �  M                                      N     O     P  (   N   A     I        �t�bhhK ��h��R�(KK
��h�C(Q  y           �      I         �t�bhhK ��h��R�(KK��h�C<   �      $  �      �  i                       �t�bhhK ��h��R�(KK��h�C8      )   P   ^     �      ^   q   R  F         �t�bhhK ��h��R�(KK��h�C`   �      e     �  i   #  �     !  �  	  S     z     �        �   w         �t�bhhK ��h��R�(KK��h�CP      �     �  5         �           >   a                    �t�bhhK ��h��R�(KK��h�C4
   �     �     F   '      H     �        �t�bhhK ��h��R�(KK��h�C  �   �  �  �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�   v            �t�bhhK ��h��R�(KK��h�C<M      \  L     
   *         =         �        �t�bhhK ��h��R�(KK��h�C4h  �  O   >   )  C   �  G   |      �         �t�bhhK ��h��R�(KK��h�CT   �            �t�bhhK ��h��R�(KK��h�C47     ;      w   5     �   J   �   8        �t�bhhK ��h��R�(KK	��h�C$T      9        �   �         �t�bhhK ��h��R�(KK��h�C\   �   �  r      �t�bhhK ��h��R�(KK��h�C0         \     (         �           �t�bhhK ��h��R�(KK��h�C@1   #      f        
   3   6     �   �               �t�bhhK ��h��R�(KK��h�C �  T     
     U        �t�bhhK ��h��R�(KK��h�C@   t     /   9   -  (   2   <           �           �t�bhhK ��h��R�(KK	��h�C$                 �         �t�bhhK ��h��R�(KK��h�C<
   V  F         �  �    �     /      {        �t�bhhK ��h��R�(KK��h�C:  �  �   �          �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C�             �t�bhhK ��h��R�(KK��h�C`"   W       X    p      Y  �  h   �     �          Z     [     \        �t�bhhK ��h��R�(KK��h�C\]     �  ^        �         �         _        :      S   Y      Q         �t�bhhK ��h��R�(KK��h�CD*      �  +                   ;  +      `  <        �t�bhhK ��h��R�(KK��h�CD   '   �  �     �  
   a                            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C<      �   %   �                 k               �t�bhhK ��h��R�(KK��h�CP
   3   6   7  }     o   ?      !      \   2   |     o               �t�bhhK ��h��R�(KK��h�C0   b  �  5         �        Z        �t�bhhK ��h��R�(KK��h�Cc     �t�bhhK ��h��R�(KK��h�C  
         �t�bhhK ��h��R�(KK��h�CD-     b        S  u  �     �     l      �  b        �t�bhhK ��h��R�(KK	��h�C$p      :          �        �t�bhhK ��h��R�(KK��h�C0�  ;  d        <                    �t�bhhK ��h��R�(KK��h�C@�   q   7  &   I     �  �  }     C  �             �t�bhhK ��h��R�(KK��h�C<   d  �     �  �     ~     l      5            �t�bhhK ��h��R�(KK��h�C<      M   �   �         �           <           �t�bhhK ��h��R�(KK��h�C1   #          �t�bhhK ��h��R�(KK��h�C�     �   e           �t�bhhK ��h��R�(KK
��h�C(,   �          	      	         �t�bhhK ��h��R�(KK��h�CD$   �     T           �           �   o               �t�bhhK ��h��R�(KK��h�C<      
   _          |  �     7  J          �t�bhhK ��h��R�(KK��h�C         e  
   c        �t�bhhK ��h��R�(KK	��h�C$�       ^     B   �        �t�bhhK ��h��R�(KK
��h�C(   (   �  �          �        �t�bhhK ��h��R�(KK��h�Cf  �   �   �         �t�bhhK ��h��R�(KK
��h�C(     �           ;   g        �t�bhhK ��h��R�(KK��h�C   J  C      !     �t�bhhK ��h��R�(KK��h�Ch  �     $   �         �t�bhhK ��h��R�(KK	��h�C$#   !   ?      
   �   F         �t�bhhK ��h��R�(KK��h�C=  	         �t�bhhK ��h��R�(KK��h�C�        o  <     �t�bhhK ��h��R�(KK��h�C<"   e   �
     �           /      ^  z           �t�bhhK ��h��R�(KK	��h�C$      3  �     k            �t�bhhK ��h��R�(KK��h�C   4  '   �   i        �t�bhhK ��h��R�(KK��h�C,%   �     j  :   @      X   �        �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6   k        �t�bhhK ��h��R�(KK��h�C8      �  c   �            l     
            �t�bhhK ��h��R�(KK��h�CL   ?   m  *      �  "  n  o  "     u  �         p           �t�bhhK ��h��R�(KK	��h�C$H  �  +            q        �t�bhhK ��h��R�(KK��h�C8%   >  r     �   �            s               �t�bhhK ��h��R�(KK��h�C<            z   
   ,            �  
            �t�bhhK ��h��R�(KK��h�C0v  �        .   s     t              �t�bhhK ��h��R�(KK��h�C0w     ;     u          "   5        �t�bhhK ��h��R�(KK��h�CD*            k         �   Q  R      �     .   �        �t�bhhK ��h��R�(KK��h�CK         Z   �     �t�bhhK ��h��R�(KK��h�C   k  j     /        �t�bhhK ��h��R�(KK��h�CX         8        �   O      ~               0   4   
   _      �        �t�bhhK ��h��R�(KK
��h�C(      )   M   +                 �t�bhhK ��h��R�(KK��h�C@a           �  	      	      	   K   	   U  	   /     �t�bhhK ��h��R�(KK��h�CP   n      �t�bhhK ��h��R�(KK��h�Cv  M             �t�bhhK ��h��R�(KK��h�C0�   7  (   �       .      �   ?         �t�bhhK ��h��R�(KK��h�C   =      �      �t�bhhK ��h��R�(KK��h�C4   (   #   !      �     $   x  
           �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C0  �      �  �   �        O  �        �t�bhhK ��h��R�(KK$��h�C�*   H     w     �  �   
   $   E         
   _      �          K       x     `         �     �   �      �  �        �t�bhhK ��h��R�(KK��h�C8V                 �     $  �              �t�bhhK ��h��R�(KK��h�Cq     �t�bhhK ��h��R�(KK��h�CT   �  �  �  �  �  h      �   L     �          v  ;      y        �t�bhhK ��h��R�(KK��h�C       z   ,               �t�bhhK ��h��R�(KK��h�C8T   �                                    �t�bhhK ��h��R�(KK��h�C   �     8   �        �t�bhhK ��h��R�(KK��h�C4
     �      u   p        �   
           �t�bhhK ��h��R�(KK��h�Cg  �           e      �t�bhhK ��h��R�(KK��h�CG     u        �t�bhhK ��h��R�(KK
��h�C(   �  &   `     �  �  �        �t�bhhK ��h��R�(KK��h�C,Z      �               �            �t�bhhK ��h��R�(KK��h�CH^  u            Y  �  :   �   �   Q      �   O  
   �        �t�bhhK ��h��R�(KK��h�C,      �  �  0  �        z        �t�bhhK ��h��R�(KK��h�Ch{        Y           �            �       �      �      �  �      h     �         �t�bhhK ��h��R�(KK��h�CT|           �     I   /   �           ;      }        �           �t�bhhK ��h��R�(KK��h�C     	      	         �t�bhhK ��h��R�(KK��h�C<�      �  �     R            �     v   �        �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK
��h�C(~    @  '   9     ]          �t�bhhK ��h��R�(KK��h�C@"   �           e      @         z   h   H   �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C      �   f     �t�bhhK ��h��R�(KK��h�C,:  
      �     M     {  7         �t�bhhK ��h��R�(KK��h�CP   �      $     �  �   Y  +      �  +      �      U      �        �t�bhhK ��h��R�(KK��h�C!  �     0   <         �t�bhhK ��h��R�(KK��h�C8            �     "     ]  �     Z        �t�bhhK ��h��R�(KK��h�Cp         �   �  �  
   #           �          $  %     >      v            �            �t�bhhK ��h��R�(KK��h�CP      &        �  �   �     '  �     �  �  
         �        �t�bhhK ��h��R�(KK��h�C<   i  �  R         /   9     7         �         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C,.  M        
        �            �t�bhhK ��h��R�(KK��h�CD            �     M   T   �   �           i           �t�bhhK ��h��R�(KK��h�C         �           �t�bhhK ��h��R�(KK��h�C   �      �t�bhhK ��h��R�(KK��h�C<�  N  
   8     ^   &  �     
      �  �        �t�bhhK ��h��R�(KK��h�C   �  
   �     �t�bhhK ��h��R�(KK��h�C<      5  �      \   �        &     
   U        �t�bhhK ��h��R�(KK��h�C              �t�bhhK ��h��R�(KK��h�Cq            �t�bhhK ��h��R�(KK��h�C\
   3   6   �  ?      !      #        �      $   �  �  �      �     �         �t�bhhK ��h��R�(KK��h�C0   >   �       �   *   �  �  V         �t�bhhK ��h��R�(KK��h�C4�  9     W     (           )  �
        �t�bhhK ��h��R�(KK��h�C@�     �           �
  :   �  
   _      �  �        �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�CD      P           *         E  �        �   �         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C1   #       +        �t�bhhK ��h��R�(KK��h�Ct   $   V  �     �     C   w         A              
      A     Z        �         �        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C �        	      	         �t�bhhK ��h��R�(KK��h�C8   �     �      *  L     �         �        �t�bhhK ��h��R�(KK��h�C4#   !      �        (      ^   Q           �t�bhhK ��h��R�(KK/��h�C�   R  %     �                             �  u      �     �     A   �     X         J   a   !         .   �      �     {      _     B     �  �         �t�bhhK ��h��R�(KK��h�Cd         0   �     �  �        (   �     �      �     w   �   �      `   /         �t�bhhK ��h��R�(KK��h�C4   W     :   �  �  �        ^            �t�bhhK ��h��R�(KK��h�C4�   ,   9  �     �      �  )      u         �t�bhhK ��h��R�(KK��h�CP        �   f     �         1   #   
   3   6     �   �            �t�bhhK ��h��R�(KK��h�C!      ,         �t�bhhK ��h��R�(KK��h�C0
        �     e  �                 �t�bhhK ��h��R�(KK��h�C�              �t�bhhK ��h��R�(KK��h�Cl�     �     +  �        �                       �      �     +  �     �   �         �t�bhhK ��h��R�(KK��h�C@,  L  �            �  &      H  �    
   �        �t�bhhK ��h��R�(KK��h�C>   �   v   r      �t�bhhK ��h��R�(KK��h�C,      )   b      #   !      �        �t�bhhK ��h��R�(KK��h�C          	      	         �t�bhhK ��h��R�(KK��h�Cb      x   
   �     �t�bhhK ��h��R�(KK	��h�C$`   b           �  �        �t�bhhK ��h��R�(KK��h�CW      �t�bhhK ��h��R�(KK��h�C    W  �   '      e         �t�bhhK ��h��R�(KK��h�CL2      =      �     �     �  �   �  7      �     J  /         �t�bhhK ��h��R�(KK��h�C0�        -  p         �      �        �t�bhhK ��h��R�(KK��h�C�     A   �     �t�bhhK ��h��R�(KK��h�C4Z         �     �  �      �     �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C8
   �   F   ?      -   1     \        +        �t�bhhK ��h��R�(KK��h�C0o  �      /      �      	      	         �t�bhhK ��h��R�(KK��h�C5     �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK	��h�C$�        .                 �t�bhhK ��h��R�(KK��h�C4*      �   F  &      U        8   �        �t�bhhK ��h��R�(KK��h�C      	      	   K      �t�bhhK ��h��R�(KK��h�Cp   �   :      Q   �  Y   �   Q     a   ;      f      �   �        .   %   �          f        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C 1   #       �              �t�bhhK ��h��R�(KK��h�C[      �     �t�bhhK ��h��R�(KK��h�C8                         <               �t�bhhK ��h��R�(KK
��h�C(�      �  	      	   K   	   �      �t�bhhK ��h��R�(KK��h�C%   �  O     �t�bhhK ��h��R�(KK
��h�C(         '  �  �   B   �        �t�bhhK ��h��R�(KK��h�C�      	      	         �t�bhhK ��h��R�(KK��h�C0�  �  .        5      �  
   6        �t�bhhK ��h��R�(KK��h�C/  q   0         �t�bhhK ��h��R�(KK��h�Cd�  �   |      �      �     �        1     �            J   �     �     W         �t�bhhK ��h��R�(KK��h�Cd      J   a   �  �       y              c  p            =      �     �         �t�bhhK ��h��R�(KK��h�Cd-      �     �     2   (   /         �  �  �   �      2   5   [         !  #        �t�bhhK ��h��R�(KK��h�C`      0   [                        ~            :     �     "              �t�bhhK ��h��R�(KK��h�C,b   #   "      �  V      J   z         �t�bhhK ��h��R�(KK��h�C2  R      �        �t�bhhK ��h��R�(KK��h�CT         �  G      �        =      [      C     "   $   �   �        �t�bhhK ��h��R�(KK��h�Cp9   �  (         j  <         �  �   |     x      "   >  D     �   �  V   2      0   <         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C0   Y      O   5      7                 �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK	��h�C$#     �   z      c  X  r      �t�bhhK ��h��R�(KK��h�C�   �     �     �t�bhhK ��h��R�(KK��h�C4V     3  &   N   
   ,                     �t�bhhK ��h��R�(KK��h�C1   #       	  l         �t�bhhK ��h��R�(KK��h�C          I   �  C         �t�bhhK ��h��R�(KK
��h�C(   E  j        k  j  /        �t�bhhK ��h��R�(KK��h�C<      b   "   W  W      �  \         0           �t�bhhK ��h��R�(KK��h�C,�     S     '   
   �   B   }         �t�bhhK ��h��R�(KK��h�C8   �  �     �   �  �  �  �  �  0  ;        �t�bhhK ��h��R�(KK
��h�C(�     I     �        �         �t�bhhK ��h��R�(KK��h�CL�      \  �   �      4     
   F  F      �   �  $     �        �t�bhhK ��h��R�(KK��h�C�     �  	         �t�bhhK ��h��R�(KK��h�Cl�   &   �     �      G       %   H  �     �   "   �  �  �  �   �     Y  �      �        �t�bhhK ��h��R�(KK��h�CD      �                    �  �          �        �t�bhhK ��h��R�(KK��h�C8?         �  �   I  V         =      n         �t�bhhK ��h��R�(KK��h�C�     A   �      �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6   t        �t�bhhK ��h��R�(KK��h�C�  4   �     �t�bhhK ��h��R�(KK��h�C1   #       i        �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�C�  5     �t�bhhK ��h��R�(KK��h�C4   &   a      +   J  
   �   $     k        �t�bhhK ��h��R�(KK	��h�C$6  �           �           �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C7  �  
   �     �t�bhhK ��h��R�(KK��h�C0      �   �         )  +   
   &        �t�bhhK ��h��R�(KK��h�C4      6  +      �  �        d  G        �t�bhhK ��h��R�(KK��h�Cd      V  �  �        5   [         U   @     �     e      �      �      �        �t�bhhK ��h��R�(KK��h�C`      D   &   D  0   4   >   P  �   �  �        N   �        .   �     �        �t�bhhK ��h��R�(KK��h�CH      �     o  ~             ?      8  
   8           �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�C�  R      �t�bhhK ��h��R�(KK��h�C,   �                            �t�bhhK ��h��R�(KK��h�C4�  �          �        �        �     �t�bhhK ��h��R�(KK��h�C   �  
   �     �t�bhhK ��h��R�(KK��h�C[   "   �     �t�bhhK ��h��R�(KK��h�C�      D      �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�C@      ]  �     �  Q     �  &   �   �             �t�bhhK ��h��R�(KK��h�C0   �  I    	     Y      O   �  �         �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   6   �     �        �t�bhhK ��h��R�(KK��h�C@   &   T   �     E      	     �           
        �t�bhhK ��h��R�(KK��h�C@�     �      N   �     �   �     %   �      I         �t�bhhK ��h��R�(KK��h�C0�   �     �   9  �     �  i   �         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK	��h�C$~     l      :        �     �t�bhhK ��h��R�(KK��h�C E      �  	      	         �t�bhhK ��h��R�(KK��h�C   
   �     �t�bhhK ��h��R�(KK��h�C
      5     �        �t�bhhK ��h��R�(KK��h�C<
   �   F   ?      �     �     #   !      P        �t�bhhK ��h��R�(KK��h�C4   .   (   �     a   �   <       <        �t�bhhK ��h��R�(KK��h�C8�
     )   N      �
                 �        �t�bhhK ��h��R�(KK��h�C<�   �        >   ;  �       %   &             �t�bhhK ��h��R�(KK��h�C0d  
   \   8   �  �  �  �     �        �t�bhhK ��h��R�(KK��h�CL
   Z        R  �     �          �     	     �   S         �t�bhhK ��h��R�(KK��h�CJ     /      �t�bhhK ��h��R�(KK��h�C    �  �   0  B   [        �t�bhhK ��h��R�(KK
��h�C(�  a  �     �  9   �  �        �t�bhhK ��h��R�(KK��h�C@      �  #      S     �  
   3   6   �             �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C`   �           %                    �
     8   �     $   A     $   p         �t�bhhK ��h��R�(KK��h�CT�        �  �            �  K  G   /      T  �   D   %   �  	        �t�bhhK ��h��R�(KK��h�C0  �     >     U     �   �   B         �t�bhhK ��h��R�(KK��h�C4   (   #   !      �     $   x  
   k        �t�bhhK ��h��R�(KK��h�C@a     G  P     $   �   �  s   �   y      �   <        �t�bhhK ��h��R�(KK��h�C�  �      �t�bhhK ��h��R�(KK��h�C@k     e      �  �     �     �   
   H   B           �t�bhhK ��h��R�(KK��h�C�  �     �  �  �     �t�bhhK ��h��R�(KK��h�C   (   �  9   �        �t�bhhK ��h��R�(KK��h�C      @          �t�bhhK ��h��R�(KK��h�C�  �          �     �t�bhhK ��h��R�(KK��h�C01   #   
   3   6   �     �     �        �t�bhhK ��h��R�(KK(��h�C��           P     2      �            �      �     �     =  i   A      .   
   _      L  �     >     �          X     d        �t�bhhK ��h��R�(KK��h�C8�  	  �   	  9   �            �
              �t�bhhK ��h��R�(KK��h�Cx   D         �     �   S        #     D      �   �           V     �      �   	  V              �t�bhhK ��h��R�(KK��h�C\               k         &        W   �  $   ;         �        �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C4      �  
         �  )   
   A   }         �t�bhhK ��h��R�(KK��h�Ce         �t�bhhK ��h��R�(KK
��h�C(#   !   '   
   �   �  ?  F         �t�bhhK ��h��R�(KK��h�C<�      �  v   �        �     ,      $   @        �t�bhhK ��h��R�(KK��h�C�      /              �t�bhhK ��h��R�(KK��h�C0      �      A     �   �     "        �t�bhhK ��h��R�(KK��h�C8�  	  +            �     �         �        �t�bhhK ��h��R�(KK��h�CL      q   B  �     �     ,        �  �  C  �     �        �t�bhhK ��h��R�(KK��h�CD   (   z         A     _  *      a          �
        �t�bhhK ��h��R�(KK��h�CX      -   P   n   ^   %  �  	     �     �  	     �                    �t�bhhK ��h��R�(KK��h�C0�        �  �            ;   �        �t�bhhK ��h��R�(KK��h�C4   5   &        �      		     $   �         �t�bhhK ��h��R�(KK��h�C,D        �           �            �t�bhhK ��h��R�(KK��h�CH*         E  H        ;      G        �  $   E   �        �t�bhhK ��h��R�(KK��h�C4�     T   a   e  �     l  �     D         �t�bhhK ��h��R�(KK��h�CH   `   b  �   �     e  9   y     &      
     �          �t�bhhK ��h��R�(KK��h�CB  �     �  �        �t�bhhK ��h��R�(KK��h�C@         �      �      7      �  F     +  �        �t�bhhK ��h��R�(KK��h�C   �  �             �t�bhhK ��h��R�(KK��h�Cd\      j     	      	      	   K   	   �   	   �   	     	   �   	   �  	   �  	   /     �t�bhhK ��h��R�(KK��h�C4E   &   �  y         �  �   �   s   7         �t�bhhK ��h��R�(KK��h�C,�     \   �         �     :        �t�bhhK ��h��R�(KK��h�C�   ]  �               �t�bhhK ��h��R�(KK��h�C   �              �t�bhhK ��h��R�(KK��h�C
	  =     �     �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C,^   �   �  �     R      �   �         �t�bhhK ��h��R�(KK��h�C@�      (  �  u      �      ,   �                    �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C4]   P        �                 G        �t�bhhK ��h��R�(KK��h�C8#   !      �  '   
   3   6   �  t              �t�bhhK ��h��R�(KK��h�C\      r  '  (      !      p      ,                  p      R      X         �t�bhhK ��h��R�(KK��h�C �     m  �                �t�bhhK ��h��R�(KK��h�C,m  �  �     �           X        �t�bhhK ��h��R�(KK��h�C<1   #      ,   �       �  
   3   6   	  �         �t�bhhK ��h��R�(KK��h�Cd   �      $     �  �   Y  +      �  +      �            U      �     	           �t�bhhK ��h��R�(KK
��h�C(   '      �     	     H        �t�bhhK ��h��R�(KK��h�C0�        �     y     �      �        �t�bhhK ��h��R�(KK��h�C�   p      �t�bhhK ��h��R�(KK��h�CI               �t�bhhK ��h��R�(KK��h�C0      h  �  �  �     S      5        �t�bhhK ��h��R�(KK��h�C,*        �  &      �     E          �t�bhhK ��h��R�(KK��h�CP�          �                 W       b  �      �  	        �t�bhhK ��h��R�(KK��h�C	  J  
            �t�bhhK ��h��R�(KK��h�C K     	                 �t�bhhK ��h��R�(KK��h�C	     �      �         �t�bhhK ��h��R�(KK
��h�C(         L  +         �        �t�bhhK ��h��R�(KK��h�C,-   n  �  7      :   M     @         �t�bhhK ��h��R�(KK��h�CH�   =  �  >     ,      A   �         E  9      �            �t�bhhK ��h��R�(KK��h�CP   @   '      -   �   e     �   
   �        /     �      K         �t�bhhK ��h��R�(KK��h�CX:   Q     z  (      M      +      j  �     �   �
     �     �  �
        �t�bhhK ��h��R�(KK��h�CP)   A   6        �            4   
   _      X  �     R  4         �t�bhhK ��h��R�(KK��h�C�  �     %   �         �t�bhhK ��h��R�(KK��h�C   +     �t�bhhK ��h��R�(KK��h�C�  
   ,      �t�bhhK ��h��R�(KK��h�C8     
   \   �             Y              �t�bhhK ��h��R�(KK
��h�C(�  �           M     	        �t�bhhK ��h��R�(KK��h�C,f         �  h        g            �t�bhhK ��h��R�(KK��h�CP      R  H           �          �   �     8   E  
   _         �t�bhhK ��h��R�(KK��h�C,j   �    �   �     �  
   �  N     �t�bhhK ��h��R�(KK��h�C,E      f   O  (  �      �  E         �t�bhhK ��h��R�(KK��h�CL�   v              �  $   k            �   s   7               �t�bhhK ��h��R�(KK	��h�C$�  (   �                    �t�bhhK ��h��R�(KK��h�C4         �  +      �     �  $           �t�bhhK ��h��R�(KK��h�C	  	         �t�bhhK ��h��R�(KK��h�C)     �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�Cl         .         D   ~   G      �  �           A   �  �
  �     �   f   Z  9            �t�bhhK ��h��R�(KK��h�CPB   P          �     �     �     �           	     �        �t�bhhK ��h��R�(KK��h�CD              �           (      v     �           �t�bhhK ��h��R�(KK��h�C\y      �  $   �     1   Q  S     d  
            �  �      R  g         �t�bhhK ��h��R�(KK��h�C        �  �        �t�bhhK ��h��R�(KK	��h�C$/   9   �  7   5      �
        �t�bhhK ��h��R�(KK��h�C             �t�bhhK ��h��R�(KK��h�C�     S  �     �t�bhhK ��h��R�(KK��h�CH   <               *  3   �  
   A   _     �  B            �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C0!      .  '   
   T     u      X         �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C@   �     �t�bhhK ��h��R�(KK��h�C�  �      N      .      �t�bhhK ��h��R�(KK��h�CD   �   �     	  	        v  �  �  u  c   �           �t�bhhK ��h��R�(KK��h�CP.  "   �     �          <     �     /     ~   �               �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C8   @   '   H   �   	     )   �   �      /         �t�bhhK ��h��R�(KK��h�C8               �  6     �     8   �        �t�bhhK ��h��R�(KK��h�CP1   #      �             �   f  
   3   6     �   �               �t�bhhK ��h��R�(KK��h�C   y     �t�bhhK ��h��R�(KK��h�C�   	  	         �t�bhhK ��h��R�(KK��h�C�  Y  �         �t�bhhK ��h��R�(KK��h�Cl     �  Q  p      u      �     �     �   �  �     A        �        z   "           �t�bhhK ��h��R�(KK��h�C<
   3   6   �     j   4   '      #   !      �        �t�bhhK ��h��R�(KK��h�CL      0   [         
   _      8   �     $   \  5   0  <         �t�bhhK ��h��R�(KK��h�CR      T     �t�bhhK ��h��R�(KK��h�C�   =     �t�bhhK ��h��R�(KK��h�CL              /               b   x   "                     �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C       �  �   7  �        �t�bhhK ��h��R�(KK��h�Cm      �         :     �t�bhhK ��h��R�(KK��h�C
   �  �  [  �        �t�bhhK ��h��R�(KK��h�C<N  7  P   �  :      	      	      	   K   	   �      �t�bhhK ��h��R�(KK��h�C	  �     �t�bhhK ��h��R�(KK��h�C@7         !  �     @      4        n  U  o        �t�bhhK ��h��R�(KK��h�Ch      \  	           �  c         ]     (        ^  )      $   k         X         �t�bhhK ��h��R�(KK��h�CH   &   �  "   �        	  u     �   "   q   �     u        �t�bhhK ��h��R�(KK��h�C`      �                  V     �          �                     �         �t�bhhK ��h��R�(KK��h�CK         �      �     �t�bhhK ��h��R�(KK��h�C�     x  �           �t�bhhK ��h��R�(KK	��h�C$�      �   9   z  q   .        �t�bhhK ��h��R�(KK��h�C O     	  �      ?        �t�bhhK ��h��R�(KK
��h�C(            �        N  �     �t�bhhK ��h��R�(KK��h�C,_        �  �     �      �        �t�bhhK ��h��R�(KK��h�C4     G  �   [      �      G     �        �t�bhhK ��h��R�(KK��h�C[      �      �t�bhhK ��h��R�(KK��h�C8   (   !      \      ]  �  
   3   6   	        �t�bhhK ��h��R�(KK��h�C�   >   5  �        �t�bhhK ��h��R�(KK��h�C !      �  	      	         �t�bhhK ��h��R�(KK��h�CHk  �  	  
   N              V  �      O     9           �t�bhhK ��h��R�(KK��h�C   �  	      	         �t�bhhK ��h��R�(KK��h�C	  �          �t�bhhK ��h��R�(KK��h�C8
   �     5     -   \   '     $   E   W        �t�bhhK ��h��R�(KK��h�C<         .   �     �  >      w   v   �           �t�bhhK ��h��R�(KK��h�C8      '   P  �     �        �              �t�bhhK ��h��R�(KK��h�C,     &      �         �   	  r      �t�bhhK ��h��R�(KK��h�C X     �  
   ]  L         �t�bhhK ��h��R�(KK��h�C1   #       �  4         �t�bhhK ��h��R�(KK��h�C@   �                  �     Q     �  �  �        �t�bhhK ��h��R�(KK��h�C0b     �     =  �  >         �        �t�bhhK ��h��R�(KK��h�C    E  j     j  /        �t�bhhK ��h��R�(KK��h�C4*   r  $  �     0     D     +  2        �t�bhhK ��h��R�(KK	��h�C$   �  +  '   �  �           �t�bhhK ��h��R�(KK��h�C#  �     p  r      �t�bhhK ��h��R�(KK
��h�C(�     !	     -      P           �t�bhhK ��h��R�(KK��h�C"	  �     �t�bhhK ��h��R�(KK��h�Cl�   q   7  &   �  Y  �   �           �   O      +  l           q     +   '      �        �t�bhhK ��h��R�(KK��h�C02      �   �   >  �  y                  �t�bhhK ��h��R�(KK��h�C<      '   H   �     �             #	           �t�bhhK ��h��R�(KK��h�C�  	         �t�bhhK ��h��R�(KK	��h�C$   @   '   �       `        �t�bhhK ��h��R�(KK��h�C@$	  �         �      �  �        �  �     `        �t�bhhK ��h��R�(KK��h�C8�   ^                        �     Y        �t�bhhK ��h��R�(KK��h�C,1   #   
   3   6   �  t              �t�bhhK ��h��R�(KK��h�C4*   �     a     2   =      Z     �        �t�bhhK ��h��R�(KK	��h�C$     �  Y  �      7         �t�bhhK ��h��R�(KK��h�C<
   �   F   ?      �     �     #   !      P        �t�bhhK ��h��R�(KK��h�C\   f   s  �      2   [  :   %	        '   �  �          d   b  (  ]         �t�bhhK ��h��R�(KK��h�C <         0   �  
   �      �t�bhhK ��h��R�(KK��h�CD1   #      b     ,     �   p   
   3   6   �     /         �t�bhhK ��h��R�(KK��h�C2   >   2     �        �t�bhhK ��h��R�(KK
��h�C(   >   =      \  �  :   W         �t�bhhK ��h��R�(KK
��h�C(q     �     �  	      	         �t�bhhK ��h��R�(KK��h�CH�     )   �     �  �     \   �  &         �
    ]        �t�bhhK ��h��R�(KK*��h�C�         O         Y      Q      �     x     J   �                �        .   
   �     
               \  �     5      7  L        �t�bhhK ��h��R�(KK��h�C1   #               �t�bhhK ��h��R�(KK��h�C0            �     �        K        �t�bhhK ��h��R�(KK��h�C        �t�bhhK ��h��R�(KK��h�C�
  	      	         �t�bhhK ��h��R�(KK��h�CL      ,  %   �                    k      l                 �t�bhhK ��h��R�(KK��h�Cd      -   �  �      �   �     �  �  '  G   C         &	     �     8   �   S        �t�bhhK ��h��R�(KK��h�C8      -   �  ^  
        "   �     �        �t�bhhK ��h��R�(KK��h�C �      '	        	         �t�bhhK ��h��R�(KK
��h�C(�     �        �  �  �        �t�bhhK ��h��R�(KK
��h�C(!         N  �  	      	         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CtY      �       X     -  J  C      �   h   �  �     X     �     �  �      (	     Y      �     �t�bhhK ��h��R�(KK��h�C8)   �  �  =     %      �   �  i   A   =        �t�bhhK ��h��R�(KK��h�C4        J  �     K     X               �t�bhhK ��h��R�(KK��h�C    (   [      �            �t�bhhK ��h��R�(KK��h�C4[      C     	      	      	   �  	   �      �t�bhhK ��h��R�(KK��h�C,N     �      d      	      	         �t�bhhK ��h��R�(KK��h�C   �  g   �            �t�bhhK ��h��R�(KK��h�C@              0   L   G      �  Z        J         �t�bhhK ��h��R�(KK
��h�C($  �  �   .        O  �        �t�bhhK ��h��R�(KK��h�C      �  �        �t�bhhK ��h��R�(KK��h�C`   `   �            .   Y  �  i   s   7      &   �  �  �  �      �      �        �t�bhhK ��h��R�(KK
��h�C(�    
         $   �            �t�bhhK ��h��R�(KK��h�C,      B   �     �  	      	         �t�bhhK ��h��R�(KK��h�C|      �      R          /  �       �     �      -  �     _     �        �     /   �   )	        �t�bhhK ��h��R�(KK��h�C4             0                       �t�bhhK ��h��R�(KK��h�CLq   �  �  �         �  x                 *   �   
  4         �t�bhhK ��h��R�(KK��h�CP      �        /  i        f   ?     /  i  �  +               �t�bhhK ��h��R�(KK��h�Cb   #   G   W         �t�bhhK ��h��R�(KK��h�CH*      �         �     C  W            ;      �   �        �t�bhhK ��h��R�(KK
��h�C(      c     +     �  �         �t�bhhK ��h��R�(KK��h�C?      �     �        �t�bhhK ��h��R�(KK
��h�C(      -   P         �  *	        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C4   (   1     \   ]   /  8   @     �        �t�bhhK ��h��R�(KK��h�C4   �        `  N               a        �t�bhhK ��h��R�(KK��h�C8#   !         =      �   ?      
   �  F         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C,      �   >      a      �          �t�bhhK ��h��R�(KK��h�C8   &   =      �  4   y   8   3  4     c         �t�bhhK ��h��R�(KK��h�C �   �  ^   �  �           �t�bhhK ��h��R�(KK��h�C<1   #         U        
   3   6   �
              �t�bhhK ��h��R�(KK��h�C<   X   '   )               �   p      B            �t�bhhK ��h��R�(KK��h�C4�     �  �      ,      A   �      �        �t�bhhK ��h��R�(KK��h�C E         	      	         �t�bhhK ��h��R�(KK��h�CH   .   W      b     �     �     f   �      &     �        �t�bhhK ��h��R�(KK��h�C,Y      O   &   -   F  C   
   H        �t�bhhK ��h��R�(KK��h�CS            �t�b�&      hhK ��h��R�(KK��h�CT         m      �     A   �     +	        M   �      �              �t�bhhK ��h��R�(KK��h�CP        i          $   n            �             ]         �t�bhhK ��h��R�(KK��h�C�  	      	         �t�bhhK ��h��R�(KK��h�C   x         �t�bhhK ��h��R�(KK��h�C    	      	      	   K      �t�bhhK ��h��R�(KK��h�C�  	      	         �t�bhhK ��h��R�(KK��h�Cd      "        s  �   [  :   %	           '   �  �          d   b  (  ]         �t�bhhK ��h��R�(KK��h�CD%     m  �            �  c           �     u         �t�bhhK ��h��R�(KK��h�C,      N   :      �     �   �         �t�bhhK ��h��R�(KK��h�CX!               	      	   K   	   �   	   I  	   U  	   /  	   �  	   �     �t�bhhK ��h��R�(KK��h�CdT      d     (   �      �   �   �     d  �   �  
   _      L  �     d     �        �t�bhhK ��h��R�(KK��h�CD$  �  �  �     >   �  $   0     *  �   �     �        �t�bhhK ��h��R�(KK��h�C0I   u      ;      0   �   !               �t�bhhK ��h��R�(KK��h�C  p      u      �t�bhhK ��h��R�(KK��h�CHw  �  (   #   !      ]   �   s     
   �  F         e        �t�bhhK ��h��R�(KK��h�C0�  "        Q     /   9     7         �t�bhhK ��h��R�(KK��h�C,1   #   
   3   6   �     �  �         �t�bhhK ��h��R�(KK��h�C0�  �       6     �     
            �t�bhhK ��h��R�(KK	��h�C$         f     M   ,	        �t�bhhK ��h��R�(KK��h�C0�     2     :     �   +     -	        �t�bhhK ��h��R�(KK��h�CX      '   -   �        �      �        .         M  �        �        �t�bhhK ��h��R�(KK��h�C,�   �   2      T          <        �t�bhhK ��h��R�(KK��h�C C  �     M     {        �t�bhhK ��h��R�(KK��h�C!           �        �t�bhhK ��h��R�(KK��h�CL�  g     �        ;            /      ;      )	  h   �         �t�bhhK ��h��R�(KK��h�Ch      )        <      x   "   Q  	     �           "   <              .            �t�bhhK ��h��R�(KK	��h�C$4   
   A      	      	         �t�bhhK ��h��R�(KK��h�C4      ]  I        �  �   !      �         �t�bhhK ��h��R�(KK��h�C�  �         �t�bhhK ��h��R�(KK��h�C   �               �t�bhhK ��h��R�(KK
��h�C(�     W  .	     N       r      �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C4*               :      n         �          �t�bhhK ��h��R�(KK��h�C4!         ?      
   �  F      
            �t�bhhK ��h��R�(KK��h�C@*   h     �  /  `        $   /	     �  b           �t�bhhK ��h��R�(KK��h�CTN  �     �  	      	      	   K   	   �   	     	   �  	   �   	   �     �t�bhhK ��h��R�(KK��h�C@1   #         �  `   �  
   3   6   �  g  �   �        �t�bhhK ��h��R�(KK��h�C<   @   '      �   5     ]     4     �   5        �t�bhhK ��h��R�(KK��h�Cq     �t�bhhK ��h��R�(KK
��h�C(   �           0	  �           �t�bhhK ��h��R�(KK��h�C      1	  2	        �t�bhhK ��h��R�(KK	��h�C$�     I  �     3	           �t�bhhK ��h��R�(KK	��h�C$T      D   4	  �  �   �        �t�bhhK ��h��R�(KK��h�C   �  �         �t�bhhK ��h��R�(KK��h�Ci     �  5	  	         �t�bhhK ��h��R�(KK��h�C�     �  �      �t�bhhK ��h��R�(KK��h�C8   �      �     %   �  6	  7	  �      D         �t�bhhK ��h��R�(KK��h�C,   B        �      �     U        �t�bhhK ��h��R�(KK��h�C   �  T     j        �t�bhhK ��h��R�(KK
��h�C(_        	      	     	   �      �t�bhhK ��h��R�(KK��h�C01   #   
   3   6         �     �         �t�bhhK ��h��R�(KK��h�CZ      �      �     �t�bhhK ��h��R�(KK��h�C   �      �  �     �t�bhhK ��h��R�(KK��h�Ck          1        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C /  ^  @     �  �         �t�bhhK ��h��R�(KK��h�C<   �        
      \        �        ?        �t�bhhK ��h��R�(KK��h�C<�   	  V  �     D   ~   �   e  i   G   �   8        �t�bhhK ��h��R�(KK��h�CK             �     �t�bhhK ��h��R�(KK��h�C4      ,  ?      �  �      �  �  �        �t�bhhK ��h��R�(KK��h�CH      G        j   4         �  �  V     v      	        �t�bhhK ��h��R�(KK	��h�C$#  �   �   �  8	     �        �t�bhhK ��h��R�(KK��h�C8        �  O      �t�bhhK ��h��R�(KK
��h�C(I   k  �  �     �     9	        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C,d  
     �     %        5         �t�bhhK ��h��R�(KK��h�C<#   !         �     (      G         $   k         �t�bhhK ��h��R�(KK��h�C4�  '                L   T   �   �        �t�bhhK ��h��R�(KK��h�C       �   �      I         �t�bhhK ��h��R�(KK��h�C#     �   r      �t�bhhK ��h��R�(KK��h�C{      �t�bhhK ��h��R�(KK��h�CL*         8   �   �      @      &      F  +           <        �t�bhhK ��h��R�(KK��h�CDE   &   r  �      W   �     �  y               �        �t�bhhK ��h��R�(KK��h�Cl  :	     ;	        �t�bhhK ��h��R�(KK��h�C<�     a   
  �     O     %            m        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C  n  
   4     �t�bhhK ��h��R�(KK��h�C          �      I         �t�bhhK ��h��R�(KK��h�C<            &   r     2  �     �  g   $	        �t�bhhK ��h��R�(KK��h�C  �   m     �        �t�bhhK ��h��R�(KK��h�CX              W  V   X        S   i   ,                 
   �         �t�bhhK ��h��R�(KK��h�CP�      L   G      o           .      m      p     <	              �t�bhhK ��h��R�(KK��h�C@            h  �       �  �     q     �        �t�bhhK ��h��R�(KK��h�C8
      =    +         r  �  	      	         �t�bhhK ��h��R�(KK��h�C\         m      s     �           M   �      �                x          �t�bhhK ��h��R�(KK��h�Ct      �           �        
   _      �        �     �     s        ;         r  �        �t�bhhK ��h��R�(KK��h�C �      d   8  �  �        �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�CP*      �  
   %       &   �                       t  �        �t�bhhK ��h��R�(KK��h�C0   Y     �   '      �     q           �t�bhhK ��h��R�(KK��h�C,  I        	      	   K   	   �      �t�bhhK ��h��R�(KK��h�Cb   #   "   $   �        �t�bhhK ��h��R�(KK��h�C0+     -	  �   +   =	        �  �        �t�bhhK ��h��R�(KK��h�C4     �   �      >	     �         �        �t�bhhK ��h��R�(KK	��h�C$      U     �     ?	        �t�bhhK ��h��R�(KK��h�C !        	      	         �t�bhhK ��h��R�(KK��h�C0   	        �   k     a     �        �t�bhhK ��h��R�(KK��h�C,Z      �               �            �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C<N  �        ,      	   K   	   �   	     	   �      �t�bhhK ��h��R�(KK��h�C43  �        �     '  
      �   �        �t�bhhK ��h��R�(KK��h�C  (         �        �t�bhhK ��h��R�(KK��h�CD   @	  �
     .      u  �  
               <        �t�bhhK ��h��R�(KK��h�C         b  �           �t�bhhK ��h��R�(KK��h�C,      �      �        �  �         �t�bhhK ��h��R�(KK��h�C4      �        0        �             �t�bhhK ��h��R�(KK��h�C,           T   A	  2   v           �t�bhhK ��h��R�(KK��h�CDM     
               �   A   w        D  v   �        �t�bhhK ��h��R�(KK1��h�CĦ     N   �     .   *   2      :      Q         S         m   
   �     x  �   �        m      �        �  �      x     �     �   F     *   �     
   A           �t�bhhK ��h��R�(KK
��h�C(#   !   ?      
   @   �   F         �t�bhhK ��h��R�(KK��h�C<^   �                  P   !   �   B	     �        �t�bhhK ��h��R�(KK��h�CH   @      �  u   ;      0   �     y  �   h   %   �           �t�bhhK ��h��R�(KK��h�C0W  �     �  B  8   �        t        �t�bhhK ��h��R�(KK��h�C    4  
   t         �t�bhhK ��h��R�(KK��h�C0      0   �     C	     $   �   �        �t�bhhK ��h��R�(KK��h�CZ   .     z        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�CLD   (   �  �  {   �       �              �  �      �        �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C         {         �t�bhhK ��h��R�(KK��h�C +     )   �     �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C@\      �      �     M    
        Q      ~         �t�bhhK ��h��R�(KK��h�C 5   �      �      �  r      �t�bhhK ��h��R�(KK��h�C0R      ]           S                  �t�bhhK ��h��R�(KK	��h�C$      2     c  X           �t�bhhK ��h��R�(KK��h�CL  h   �  �   :      B   ?     X     ,         �     a   �     �t�bhhK ��h��R�(KK��h�CX   5  _  D   �     �   f     _  C      ,   �              �  �        �t�bhhK ��h��R�(KK��h�Ch   D	  
   �         �  ?               ^   %        �  ?     �   �  �  
   T        �t�bhhK ��h��R�(KK��h�C�      D      V     �t�bhhK ��h��R�(KK��h�CN  7      �t�bhhK ��h��R�(KK��h�CD-   H   �    �   �      .      �     !       @        �t�bhhK ��h��R�(KK��h�CL         8   �   �           &      F  +           <        �t�bhhK ��h��R�(KK
��h�C(�  {           �             �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�CX   >   =         �  4   
   _      {   y   8   4         P   {     c         �t�bhhK ��h��R�(KK��h�CX"   X   E	     g           2      .   �  �     |     F	  �     }        �t�bhhK ��h��R�(KK��h�Cp            Z        S   Y      Q      Q     Q         x        ;      y  ^              �t�bhhK ��h��R�(KK	��h�C$"   G	        )   �   +        �t�bhhK ��h��R�(KK��h�CX     �   �     �t�bhhK ��h��R�(KK��h�C�  T     �t�bhhK ��h��R�(KK��h�Cb      	      	         �t�bhhK ��h��R�(KK��h�C<�   7        ;      �  e  ,                     �t�bhhK ��h��R�(KK��h�C,f   �     @        �  
   ~        �t�bhhK ��h��R�(KK��h�C )     T      $   �        �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C,   �   �             G   �         �t�bhhK ��h��R�(KK��h�Cp   Y        S   X  i   ,            �  �  �     T        �  P        �                �t�bhhK ��h��R�(KK��h�CP   R      �t�bhhK ��h��R�(KK��h�C0      :     �   
   ,      
            �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C
  �     �t�bhhK ��h��R�(KK	��h�C$p         M  	      	         �t�bhhK ��h��R�(KK��h�C       z   ,      X        �t�bhhK ��h��R�(KK��h�Cx     �  �   O     ;     I   %   /      �           �  �        �  C      �  h      �   �         �t�bhhK ��h��R�(KK��h�C\   w   �   �
              �     �       �        P      n      +         �t�bhhK ��h��R�(KK��h�CT
        2   �   0  p  
   z  �   7      �  �  p  
   z  s   7         �t�bhhK ��h��R�(KK��h�C1   #       �        �t�be(hhK ��h��R�(KK��h�C4      m     �t�bhhK ��h��R�(KK��h�C	     �t�bhhK ��h��R�(KK��h�C4#   !         k  �  (      
   u  F         �t�bhhK ��h��R�(KK��h�CH         �     7         0   �  �  �  �   $               �t�bhhK ��h��R�(KK��h�C,      �  �   �  G     �  �         �t�bhhK ��h��R�(KK	��h�C$�   �   E           �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK	��h�C$T   >      v      [  w         �t�bhhK ��h��R�(KK��h�Ch  =     �t�bhhK ��h��R�(KK��h�CH7  �  �   H	          �      z  M     {  �     U        �t�bhhK ��h��R�(KK
��h�C(j                   /        �t�bhhK ��h��R�(KK��h�C0�     `        �  d         �        �t�bhhK ��h��R�(KK��h�CL         4      k                  ;      Q  R      	        �t�bhhK ��h��R�(KK��h�C<'  �  
      
   �   }       ,                     �t�bhhK ��h��R�(KK��h�C4�  $   �        �  s   �   y      l        �t�bhhK ��h��R�(KK��h�CD   �   b     �      �        �     ,   	      	         �t�bhhK ��h��R�(KK��h�C,�      (     �  )   �      �         �t�bhhK ��h��R�(KK��h�CD                 &      U   |      �   y      �         �t�bhhK ��h��R�(KK��h�CH
   �  F   '   \     B   I  V         z   ,   
   �   �         �t�bhhK ��h��R�(KK��h�C@�  ]  �  I	  �     �  �   J	  
   _      d   �         �t�bhhK ��h��R�(KK��h�Cb        �      �t�bhhK ��h��R�(KK��h�C h  �  K	  "              �t�bhhK ��h��R�(KK��h�C0g   �     2   �   E         d  E         �t�bhhK ��h��R�(KK��h�C0   "   >  0   <      �                 �t�bhhK ��h��R�(KK
��h�C(T            ;      �   �        �t�bhhK ��h��R�(KK��h�C8      v            �              �        �t�bhhK ��h��R�(KK
��h�C(1   #      �  
   3   6            �t�bhhK ��h��R�(KK��h�C8         5   �       �  g   �      �        �t�bhhK ��h��R�(KK��h�C   i     �t�bhhK ��h��R�(KK��h�C4      �
  8  �
     Z       �  �        �t�bhhK ��h��R�(KK��h�C�  >      
   c        �t�bhhK ��h��R�(KK��h�C         
   s            �t�bhhK ��h��R�(KK��h�C 1  ^     /        �     �t�bhhK ��h��R�(KK	��h�C$�  �   L	  �   +     "        �t�bhhK ��h��R�(KK��h�C8   �   �  �   C      8   S     �  j  /        �t�bhhK ��h��R�(KK��h�C �        k               �t�bhhK ��h��R�(KK��h�C,            �     �   �   /         �t�bhhK ��h��R�(KK��h�C@      �     �           >      F  +              �t�bhhK ��h��R�(KK��h�CP            �     i  �   �     �     �  �   �     �  �        �t�bhhK ��h��R�(KK��h�Cx            M	  \  &      M      `   .  �     �
  �      �  R  �   *   �      �   �  c      �        �t�bhhK ��h��R�(KK��h�C0      f  '            �  
   �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6   N	        �t�bhhK ��h��R�(KK��h�Cj  g  k     �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�  O	  �         �t�bhhK ��h��R�(KK��h�C@      )   M   �   
      �   �     
   �               �t�bhhK ��h��R�(KK��h�C8!              	      	      	   K   	   ^     �t�bhhK ��h��R�(KK��h�CH:   �   �  '   �   �     @      A        u                 �t�bhhK ��h��R�(KK��h�C,.     �  �      B        u        �t�bhhK ��h��R�(KK��h�Cd      P	          �  V   X     ,   :  D   -         �  }   �      %   6  �        �t�bhhK ��h��R�(KK	��h�C$      �   5           Q	     �t�bhhK ��h��R�(KK��h�C_     (         �t�bhhK ��h��R�(KK��h�C  2       x     �t�bhhK ��h��R�(KK��h�Ch         �  �         o  O         l              0   4         
   _      �        �t�bhhK ��h��R�(KK��h�C4!        h  �     �                   �t�bhhK ��h��R�(KK��h�CD     .     7  R	  
     l      S	           7        �t�bhhK ��h��R�(KK��h�Cm      4      �t�bhhK ��h��R�(KK��h�Ct-      /      �  8     �           0   o  �         �     (   �      �   S   Q      �   8        �t�bhhK ��h��R�(KK
��h�C(2      0         �              �t�bhhK ��h��R�(KK��h�C0"  #  \   I  �        �               �t�bhhK ��h��R�(KK��h�C`      �   �  i   d        �  �      4   >   l  T	     .   �            U	        �t�bhhK ��h��R�(KK��h�CT      �  =      �  &      U   �      (        �   �  �     "        �t�bhhK ��h��R�(KK��h�C,   ?   #   !         
   $  F         �t�bhhK ��h��R�(KK��h�C@      �      �  L      ]   S     �     B   ?        �t�bhhK ��h��R�(KK��h�C\      �         T     �   5     &      �  �   $   E   �   �  �   �            �t�bhhK ��h��R�(KK��h�CD      �      �  �         �   �      �  *   %  ]        �t�bhhK ��h��R�(KK��h�C4&  �   �   �  O      '                    �t�bhhK ��h��R�(KK��h�C4      �     �  V	        �  �   �        �t�bhhK ��h��R�(KK��h�CX   �   R      u   �     �t�bhhK ��h��R�(KK��h�C,      )  8   /      �      �        �t�bhhK ��h��R�(KK��h�C,#   !      P  '   
   �     F         �t�bhhK ��h��R�(KK��h�CW	     �t�bhhK ��h��R�(KK��h�C8(  )  *  �  0  �     +           �        �t�bhhK ��h��R�(KK��h�C01     �   	  ?         .   
           �t�bhhK ��h��R�(KK��h�C   5   ,     8   �     �t�bhhK ��h��R�(KK��h�C@      0   -  
   �   |  -   *   $   k   �   $   �         �t�bhhK ��h��R�(KK��h�CT            v  �     5      -               �  
   �     @        �t�bhhK ��h��R�(KK	��h�C$      �  �     �
  �
        �t�bhhK ��h��R�(KK��h�C@d  
   \      &   �  ^  8   �     $         �        �t�bhhK ��h��R�(KK��h�C8*      �       �     C      )   �  X	        �t�bhhK ��h��R�(KK��h�C0   %   �  .     X  �  ,               �t�bhhK ��h��R�(KK��h�C�  "   �     �t�bhhK ��h��R�(KK��h�C<*   �  �     �     �        \   �     �        �t�bhhK ��h��R�(KK��h�C @     /  	      	         �t�bhhK ��h��R�(KK��h�C@   �        �  +      &      U   Y	  �     Z	        �t�bhhK ��h��R�(KK��h�C�   �     �t�bhhK ��h��R�(KK��h�C,   @         �   `     H   3        �t�bhhK ��h��R�(KK��h�CH   2   �     �     2   �       <     �  �   �   {         �t�bhhK ��h��R�(KK��h�C0�  �  
   ,            K      �         �t�bhhK ��h��R�(KK��h�C f   ?  �   �   �  �        �t�bhhK ��h��R�(KK��h�CL   i  7   v        �   -         �   [	     �  �  0           �t�bhhK ��h��R�(KK��h�C<        �  �        :   z  7      �            �t�bhhK ��h��R�(KK��h�C`         �         =         +  ^   =  b  *     �  �  	     �  *           �t�bhhK ��h��R�(KK��h�C,q     	  /      a  	      	         �t�bhhK ��h��R�(KK��h�C �     1  	      	         �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   6   �  :            �t�bhhK ��h��R�(KK��h�C\	  4  '  O  7         �t�bhhK ��h��R�(KK	��h�C$      ~     2     2        �t�bhhK ��h��R�(KK��h�C�   !         	         �t�bhhK ��h��R�(KK��h�C -   $   �      �   P        �t�bhhK ��h��R�(KK��h�C�  
   =     �        �t�bhhK ��h��R�(KK��h�Cd                        �     �     %   �   �     $     �        �   �        �t�bhhK ��h��R�(KK��h�C02         .   c     �  |              �t�bhhK ��h��R�(KK��h�C,O      I   ?     �  C               �t�bhhK ��h��R�(KK��h�C�  g        3        �t�bhhK ��h��R�(KK��h�C0
   K  '   �   4     5     �  6        �t�bhhK ��h��R�(KK��h�C<S     �     .   
   7     "   �     G            �t�bhhK ��h��R�(KK��h�CPW  �     =      �  m  G   W   h   �  �   :      �     �  �         �t�bhhK ��h��R�(KK��h�C0�     8              F      �        �t�bhhK ��h��R�(KK��h�C`�   �  �     �   D      V  w  9   b        J   �  �  D      4	  �  �   �        �t�bhhK ��h��R�(KK��h�C          	      	         �t�bhhK ��h��R�(KK��h�C4D      a   o  �      �      �   S   Q         �t�bhhK ��h��R�(KK��h�CD�   =     �   �  i   %   *     �  c      o      n        �t�bhhK ��h��R�(KK��h�C89      �     �     �  �      �  h   �        �t�bhhK ��h��R�(KK��h�C01   #      �     �  
   3   6   �        �t�bhhK ��h��R�(KK��h�C,         �         �  �
     �     �t�bhhK ��h��R�(KK
��h�C(�       9     ]	     �        �t�bhhK ��h��R�(KK��h�C !      �  
   :  	         �t�bhhK ��h��R�(KK��h�Cl"   �   -        z      �  +   c  ;     c     I   ^	  �  h   _	     �     <     =        �t�bhhK ��h��R�(KK��h�C<
   _      8   �        )   0   �  
   �  >        �t�bhhK ��h��R�(KK��h�C8      ?  '        j      �     �   o         �t�bhhK ��h��R�(KK��h�C ]     /     8   �        �t�bhhK ��h��R�(KK��h�C8g            �      �        �              �t�bhhK ��h��R�(KK��h�C4   �      	           `	     a	           �t�bhhK ��h��R�(KK ��h�C�
   �  [  '      �   �  q        ;        u      �         `        l      J   %  C      !  �        �t�bhhK ��h��R�(KK��h�C+              �t�bhhK ��h��R�(KK��h�C@      �  �  "      ^   |      �      �              �t�bhhK ��h��R�(KK��h�C\      P         �        �      B     T         E  �  �      �   �         �t�bhhK ��h��R�(KK��h�C4X   �   =  �     �  c      @  �  �        �t�bhhK ��h��R�(KK��h�C ]   �                    �t�bhhK ��h��R�(KK"��h�C�      6     �  "   �  �  V            d     �   �  
   �      v  �         .                        �        �t�bhhK ��h��R�(KK��h�C<T   �     ;      2   �   b	           !  �        �t�bhhK ��h��R�(KK��h�C0     �  �  �     �  B   �          �t�bhhK ��h��R�(KK��h�C0      )   b      x   "   �     �        �t�bhhK ��h��R�(KK��h�C\
   3   6   �     �      �  ?      !      �         P   <      m               �t�bhhK ��h��R�(KK��h�C<      -   b      $   �   |  "   �   c	     �        �t�bhhK ��h��R�(KK	��h�C$   A  �                     �t�bhhK ��h��R�(KK��h�C8        �  B     �     8        �        �t�bhhK ��h��R�(KK��h�Cp      �     
      �    �  �  !      �     u            �         
      �              �t�bhhK ��h��R�(KK��h�CHy      @  t         }           !     '   
   �  C        �t�bhhK ��h��R�(KK
��h�C(�        '   
   @   �   F         �t�bhhK ��h��R�(KK��h�C D  E           F  �     �t�bhhK ��h��R�(KK��h�C�  7      �t�bhhK ��h��R�(KK��h�C'  G  	      	         �t�bhhK ��h��R�(KK��h�C�     	      	         �t�bhhK ��h��R�(KK��h�C1   #       �           �t�bhhK ��h��R�(KK��h�C<   H  %     ^  8   �     `        `   �        �t�bhhK ��h��R�(KK��h�CT   "  c      �      �         �   �         ]               �        �t�bhhK ��h��R�(KK��h�CXT         P   �               d	           ;     �      �  E  �         �t�bhhK ��h��R�(KK
��h�C(F     e	     �         I        �t�bhhK ��h��R�(KK��h�C<1   #      f	     4      3   �     Y      O         �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C0   �         �   #          �        �t�bhhK ��h��R�(KK	��h�C$   A  &      �  g	  J        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C�  �            �t�bhhK ��h��R�(KK��h�CD�      w   5              B     $   �  �     ;         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C 1   #       �      D         �t�bhhK ��h��R�(KK��h�CK  >   3	  r        �t�bhhK ��h��R�(KK��h�CLB     �         �        �   L     +      &   }     o         �t�bhhK ��h��R�(KK��h�Ch	  9     �t�bhhK ��h��R�(KK��h�C0u  R   "   e   �   ?      
   �   F         �t�bhhK ��h��R�(KK��h�C,j  S  �     �      7      �        �t�bhhK ��h��R�(KK��h�C`�   �   &   �   �  �  *      $  2     �           p      �     M              �t�bhhK ��h��R�(KK��h�CHM   �      |      �   �   �     "        N  =      �        �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�CH      =         �     �   �     I     '   
   �   F         �t�bhhK ��h��R�(KK
��h�C(W   �      �  D   �  9  7         �t�bhhK ��h��R�(KK��h�C!         l      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C D      �   �   �   �        �t�bhhK ��h��R�(KK��h�C<   f   �   �  �       �      �     �   ^        �t�bhhK ��h��R�(KK��h�C      O  �  �        �t�bhhK ��h��R�(KK��h�CL   f     (      �   .  "   �  )         G        j   4         �t�bhhK ��h��R�(KK��h�CP  	      	         �t�bhhK ��h��R�(KK��h�C\           r      �t�bhhK ��h��R�(KK��h�C@   (   �         �        �   �   i	                 �t�bhhK ��h��R�(KK��h�CZ      �      Q     �t�bhhK ��h��R�(KK	��h�C$   �     9     �  R        �t�bhhK ��h��R�(KK��h�Ch�        �     �   E      )   r  �   h  Z        �      .         X   o  9   y        �t�bhhK ��h��R�(KK��h�CT      "     0      �  �        �           �  S  {      �        �t�bhhK ��h��R�(KK��h�C             v   $   "     �t�bhhK ��h��R�(KK��h�C\   �                 �  �  �               /            �     7         �t�bhhK ��h��R�(KK��h�C0$  �  "     �   .        O  �        �t�bhhK ��h��R�(KK��h�C8�   &   a      �  �        �  �      �        �t�bhhK ��h��R�(KK��h�CX,   O      �     j	  �  -   �  �       �     !  �                    �t�bhhK ��h��R�(KK��h�C@�  �  &   k	  h   s   �   g         l  �   
   �        �t�bhhK ��h��R�(KK	��h�C$M	  \     �         e  /      �t�bhhK ��h��R�(KK��h�C0l	  T  �
  �  U     V     l	           �t�bhhK ��h��R�(KK��h�Ch      f     W     �           m	           �              X  �  Y  Y  h        �t�bhhK ��h��R�(KK
��h�C(   Z  w  &      �   j  /        �t�bhhK ��h��R�(KK��h�C�  T     �t�bhhK ��h��R�(KK��h�C1   #          �t�bhhK ��h��R�(KK��h�C01   �  
   3   6   �     :             �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C8!         =        ?      
   3   6   �        �t�bhhK ��h��R�(KK��h�CD
   3   6         �   '   #   !      m                    �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�C\      �   ]   �        5   �      '        \     J   �      [     n	        �t�bhhK ��h��R�(KK
��h�C(/   (      .                     �t�bhhK ��h��R�(KK��h�CH�  \     C         �        .   ^  �     �     ]        �t�bhhK ��h��R�(KK��h�CT
   �   F   '                  �         �        �  ^     �         �t�bhhK ��h��R�(KK
��h�C(&  �   p  &   q     "            �t�bhhK ��h��R�(KK��h�C4   G   /   9   -       T     �           �t�bhhK ��h��R�(KK	��h�C$I   _  o	  �      �  �         �t�bhhK ��h��R�(KK��h�CX�               �           �      
   �  �        �  `              �t�bhhK ��h��R�(KK��h�CX!      �   ?      
         a     �        
   ,            
            �t�bhhK ��h��R�(KK��h�C0   �      �  
   ,                     �t�bhhK ��h��R�(KK��h�C0�  [   x  /      �  h   p     �         �t�bhhK ��h��R�(KK��h�C    �           b  �     �t�bhhK ��h��R�(KK��h�C8   �     �     g  �      p	     c  E        �t�bhhK ��h��R�(KK��h�C@      -   b      �     �      �      {      �        �t�bhhK ��h��R�(KK��h�C8   (   �   
   �   |        �         �        �t�bhhK ��h��R�(KK	��h�C$   �     �   �              �t�bhhK ��h��R�(KK��h�CXW  )   �        d        �  �     1   S  �  I   q	  y      r	  �         �t�bhhK ��h��R�(KK��h�CD�      (     |      s	        �  +      �     �         �t�bhhK ��h��R�(KK��h�CL�      -   r     �   %   �         Y	        6  �   �           �t�bhhK ��h��R�(KK+��h�C�         k               =      �  �        e        �      /   9   �   7      �  �        e        �      f     �  M     {  G   W         �t�bhhK ��h��R�(KK��h�CLH  C  $   0                 �           R  H              �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�Ch   .   �  �  �     $  [  �     g                    E  
   ,         "   n        �t�bhhK ��h��R�(KK��h�C0
   �  �   �   -   �  h  
   B   }         �t�bhhK ��h��R�(KK��h�CH   �   i  j                 '   !      3  �  �   �        �t�bhhK ��h��R�(KK��h�C4   t	           �   f     )      �        �t�bhhK ��h��R�(KK��h�C      �   �        �t�bhhK ��h��R�(KK��h�C�   �   k     �t�bhhK ��h��R�(KK��h�C<      =      �     �  J  E   
        �        �t�bhhK ��h��R�(KK��h�CX*      @          �  $   0  &      M      +   8   3     �     �        �t�bhhK ��h��R�(KK
��h�C(�  �   �  �          �        �t�bhhK ��h��R�(KK��h�CTl                 m     �     h  �     �   '      n  
   y        �t�bhhK ��h��R�(KK��h�CX   2      �  �  &      �   w   *        �      �   ,     L      o        �t�bhhK ��h��R�(KK��h�CL      5   �   9   �   �  &      U     �   
   �  *      �        �t�bhhK ��h��R�(KK��h�CXg   �     e  �     �  H  '        M   �      D      b  Y     a        �t�bhhK ��h��R�(KK��h�C4   �      �   �      �   ]   )   d   �         �t�bhhK ��h��R�(KK	��h�C$      �  3     p     u	     �t�bhhK ��h��R�(KK��h�C0�  �     �        ,                 �t�bhhK ��h��R�(KK��h�C8         �       ]         0      �        �t�bhhK ��h��R�(KK��h�CH      �        �       $   �     %           	        �t�bhhK ��h��R�(KK��h�CX   �  �       8  �  )   �  �   T   5            :   �     �           �t�bhhK ��h��R�(KK��h�CT   A   �  (   �   s     	     ~     D   *   D      G   �     v	        �t�bhhK ��h��R�(KK��h�Cq     r     �t�bhhK ��h��R�(KK��h�C`     t        �t�bhhK ��h��R�(KK��h�C                �t�bhhK ��h��R�(KK��h�Co  �   �   P     �t�bhhK ��h��R�(KK��h�CP9      ]  �  �              �     �  �  �  s     H   �        �t�bhhK ��h��R�(KK��h�C0T   5            �  4         �         �t�bhhK ��h��R�(KK��h�C �  ?   
   $   �           �t�bhhK ��h��R�(KK��h�C         p            �t�bhhK ��h��R�(KK��h�C,B  >   k	  h   �   �   :   d   t        �t�bhhK ��h��R�(KK��h�C<      �     s     �t�bhhK ��h��R�(KK��h�C0      �      �        (      v        �t�bhhK ��h��R�(KK	��h�C$'  
   �     �              �t�bhhK ��h��R�(KK��h�Cm      �  r      �t�bhhK ��h��R�(KK��h�C 2   �      �      �        �t�bhhK ��h��R�(KK��h�C      �        �        �t�bhhK ��h��R�(KK��h�C O        	      	         �t�bhhK ��h��R�(KK��h�C   J  C      �t�bhhK ��h��R�(KK��h�C,@     �       �  �  �   �        �t�bhhK ��h��R�(KK��h�C4]   �  '      
      }                     �t�bhhK ��h��R�(KK��h�C�  4      �      �t�bhhK ��h��R�(KK	��h�C$F	     �                    �t�bhhK ��h��R�(KK��h�C�        	         �t�bhhK ��h��R�(KK��h�C@s     O        w	  �  M     �        x	  �        �t�bhhK ��h��R�(KK��h�C    �  �   $   �           �t�bhhK ��h��R�(KK��h�CZ   t     �t�bhhK ��h��R�(KK��h�C<   0   u     �   h        �                    �t�bhhK ��h��R�(KK��h�C%   �  �     �        �t�bhhK ��h��R�(KK��h�C1   #                 �t�bhhK ��h��R�(KK��h�CX   y	  L           z	              S   Y      Q      5   y	     {	        �t�bhhK ��h��R�(KK
��h�C(z    �  �  
   �     �        �t�bhhK ��h��R�(KK��h�Cv     �t�bhhK ��h��R�(KK
��h�C(   �  �            �           �t�bhhK ��h��R�(KK��h�C<1   #      ]   
   3   6   �     /   �              �t�bhhK ��h��R�(KK��h�C<2   5   �     d  �  �  
   #  �      a  c         �t�bhhK ��h��R�(KK��h�C �        	      	         �t�bhhK ��h��R�(KK��h�C �     j  "   �           �t�bhhK ��h��R�(KK��h�C,   �  "   �      (  a     r  '     �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C`            v   �  
      :     &      U   w     �           x     �        �t�bhhK ��h��R�(KK��h�C     k  5	     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C�  ;     �t�bhhK ��h��R�(KK��h�C<   �  �   )   �  �   �   6     �  �     u         �t�bhhK ��h��R�(KK��h�Ci     �      �t�bhhK ��h��R�(KK��h�C4j  �      ?     �      y     H   �        �t�bhhK ��h��R�(KK��h�C0$   �     s           �  A            �t�bhhK ��h��R�(KK��h�C0p     )   P   n   ^   z  {  |  �        �t�bhhK ��h��R�(KK	��h�C$d   �  8     �             �t�bhhK ��h��R�(KK��h�C,*         �         �   V      �     �t�bhhK ��h��R�(KK��h�C<   �    
   \   �  L      5   [      $   �        �t�bhhK ��h��R�(KK��h�C   �   ]   ,   O      �t�bhhK ��h��R�(KK��h�C\�     �  +      u     !                 $   0        
      }          �t�bhhK ��h��R�(KK��h�CX      5   <         �     �  �                    U   $   W  N        �t�bhhK ��h��R�(KK��h�CL�     -   l                 �   f  a   ;      �  :   W         �t�bhhK ��h��R�(KK��h�Cx   �   �  �   Y     /                 �  P   <      .   G   /  i     "   C          �  O        �t�bhhK ��h��R�(KK��h�C [      �  	      	         �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�CH�  "   T  �   x      �      -  �  �  �      |	              �t�bhhK ��h��R�(KK��h�Ch�      L   G      Z     i        5   �                       1  8                 �t�bhhK ��h��R�(KK��h�C     ^  �     �t�bhhK ��h��R�(KK��h�CD        =      �         }	  /            l           �t�bhhK ��h��R�(KK	��h�C$-      �  8     U   �
        �t�bhhK ��h��R�(KK��h�C8   &   �  �   �     $   E      4      �          �t�bhhK ��h��R�(KK��h�Cq      	      	         �t�bhhK ��h��R�(KK
��h�C(      t	  ~        �   �        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C4�        a	     �  S  �   +     "        �t�bhhK ��h��R�(KK��h�C4�       d  (      �     �  �           �t�bhhK ��h��R�(KK��h�C8      '   )             �   B   �           �t�bhhK ��h��R�(KK	��h�C$q   �     ~	  �     I         �t�bhhK ��h��R�(KK��h�C�  	         �t�bhhK ��h��R�(KK	��h�C$   k        �   
   �        �t�bhhK ��h��R�(KK��h�C�   =     �t�bhhK ��h��R�(KK��h�C�  �         �t�bhhK ��h��R�(KK	��h�C$�  R      �        	         �t�bhhK ��h��R�(KK��h�CL               �        �      ;         �   �               �t�bhhK ��h��R�(KK��h�C�     v     �t�bhhK ��h��R�(KK��h�C,1   #      �  
   3   6       �        �t�bhhK ��h��R�(KK��h�C0     	  �   *      A   E      �        �t�bhhK ��h��R�(KK
��h�C(   5   -         :   Q  �        �t�bhhK ��h��R�(KK ��h�C�         �   �	     j  
               f   �   0   [      �  �               ]   �     $   �     �	        �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C     �     �t�bhhK ��h��R�(KK��h�C<      ;      �     �     �      z               �t�bhhK ��h��R�(KK��h�C,      	      	      	   �   	   /     �t�bhhK ��h��R�(KK��h�C�  	         �t�bhhK ��h��R�(KK��h�C      �     �t�bhhK ��h��R�(KK��h�C0      b      ]   
           l        �t�bhhK ��h��R�(KK��h�CP            ,               �      &  *      �  �   G   �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�Cd�  �            �           �        �      �  �  �     �	        �           �t�bhhK ��h��R�(KK��h�Cp      G           A  #  �      $   �         �	  o      5         w     v                 �t�bhhK ��h��R�(KK��h�C,5     �   
   �  �  	      	         �t�bhhK ��h��R�(KK��h�C 8         �  
            �t�bhhK ��h��R�(KK��h�C,t  �  
             �	  +         �t�bhhK ��h��R�(KK��h�C�             �t�bhhK ��h��R�(KK��h�C4#   !         ?      
   3   6   �  4         �t�bhhK ��h��R�(KK��h�C0      -   w   �  �  $   �  �           �t�bhhK ��h��R�(KK
��h�C(      w   P   !      u  *        �t�bhhK ��h��R�(KK��h�CD   
   B   �  	      	      	   K   	   �   	   �   	   /     �t�bhhK ��h��R�(KK��h�Cd   �   "         �t�bhhK ��h��R�(KK��h�C\0     -        m        x  �        U     x          �	     &        �t�bhhK ��h��R�(KK��h�C,�   �      �	     �	  A  s   o        �t�bhhK ��h��R�(KK��h�C @     /  	      	         �t�bhhK ��h��R�(KK��h�C�     �         �t�bhhK ��h��R�(KK��h�C0�  �     .      �  �                 �t�bhhK ��h��R�(KK	��h�C$      1	  -                  �t�bhhK ��h��R�(KK��h�C      
   �     �        �t�bhhK ��h��R�(KK��h�C0   X   '   R         �  �     �        �t�bhhK ��h��R�(KK��h�Cy  �     �     �t�bhhK ��h��R�(KK��h�CD      J   4        t     ~         5         4         �t�bhhK ��h��R�(KK��h�CD        �      )  �        !          !  �         �t�bhhK ��h��R�(KK
��h�C(                 �   w        �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C0�     �  �     	      	      	   K      �t�bhhK ��h��R�(KK
��h�C(   =      o  �  	      	         �t�bhhK ��h��R�(KK��h�Cx*      �  �  �            �   �        �     `               -   �        #  �       +         �t�bhhK ��h��R�(KK
��h�C(�  
        �  
   �  �        �t�bhhK ��h��R�(KK��h�C�            �t�bhhK ��h��R�(KK��h�C<         �      �   #  �   z  $   �  N   +        �t�bhhK ��h��R�(KK��h�CT-      L              l     �   S   �     Q     Q      {           �t�bhhK ��h��R�(KK��h�C@        (                      �              �t�bhhK ��h��R�(KK+��h�C�        )   p      ,      �                    |           S   X  i   ,            ^        O  �        ,   �            �     V        �t�bhhK ��h��R�(KK��h�C0�  �  �   O  7   �                    �t�bhhK ��h��R�(KK��h�C    1     �  �           �t�bhhK ��h��R�(KK��h�CL      (   �  
   $        E      4         ;                �t�bhhK ��h��R�(KK	��h�C$   %   �    '               �t�bhhK ��h��R�(KK��h�C�     4      �t�bhhK ��h��R�(KK��h�C@d  -   
     �        
  :   `   �	     A   �        �t�bhhK ��h��R�(KK��h�CX*         �         ;      �   �  &      �   )  <     `   �     W         �t�bhhK ��h��R�(KK��h�C4   &   �     t   �        �  �   n        �t�bhhK ��h��R�(KK��h�C -   �  h  H   �  �        �t�bhhK ��h��R�(KK
��h�C(�   &   8   /   a      o  ~        �t�bhhK ��h��R�(KK��h�CL      =      �  )   �     �   T   �  �  
   �  �  
   o        �t�bhhK ��h��R�(KK��h�C�      u      �t�bhhK ��h��R�(KK��h�C@     �t�bhhK ��h��R�(KK��h�C`�        I          b     &   a   �     0         p      �       O         �t�bhhK ��h��R�(KK��h�CT'  �  �     }     �         �   �  v  3        �        �         �t�bhhK ��h��R�(KK��h�C      	      	         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C@      q   �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C<#   !      X     k   '   
   3   6   2              �t�bhhK ��h��R�(KK��h�C@      J   z   "      {  &      M   �   �      �        �t�bhhK ��h��R�(KK��h�C,   W  �     ^  '   "   ~  y        �t�bhhK ��h��R�(KK��h�C   �      �t�bhhK ��h��R�(KK	��h�C$      �  �        *        �t�bhhK ��h��R�(KK��h�Ct            �  4      {               =         0  4   *         �        s   7   j   �        �t�bhhK ��h��R�(KK��h�C4a     Z           �   m  "     �	        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C  ^  �     �t�bhhK ��h��R�(KK	��h�C$   (   �   <     $   n         �t�bhhK ��h��R�(KK
��h�C(�         0                     �t�bhhK ��h��R�(KK��h�C0
      ]  T  '   �  !      �   �        �t�bhhK ��h��R�(KK��h�C,
   K  '   4     5     �  6        �t�bhhK ��h��R�(KK��h�C<         /      &   �  +      M   �      |        �t�bhhK ��h��R�(KK&��h�C��          ,                  K      �      �                 I     �     �     U     �     �        �     �         �t�bhhK ��h��R�(KK��h�C�   �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C48   /         9   -        �   �  �        �t�bhhK ��h��R�(KK��h�C	     �      �         �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�C/         �   O      �t�bhhK ��h��R�(KK��h�C\      �   |         T      5   !      |      <  R      D     .  
   y        �t�bhhK ��h��R�(KK��h�Cp          �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�C4,   �     �  }      �                    �t�bhhK ��h��R�(KK��h�CHD   >   N   9     7   �     �     �  T        4   V        �t�bhhK ��h��R�(KK	��h�C$   T  ~   �                 �t�bhhK ��h��R�(KK��h�C81   #      �      n     �     Y      O         �t�bhhK ��h��R�(KK��h�CX!      �  	      	      	   �   	   �   	   I  	   /  	   s  	   )  	   �     �t�bhhK ��h��R�(KK��h�C   �	         �t�bhhK ��h��R�(KK��h�C8�     %   )   1     �     J        �	        �t�bhhK ��h��R�(KK��h�C@1   #   
   3   6   �     �                           �t�bhhK ��h��R�(KK��h�C`      '   �   �   |        :         C  8  (  ]      �   �      �
  �   d        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C@         �   �        	     U      "   e   �         �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   6   �  "   �         �t�bhhK ��h��R�(KK��h�C`#   !      �          ^  @     �  �  (            S            Z            �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C   �     �        �t�bhhK ��h��R�(KK��h�CL      =      �	  =  ^   �   �        
   �     �     �        �t�bhhK ��h��R�(KK��h�CD      �     �     .   %   [      W   �      �           �t�bhhK ��h��R�(KK��h�C<         �     �     �t�bhhK ��h��R�(KK��h�C�      	      	         �t�bhhK ��h��R�(KK��h�C8      �    7               �              �t�bhhK ��h��R�(KK��h�C�          �t�bhhK ��h��R�(KK��h�C0b   
   $      �         P               �t�bhhK ��h��R�(KK��h�C R      M  	      	         �t�bhhK ��h��R�(KK��h�C       �  	      	         �t�bhhK ��h��R�(KK��h�C0*              &      �      L         �t�bhhK ��h��R�(KK��h�CD   8   {   �  �   �   �   &      =            G   H        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C<   `     m     
   +	        �     P   <         �t�bhhK ��h��R�(KK��h�C      �  �            �t�bhhK ��h��R�(KK��h�C@*      l  
      �  �   &      �   8        �         �t�bhhK ��h��R�(KK��h�C4   f   w     :  "   �   �  �   N   �        �t�bhhK ��h��R�(KK
��h�C(             �  j  /        �t�bhhK ��h��R�(KK��h�CH      �	  �         z  �	     h  Y     k        �	        �t�bhhK ��h��R�(KK��h�C8�     �     
   Z     y      �      �        �t�bhhK ��h��R�(KK��h�C�      �     u      �t�bhhK ��h��R�(KK��h�C4     '   s   �                 �	        �t�bhhK ��h��R�(KK��h�C0�     �  *      &   N   �     �	        �t�bhhK ��h��R�(KK��h�C`      L        �     M     �     �  ^      �         l  �	                 �t�bhhK ��h��R�(KK��h�C4�   �   7  (   �    
   _         �        �t�bhhK ��h��R�(KK��h�C0      �     @         �               �t�bhhK ��h��R�(KK��h�C82         .   �        J  x     A   8        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK
��h�C(   p  �  
   q                  �t�bhhK ��h��R�(KK��h�C�     	      	         �t�bhhK ��h��R�(KK��h�CP   d   �           �      �   =            
   �   �  :   >        �t�bhhK ��h��R�(KK��h�C0#   !      $	  (      :                  �t�bhhK ��h��R�(KK��h�C01   #   
   3   6     �   �               �t�bhhK ��h��R�(KK��h�CH]   �     2         .   (   �        /   *   %               �t�bhhK ��h��R�(KK��h�C<"   p  C  �        '   �     �  �   q   7        �t�bhhK ��h��R�(KK��h�CH                              -   R  �     �  Z        �t�bhhK ��h��R�(KK
��h�C(�   '                 �        �t�bhhK ��h��R�(KK��h�C,   �     B            �  �         �t�bhhK ��h��R�(KK��h�CD1   #      b     ,     �   p   
   3   6      �            �t�bhhK ��h��R�(KK��h�C�        	         �t�bhhK ��h��R�(KK��h�CU  �  �   �        �t�bhhK ��h��R�(KK��h�C<      �  �          �        �        �     �t�bhhK ��h��R�(KK��h�C�   p      �t�bhhK ��h��R�(KK
��h�C(�  :                          �t�bhhK ��h��R�(KK��h�CH�  
   �  �  �  �      
   +      8   /         �   O         �t�bhhK ��h��R�(KK��h�C|A     `                u      �                             �  !                    �        �t�bhhK ��h��R�(KK ��h�C�      �     /         	  i   �   7   '        =      �  :   >     �        .   N   d   �     �   S        �t�bhhK ��h��R�(KK��h�C�  �   �  	         �t�bhhK ��h��R�(KK��h�Ct   ?   3     �     �  m   -   
   3   6   �     �  m      )  ?   �   <   *   /      �      m   r      �t�bhhK ��h��R�(KK��h�CT?  (      �  j              Z           &   �           
        �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK
��h�C(      $  )      7     8        �t�bhhK ��h��R�(KK��h�C
   2     �t�bhhK ��h��R�(KK��h�C8      �         �        D        �         �t�bhhK ��h��R�(KK��h�CT         E  �            �        �     �      (     8   �         �t�bhhK ��h��R�(KK
��h�C(�        E      `     �	        �t�bhhK ��h��R�(KK��h�C0^   �   o         )   0      D  2        �t�bhhK ��h��R�(KK��h�CP�  b     �   �     I   /      �     �    }          >        �t�bhhK ��h��R�(KK��h�C4g  �        �             P   �         �t�bhhK ��h��R�(KK��h�C l  �   �        �         �t�bhhK ��h��R�(KK��h�C8     
               \   �   �              �t�bhhK ��h��R�(KK��h�C4   '               �                     �t�bhhK ��h��R�(KK��h�C8          
   i	           h  �  |        �t�bhhK ��h��R�(KK
��h�C(   .      �            �         �t�bhhK ��h��R�(KK��h�C,   �       �     �t�bhhK ��h��R�(KK��h�CP*      �          P        *     b   #  8   t  &   J           �t�bhhK ��h��R�(KK��h�C4#   !      �      ?      -   
   �   F         �t�bhhK ��h��R�(KK��h�CT   U           �     �    
   \   H            �      �   �        �t�bhhK ��h��R�(KK��h�C@         	        J   �  �            8   �         �t�bhhK ��h��R�(KK��h�C,�           �         R           �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CT�     �  �      �        �  �     �	       )   �                  �t�bhhK ��h��R�(KK��h�CT   S  &      �   �      �	       �     t      �        $   k         �t�bhhK ��h��R�(KK��h�CL            
               &      b   x   "   $   �            �t�bhhK ��h��R�(KK��h�CHB     �   �  �     �     �      �          
   A        �t�bhhK ��h��R�(KK��h�C4                     q     �           �t�bhhK ��h��R�(KK��h�C,%     �  	  �   4                 �t�bhhK ��h��R�(KK��h�C,�           N   e                �t�bhhK ��h��R�(KK��h�C@s     O        w	  �  M     �        x	  �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�      �     	         �t�bhhK ��h��R�(KK��h�C0      '   -   H   j           u         �t�bhhK ��h��R�(KK��h�CL                                   n  I   �     R         �t�bhhK ��h��R�(KK��h�C4      	     K        )     $   �        �t�bhhK ��h��R�(KK��h�C`�   �  A   T     �  s  C         �  �   �        �      �         �          �t�bhhK ��h��R�(KK��h�C,k     �  "   L     ~     p          �t�bhhK ��h��R�(KK��h�C\�     �	  �                R  "  h                                   �t�bhhK ��h��R�(KK��h�C1   #       �         �t�bhhK ��h��R�(KK��h�CP   e   '   H   �  j     �     A   j  ^        -      �  �        �t�bhhK ��h��R�(KK	��h�C$U   �  �	     �     �        �t�bhhK ��h��R�(KK��h�C1   #       +     �t�bhhK ��h��R�(KK��h�C,           �  *        �         �t�bhhK ��h��R�(KK#��h�C�         O         Y      Q      Q     Q      
  Q      x     J   4              �     o      5      7  4         �t�bhhK ��h��R�(KK��h�C,!      �     	      	      	   K      �t�bhhK ��h��R�(KK��h�C]      �        �t�bhhK ��h��R�(KK��h�CT   f   �         �  0      �     �     4         
   _      �        �t�bhhK ��h��R�(KK��h�C!            �t�bhhK ��h��R�(KK��h�C\
   �          F   '      H     %        B  �      *         �   �         �t�bhhK ��h��R�(KK��h�CL�   �     8  >   �         �  	  C  �     0   {      p         �t�bhhK ��h��R�(KK
��h�C(  �     �                    �t�bhhK ��h��R�(KK1��h�C�*      V  �   �	        0   [      <      $      "   K     i        
   C     �                    !  h         m  �            �              �   G   �	        �t�bhhK ��h��R�(KK��h�CL�  �      N         *   2      .      :      Q         S         �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK	��h�C$   �    '   -   �            �t�bhhK ��h��R�(KK��h�C0      -   P   �                     �t�bhhK ��h��R�(KK��h�Cl*         E  c          P   +      �  �   e  h   c  �     "      �     "              �t�bhhK ��h��R�(KK��h�C80     ;      0   �     9         9   �         �t�bhhK ��h��R�(KK��h�CD!      �   �  ?      
   }  n     e      n     @         �t�bhhK ��h��R�(KK��h�C      �     �t�bhhK ��h��R�(KK*��h�C�   �  �  �                  �         �  N      <   *   2   �         {         �     S     {  �        c  
   �      2      E  �         �t�bhhK ��h��R�(KK��h�C0      �   2      �     :  �   7         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C,�     �   �  �   7        �         �t�bhhK ��h��R�(KK��h�C �        	      	         �t�bhhK ��h��R�(KK��h�C,�     �     ,            ^        �t�bhhK ��h��R�(KK��h�CT�            ;      )     �     �         �     �  �      k        �t�bhhK ��h��R�(KK��h�C,4      m        J	     I   q        �t�bhhK ��h��R�(KK��h�C0      �  	      	      	   K   	   U     �t�bhhK ��h��R�(KK��h�C4�     �      C  �     �                �t�bhhK ��h��R�(KK��h�C<   �  R   �  -               �   �  �   �        �t�bhhK ��h��R�(KK��h�C<�     7  �  �        M   �      �     V        �t�bhhK ��h��R�(KK��h�C<$        $   �     a  �                       �t�bhhK ��h��R�(KK��h�C&	     m     �t�bhhK ��h��R�(KK��h�C0         �  `     �     I           �t�bhhK ��h��R�(KK��h�C<           x      <   -               �        �t�bhhK ��h��R�(KK��h�C!            �t�bhhK ��h��R�(KK��h�C�	  	         �t�bhhK ��h��R�(KK��h�C             �           �t�bhhK ��h��R�(KK��h�C8      �     �     
   A        
   [        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK%��h�C�               t           v     �   )         �      ~            �  �        �  C   w         t                    �t�bhhK ��h��R�(KK��h�C1   #   
     �          �t�bhhK ��h��R�(KK��h�C,      �                 �        �t�bhhK ��h��R�(KK��h�CT�   �      �	     �	     A  s      g   �        J   �     �  7         �t�bhhK ��h��R�(KK��h�C\,   �      �         %   �        �     �      -                  }         �t�bhhK ��h��R�(KK��h�CL      �  
      4           (      �  :   2     �           �t�bhhK ��h��R�(KK��h�Ch   �           �      �	  
   C   w                                   �	           �t�bhhK ��h��R�(KK��h�C0
   �	  6   '      �  �   q   �  �         �t�bhhK ��h��R�(KK��h�C       �  �  �  �        �t�bhhK ��h��R�(KK��h�C,   2     N         m        .      �t�bhhK ��h��R�(KK��h�C0M      +   �          �     �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   6       g   O        �t�bhhK ��h��R�(KK��h�C,   �      ,  ~  l         �  �      �t�bhhK ��h��R�(KK��h�C8}  +            c  ,            `   �        �t�bhhK ��h��R�(KK��h�C,�      2   0   <         0   /         �t�bhhK ��h��R�(KK��h�C`      5   �  [   �  
   _      �  &      =      �   
        9   E      g        �t�bhhK ��h��R�(KK��h�C0:  "      �     �	           �        �t�bhhK ��h��R�(KK��h�C@                 @         ~  y     e            �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C,T   r  �  �  
   �     �           �t�bhhK ��h��R�(KK��h�C`            s  4      �     _               �        �  @  {  �  �        �t�bhhK ��h��R�(KK��h�C<      E     �t�bhhK ��h��R�(KK	��h�C$�         	      	   �     �t�bhhK ��h��R�(KK��h�CL         E     �               0      4         P   {         �t�bhhK ��h��R�(KK��h�C8`        .   �     �  q                   �t�bhhK ��h��R�(KK��h�C`      �  /      �             +   
   �   �         U                        �t�bhhK ��h��R�(KK��h�Cx�     �  	      	      	   K   	   �   	     	   �  	   U  	   �  	   �   	   �  	   �  	   �  	        �t�bhhK ��h��R�(KK��h�C4   �              �  
   �              �t�bhhK ��h��R�(KK��h�C1   #       9     �t�bhhK ��h��R�(KK��h�C      �     �t�bhhK ��h��R�(KK��h�C`      5   �	     [      $   �                  �  =        �	                 �t�bhhK ��h��R�(KK ��h�C�      �  r  +         
   �   �   _         a   ;      �   )               �	        4   
   _      {         �t�bhhK ��h��R�(KK��h�CH      (   4            `      =      �   
   _      �        �t�bhhK ��h��R�(KK ��h�C�              �   f     �           g                  ;      P   �           G   W      �           �t�bhhK ��h��R�(KK��h�C [         	      	         �t�bhhK ��h��R�(KK��h�C0"        2      .   �                  �t�bhhK ��h��R�(KK	��h�C$;           	      	         �t�bhhK ��h��R�(KK��h�CT�  �   �	  �     �        /   9     7      )      %      ~   �         �t�bhhK ��h��R�(KK��h�C@v                 t  
   �   :        �   "        �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C0           K  G   %  D   ~   �        �t�bhhK ��h��R�(KK��h�C8q   �  �           �        A     �	        �t�bhhK ��h��R�(KK��h�C`   Q                 '      �              V         �   B              �t�bhhK ��h��R�(KK��h�C8G                            �  �         �t�bhhK ��h��R�(KK!��h�C�  {   �     {      �     K           �         �  �  �            [      d      Q     �	     �            �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�CD!      �      �  R   ?      
   3   6   �     �   f        �t�bhhK ��h��R�(KK��h�CP        �             �         �         
   y     �        �t�bhhK ��h��R�(KK��h�C@   @   '   )   H   �     V   %   �      G  
            �t�bhhK ��h��R�(KK��h�C8�	           l      (   X  �	  	      	         �t�bhhK ��h��R�(KK��h�CH
      ]  T  �  '     �   [      �   �      �	     �	        �t�bhhK ��h��R�(KK��h�C0      '               /      �         �t�bhhK ��h��R�(KK��h�C8%      �     I      J   6  C      c  ,         �t�bhhK ��h��R�(KK��h�CD*      J   �   L      �  &      �   X  �     $   k         �t�bhhK ��h��R�(KK��h�C8     �     �t�bhhK ��h��R�(KK��h�CPy      @  t         }                      �  
   �  C        �t�bhhK ��h��R�(KK	��h�C$�	     �	                    �t�bhhK ��h��R�(KK��h�C�      R              �t�bhhK ��h��R�(KK��h�CA     �     �t�bhhK ��h��R�(KK��h�C4�        �    7                        �t�bhhK ��h��R�(KK��h�C,M      +      �     �     �        �t�bhhK ��h��R�(KK	��h�C$      E  `     p  �         �t�bhhK ��h��R�(KK��h�C   �         �t�bhhK ��h��R�(KK��h�C	         �t�bhhK ��h��R�(KK��h�CL   D      s   �     �     �	        S   �            �        �t�bhhK ��h��R�(KK��h�C X     �  
   ]  L         �t�bhhK ��h��R�(KK��h�C   	  	      	         �t�bhhK ��h��R�(KK��h�C   J  C      
     �t�bhhK ��h��R�(KK��h�C,�  �      [         	      	         �t�bhhK ��h��R�(KK��h�C4        I   Y      ?     t              �t�bhhK ��h��R�(KK
��h�C(!      p     �  	      	         �t�bhhK ��h��R�(KK��h�C<      0   �   )               G                �t�bhhK ��h��R�(KK��h�C Y  >   �   w   �          �t�bhhK ��h��R�(KK%��h�C�   D   �  �       ,               2     �     �	  �  �      �   :       �         �   �        �	  �                 �t�bhhK ��h��R�(KK��h�CH   ,      	   K   	   �   	   I  	   U  	   /  	   �  	   �     �t�bhhK ��h��R�(KK��h�C<      �   �           [  �  B   [              �t�bhhK ��h��R�(KK
��h�C(      �  s   7   �   j   �        �t�bhhK ��h��R�(KK��h�CT
   3   6      ?      !      #        �         �           �         �t�bhhK ��h��R�(KK��h�CT�        �  h      �  p  :   $   �   x  �  �  �   y      5            �t�bhhK ��h��R�(KK��h�C<      �     m  �  �           �     �        �t�bhhK ��h��R�(KK
��h�C(      -        6     _        �t�bhhK ��h��R�(KK��h�C08   /      
      �     �               �t�bhhK ��h��R�(KK��h�CH!        U          )   ;      �  �      (	             �t�bhhK ��h��R�(KK��h�CD         B           �t�bhhK ��h��R�(KK��h�Ct   d   �        ,   �         �  �      �         6  O        D   0     p                     �t�bhhK ��h��R�(KK��h�C           �	  	         �t�bhhK ��h��R�(KK��h�CZ        �t�bhhK ��h��R�(KK��h�C,1   #   
   3   6     �               �t�bhhK ��h��R�(KK��h�C       0   �  �           �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�	        �t�bhhK ��h��R�(KK��h�CL         E  �               0      �  4         P   {         �t�bhhK ��h��R�(KK	��h�C$   �      B  "   �           �t�bhhK ��h��R�(KK��h�CD   C    �      ]  '        �     _  g   d   t        �t�bhhK ��h��R�(KK��h�C    �	     &      �        �t�bhhK ��h��R�(KK��h�C,1   #   
   3   6           ?        �t�bhhK ��h��R�(KK	��h�C$   @      M  '               �t�bhhK ��h��R�(KK��h�C  M     �t�bhhK ��h��R�(KK��h�Ct         
  4   
   _      �     �     (   ;      k                  ,       $   �   x        �t�bhhK ��h��R�(KK��h�CL      b   x      �              �   L   G   �                 �t�bhhK ��h��R�(KK��h�CH      '         V                 `   3  T             �t�bhhK ��h��R�(KK��h�C@      J   �     �        &      z   ,               �t�b�
      hhK ��h��R�(KK��h�C\   (   �      r      �t�bhhK ��h��R�(KK��h�C,1   #       �  Y  �      Z          �t�bhhK ��h��R�(KK��h�Cd                          �     �     d        .        �             �t�bhhK ��h��R�(KK��h�CX            .   N         o        �   S   �                         �t�bhhK ��h��R�(KK��h�C       �      �   L         �t�bhhK ��h��R�(KK��h�C\   �	           �  �        3  �   �   �	        Q   V         E  �         �t�bhhK ��h��R�(KK��h�C4
   �             $   �  �  �           �t�bhhK ��h��R�(KK��h�C �  �     �  �     ?     �t�bhhK ��h��R�(KK��h�C0      �     �t�bhhK ��h��R�(KK��h�CP            ;      %   �              �   L   
      �   D        �t�bhhK ��h��R�(KK��h�C  	         �t�bhhK ��h��R�(KK��h�C �     s        �        �t�bhhK ��h��R�(KK��h�C   �         �t�bhhK ��h��R�(KK��h�C\   |  �      o   r      �t�bhhK ��h��R�(KK��h�C@   H  �   +      �  �   
   $        (      4         �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   �       u        �t�bhhK ��h��R�(KK��h�C0        �      $   8  �   s   7         �t�bhhK ��h��R�(KK��h�C,              �     ,   K        �t�bhhK ��h��R�(KK��h�C8      �      �  �      �        P   +        �t�bhhK ��h��R�(KK��h�C4   �   J      �   �     �  �              �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK#��h�C��	                 {                 �     `     V   %        C      �   �           �  �  �     �           �t�bhhK ��h��R�(KK��h�C8   �  C         L               B   #        �t�bhhK ��h��R�(KK��h�C �      ,   �   "   �   n     �t�bhhK ��h��R�(KK	��h�C$�     ^     �     �         �t�bhhK ��h��R�(KK��h�C   �           �t�bhhK ��h��R�(KK��h�C�  �   �        �     �t�bhhK ��h��R�(KK��h�CP   �     D      �   (   [      .      �      k  y   2   t  v        �t�bhhK ��h��R�(KK��h�CX      �      �   G     )           a      �       4     
           �t�bhhK ��h��R�(KK��h�C!        	         �t�bhhK ��h��R�(KK��h�C          5     V  �      �t�bhhK ��h��R�(KK��h�C   �     	         �t�bhhK ��h��R�(KK��h�C0�   l     
   �     �   �  
            �t�bhhK ��h��R�(KK��h�CpK        �      �            �   �        �     �            d  $   N     �              �t�bhhK ��h��R�(KK��h�C,      "     n   
      �            �t�bhhK ��h��R�(KK
��h�C(+  �             G   �
        �t�bhhK ��h��R�(KK��h�C,B    �         �       �        �t�bhhK ��h��R�(KK��h�C<$   K     �              W     +      �   �     �t�bhhK ��h��R�(KK��h�C`           �            �
     f   �   =         �  G   �     �               �t�bhhK ��h��R�(KK��h�C,      J         )   �    �        �t�bhhK ��h��R�(KK��h�C                    �t�bhhK ��h��R�(KK��h�CH�   �       &   [     �      �  �     0  `     �        �t�bhhK ��h��R�(KK��h�CX   �   �      6  C   �   
   �   �      �     B  �     !  �              �t�bhhK ��h��R�(KK��h�CL�	  �     D     ;      M      �      `   b           `        �t�bhhK ��h��R�(KK��h�C�  �      �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�CH         �	     c  X     $   �	           0      �        �t�bhhK ��h��R�(KK��h�C8   �     �                 "              �t�bhhK ��h��R�(KK��h�C,�    �  
   �        �   L         �t�bhhK ��h��R�(KK��h�C�  \     �t�bhhK ��h��R�(KK
��h�C(!      n        	      	         �t�bhhK ��h��R�(KK��h�C�  7      �t�bhhK ��h��R�(KK��h�C,   4  '   �   s         #  �        �t�bhhK ��h��R�(KK��h�CH      �     *      w   $        �   �     �    w         �t�bhhK ��h��R�(KK��h�C �       I   _  �  �     �t�bhhK ��h��R�(KK��h�C0*   '    �       �                  �t�bhhK ��h��R�(KK��h�CLl      �            E     M   �      �	  �	  "   �   �   k        �t�bhhK ��h��R�(KK��h�C`      �     E     +        p              P                 J  E         �t�bhhK ��h��R�(KK��h�C   @   '   �   �	        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C<a  �      �     �     �           �	  �  �     �t�bhhK ��h��R�(KK��h�CT      �   L  v  7  �      b     �        N   ^  T   2     �         �t�bhhK ��h��R�(KK��h�C<)   ^     e  C         �  �        �           �t�bhhK ��h��R�(KK��h�C8   &      S   F  �     v        �  �        �t�bhhK ��h��R�(KK��h�C`   �        c      =  �                       M   c      
   w  j            �t�bhhK ��h��R�(KK��h�Cx     �     �t�bhhK ��h��R�(KK��h�C4   f   e    �  
   �   S   }   i   ,         �t�bhhK ��h��R�(KK��h�CP   �      �      �     �      �  L   :                 �        �t�bhhK ��h��R�(KK
��h�C(�      %         ,               �t�bhhK ��h��R�(KK��h�C@      0   U           7      �  9   A  �   7         �t�bhhK ��h��R�(KK��h�C`�        �  �  ,            �        �	     }         �  5   [      �         �t�bhhK ��h��R�(KK
��h�C(   %     m  N   �      �          �t�bhhK ��h��R�(KK��h�C8�	  
         $   �     $   �     �           �t�bhhK ��h��R�(KK��h�C             �t�bhhK ��h��R�(KK��h�CDV         b      x      0   [      �	     ~     /         �t�bhhK ��h��R�(KK��h�CL�	  4     t      �  �  4        &        �   S   �  �        �t�bhhK ��h��R�(KK	��h�C$^   �   �	     �     �        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CP   P     2   
      I    �      e  z    i   
      �          �t�bhhK ��h��R�(KK��h�CP}       Q         O               f   �   �         j   4         �t�bhhK ��h��R�(KK��h�CL      ,     (           �   5         o                  �t�bhhK ��h��R�(KK��h�Cl   �	  �   l     �      ;        %   R   �      �   5   
   �   �     %   h  k     <        �t�bhhK ��h��R�(KK��h�C0
   �  �   Q     
   H   �     4        �t�bhhK ��h��R�(KK��h�C�      �     �t�bhhK ��h��R�(KK��h�CX      J   6     �	     X         P        �	          �     :        �t�bhhK ��h��R�(KK��h�C�
     �t�bhhK ��h��R�(KK��h�CL
   Z     o           R              �     �              �t�bhhK ��h��R�(KK��h�CD      &   �  +         ?      y  !   
   3   6            �t�bhhK ��h��R�(KK��h�C0   9   �       �      �   s   7         �t�bhhK ��h��R�(KK��h�C<y         0   �  >      2           �            �t�bhhK ��h��R�(KK��h�C,   X   �        p         �	        �t�bhhK ��h��R�(KK��h�C4               J   �           :   M     �t�bhhK ��h��R�(KK��h�C8   X     �  
   ,            K               �t�bhhK ��h��R�(KK��h�C41   #         �   �   
   3   6      p         �t�bhhK ��h��R�(KK��h�C`         O         Y      Q      �     x     5      7  4      L              �t�bhhK ��h��R�(KK��h�C8   5   �  *  �   8      *      �               �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK	��h�C$b         
   $   �            �t�bhhK ��h��R�(KK��h�C4�	     i        h                        �t�bhhK ��h��R�(KK��h�CH      ~      ,     �
     z     �     �                �t�bhhK ��h��R�(KK��h�C48   �     �                  �            �t�bhhK ��h��R�(KK��h�ChS     �        Y      O      �	        t        Y      O      �     �               �t�bhhK ��h��R�(KK��h�Cd*      m     �   o         R     �     ;  $   o  9      L   T      �  $   �        �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�Cxl         �     �     %   �  !  j   <         .   �     l      �        0   M   �      '          �t�bhhK ��h��R�(KK��h�C0�  !         ?      ^   �     �         �t�bhhK ��h��R�(KK��h�C<      G     �t�bhhK ��h��R�(KK��h�CP   f   w        K     ~      D   =      (           "   W         �t�bhhK ��h��R�(KK��h�C 4         	      	         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C1   #       �      �t�bhhK ��h��R�(KK��h�C�      	      	         �t�bhhK ��h��R�(KK��h�C 1   #       F     �        �t�bhhK ��h��R�(KK��h�C4
   2     �           $  �   "  �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�Cm     �  m     �t�bhhK ��h��R�(KK��h�Cp      :          �t�bhhK ��h��R�(KK��h�C<
   3   6   {     �  ?      !                    �t�bhhK ��h��R�(KK��h�C0B               �   
   $   �        �t�bhhK ��h��R�(KK��h�C   X   '   �   �        �t�bhhK ��h��R�(KK��h�C      �        �t�bhhK ��h��R�(KK	��h�C$�        N                  �t�bhhK ��h��R�(KK��h�CD      �  H     �        E               8   4         �t�bhhK ��h��R�(KK��h�CT   �	  �  3  *            S        �	        t        Y      O      �t�bhhK ��h��R�(KK	��h�C$#   !                         �t�bhhK ��h��R�(KK��h�C@r  )     s                  �            �         �t�bhhK ��h��R�(KK��h�C8
   �  '   �   �   ^     �   Q                 �t�bhhK ��h��R�(KK��h�C8�        �     )  C      �	     \  L         �t�bhhK ��h��R�(KK��h�C�  �     ?          �t�bhhK ��h��R�(KK��h�C@�       �      �     �     �  �      �     �     �t�bhhK ��h��R�(KK��h�C4         {      &   �  /        �         �t�bhhK ��h��R�(KK��h�C�     	      	         �t�bhhK ��h��R�(KK��h�C4�         t      �     \  L               �t�bhhK ��h��R�(KK��h�CPX   �   h  B   R      �     �   �      0   �      �     �  �         �t�bhhK ��h��R�(KK��h�C �      )     
            �t�bhhK ��h��R�(KK��h�C\
   3   6      �      4   ?      !      #        �         (      *  �         �t�bhhK ��h��R�(KK��h�C D  E           F  M     �t�bhhK ��h��R�(KK��h�CL      b   x      �      -  �	     �  "   $   �   |      �        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C<  R      |        �t�bhhK ��h��R�(KK��h�C�     �	     �t�bhhK ��h��R�(KK��h�C+     �t�bhhK ��h��R�(KK��h�C<�  �   +            !  �     �  �     �         �t�bhhK ��h��R�(KK
��h�C(      -   �	  `   �  
   &        �t�bhhK ��h��R�(KK��h�C �     �  	      	         �t�bhhK ��h��R�(KK��h�CP[      <      `     �  �                  %   �      �            �t�bhhK ��h��R�(KK��h�CP      ;      *  �           �        �     0         ]         �t�bhhK ��h��R�(KK��h�CH      0   �        
        �	     {      �      x        �t�bhhK ��h��R�(KK��h�C0�     �  X     "   >  ;      �        �t�bhhK ��h��R�(KK��h�CP   f   ?     D   ;      W    �  �   �        �  �     '        �t�bhhK ��h��R�(KK��h�C,      -   �     �      �  �         �t�bhhK ��h��R�(KK
��h�C(      L              �        �t�bhhK ��h��R�(KK��h�CD   v  )                        (   :   t               �t�bhhK ��h��R�(KK
��h�C([  (      �     #     C         �t�bhhK ��h��R�(KK��h�Cq     r     �t�bhhK ��h��R�(KK��h�C�      �     �t�bhhK ��h��R�(KK��h�C�     E      �        �t�bhhK ��h��R�(KK��h�Ch               "      �      ,     �        E   
   �     �   �      
   �  �        �t�bhhK ��h��R�(KK��h�C�  :   Y      �     �t�bhhK ��h��R�(KK��h�C`�	  }     �   @                              )   �     /     �     4        �t�bhhK ��h��R�(KK��h�C�            �t�bhhK ��h��R�(KK��h�C<         �     s                 k            �t�bhhK ��h��R�(KK
��h�C(|         	      	      	   K      �t�bhhK ��h��R�(KK��h�C0   8   /   \  &      U     "   >        �t�bhhK ��h��R�(KK��h�CH   %   .          M   �   �     �   y   2   (      n         �t�bhhK ��h��R�(KK��h�Cp      =      �  h   p     8   /   =  ^   �                 
   �   F      E      �           �t�bhhK ��h��R�(KK��h�Cl   �      @      �     t      ~     �     W      $           ~     �     =           �t�bhhK ��h��R�(KK��h�C�  �         �t�bhhK ��h��R�(KK
��h�C(�   �   )   �  q     �  /         �t�bhhK ��h��R�(KK��h�CH|      �      W      <  C  $   ;            @  9   �        �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�CH%         �     7      P   C              �   �   �        �t�bhhK ��h��R�(KK��h�CD�     �   �     -                 �      �   �	        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C�     1  	         �t�bhhK ��h��R�(KK��h�CL  �        �t�bhhK ��h��R�(KK��h�Cx            �     J  C      !  *      d  �       +      .     $         `   �     �  1        �t�bhhK ��h��R�(KK��h�C!      �     �t�bhhK ��h��R�(KK��h�Cq      	      	         �t�bhhK ��h��R�(KK��h�C�     %           �t�bhhK ��h��R�(KK��h�CT�        .      ;      �   �       J  S                �	        �t�bhhK ��h��R�(KK��h�C!                  �t�bhhK ��h��R�(KK��h�C4   %   h  �  ?      !   
   X   �   F         �t�bhhK ��h��R�(KK��h�C �   [  �       &         �t�bhhK ��h��R�(KK	��h�C$6  �                       �t�bhhK ��h��R�(KK��h�C0/     )     ^   &  
        V        �t�bhhK ��h��R�(KK��h�C�  �            �t�bhhK ��h��R�(KK��h�CX-      .      S                 �                G     6  +         �t�bhhK ��h��R�(KK��h�Cz  +      f  �     �t�bhhK ��h��R�(KK��h�CD^   �      '	     2      .   P      �         ,   �         �t�bhhK ��h��R�(KK��h�C  -   '  �        �t�bhhK ��h��R�(KK��h�C          	      	         �t�bhhK ��h��R�(KK��h�Ch�  R      �  �            �        b           0   0     {  Q  �  :     k        �t�bhhK ��h��R�(KK��h�C41   #   
   3   6   Y      O      (  O         �t�bhhK ��h��R�(KK��h�C)         �t�bhhK ��h��R�(KK��h�C �   �                   �t�bhhK ��h��R�(KK��h�C 
   .  c    �   �        �t�bhhK ��h��R�(KK��h�C81   #           �  
   3   6   1     	        �t�bhhK ��h��R�(KK��h�C4�   �   �  �      �             �         �t�bhhK ��h��R�(KK��h�C      	      	         �t�bhhK ��h��R�(KK��h�C�   k  �     �t�bhhK ��h��R�(KK��h�Cd   �      $     �  �   Y  +      �  +      �            U   �   i     i           �t�bhhK ��h��R�(KK��h�C
       $   |        �t�bhhK ��h��R�(KK��h�C,   �     �  �                    �t�bhhK ��h��R�(KK��h�C82   �        �      �  9   �  
      *        �t�bhhK ��h��R�(KK��h�C<            �   2               t  �   �        �t�bhhK ��h��R�(KK��h�C@1   #         P   �         
   T  )  ?   �   �   r      �t�bhhK ��h��R�(KK
��h�C(!         	      	   �   	   �      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CD        I   ,   O      �    7   ;      �  "   �        �t�bhhK ��h��R�(KK��h�C`  (  
   ,         �t�bhhK ��h��R�(KK	��h�C$               y   �	        �t�bhhK ��h��R�(KK��h�Ca        	         �t�bhhK ��h��R�(KK	��h�C$      �	  +  �  
   y        �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�Cd9   ,     0  -     �      C      �     v	     �      -     0          �         �t�bhhK ��h��R�(KK��h�CP      J   =      o  �   >      D  ,                  ,            �t�bhhK ��h��R�(KK��h�C4!      �      	   I  	   U  	   /  	   s     �t�bhhK ��h��R�(KK��h�CH      �   �  �  �  &      �  )  �     �        Z        �t�bhhK ��h��R�(KK	��h�C$$  
   2     �              �t�bhhK ��h��R�(KK	��h�C$#  a  �   *            r      �t�bhhK ��h��R�(KK��h�C<1   #         r  '     �  
   3   F   3           �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C<7      �  e           �  7   �  �             �t�bhhK ��h��R�(KK	��h�C$   .      d   ]  U            �t�bhhK ��h��R�(KK��h�C`   /   (   o  �   -      �  �              (   �      �   �   Q      �   8        �t�bhhK ��h��R�(KK��h�CD�     s        �     �            .                 �t�bhhK ��h��R�(KK��h�CD     �  
   B     P     �            b              �t�bhhK ��h��R�(KK
��h�C(      0   /  
   ,               �t�bhhK ��h��R�(KK��h�C       �         �	        �t�bhhK ��h��R�(KK��h�C0�  
   �  }      �         �           �t�bhhK ��h��R�(KK��h�C4�	  
         k  �                       �t�bhhK ��h��R�(KK��h�C44        �        %   �                �t�bhhK ��h��R�(KK
��h�C(�  �     �     5  
            �t�bhhK ��h��R�(KK��h�CD         �  �          c   �      �   �               �t�bhhK ��h��R�(KK��h�C          �     �        �t�bhhK ��h��R�(KK��h�CP#   !      d        B     '   
   3   6   �             �        �t�bhhK ��h��R�(KK��h�CH      �     Y     7   &      �  a      �     /  �        �t�bhhK ��h��R�(KK��h�CHj   �   (         �   �  <     )         �       w         �t�bhhK ��h��R�(KK��h�C,�  �	     �   �  �     �  P        �t�bhhK ��h��R�(KK��h�C0H   �  �   )   p      �      B           �t�bhhK ��h��R�(KK��h�C/         �  O      �t�bhhK ��h��R�(KK��h�CD      '      �        0        9   �	                 �t�bhhK ��h��R�(KK��h�C,         9   N     �      7   v     �t�bhhK ��h��R�(KK��h�C2     �
     �t�bhhK ��h��R�(KK��h�C    �  (      
   Z        �t�bhhK ��h��R�(KK
��h�C(�        �           �         �t�bhhK ��h��R�(KK��h�C@   �        �   �  R   )      e         $   k         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C      �	     ?        �t�bhhK ��h��R�(KK
��h�C(      �   �                    �t�bhhK ��h��R�(KK��h�CL         Y        $   E               .   
   _               �t�bhhK ��h��R�(KK��h�C�     �	     e         �t�bhhK ��h��R�(KK��h�C   �	        �t�bhhK ��h��R�(KK��h�Cd^            0               !  +         g   {      _           �  �   o         �t�bhhK ��h��R�(KK��h�C,   �   
      �     �      �        �t�bhhK ��h��R�(KK��h�C�	     6     �t�bhhK ��h��R�(KK
��h�C(      �	  $   �     &           �t�bhhK ��h��R�(KK��h�CD   -            1        $   V  �      �  C   w         �t�bhhK ��h��R�(KK��h�C<I      �         �	  &   �   �      E      ,        �t�bhhK ��h��R�(KK��h�C<'        0   *                       ~        �t�bhhK ��h��R�(KK��h�C@      �     �   "     0      �  
      �   �        �t�bhhK ��h��R�(KK��h�C,   �    
     Q                  �t�bhhK ��h��R�(KK��h�C4�     �      7     h     �  
            �t�bhhK ��h��R�(KK��h�C@�        h              V     +   �        h     �t�bhhK ��h��R�(KK��h�C,  �   �     �     �t�bhhK ��h��R�(KK��h�CP�	  2  �      $   �     �  �  *   �   �      A     �  Y  �         �t�bhhK ��h��R�(KK��h�C 
      I  '               �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�CD�  �  $         �        0             H  �         �t�bhhK ��h��R�(KK��h�C\      /   9   q  7   \       d            H  '        M   �      D         �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�Cl)      0     
  p      v        �  *   x  ]        H   �   �   �      �  C   #   p         �t�bhhK ��h��R�(KK��h�C      �           �t�bhhK ��h��R�(KK
��h�C(8  �  ;  S  y      |  �        �t�bhhK ��h��R�(KK��h�CX      0      �           �                 �     \     (  �         �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CH      B            �     n  I   c  O  h         �        �t�bhhK ��h��R�(KK��h�C   (      k  �	     �t�bhhK ��h��R�(KK��h�C<      �  c   8   �        o  �  
      �        �t�bhhK ��h��R�(KK��h�C01   #   
   3   6   �     �     �        �t�bhhK ��h��R�(KK��h�C`!      �        	      	      	   �   	   �   	   I  	   /  	   s  	   )  	   �     �t�bhhK ��h��R�(KK��h�C 1   #          }     o      �t�bhhK ��h��R�(KK��h�Cl�  �     �        %  �      �   �	           '      �  �     $   n   O     d  �        �t�bhhK ��h��R�(KK��h�CD   �  <         �  �            B   �  �	     4        �t�bhhK ��h��R�(KK��h�C<!           8  ?      
   3   6                 �t�bhhK ��h��R�(KK	��h�C$�           g              �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C4{      �  +   �  ;      �  �              �t�bhhK ��h��R�(KK��h�CT            3                                              �t�bhhK ��h��R�(KK��h�C<$   ;      �     @        0     
   G   W         �t�bhhK ��h��R�(KK��h�C\     |            9  
   ,      �	  
         �	  
         4  
   K         �t�bhhK ��h��R�(KK��h�C0H   �     -  5  
      R              �t�bhhK ��h��R�(KK��h�CHW  �     )  +   -   �   g   �      X        �              �t�bhhK ��h��R�(KK��h�C,6     7  "     N  �     �         �t�bhhK ��h��R�(KK��h�C8W      )   �  �         �                     �t�bhhK ��h��R�(KK��h�CH   �  {  
   _            �  8  �        �
     �        �t�bhhK ��h��R�(KK��h�C�	           �t�bhhK ��h��R�(KK��h�Ch   3  h      �   L     x     [	     v  �   �   
      ]  �        .      �  p        �t�bhhK ��h��R�(KK��h�Cp        /      9   �   7         d   K  0   �        :     *   �      �   �  D      V        �t�bhhK ��h��R�(KK��h�C@#   !                 �     �       �            �t�bhhK ��h��R�(KK	��h�C$�   p         	      	         �t�bhhK ��h��R�(KK��h�CD         k      l                 ,  %   �            �t�bhhK ��h��R�(KK��h�CP*            k         ;      �   �  �  R   �     .   �   �        �t�bhhK ��h��R�(KK��h�CxY         	      	      	   �   	   �   	   I  	   /  	   s  	   )  	   �  	   �	  	   �  	   �  	   �     �t�bhhK ��h��R�(KK$��h�C�      >   $  �      [     �         ,                    '   �   S   }      �        D             �               �t�bhhK ��h��R�(KK��h�C0   @   '      �	          �  �        �t�bhhK ��h��R�(KK��h�CH                 e  b  2            #     �   2         �t�bhhK ��h��R�(KK	��h�C$
   �	  �  ;  )   A   |        �t�bhhK ��h��R�(KK��h�C4     �   �      ,              �        �t�bhhK ��h��R�(KK��h�C  �      �t�bhhK ��h��R�(KK��h�C4�	     ;      �     �   �  T   �	  �        �t�bhhK ��h��R�(KK��h�C �        	      	         �t�bhhK ��h��R�(KK��h�CH�  �    
        %   9  �     O    2   �	  
   c        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C        �t�bhhK ��h��R�(KK��h�C   �	     �t�bhhK ��h��R�(KK��h�CZ             �t�bhhK ��h��R�(KK
��h�C(  �     �           ,         �t�bhhK ��h��R�(KK��h�CD   '   )   f   A   �   V         =      �   �   q   7        �t�bhhK ��h��R�(KK��h�C1   #       �        �t�bhhK ��h��R�(KK��h�C`   �     �
        8     �
     9  V      {  $   �     $   :     �  �        �t�bhhK ��h��R�(KK��h�C8         �     ,   K  �            Y        �t�bhhK ��h��R�(KK��h�C,*      ,        >      v   �        �t�bhhK ��h��R�(KK��h�C:  �     �t�bhhK ��h��R�(KK��h�C<         h      5      -      y                 �t�bhhK ��h��R�(KK��h�C0      �     �	  �         I           �t�bhhK ��h��R�(KK��h�CD      �  �   E      <    �   s     ^   �     s        �t�bhhK ��h��R�(KK��h�C@
   ;     2               �      A   �              �t�bhhK ��h��R�(KK��h�C1   #       m  �         �t�bhhK ��h��R�(KK
��h�C(G     �       Q      �        �t�bhhK ��h��R�(KK��h�CH
   T  '   )   !         �      +        �     -          �t�bhhK ��h��R�(KK��h�C<     �t�bhhK ��h��R�(KK��h�C%   �   -           �t�bhhK ��h��R�(KK	��h�C$   �  �               �      �t�bhhK ��h��R�(KK��h�C�  
   ,      �t�bhhK ��h��R�(KK��h�C4   
        	      	      	   K   	   �      �t�bhhK ��h��R�(KK��h�C�   !      �t�bhhK ��h��R�(KK��h�CP                 >     �     �  �         C  V              �t�bhhK ��h��R�(KK��h�Cp      �t�bhhK ��h��R�(KK��h�C<�     �   �   �   �  �               �   �        �t�be(hhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�C|   f   �      P  )   �  A   =                             $   �	     �     $   0           =        �t�bhhK ��h��R�(KK��h�C,V   '   �  
     i   9  B   }         �t�bhhK ��h��R�(KK��h�C0-   H        ;      �  c   f   �        �t�bhhK ��h��R�(KK��h�C0#   !   (      
   �     �     F         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK
��h�C(1   #   9          �           �t�bhhK ��h��R�(KK��h�C �     >  	      	         �t�bhhK ��h��R�(KK	��h�C$   O  :  �  H   �	  �        �t�bhhK ��h��R�(KK��h�C,   '   -   A   #  i   �     +        �t�bhhK ��h��R�(KK"��h�C�                              %   �                 �     �      O           �	                          �t�bhhK ��h��R�(KK��h�C   @   '   H   �        �t�bhhK ��h��R�(KK��h�C,   �        �	     �   "   t         �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK	��h�C$�   _              �        �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C0*     2                            �t�bhhK ��h��R�(KK
��h�C(�          ?        �        �t�bhhK ��h��R�(KK
��h�C("   K  r  )   �                 �t�bhhK ��h��R�(KK��h�C|n  I   �	        �     f     g  (  �   2      0         )      2         G        f     g  )        �t�bhhK ��h��R�(KK��h�CT                                    >        �   )   �           �t�bhhK ��h��R�(KK��h�C<                              �  o           �t�bhhK ��h��R�(KK��h�C,   .        �   �  B  h   �         �t�bhhK ��h��R�(KK��h�C`     0   [      x      @                   �	                            �t�bhhK ��h��R�(KK��h�C8         �       A        0      �        �t�bhhK ��h��R�(KK
��h�C(   >   �  �  v   "             �t�bhhK ��h��R�(KK��h�C4%   _  C   -         A   Y  }      �        �t�bhhK ��h��R�(KK	��h�C$1  �    
                  �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�CP      n     *     %   �           �              
   &        �t�bhhK ��h��R�(KK��h�C8      �  8   �  "     �	          �        �t�bhhK ��h��R�(KK��h�C B  �   �   �      u         �t�bhhK ��h��R�(KK��h�C       A   6     N          �t�bhhK ��h��R�(KK��h�CH
        '  ,      �         �         �       ,         �t�bhhK ��h��R�(KK��h�C0T         P      �         C  E         �t�bhhK ��h��R�(KK��h�C �        	      	         �t�bhhK ��h��R�(KK��h�CD               �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�Cn     !        �t�bhhK ��h��R�(KK��h�CT%         .   �     �	     s   `     s   �  �   �       i   s   8     �t�bhhK ��h��R�(KK��h�C<�         v        �   E  �           �        �t�bhhK ��h��R�(KK��h�CL      9   %   Z  T   �  �   �   "   �     �   9                  �t�bhhK ��h��R�(KK��h�C�   -     �t�bhhK ��h��R�(KK��h�CH   o   �   F           �t�bhhK ��h��R�(KK��h�CH   8   S       i      �	  >            �     �   �	        �t�bhhK ��h��R�(KK��h�C    R        �   h        �t�bhhK ��h��R�(KK��h�C   �               �t�bhhK ��h��R�(KK	��h�C$�  �        i  "            �t�bhhK ��h��R�(KK��h�C\�                   B         �  +      �             0   !          �t�bhhK ��h��R�(KK��h�CH�     �      
   �           -   N      S        �        �t�bhhK ��h��R�(KK��h�C,%   '           �        ?        �t�bhhK ��h��R�(KK��h�CP      <               .            C      �	  
   C      	        �t�bhhK ��h��R�(KK	��h�C$      	      	      	   K      �t�bhhK ��h��R�(KK��h�CT   &        �   j        J   b   �              .                  �t�bhhK ��h��R�(KK��h�CP      5   <      [      �     �            �   L                  �t�bhhK ��h��R�(KK��h�C       �	  s      �   �      �t�bhhK ��h��R�(KK��h�C    ?     
   �            �t�bhhK ��h��R�(KK��h�C       0        �        �t�bhhK ��h��R�(KK��h�CTo  S        ,     �        �     ,   	      	   K   	     	   �      �t�bhhK ��h��R�(KK��h�C G     �      �          �t�bhhK ��h��R�(KK��h�C<;     	      	      	   K   	   I  	   /  	   �     �t�bhhK ��h��R�(KK��h�C4*         H     �         =      4         �t�bhhK ��h��R�(KK��h�CP*      &   $  �   "   F              �   L   
   c  
   F  F         �t�bhhK ��h��R�(KK��h�CI     !  �      �t�bhhK ��h��R�(KK��h�C,`           Q          I         �t�bhhK ��h��R�(KK��h�C@      	      	         �t�bhhK ��h��R�(KK��h�C,�     q   �  :   �        �
        �t�bhhK ��h��R�(KK��h�C0!      �	  �     R   '   
   �  F         �t�bhhK ��h��R�(KK��h�C@         O      �   S   Q   5         4      �         �t�bhhK ��h��R�(KK	��h�C$�  �   +   !      B   J        �t�bhhK ��h��R�(KK��h�C,f           �     p   �   :        �t�bhhK ��h��R�(KK��h�C<   f   �         0   	  )   y      �    7         �t�bhhK ��h��R�(KK��h�C@  �     �        �t�bhhK ��h��R�(KK��h�C1   #       �   p         �t�bhhK ��h��R�(KK��h�CH   �   �           v               �   �        �        �t�bhhK ��h��R�(KK��h�Clw       ]     p      �     �           y     K  z  �       �     �   /  A        �t�bhhK ��h��R�(KK��h�C L  �  �   M     �        �t�bhhK ��h��R�(KK��h�CT      �     N        S   Q      5         g  
  �      �   �        �t�bhhK ��h��R�(KK��h�C\      -   �   k  
              b      �            5   B  <      �        �t�bhhK ��h��R�(KK
��h�C(�  ?   2   �  H  �              �t�bhhK ��h��R�(KK��h�C@   $   �           !     W  
   \   �  �  Y        �t�bhhK ��h��R�(KK��h�Cx     �t�bhhK ��h��R�(KK��h�C0   P   4   
   _         	      	         �t�bhhK ��h��R�(KK��h�CT]     
        \   �	  �        �   :     Q         �              �t�bhhK ��h��R�(KK	��h�C$1   #       *      �  /         �t�bhhK ��h��R�(KK��h�C0"      '   H   B   �           z         �t�bhhK ��h��R�(KK��h�CT*      �       5         �        u     !     �   �   	  �        �t�bhhK ��h��R�(KK��h�C�      {      �     �t�bhhK ��h��R�(KK
��h�C(j  /  �     I   Y      ?        �t�bhhK ��h��R�(KK��h�C,O  �       �      i     �        �t�bhhK ��h��R�(KK��h�C<�  P     �  P     �   �	        m      �         �t�bhhK ��h��R�(KK��h�C Q        	      	         �t�bhhK ��h��R�(KK��h�C0S        	      	      	   K   	   �      �t�bhhK ��h��R�(KK��h�C@  �  2   �  )                        �  )        �t�bhhK ��h��R�(KK��h�C0�  &   N   �  9   �  $   �              �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�C<�     Z  R      �     l         �    7         �t�bhhK ��h��R�(KK��h�C<9        R  (      �   �     *         f        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C<
   T  �	  ?      �     '      �  
               �t�bhhK ��h��R�(KK��h�C4�  {     .        >	  T   D   �  N        �t�bhhK ��h��R�(KK
��h�C(�             	      	         �t�bhhK ��h��R�(KK��h�CS     �t�bhhK ��h��R�(KK��h�C4   R  )      �      ]           C        �t�bhhK ��h��R�(KK��h�C`   5   7        g              �  �	     �        �        Y      Q         �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�CL   	     l      T  C   :   �  m   x  *             >        �t�bhhK ��h��R�(KK��h�C4   (   �  �     �        ]  j   �        �t�bhhK ��h��R�(KK	��h�C$      -   N   U  
   �        �t�bhhK ��h��R�(KK��h�C,/      �   �
  �     5     e        �t�bhhK ��h��R�(KK��h�C\*   2         �   �     C   �  %   �      �      I   a     2   �             �t�bhhK ��h��R�(KK	��h�C$�   �     �      �  �         �t�bhhK ��h��R�(KK��h�C   �  �           �t�bhhK ��h��R�(KK��h�C\   (        x         =      �	     �  �     	  �         }              �t�bhhK ��h��R�(KK��h�CP   #  (           ;      \    h   �   a  g                    �t�bhhK ��h��R�(KK��h�C`      ]  �     '     %              >   M   �      *         �              �t�bhhK ��h��R�(KK��h�C`        I                     �   �           �
     /      p     �        �t�bhhK ��h��R�(KK��h�C,      l   �     7   �	  "            �t�bhhK ��h��R�(KK��h�C             �t�bhhK ��h��R�(KK��h�C �         7     	         �t�bhhK ��h��R�(KK��h�C�       �t�bhhK ��h��R�(KK��h�C�	       �  �   _     �t�bhhK ��h��R�(KK��h�Cd
   �  !        c  
   ,                  �                  &  
   8   X        �t�bhhK ��h��R�(KK��h�C,      �     V  D  �   �   �        �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   �        �        �t�bhhK ��h��R�(KK��h�C<     �	                      p     �        �t�bhhK ��h��R�(KK��h�C,V      2   )   z   ,      A   }         �t�bhhK ��h��R�(KK��h�CH�         /         9      7   �  �     T  �   �  o        �t�bhhK ��h��R�(KK��h�C8      �	     �      $   �	     �      (        �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C1   #       �        �t�bhhK ��h��R�(KK
��h�C(      �  �     `             �t�bhhK ��h��R�(KK	��h�C$1  '   
        @   �         �t�bhhK ��h��R�(KK��h�C0�  )                .  3  �        �t�bhhK ��h��R�(KK	��h�C$      -   a   �      �        �t�bhhK ��h��R�(KK��h�C,H   3  �     E     e      @         �t�bhhK ��h��R�(KK��h�C�  �         �t�bhhK ��h��R�(KK��h�C@�              J   �  ;               �           �t�bhhK ��h��R�(KK��h�Ct      �  l  �         S   Q      F  �      �      7         $   ;         �   �                  �t�bhhK ��h��R�(KK��h�CP   e   �   �     ,            e        e   {                    �t�bhhK ��h��R�(KK��h�C,"     ,  �     .      �             �t�bhhK ��h��R�(KK��h�C�  q     �t�bhhK ��h��R�(KK��h�C4         x      �     �  
   �   �        �t�bhhK ��h��R�(KK��h�C0   @   '      �              �        �t�bhhK ��h��R�(KK��h�Cv  �  �     G  w     �t�bhhK ��h��R�(KK��h�C,            K        �   O         �t�bhhK ��h��R�(KK��h�C0�  �      =      B   �	     �   �        �t�bhhK ��h��R�(KK��h�C<b   #      ?  
                 l     W        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C@      (               �   �         9   �  �        �t�bhhK ��h��R�(KK��h�CL�  (   �     D      �        �     l  �     C             �t�bhhK ��h��R�(KK��h�C0                           �        �t�bhhK ��h��R�(KK��h�C<*      �	     �      M               �	           �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C,a     E   y   8      4     c         �t�bhhK ��h��R�(KK��h�C,                  $              �t�bhhK ��h��R�(KK��h�C0                                    �t�bhhK ��h��R�(KK��h�C_     �         �t�bhhK ��h��R�(KK��h�Cd      P         �  T         E           �     �                 S   Q         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C�   �   E  	         �t�bhhK ��h��R�(KK��h�CD      �   X     M   T   �      �       
   8   �        �t�bhhK ��h��R�(KK��h�C,!         �         	      	         �t�bhhK ��h��R�(KK��h�Ch   $   n      �	        .      H          �             f   �     %   I  �        �t�bhhK ��h��R�(KK
��h�C(2  �           �  �  {        �t�bhhK ��h��R�(KK��h�Ct            �  4   
   _      �        =         0  4   *      t     +   �         0  4         �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C K  �   Y  	      	         �t�bhhK ��h��R�(KK
��h�C(      
   c  b   D     ]         �t�bhhK ��h��R�(KK��h�C   m        �t�bhhK ��h��R�(KK��h�C,1   #      �   "   �   
   T  �	        �t�bhhK ��h��R�(KK��h�C<�  q  �      .      B         �   ]     �        �t�bhhK ��h��R�(KK��h�C<%            %   �        `   �     A   [        �t�bhhK ��h��R�(KK��h�C8[  L  
   y       �   �   M     {  _        �t�bhhK ��h��R�(KK��h�CZ   Z     �t�bhhK ��h��R�(KK��h�Ch         O      �   S   Q            8   4      �   ;      �      �  �        �         �t�bhhK ��h��R�(KK��h�C,   w  J  2   C   ^   e   �   F         �t�bhhK ��h��R�(KK��h�C@         O         
  Q   5         4               �t�bhhK ��h��R�(KK��h�C4   5   4      m        ,     .             �t�bhhK ��h��R�(KK��h�CD
   �        -         S  [    D	  3  i   
   �        �t�bhhK ��h��R�(KK��h�C<f           �              ,   	      	         �t�bhhK ��h��R�(KK��h�C<�   f     g        �              �   �        �t�bhhK ��h��R�(KK��h�CT*   �  '   
   �     �     �      �   B     A  #  2        �	        �t�bhhK ��h��R�(KK'��h�C�<      !      l                  	      	      	   K   	   �   	   �   	     	   I  	   �  	   U  	   �   	   �  	   �  	   �  	        �t�bhhK ��h��R�(KK
��h�C(     �  "     @               �t�bhhK ��h��R�(KK��h�C0�     W     ?      
   $   \  F         �t�bhhK ��h��R�(KK��h�C      &      w  ]     �t�bhhK ��h��R�(KK��h�C ?  �     �   S   X        �t�bhhK ��h��R�(KK
��h�C(      �     2   �  �  \        �t�bhhK ��h��R�(KK��h�C4^        #  !     .  �  :   �           �t�bhhK ��h��R�(KK��h�C8�   '      �      V         �  
            �t�bhhK ��h��R�(KK��h�C8      �  u  C  h                  +         �t�bhhK ��h��R�(KK��h�C/  ^            �t�bhhK ��h��R�(KK��h�C8�  J  )     
   _      �
                   �t�bhhK ��h��R�(KK��h�CD!      |      <  R   ?      
   3   6   �     �   f        �t�bhhK ��h��R�(KK&��h�C�         E  H     �     �   S   Y      Q            x     #     $     �     y      W           �  $   E                  �t�bhhK ��h��R�(KK
��h�C(#   !   ?      
   X   �   F         �t�bhhK ��h��R�(KK��h�C0�     ;     w  V   2   5   B  �         �t�bhhK ��h��R�(KK
��h�C(b         "   �	                 �t�bhhK ��h��R�(KK	��h�C$   ]   �      H  d   �         �t�bhhK ��h��R�(KK��h�C   y     �t�bhhK ��h��R�(KK��h�C,      c  
         	      	         �t�bhhK ��h��R�(KK��h�C                     �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CP      �     $  `   �      [     5  _     0   !                �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK	��h�C$1   A  S  y      r	           �t�bhhK ��h��R�(KK	��h�C$q   l  }      ,               �t�bhhK ��h��R�(KK��h�CPY      O               ,        -   �  �      (	     q   �	        �t�bhhK ��h��R�(KK��h�C@         4                       '   `          �t�bhhK ��h��R�(KK��h�C,               �  �               �t�bhhK ��h��R�(KK��h�C    ?   �  
   �	  F         �t�bhhK ��h��R�(KK��h�CR      �     �t�bhhK ��h��R�(KK��h�CE      4           �t�bhhK ��h��R�(KK	��h�C$�     �  K  	      	         �t�bhhK ��h��R�(KK��h�C       M  	      	         �t�bhhK ��h��R�(KK��h�CL      �  o   �  8            �           0   `     �        �t�bhhK ��h��R�(KK��h�CX      \       �  c         ]           d  �    �     U   �        �t�bhhK ��h��R�(KK��h�C8   %   �  :           �         o  �         �t�bhhK ��h��R�(KK��h�C*         %     �t�bhhK ��h��R�(KK��h�C@b   $   �   �        $  
      �        J   P         �t�bhhK ��h��R�(KK
��h�C(   �        /      9  7         �t�bhhK ��h��R�(KK��h�C�  '   9               �t�bhhK ��h��R�(KK��h�CH
   �  F   '   \     B   I  V         z   ,   
   �   �         �t�bhhK ��h��R�(KK��h�Cl   4        �  B   �  a        .         S   X        �        d  i         �        �t�bhhK ��h��R�(KK��h�C@  �     �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK
��h�C(b   #   G   �   �     R  �         �t�bhhK ��h��R�(KK��h�C8   �     L  h   �  L   >   p  �  
   �        �t�bhhK ��h��R�(KK��h�C,   �  �       F        b        �t�bhhK ��h��R�(KK��h�C`
   �              �                     �                                �t�bhhK ��h��R�(KK��h�C8      K     W   C  $   ;      %   �           �t�bhhK ��h��R�(KK��h�Cl   X   M     
   ,   -   
                                          �                 �t�bhhK ��h��R�(KK��h�CD*   D   l     5  �  2   �      �      I        P	        �t�bhhK ��h��R�(KK��h�C &        �   p  �        �t�bhhK ��h��R�(KK��h�CL   @   '   �  "     V   l      G        j   �      0            �t�bhhK ��h��R�(KK��h�C8U  4     A   F     �     �
  +      n         �t�bhhK ��h��R�(KK��h�C\R    
   %     �        b         :     Q      �      +   �              �t�bhhK ��h��R�(KK	��h�C$�     o  �  	      	         �t�bhhK ��h��R�(KK��h�C]   �              �t�bhhK ��h��R�(KK��h�C �     M  	      	         �t�bhhK ��h��R�(KK
��h�C("   �      2      �     �         �t�bhhK ��h��R�(KK
��h�C(1   #       �	     /      �         �t�bhhK ��h��R�(KK
��h�C(   �        �   �   �  7         �t�bhhK ��h��R�(KK��h�C,      �  
   ,                     �t�bhhK ��h��R�(KK��h�C8        �    �      ,         Y  �        �t�bhhK ��h��R�(KK��h�C8*      �  B  7   �  �  @   �                 �t�bhhK ��h��R�(KK��h�CHB     `   �  "                �  )         !  �         �t�bhhK ��h��R�(KK��h�CL*      �     �     W  �     5  8   t     �        �         �t�bhhK ��h��R�(KK��h�C      Y        �t�bhhK ��h��R�(KK��h�CD      �            2   (   H     j   �   �   �  �        �t�bhhK ��h��R�(KK
��h�C(   `        z   h   H   �        �t�bhhK ��h��R�(KK	��h�C$u      ;         r  �        �t�bhhK ��h��R�(KK��h�CZ     L           �t�bhhK ��h��R�(KK��h�CX   H     ?      �  
         /     �      �     I     �      K         �t�bhhK ��h��R�(KK��h�C �  @     m	              �t�bhhK ��h��R�(KK��h�Ch      �     $      �  =     �      L            
        8   �     G      �	        �t�bhhK ��h��R�(KK��h�Ct*               �  W   �   �      $   �           �   �               �     @     �  �        �t�bhhK ��h��R�(KK��h�C<   �  (            �  
   _      F              �t�bhhK ��h��R�(KK��h�C  �         �t�bhhK ��h��R�(KK��h�C<      0   +  4                  m              �t�bhhK ��h��R�(KK��h�C0�   c  �   I   �     c  �   I   �         �t�bhhK ��h��R�(KK��h�CX   �      $     �  �   Y  +      �  +      �            U      �        �t�bhhK ��h��R�(KK��h�C|      �	          .            o  9               S   Y   �   Q     Q      x     �  i      7         �t�bhhK ��h��R�(KK��h�C\9   �     �  '   �     /   9   9  7   "   ~  y     e      
   d     @         �t�bhhK ��h��R�(KK��h�CD         :   n     �  �     %     �      e           �t�bhhK ��h��R�(KK��h�C\      �  �     �  �     D            �  �  s    N  D   &   O           �t�bhhK ��h��R�(KK��h�CC                �t�bhhK ��h��R�(KK��h�C1   #          �t�bhhK ��h��R�(KK��h�C	  	      	         �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�C4      �      �t�bhhK ��h��R�(KK	��h�C$�     �   �     �   �        �t�bhhK ��h��R�(KK��h�CH
        @   �         V   2      �	  C         c  ,         �t�bhhK ��h��R�(KK��h�C\   $   8     4            ~               0   4         
   _      �        �t�bhhK ��h��R�(KK��h�C8     T  C   :   m         �                �t�bhhK ��h��R�(KK��h�C8
   3   6   �  '   !         �     W   �         �t�bhhK ��h��R�(KK��h�C   �     $  �        �t�bhhK ��h��R�(KK��h�C@  K	  G   W         �t�bhhK ��h��R�(KK��h�CL      P         �        �   
      �  }         �  E         �t�bhhK ��h��R�(KK��h�C<�  �           .   @            �   -  5        �t�bhhK ��h��R�(KK��h�C<�   '      .   
                    (           �t�bhhK ��h��R�(KK��h�C   �            �t�bhhK ��h��R�(KK
��h�C(�  ~   H   z        �  *        �t�bhhK ��h��R�(KK��h�C   �  �      �t�bhhK ��h��R�(KK��h�C8         1  �  �     c        
           �t�bhhK ��h��R�(KK��h�C@�  l     w  �   :   .        �  T   A     �         �t�bhhK ��h��R�(KK��h�C0       .   "   H                     �t�bhhK ��h��R�(KK��h�C,      �  &         .     �        �t�bhhK ��h��R�(KK��h�C8   X   '   s   `     �	                       �t�bhhK ��h��R�(KK��h�CD   @      u     w       �   &  �  �   0  B   �        �t�bhhK ��h��R�(KK��h�CX�   �      �     I     �   �     �           �  �     )   �   <         �t�bhhK ��h��R�(KK��h�C�                     �t�bhhK ��h��R�(KK	��h�C$M   �      �  
   $   �        �t�bhhK ��h��R�(KK��h�C      �           �t�bhhK ��h��R�(KK��h�CDO     �          �   l     �  M     �     �  �        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK
��h�C(I      ]  �     R               �t�bhhK ��h��R�(KK	��h�C$�  ;              P        �t�bhhK ��h��R�(KK��h�CD�         b      x      0   [      �	     ~     /         �t�bhhK ��h��R�(KK��h�CL   [  �     .   �     W      �      (        "   e   �         �t�bhhK ��h��R�(KK��h�C9  7      �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C8f  �  �  M     �     �  �  �     �        �t�bhhK ��h��R�(KK��h�CD      A   g     %   s         �        "     g        �t�bhhK ��h��R�(KK��h�C0        '      h     \               �t�bhhK ��h��R�(KK��h�C   �         �t�bhhK ��h��R�(KK��h�C4   >  v           '                    �t�bhhK ��h��R�(KK��h�C8         Y      O   5         4               �t�bhhK ��h��R�(KK��h�C,�	          �     M  �     ,      �t�bhhK ��h��R�(KK	��h�C$      i     i  
   w        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C\         �  "   �      (        b      �     ,         "   �      (        �t�bhhK ��h��R�(KK��h�C�     �      �        �t�bhhK ��h��R�(KK��h�C    @   '   )   #  W        �t�bhhK ��h��R�(KK��h�C j  &   a   �     �        �t�bhhK ��h��R�(KK
��h�C(1   #       �     �	              �t�bhhK ��h��R�(KK��h�C<      �  $   0  "   �  �     �   "   q   �        �t�bhhK ��h��R�(KK��h�Cd         �      G  :      Q   �  Q     �  5      -         y         �   >        �t�bhhK ��h��R�(KK��h�C"           �t�bhhK ��h��R�(KK��h�C,.  M     �  
   �    
   ,         �t�bhhK ��h��R�(KK��h�C@     C         �  �  %        �                 �t�bhhK ��h��R�(KK��h�C
   y     �t�bhhK ��h��R�(KK��h�CH�         �   ,                      �   �               �t�bhhK ��h��R�(KK��h�CHq   k  �	        �	     l  g      �  %   �   m     E        �t�bhhK ��h��R�(KK	��h�C$�  �        	      	         �t�bhhK ��h��R�(KK��h�Cn        �t�bhhK ��h��R�(KK#��h�C�         �           .      0      n	  �  g	     &      �        $                       \      �  $            �t�bhhK ��h��R�(KK��h�CL      �   E   &      �  #           �  3     �  D  �        �t�bhhK ��h��R�(KK��h�C8#   !      t        (      
   3   6   n        �t�bhhK ��h��R�(KK��h�CT      �   f  &      )  +   G   |      �   �       �     $            �t�bhhK ��h��R�(KK
��h�C(%   �   &   -   �  �	     �        �t�bhhK ��h��R�(KK��h�C0   f   ,  '      -                     �t�bhhK ��h��R�(KK	��h�C$�  "  S       �            �t�bhhK ��h��R�(KK��h�C04     (     9       
   8   �	        �t�bhhK ��h��R�(KK��h�C0+  �     Y      O   �	  �  :   H        �t�bhhK ��h��R�(KK��h�C4      H   A   ?     m        �  n        �t�bhhK ��h��R�(KK(��h�C�
   t            9         �     ]   �	     )   0      �   ~              �  �     
  T      o  4      $   �     Y      O            �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   6         �        �t�bhhK ��h��R�(KK��h�C�   =  	         �t�bhhK ��h��R�(KK
��h�C(   �  �	  �	     Q  $   �        �t�bhhK ��h��R�(KK��h�C<K  �  �      �  �      6     �        �        �t�bhhK ��h��R�(KK��h�Cd�      �   �              �     4          b       �   p  q  �  7            �t�bhhK ��h��R�(KK��h�C0]           %     �        �        �t�bhhK ��h��R�(KK��h�CX*               
   _      �              ;      �      z               �t�bhhK ��h��R�(KK��h�C07      �  @      �   �  �  
            �t�bhhK ��h��R�(KK��h�Cx4  �         0  s   �                             �           X  E                 p         �t�bhhK ��h��R�(KK��h�C02      )      �               y        �t�bhhK ��h��R�(KK��h�CH      0   c  �            v           +   :      �         �t�bhhK ��h��R�(KK��h�C         	         �t�bhhK ��h��R�(KK
��h�C(�  �     R     	      	         �t�bhhK ��h��R�(KK��h�C�   �   p     �t�bhhK ��h��R�(KK��h�CD           %             H  �                     �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C8   �              r  s     %               �t�bhhK ��h��R�(KK	��h�C$   �	     	                 �t�bhhK ��h��R�(KK��h�C4*         &      �  $   !       Z        �t�bhhK ��h��R�(KK��h�C@1   #      �     �   
   3   6   �     :             �t�bhhK ��h��R�(KK��h�CH     t     �	  �            
   _      �   u  �        �t�bhhK ��h��R�(KK��h�CD%  �        �	              G     �        �         �t�bhhK ��h��R�(KK��h�C@   (   #   !      [        "   �  
   $   �   �        �t�bhhK ��h��R�(KK��h�CL�	  �   �                          O         Y      Q         �t�bhhK ��h��R�(KK��h�C0M      +   3        &   i  �  �        �t�bhhK ��h��R�(KK��h�CH!           �   (      "   k     �  "   �  v  �          �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�Cb   #   G   W         �t�bhhK ��h��R�(KK��h�CD*           �           &      n  �   v               �t�bhhK ��h��R�(KK��h�Cw     x        �t�bhhK ��h��R�(KK��h�C01   #       q         �
     �
           �t�bhhK ��h��R�(KK��h�CdX     y  =  i     z        �  �                          �   �	     T        �t�bhhK ��h��R�(KK��h�C<"   �  �  (      x      <         �     o         �t�bhhK ��h��R�(KK��h�C l     �        �         �t�bhhK ��h��R�(KK��h�C f   �	           [         �t�bhhK ��h��R�(KK��h�C\      J     `   �            %   �         E  �         <      {  b        �t�bhhK ��h��R�(KK��h�C8   ]   �         =      L     ]   �  �        �t�bhhK ��h��R�(KK��h�Ct                        w      �        |  =      4   h   �   �            �  =      �        �t�bhhK ��h��R�(KK��h�C<>        ?      �         
     
               �t�bhhK ��h��R�(KK��h�Cd      >     �        $   n         �       �         0   �     �      <        �t�bhhK ��h��R�(KK��h�C �        	      	         �t�bhhK ��h��R�(KK��h�C`   $   n      �	     .      H          �          f   �     %   I  �        �t�bhhK ��h��R�(KK
��h�C(8        �    	      	         �t�bhhK ��h��R�(KK��h�C�  �      S     �t�bhhK ��h��R�(KK��h�CH
      ]  T  '   !            �   �      �     �            �t�bhhK ��h��R�(KK��h�C,�     j                 �        �t�bhhK ��h��R�(KK��h�CD      '   �   �     ,        �  	  C  �     �        �t�bhhK ��h��R�(KK��h�C<
   @   �   F   '   #   !      �         i  }        �t�bhhK ��h��R�(KK��h�C\         .   0         F     �                 D  �   �     8   S        �t�bhhK ��h��R�(KK��h�C�              �t�bhhK ��h��R�(KK��h�C    �  �  �     c         �t�bhhK ��h��R�(KK��h�CP      -   �   L   G        �     ~        Z  
   $   �   N        �t�bhhK ��h��R�(KK��h�C4   f   �      �  N      �      $   L        �t�bhhK ��h��R�(KK��h�C4      �     �  "   �     T     C        �t�bhhK ��h��R�(KK��h�C�  J  �         �t�bhhK ��h��R�(KK��h�C@`     �  �	  N           �              a        �t�bhhK ��h��R�(KK��h�C1   #       �         �t�bhhK ��h��R�(KK��h�C'  �  �      `     �t�bhhK ��h��R�(KK��h�C�     C     �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C#  a    r      �t�bhhK ��h��R�(KK��h�CP1   #      �      A   �  �         �   �  �	  
   3   6      �        �t�bhhK ��h��R�(KK��h�C`      �     I        i              Z                                   �t�bhhK ��h��R�(KK��h�Ch�      �                 .  &                                                  �t�bhhK ��h��R�(KK��h�Ct"   m      �      �  (      <        ^  �
           �   �  ?       ^  @     �   
  T        �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�Ch"   �  B  h   �         U   @     �     �  �  �                �  �  �   �        �t�bhhK ��h��R�(KK��h�C�     �  �   r      �t�bhhK ��h��R�(KK��h�Ct   ]  T     ;     +         O      �   S   Q         Y      Q      #     $     x     �        �t�bhhK ��h��R�(KK��h�CH      L             ?        2   
         �	  �        �t�bhhK ��h��R�(KK��h�C`      J      8   /   &   �     �  �           �     b      �     $   k         �t�bhhK ��h��R�(KK��h�C,         Y      O         O          �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C4   f     '            �  V   �  �        �t�bhhK ��h��R�(KK��h�C1   #       +     �t�bhhK ��h��R�(KK��h�Cd   B  (   2   )   <   "   X   �   @     �     �  �  �                �  �        �t�bhhK ��h��R�(KK��h�C8#   !      \      a  u	  ?      
   �  F         �t�bhhK ��h��R�(KK��h�Cd      -   v      
   &           X	                                            �t�bhhK ��h��R�(KK��h�C
  �     �      �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C,         &      
     �          �t�bhhK ��h��R�(KK��h�C1   #       9        �t�bhhK ��h��R�(KK��h�C,U     *      �           %        �t�bhhK ��h��R�(KK��h�CH�           �   H         �          �  /      �         �t�bhhK ��h��R�(KK��h�C,G        6  C   I  ,      |        �t�bhhK ��h��R�(KK ��h�C�M      +   `      	      	      	   �   	   �   	   I  	   /  	   s  	   )  	   �  	   �	  	   �  	   �  	   �     �t�bhhK ��h��R�(KK��h�CD      J      `            �   �  B                    �t�bhhK ��h��R�(KK��h�C            B            �t�bhhK ��h��R�(KK��h�C|  �      �     �     �t�bhhK ��h��R�(KK!��h�C�   5   �      �  �   `   �          �      �         �      M      �               �      �   J   *  �         �t�bhhK ��h��R�(KK��h�CL     '      f        &     s   (        �
        �        �t�bhhK ��h��R�(KK
��h�C(�           P  
     �         �t�bhhK ��h��R�(KK��h�C�      {      �t�bhhK ��h��R�(KK��h�CX�     �  �  >   N            2   �  :   �   &   D  �  �   U             �t�bhhK ��h��R�(KK��h�CD*            �  &      U                  $            �t�bhhK ��h��R�(KK��h�C@      �  �   $   b   ^      
   ,                     �t�bhhK ��h��R�(KK��h�C82         =         �  �  ^   �              �t�bhhK ��h��R�(KK��h�Ch  �     �t�bhhK ��h��R�(KK��h�C �  a  �           �     �t�bhhK ��h��R�(KK��h�CH�  
      �   x      �      $  �  �  �      
              �t�bhhK ��h��R�(KK��h�C,      W	     @      z  �          �t�bhhK ��h��R�(KK��h�C@           �      �  �      �   U   U  ^   �         �t�bhhK ��h��R�(KK��h�C0�	  �  �  �     $   E      �  �         �t�bhhK ��h��R�(KK��h�C8)      /      �        5      4               �t�bhhK ��h��R�(KK	��h�C$�	  �  7  h     q   �        �t�bhhK ��h��R�(KK��h�CX      X   '      �     �
  X   "      �     "      9        �	           �t�bhhK ��h��R�(KK��h�Cd        �   O         �t�bhhK ��h��R�(KK��h�Cc  �  	      	         �t�bhhK ��h��R�(KK"��h�C�V  �      ;         D	     !     �  �           �     �                �  j      �        �  �           �t�bhhK ��h��R�(KK��h�C4   X   '   s                               �t�bhhK ��h��R�(KK��h�CT      )  +         �      �     y           �      .     �        �t�bhhK ��h��R�(KK��h�C�      �     �t�bhhK ��h��R�(KK��h�C8      N      U  �  D      a  c   �  s         �t�bhhK ��h��R�(KK	��h�C$        �                  �t�bhhK ��h��R�(KK��h�C\�   N        �   �     �        2      �         �   L           Z        �t�bhhK ��h��R�(KK��h�CT   $   �  �      
      
    �  Y  �           U   �     �        �t�bhhK ��h��R�(KK��h�C@            0   �  )   "   t      2  
   $   �        �t�bhhK ��h��R�(KK��h�C,1   #      >  
   3   6      [        �t�bhhK ��h��R�(KK��h�C<8        l  �  [  �      H   �     �      d      �t�bhhK ��h��R�(KK��h�CPT   �  �     .   \   �  �     �         \   2         :   �         �t�bhhK ��h��R�(KK��h�C�     W     �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�CP
               F         P   !         
   $   �     C  �        �t�bhhK ��h��R�(KK��h�C      U             �t�b�      hhK ��h��R�(KK��h�C,v        .   �           
        �t�bhhK ��h��R�(KK��h�CD     X         �t�bhhK ��h��R�(KK��h�Ct     �	     �t�bhhK ��h��R�(KK��h�C`   �  C      ;  C         <     S     Y  
     e  i      �  �	     �        �t�bhhK ��h��R�(KK��h�C4      J   4        5      �      4         �t�bhhK ��h��R�(KK
��h�C(�              -   
           �t�bhhK ��h��R�(KK��h�C "   >  �        �        �t�bhhK ��h��R�(KK��h�C             �t�bhhK ��h��R�(KK��h�C�  !      �          �t�bhhK ��h��R�(KK��h�Cl   C          D   �        T   �  �  �     �     �      D      )      �   ~   �         �t�bhhK ��h��R�(KK	��h�C$
        �      
   �        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�CB  q     �        �t�bhhK ��h��R�(KK��h�C   9     �  7      �t�bhhK ��h��R�(KK��h�Ch      �     �	       
         �     �        �     ,      K                     �t�bhhK ��h��R�(KK��h�C<      =      
  G   �        �     �           �t�bhhK ��h��R�(KK��h�C�              �t�bhhK ��h��R�(KK��h�C0v  w        .   �                    �t�bhhK ��h��R�(KK
��h�C(W   �   �      
   8   t           �t�bhhK ��h��R�(KK��h�C,M         �          8   4         �t�bhhK ��h��R�(KK��h�C`�   �   �  A  :   �   �     $   �               $   A  g            E  �         �t�bhhK ��h��R�(KK��h�C<1   #           o     �  
   3   6      l         �t�bhhK ��h��R�(KK��h�Cpq         �                 #                 �                                      �t�bhhK ��h��R�(KK��h�C8\   �  [      (     
   \   �   <      5         �t�bhhK ��h��R�(KK��h�C-	              �t�bhhK ��h��R�(KK��h�C8"   6    )         5   �      Z     i        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C1        	         �t�bhhK ��h��R�(KK��h�C1   #       �          �t�bhhK ��h��R�(KK��h�C,   �  �   )                       �t�bhhK ��h��R�(KK��h�C	     �t�bhhK ��h��R�(KK��h�C8           �  	      	   K   	     	   �      �t�bhhK ��h��R�(KK��h�C1   #       �         �t�bhhK ��h��R�(KK��h�C	  �  �     �t�bhhK ��h��R�(KK��h�CL         '   �                      �  h      �   t        �t�bhhK ��h��R�(KK
��h�C(o  �         �   �     4         �t�bhhK ��h��R�(KK��h�C42   	
  (     �                         �t�bhhK ��h��R�(KK
��h�C(      I  ,                     �t�bhhK ��h��R�(KK��h�C,
   )  &   2   �	  C                  �t�bhhK ��h��R�(KK��h�C0   �     S                           �t�bhhK ��h��R�(KK��h�C01   #   
   3   6   �           �         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CL      -   �   L   G      �   

        R      9  �     �        �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C�      '	        �t�bhhK ��h��R�(KK��h�CP      �     .   J   �	        9      &   ]   �  9   %               �t�bhhK ��h��R�(KK��h�C<      �              �  :   I   �              �t�bhhK ��h��R�(KK��h�C1         �t�bhhK ��h��R�(KK��h�C      �           �t�bhhK ��h��R�(KK��h�CH         Y     l      +	     C  V     A         +	        �t�bhhK ��h��R�(KK��h�CD   �    �      .         *      &   N   �     �	        �t�bhhK ��h��R�(KK
��h�C(      0   <   
   �   B   }         �t�bhhK ��h��R�(KK��h�CG  	         �t�bhhK ��h��R�(KK	��h�C$   5      �   L   
   �        �t�bhhK ��h��R�(KK��h�C   s  �        �t�bhhK ��h��R�(KK��h�C�          �           �t�bhhK ��h��R�(KK��h�C0   �     �        �       �        �t�bhhK ��h��R�(KK��h�C       P   �  G   W         �t�bhhK ��h��R�(KK��h�CX         F     �  L   &      M     
      �      N           +         �t�bhhK ��h��R�(KK��h�C �              �         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK
��h�C(f   _     k  u  _              �t�bhhK ��h��R�(KK��h�C <      a  	      	         �t�bhhK ��h��R�(KK
��h�C(   (   �   )   "      M	  \        �t�bhhK ��h��R�(KK��h�CD            o      X            �  G     X   �        �t�bhhK ��h��R�(KK��h�C      �     �t�bhhK ��h��R�(KK��h�C8�	     v         �           T   �	           �t�bhhK ��h��R�(KK��h�C4
   3   6   {     �  ?      !               �t�bhhK ��h��R�(KK��h�C�     �      �t�bhhK ��h��R�(KK��h�C4      �
  8  �
     Z       �  �        �t�bhhK ��h��R�(KK��h�C0�         R      �     �  �        �t�bhhK ��h��R�(KK��h�C@   �  �      S         �     �        =   �        �t�bhhK ��h��R�(KK
��h�C(�  !   ?      
   �    _        �t�bhhK ��h��R�(KK��h�C�      �     �t�bhhK ��h��R�(KK��h�CL
   X     M                 V   2      �	  
      c  ,         �t�bhhK ��h��R�(KK��h�CH�           <      q  �  �     Q          �	           �t�bhhK ��h��R�(KK��h�C 1   #       �     _        �t�bhhK ��h��R�(KK��h�C<;     )   =         0  �  �      C  J  <        �t�bhhK ��h��R�(KK��h�Ct]   �        9           N  Y                                  �   w         
  8        �t�bhhK ��h��R�(KK��h�C   �  7   �           �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C8   (   #   !   
   3   6   9     �              �t�bhhK ��h��R�(KK��h�C@     q            �t�bhhK ��h��R�(KK��h�C             m  ;          �t�bhhK ��h��R�(KK��h�C,)         q   k  �         u         �t�bhhK ��h��R�(KK��h�C
  �  �     A   �      �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK	��h�C$1   #       �  �      S        �t�bhhK ��h��R�(KK��h�C,Z      �               �            �t�bhhK ��h��R�(KK��h�C0     �     S     
   �   B   }         �t�bhhK ��h��R�(KK��h�C@E      -     �         d     `   U  &   q           �t�bhhK ��h��R�(KK��h�Ca  P           �     �t�bhhK ��h��R�(KK��h�C \   �  
  Z  �  
   }     �t�bhhK ��h��R�(KK��h�C�   �     
     �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�C@        �        �t�bhhK ��h��R�(KK��h�C %      �      A   R         �t�bhhK ��h��R�(KK��h�C`      M     
            "     F     k            +   "   t   
   $   �        �t�bhhK ��h��R�(KK��h�C �  	  *  �        r      �t�bhhK ��h��R�(KK��h�C        
   K        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�Cx         @  
   �  }      
   ,               A   �     2   -   �  
   �   
         �              �t�bhhK ��h��R�(KK��h�C8   �                 �   �     �           �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C,%   �   +      �        8           �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C 
                      �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�CL   �      c  X  e     �      (           �    
           �t�bhhK ��h��R�(KK��h�C0                     �  �   �         �t�bhhK ��h��R�(KK��h�C4        a   /      �           �        �t�bhhK ��h��R�(KK��h�C�      0   !  �     �t�bhhK ��h��R�(KK!��h�C�         Y     A   ?                          >      w   M     
            ;      0   �  :   �   ?        �t�bhhK ��h��R�(KK��h�C,$   �  5      N   �     �   �          �t�bhhK ��h��R�(KK��h�C�      ,      /      �t�bhhK ��h��R�(KK	��h�C$#   !   ?      
   �  F         �t�bhhK ��h��R�(KK��h�C0b   #      �           W  �           �t�bhhK ��h��R�(KK	��h�C$
   )        �      R        �t�bhhK ��h��R�(KK��h�C<�  g  k              
     �  k     X         �t�bhhK ��h��R�(KK��h�C       �      c    e     �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C@�   �     �     l             �   �               �t�bhhK ��h��R�(KK��h�Cb   #   
   W         �t�bhhK ��h��R�(KK��h�C0!      0     x   "      	      	         �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK	��h�C$E      �   L     s            �t�bhhK ��h��R�(KK��h�C   =  �  �     �t�bhhK ��h��R�(KK
��h�C(�     )   �          �        �t�bhhK ��h��R�(KK��h�CLy      J  +      �   &      �   +            
   %   B            �t�bhhK ��h��R�(KK��h�C8      X                    �               �t�bhhK ��h��R�(KK!��h�C�   &   �     �           �                                   �     �              
     %   �         �t�bhhK ��h��R�(KK
��h�C(!         	   K   	   �   	   ^     �t�bhhK ��h��R�(KK��h�CX   K     D         l        >   N   d   �        D   &   D  0   4         �t�bhhK ��h��R�(KK
��h�C(   (   �  3  -   :   �   �        �t�bhhK ��h��R�(KK��h�CP      M   c   A    _     $   
       d              �        �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK��h�C8�   >      �      L   G   �                  �t�bhhK ��h��R�(KK��h�C8      ;     l         �   �      
           �t�bhhK ��h��R�(KK��h�C\
     '            �                 �   y  !            R      	        �t�bhhK ��h��R�(KK��h�C@�  (      9   �   _     �   �            8            �t�bhhK ��h��R�(KK��h�C4   "   �     �   �      ,   �   
            �t�bhhK ��h��R�(KK
��h�C(%   �   +         +               �t�bhhK ��h��R�(KK��h�C       0   �  :   W         �t�bhhK ��h��R�(KK��h�C D     [      a  	         �t�bhhK ��h��R�(KK��h�C<      ~     /      �t�bhhK ��h��R�(KK	��h�C$�	             l  �        �t�bhhK ��h��R�(KK��h�Ch        �   o         `      :      Q         S      -         `   �                 �t�bhhK ��h��R�(KK��h�C<
   3   6   1     	  ?      !      R      	        �t�bhhK ��h��R�(KK��h�C  
   �     �t�bhhK ��h��R�(KK��h�C4      '   H   o      �   B   
              �t�bhhK ��h��R�(KK��h�CD%                       X   V   2   (   [      x         �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK
��h�C(   @          H   3  �        �t�bhhK ��h��R�(KK��h�Cl*      d  �
  &      R     S   1        �                �        �   ;     +        �t�bhhK ��h��R�(KK��h�C0"   �  �  �     p   �       u         �t�bhhK ��h��R�(KK��h�C8   (   #   !      k   
   3   6   2              �t�bhhK ��h��R�(KK��h�C@   J  E   �   s   o  �   7      
        
   �        �t�bhhK ��h��R�(KK��h�Cl   &     �        �        Y      Q              Y   
  �         5   &     �        �t�bhhK ��h��R�(KK��h�C0B  
   c  %  
          �   ~        �t�bhhK ��h��R�(KK	��h�C$(       �  :   1          �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK
��h�C(*      J      $   �     `   �     �t�bhhK ��h��R�(KK��h�CD   >   �   a   L     ;      G        �   �   j   L        �t�bhhK ��h��R�(KK��h�C,#   !         ?      
   T           �t�bhhK ��h��R�(KK��h�CD�           �   R  �  �      �     E     A   !        �t�bhhK ��h��R�(KK��h�C<�        P   <   "   @       '   
   H   [        �t�bhhK ��h��R�(KK��h�C�   
           �t�bhhK ��h��R�(KK��h�C8      �               �   5         4         �t�bhhK ��h��R�(KK	��h�C$<      �          �  �     �t�bhhK ��h��R�(KK��h�C,!         i     �  	      	         �t�bhhK ��h��R�(KK��h�C0*      /   �        �        �  0      �t�bhhK ��h��R�(KK��h�C   ?   �  
   �        �t�bhhK ��h��R�(KK	��h�C$   p       d              �t�bhhK ��h��R�(KK��h�C8   �         �        �  ;  �     �        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C&     .  �  �         �t�bhhK ��h��R�(KK��h�C\1   #      l     /   
   3   �  �	     �        K                r         �t�bhhK ��h��R�(KK��h�CLT   �  2   [     �  �     �  I  z     �  �  �  
            �t�bhhK ��h��R�(KK	��h�C$  	  �  A   3  �  �        �t�bhhK ��h��R�(KK��h�C@�      *     �     g  �    7   g      x  �        �t�bhhK ��h��R�(KK��h�CD         m      s     �     &      M   �      b        �t�bhhK ��h��R�(KK��h�C`              �   f     �     �  W      �        �      �     H   �        �t�bhhK ��h��R�(KK
��h�C(         �     )  ^            �t�bhhK ��h��R�(KK��h�C�     �      �t�bhhK ��h��R�(KK��h�C1     3   T         �t�bhhK ��h��R�(KK��h�C,d   �     �   O      �      �        �t�bhhK ��h��R�(KK��h�C,,      V     z  �  �     �        �t�bhhK ��h��R�(KK��h�C �  �  �     ,   O         �t�bhhK ��h��R�(KK��h�C0�  �
           �	     �     v	        �t�bhhK ��h��R�(KK��h�CD      �        �      �  4   y   8   3  4     c         �t�bhhK ��h��R�(KK��h�Cp*   �   1     �     5   <         �        �        �   =                                 �t�bhhK ��h��R�(KK��h�C@   �  �  u            4      u            Z        �t�bhhK ��h��R�(KK��h�Cl   $   \     M	              �   '      #   !      �      
   3   6     *         F        �t�bhhK ��h��R�(KK��h�C0�  �  �   
  
   ,            K         �t�bhhK ��h��R�(KK��h�C8        >                    D  �        �t�bhhK ��h��R�(KK
��h�C(�  �     �   �        8   �      �t�bhhK ��h��R�(KK	��h�C$�  4      K  	      	         �t�bhhK ��h��R�(KK��h�C46  �        �  F     G     C  /         �t�bhhK ��h��R�(KK��h�C,%          @      �              �t�bhhK ��h��R�(KK	��h�C$   �      w   �     �        �t�bhhK ��h��R�(KK��h�C %	        f   �            �t�bhhK ��h��R�(KK��h�C       ;      �           �t�bhhK ��h��R�(KK��h�C b   #   "   $   �   N        �t�bhhK ��h��R�(KK
��h�C(�  W     �   �  j      
        �t�bhhK ��h��R�(KK��h�CL%   .  �  g   ,            K      �                 �         �t�bhhK ��h��R�(KK��h�CT        /      	  i   �   7      �  0   �     �      D      V        �t�bhhK ��h��R�(KK��h�C4�     �   G   Q     y      �     �
        �t�bhhK ��h��R�(KK��h�CL   �     #        !     u  V   �  �   [  �   S     "        �t�bhhK ��h��R�(KK��h�CX         m         v         `     U   O              �              �t�bhhK ��h��R�(KK��h�CH         E  O     �  �      �
             �   A        �t�bhhK ��h��R�(KK��h�C0�           �   �   �      "           �t�bhhK ��h��R�(KK��h�C@      J   4        >      a      4      �   >         �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6            �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C0      =      �  "   �     $   k         �t�bhhK ��h��R�(KK��h�C�     �  r      �t�bhhK ��h��R�(KK��h�CH         $   k                 ,  %   �        
        �t�bhhK ��h��R�(KK
��h�C(      P   
  +  -      �        �t�bhhK ��h��R�(KK��h�CD
   3   6      ?      #   !   ;     l            
        �t�bhhK ��h��R�(KK��h�C0
      �   D  >      v     �  w         �t�bhhK ��h��R�(KK��h�Cv  	         �t�bhhK ��h��R�(KK��h�C
   �   |         �t�bhhK ��h��R�(KK��h�C,1   #      �   _  
   T  
  �	        �t�bhhK ��h��R�(KK��h�CD           <      �      -           o   G            �t�bhhK ��h��R�(KK��h�CT      6  +         <      �
             �     $   �               �t�bhhK ��h��R�(KK	��h�C$!      5  ,   	      	         �t�bhhK ��h��R�(KK��h�C,   (   -      
  *                 �t�bhhK ��h��R�(KK��h�CD      -     
  �  �  x     p      �  w  
   �         �t�bhhK ��h��R�(KK��h�Cd
                   �   �               ;      �   �        ~   �               �t�bhhK ��h��R�(KK	��h�C$      �     
  �      �      �t�bhhK ��h��R�(KK��h�C8      P      H            J  E      �        �t�bhhK ��h��R�(KK��h�C4�  �     w  �    a        "  �        �t�bhhK ��h��R�(KK��h�C@#   !      ,  '   
   �                             �t�bhhK ��h��R�(KK��h�CD     `     �t�bhhK ��h��R�(KK��h�C@�   >   %      ,        v     
   �                 �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK	��h�C$�  ;               �        �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�C<?                 	   �   	   I  	   /  	   s     �t�bhhK ��h��R�(KK��h�CT     [  
        �t�bhhK ��h��R�(KK��h�C      �     �t�bhhK ��h��R�(KK��h�Cp            �
     �   
   _      \     �        =      �              X                 �t�bhhK ��h��R�(KK��h�C       j      
            �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   6   {     �        �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CA  {     �     �t�bhhK ��h��R�(KK��h�C/      �      �t�bhhK ��h��R�(KK��h�C�  �  #        �t�bhhK ��h��R�(KK��h�C<      �   T                  C   q              �t�bhhK ��h��R�(KK��h�C   :     �     �t�bhhK ��h��R�(KK��h�C<T   A	  2   %   �            W                    �t�bhhK ��h��R�(KK��h�C<1   #      d   �   
   T  �     /   �              �t�bhhK ��h��R�(KK��h�C,   ?  �     �  �	        �        �t�bhhK ��h��R�(KK��h�CL   �         �     C      M     
      �     �  �            �t�bhhK ��h��R�(KK��h�C4�                    �      �           �t�bhhK ��h��R�(KK��h�CL�  v  �       q   .    V   2      e  C   h   H   B   3        �t�bhhK ��h��R�(KK��h�C01   #   
   3   6         �  Y  �         �t�bhhK ��h��R�(KK��h�CH   �        .   !
     A     n                �        �t�bhhK ��h��R�(KK��h�C\�  �	        �        "
              Y      Q      Q     Q      x        �t�bhhK ��h��R�(KK
��h�C(U   \        J   a      �        �t�bhhK ��h��R�(KK��h�CH�  L     %   ?  V      G     �               �  �        �t�bhhK ��h��R�(KK��h�C[                 �t�bhhK ��h��R�(KK��h�CH$   �           �                 #
  �            +      �t�bhhK ��h��R�(KK
��h�C(#   !   ?      
   e   �   F         �t�bhhK ��h��R�(KK��h�CL
   Z        )   R  q     �     �  �                        �t�bhhK ��h��R�(KK��h�C4!      s  
  '      S   
   q      F         �t�bhhK ��h��R�(KK��h�C,D      0            �     �         �t�bhhK ��h��R�(KK%��h�C��      v                  �  �     �           �  �   �        �  (   2   ;      �  �   �                     �        �t�bhhK ��h��R�(KK��h�Ct         F     �  L      $   �      
  �   +     9   �        P   �   �  *   U     
  �        �t�bhhK ��h��R�(KK��h�C0%   >   v   �   �     	     h          �t�bhhK ��h��R�(KK��h�C0!         �  "        	      	         �t�bhhK ��h��R�(KK��h�C*     �        �t�bhhK ��h��R�(KK
��h�C(d   �           l        /      �t�bhhK ��h��R�(KK��h�C       �   k  
           �t�bhhK ��h��R�(KK	��h�C$!  -  �  �  �      I         �t�bhhK ��h��R�(KK��h�C<            �        
   �  j      �  �         �t�bhhK ��h��R�(KK��h�C0      =      (  :   >     �   w         �t�bhhK ��h��R�(KK��h�CH   (   <   
   ,               
   %   �     )   
            �t�bhhK ��h��R�(KK��h�CD*      �           %     U   �     $
     $   k         �t�bhhK ��h��R�(KK��h�C   �     �      �t�bhhK ��h��R�(KK
��h�C(         f       d   d        �t�bhhK ��h��R�(KK��h�C<H  %
  +   �  4      �        3  �  �  �        �t�bhhK ��h��R�(KK��h�CH      �           �  �                  .      &
        �t�bhhK ��h��R�(KK
��h�C(�   �   7     `     �  �
        �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�CD   H  5   �  =     +      �  ]      �        �         �t�bhhK ��h��R�(KK��h�C q   �     	      	         �t�bhhK ��h��R�(KK	��h�C$K      �   �                 �t�bhhK ��h��R�(KK��h�C\?     �                �            2      0      �   �  �              �t�bhhK ��h��R�(KK	��h�C$  ?  '   
                  �t�bhhK ��h��R�(KK��h�CP   �	     ;      #     �  �        .   z      �      �          �t�bhhK ��h��R�(KK��h�C    0     	      	         �t�bhhK ��h��R�(KK��h�CL   P  -              w   (   s  �              8   S        �t�bhhK ��h��R�(KK��h�C,      �         s   o     �        �t�bhhK ��h��R�(KK	��h�C$�  (     �         ]        �t�bhhK ��h��R�(KK��h�C`   5   �  �     �  -      u     �                    �     8   E  �        �t�bhhK ��h��R�(KK��h�Ch�  �  �   �      ,               �         +         �   �     �        �   f        �t�bhhK ��h��R�(KK��h�C   9     �t�bhhK ��h��R�(KK��h�C4     '               4  '   H   i        �t�bhhK ��h��R�(KK��h�Cx     H  ?             �  �  t           �     �  
      h  N        2   >   w   v            �t�bhhK ��h��R�(KK��h�C�      �      �     �t�bhhK ��h��R�(KK��h�C,         6     �  j               �t�bhhK ��h��R�(KK��h�C       
   _      $   \     �t�bhhK ��h��R�(KK��h�C �  �   u     B   J        �t�bhhK ��h��R�(KK��h�C�   
   B   }          �t�bhhK ��h��R�(KK��h�C,�     �   '
        	      	         �t�bhhK ��h��R�(KK��h�C@�     "   >  �     �        �        �           �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C<�     `  &   �  �  "   2        �              �t�bhhK ��h��R�(KK	��h�C$�      
                  �t�bhhK ��h��R�(KK��h�C,�           	      	      	   K      �t�bhhK ��h��R�(KK��h�C4      J   �  �   &      �  ]      t         �t�bhhK ��h��R�(KK��h�C1        	         �t�bhhK ��h��R�(KK��h�C   =      �     �t�bhhK ��h��R�(KK��h�C0u      )   $  �   "   �        �        �t�bhhK ��h��R�(KK��h�C,4      �   ]   ,     	      	         �t�bhhK ��h��R�(KK��h�C,      �  0   [         :   W         �t�bhhK ��h��R�(KK��h�C8�     �  	      	      	   K   	   U  	   /     �t�bhhK ��h��R�(KK��h�CD*        E      �      �  �   l     #  �   �  �        �t�bhhK ��h��R�(KK��h�Cb     �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C,      �   �   
   B   [              �t�bhhK ��h��R�(KK��h�C      R          �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�CHH         )            T   2      �      �   j      �        �t�bhhK ��h��R�(KK��h�C<      5   �  <      �     E     �  j  /        �t�bhhK ��h��R�(KK
��h�C(!      �         	      	         �t�bhhK ��h��R�(KK��h�C,u  
     �      �   �              �t�bhhK ��h��R�(KK��h�CH�     (
             �	     �               �   l         �t�bhhK ��h��R�(KK��h�C<
   )
           .   0   <      �  m      �        �t�bhhK ��h��R�(KK
��h�C(�        �   -      H   �        �t�bhhK ��h��R�(KK��h�C^     b     �t�bhhK ��h��R�(KK��h�C�      4      �t�bhhK ��h��R�(KK��h�C M   �         �   D        �t�bhhK ��h��R�(KK��h�C0      =      �      	     �           �t�bhhK ��h��R�(KK	��h�C$�   &   �        !  �         �t�bhhK ��h��R�(KK��h�C  �     z      r      �t�bhhK ��h��R�(KK��h�C8M         g  �                 �   f        �t�bhhK ��h��R�(KK��h�C`     �      ;     �      ^           $           J   �  �   �     ,   *
     �t�bhhK ��h��R�(KK��h�C@   .                  �                          �t�bhhK ��h��R�(KK��h�Cb     �t�bhhK ��h��R�(KK	��h�C$      '                     �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�ClW  �  �     �         =      4      +      j   �     $   E      �   �      �   �           �t�bhhK ��h��R�(KK��h�C�  "   ~  y     �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C`�        �        �     6  �  !             �                  �        �t�bhhK ��h��R�(KK��h�C      	      	         �t�bhhK ��h��R�(KK��h�C          
   �  *        �t�bhhK ��h��R�(KK��h�C,   �  �    �  :   q     �        �t�bhhK ��h��R�(KK��h�Cp           �   �   J   0      r  '        L        &      U   +  "   @   �   @     �        �t�bhhK ��h��R�(KK
��h�C(  �   )   �         �          �t�bhhK ��h��R�(KK��h�C4      �      �      L   
                �t�bhhK ��h��R�(KK��h�C               �t�bhhK ��h��R�(KK	��h�C$�     �	  �      �     9     �t�bhhK ��h��R�(KK��h�C@O         
  Q           l        %   �  �  	     �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�Cd
   k  r     /      \  	     �              x   ^      �  �     �              �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�C{      �t�bhhK ��h��R�(KK��h�C0      !      k     �   �     �        �t�bhhK ��h��R�(KK��h�Ct   Y      O         �                     �        �                      �              �t�bhhK ��h��R�(KK	��h�C$[      �  M  	      	         �t�bhhK ��h��R�(KK��h�Ct     �t�bhhK ��h��R�(KK��h�C �      ,   �   "   �   n     �t�bhhK ��h��R�(KK��h�CH   y             V         0   �        
   B   }         �t�bhhK ��h��R�(KK��h�C+
  �         �t�bhhK ��h��R�(KK��h�C=  	         �t�bhhK ��h��R�(KK��h�C<�     t        �  +      �  +   �     "        �t�bhhK ��h��R�(KK!��h�C�                        D     �     $     (      �        *         a  #  �   �     �	  �   $           �t�bhhK ��h��R�(KK��h�C@*              {           
   8   ,
              �t�bhhK ��h��R�(KK��h�C      �  	         �t�bhhK ��h��R�(KK��h�C4      N   �   �   �      A  s   7   �        �t�bhhK ��h��R�(KK��h�C\   �  �  2   �   �           �   �         �     #   %     :  #   �        �t�bhhK ��h��R�(KK��h�C\   �
     8   -
  �  �  S     
   _      	     8   /         2              �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C@   �       S   
     b     <     �   ~            �t�bhhK ��h��R�(KK��h�C d  S  
      ?  �        �t�bhhK ��h��R�(KK��h�C<      )   0   �  
   �  B   .
     q             �t�bhhK ��h��R�(KK��h�C4�     �     �  �   *         �  �        �t�bhhK ��h��R�(KK��h�C,m      @     �                    �t�bhhK ��h��R�(KK��h�C      �  �      �t�bhhK ��h��R�(KK��h�C4        %     �  k  }     $   k         �t�bhhK ��h��R�(KK��h�C0!         �   �      K  	      	         �t�bhhK ��h��R�(KK	��h�C$D       �        �        �t�bhhK ��h��R�(KK��h�CZ         Z         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK	��h�C$      �      	      	         �t�bhhK ��h��R�(KK��h�C �   E      P     �         �t�bhhK ��h��R�(KK1��h�C�   �              _  C   :        &  
   �                 '   �        �   R     w     �  H          �         �     �     �         /
                 �t�bhhK ��h��R�(KK��h�C     	      	         �t�bhhK ��h��R�(KK��h�C0   >  �  0
     �   �                 �t�bhhK ��h��R�(KK��h�CX�     �           $   k   �  �      +         5   �         $   n         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CL-                  �                 k  t                 �t�bhhK ��h��R�(KK��h�CW           �t�bhhK ��h��R�(KK��h�C4      �           1     �     $	        �t�bhhK ��h��R�(KK��h�C5         1  r      �t�bhhK ��h��R�(KK��h�C`   �   '             �      f                          �        �        �t�bhhK ��h��R�(KK��h�CH      -   a   ;         �   �               ,              �t�bhhK ��h��R�(KK��h�CD�      ;     l            �     ,                     �t�bhhK ��h��R�(KK��h�C'  �  �         �t�bhhK ��h��R�(KK��h�C,8   4         %  �      (   �         �t�bhhK ��h��R�(KK��h�CXW   �  �      
   �   �     �   �      s  �   ^   �     '   
   �            �t�bhhK ��h��R�(KK��h�CD   <      �         
   c  �	           v   (          �t�bhhK ��h��R�(KK��h�Che   �   �   �        %   8     �  /      V        '      .   �     �   5             �t�bhhK ��h��R�(KK��h�C;      0   �            �t�bhhK ��h��R�(KK��h�C !         �     	         �t�bhhK ��h��R�(KK��h�C@#   !            C        e   ?      
      F         �t�bhhK ��h��R�(KK	��h�C$E     F  ,   	      	         �t�bhhK ��h��R�(KK��h�C0      �  ]  g                        �t�bhhK ��h��R�(KK	��h�C$   >      =         �        �t�bhhK ��h��R�(KK��h�C\   (   G           �   S   Q        j   4   �   �     8   L        Z        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CX%   �  k     �   �  �   n      %         �        �   n   
   A           �t�bhhK ��h��R�(KK��h�Ch         1
     L   G   �     �         �   
      L   &      �   �     [  $   L         �t�bhhK ��h��R�(KK��h�C@g  
   �                        E  "        .     �t�bhhK ��h��R�(KK��h�C
                  �t�bhhK ��h��R�(KK��h�CXH  �      �                    �     9      �            �   '        �t�bhhK ��h��R�(KK��h�Cx/      �     /   :     �     0   )                    �  H   /   J  C      �          �         �t�bhhK ��h��R�(KK��h�C ,     N   A  #  �         �t�bhhK ��h��R�(KK��h�Cv     -               �t�bhhK ��h��R�(KK��h�C0   �   !  <            /   
            �t�bhhK ��h��R�(KK��h�C�     	         �t�bhhK ��h��R�(KK��h�C\     &  �	  T   s        l   �           }     &  �      �              �t�bhhK ��h��R�(KK��h�C`     �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C   �  �  �         �t�bhhK ��h��R�(KK��h�CT2
             �     `   A   b     $   |        �  /  �          �t�bhhK ��h��R�(KK	��h�C$                           �t�bhhK ��h��R�(KK��h�CH
      '      S   �
     �            �     !      a        �t�bhhK ��h��R�(KK
��h�C(�        �  �      h  |        �t�bhhK ��h��R�(KK��h�C   m     r        �t�bhhK ��h��R�(KK��h�C �   �     U	     �	        �t�bhhK ��h��R�(KK	��h�C$   �  
   �     �  *        �t�bhhK ��h��R�(KK��h�C8!      B        2     �  '   
   �   F         �t�bhhK ��h��R�(KK
��h�C(T         K        "   U        �t�bhhK ��h��R�(KK	��h�C$"    �      :  �   �        �t�bhhK ��h��R�(KK��h�Ct      J   "     �   +  &      U         �  c   �      W       *         6     �  
   �         �t�bhhK ��h��R�(KK
��h�C(   =      o     	      	         �t�bhhK ��h��R�(KK��h�C<      �     �t�bhhK ��h��R�(KK��h�CE      4      �        �t�bhhK ��h��R�(KK��h�CL
   �  F   '            ,   �   V         z   ,   
   �   �         �t�bhhK ��h��R�(KK��h�CP                     q   �
          �          �          �t�bhhK ��h��R�(KK	��h�C$�  �         	      	         �t�bhhK ��h��R�(KK��h�C4b   $   �      �  �  �   �        �         �t�bhhK ��h��R�(KK��h�CX)	  h   �   �     �  �   $     �   /	  �   �  /      �   �  d   A   K        �t�bhhK ��h��R�(KK
��h�C(           �   �               �t�bhhK ��h��R�(KK��h�CTB  �   �   s   B   �  �                     �                       �t�bhhK ��h��R�(KK!��h�C�                  V  �            �      �      N      >     <                  .   �     �  "            �t�bhhK ��h��R�(KK��h�C8   �       &      �   D     �      �        �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�CT�   �  �     .            �           e                           �t�bhhK ��h��R�(KK��h�C(  �   �         �t�bhhK ��h��R�(KK��h�C          	      	         �t�bhhK ��h��R�(KK��h�C*   &   �   v   �  r      �t�bhhK ��h��R�(KK	��h�C$V   ?      )   �     &        �t�bhhK ��h��R�(KK	��h�C$1   #   
   3   6      m         �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�C  b     �t�bhhK ��h��R�(KK��h�C �	        	      	         �t�bhhK ��h��R�(KK	��h�C$�       �              3
     �t�bhhK ��h��R�(KK��h�C0�  "        R     /   9     7         �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�C   (          �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CL
      �  2   
   ,      �         �         �       ,         �t�bhhK ��h��R�(KK��h�C0G      �   �  >      v     �  w         �t�bhhK ��h��R�(KK��h�C8   4  '   )   �     �  �     �	              �t�bhhK ��h��R�(KK��h�CDM            �                    
   �  N  j   �      �t�bhhK ��h��R�(KK��h�C   �         �         �t�bhhK ��h��R�(KK��h�C\      J   a   �         �                   <   "      "   q   �  �        �t�bhhK ��h��R�(KK��h�CT�   �      �     �  :                                             �t�bhhK ��h��R�(KK��h�C0         �     
  Y  �  �  7         �t�bhhK ��h��R�(KK��h�C@   �       �  r  
         �        �           �t�bhhK ��h��R�(KK��h�Cl
        %     �        K              �	  �     '   !      x      8     1  �         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CX   �     /   9   -  (      !   
   T     �        "                     �t�bhhK ��h��R�(KK��h�CH*      �     P     W  �     5  8   t     �   �           �t�bhhK ��h��R�(KK��h�C #   !   '   
   �            �t�bhhK ��h��R�(KK��h�C@   �           P  *         
  �   �               �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C4N  c   I  
   �  F      �                �t�bhhK ��h��R�(KK��h�C4g   �                    M   c   �        �t�bhhK ��h��R�(KK��h�C@
   %   .     '   �   �	     
      [  -   �   +        �t�bhhK ��h��R�(KK��h�C         �   �      �t�bhhK ��h��R�(KK��h�C   }          �t�bhhK ��h��R�(KK��h�C0   @   '   H     
   B   �     4        �t�bhhK ��h��R�(KK��h�C0�  �  �      
   ,            K         �t�bhhK ��h��R�(KK��h�C:   �      �     �t�bhhK ��h��R�(KK��h�CX      :  "   9          �             P   n   G                   �t�bhhK ��h��R�(KK��h�CL-   `         a   ;      �   R      %            �      +         �t�bhhK ��h��R�(KK7��h�C�                        �   "   �              "     ^  @     �  �     �  9     W        �        M     �               �      �     �  �   �     �	  �      �     �        �t�bhhK ��h��R�(KK ��h�C�        �  �     i  7      0   <   "      2     �     m      .         �             �              �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�CLV   �      +      �        �            �        �  4
        �t�bhhK ��h��R�(KK��h�C4T   �	        ,  �  �   �     `            �t�bhhK ��h��R�(KK��h�CL          
   8   �        
          J   a      +         �t�bhhK ��h��R�(KK��h�CH   .   h   @        V       �        h         �        �t�bhhK ��h��R�(KK��h�C,      �     D  �     h   �         �t�bhhK ��h��R�(KK��h�C4      -      8   �   �      M               �t�bhhK ��h��R�(KK��h�C,      �     ;  a        �         �t�bhhK ��h��R�(KK��h�CT   �                     �      
        �     "      �           �t�bhhK ��h��R�(KK��h�C0   s  �  (         �   9   �           �t�bhhK ��h��R�(KK��h�C      O  �     �t�bhhK ��h��R�(KK��h�C    �     z  s   7         �t�bhhK ��h��R�(KK	��h�C$      -   P   T  ^   &        �t�bhhK ��h��R�(KK��h�CX*      a  g      n         �                  �            �   �         �t�bhhK ��h��R�(KK��h�C 1   #       F     �        �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�Ct      �     �t�bhhK ��h��R�(KK��h�C!      �           �t�bhhK ��h��R�(KK��h�Ch	       p      u      �t�bhhK ��h��R�(KK	��h�C$!      �     	      	         �t�bhhK ��h��R�(KK	��h�C$     e  �   
   8           �t�bhhK ��h��R�(KK��h�C1   #             �t�bhhK ��h��R�(KK��h�C(                 �t�bhhK ��h��R�(KK��h�CHT         �      b           ;      5     �   �   �        �t�bhhK ��h��R�(KK��h�C 1   #          }     o      �t�bhhK ��h��R�(KK��h�C        �     �t�bhhK ��h��R�(KK��h�C-     .  /  *     �t�bhhK ��h��R�(KK��h�CP            %   b  z           2   J   *  !	                    �t�bhhK ��h��R�(KK��h�C0�      N      .   �      ,              �t�bhhK ��h��R�(KK��h�C\   M   C      �                              �       0      �           �t�bhhK ��h��R�(KK��h�C4%   ^     �      N      �      B           �t�bhhK ��h��R�(KK��h�C<�          N      .   L  �     �     d        �t�bhhK ��h��R�(KK��h�C�  h         �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C<�     �     �     V  �     �  7     �        �t�bhhK ��h��R�(KK��h�C4%   �        �  
   `   b  :   �     y     �t�bhhK ��h��R�(KK��h�CX      �     �  G      �     8   E     b           �  G   R  �        �t�bhhK ��h��R�(KK��h�C,#   !      v  w  (      "   W         �t�bhhK ��h��R�(KK	��h�C$
   f   [  �  )   #  �        �t�bhhK ��h��R�(KK��h�CD`   �     0      n   �     8   5
     `   6
     b        �t�bhhK ��h��R�(KK��h�C@�     0     m  G   W   �  s   �   �      "  �        �t�be(hhK ��h��R�(KK��h�C<q   c              �   ,  *   %                  �t�bhhK ��h��R�(KK��h�CH   �   '   �  
            B   �
  �   j        �  q        �t�bhhK ��h��R�(KK��h�Ch  d     �t�bhhK ��h��R�(KK��h�C,�  �      )         �     �         �t�bhhK ��h��R�(KK��h�C4�   3     %   l         ;      �            �t�bhhK ��h��R�(KK
��h�C(   	      	      	   K   	   U     �t�bhhK ��h��R�(KK��h�Cx      �   F                 ;      �  �   h      �        �        .   
      N        y        �t�bhhK ��h��R�(KK��h�Cd   �  �     .   %   �   m     I         �        �   x     \      ,   K  �        �t�bhhK ��h��R�(KK��h�C�  d  2   �           �t�bhhK ��h��R�(KK��h�C"   �     :           �t�bhhK ��h��R�(KK	��h�C$   ?      
   �              �t�bhhK ��h��R�(KK��h�CZ            �t�bhhK ��h��R�(KK��h�C0         k         (      �  �        �t�bhhK ��h��R�(KK
��h�C(U   8   �  �   *                  �t�bhhK ��h��R�(KK��h�C0      (      #   !   
   3   6   �        �t�bhhK ��h��R�(KK��h�CD   �         �     (   D   o  �      �   �  �   �          �t�bhhK ��h��R�(KK��h�C�     �   o            �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK
��h�C(      -   �         �          �t�bhhK ��h��R�(KK��h�CI      ;      �     �t�bhhK ��h��R�(KK��h�C0   �   S   �  �        �              �t�bhhK ��h��R�(KK��h�C!         	         �t�bhhK ��h��R�(KK��h�CT�  !      �      ,               ?      
   3   6   �        �         �t�bhhK ��h��R�(KK
��h�C()      �     �  C               �t�bhhK ��h��R�(KK
��h�C(
   ]   1                 :      �t�bhhK ��h��R�(KK��h�C@         .               N      0   `   %  (        �t�bhhK ��h��R�(KK��h�C@      �   L     �   w   -  4     e  �  �            �t�bhhK ��h��R�(KK	��h�C$7
          �             �t�bhhK ��h��R�(KK��h�C       P   �               �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C<*      ]     n   >      -   v   8
                 �t�bhhK ��h��R�(KK	��h�C$                 S   Q      �t�bhhK ��h��R�(KK��h�CD%      �     -   
         �  (   2         L   V         �t�bhhK ��h��R�(KK��h�C�  �              �t�bhhK ��h��R�(KK��h�C �     -   �   �   �         �t�bhhK ��h��R�(KK��h�C�  �                �t�bhhK ��h��R�(KK��h�C    8   �      �  �  {     �t�bhhK ��h��R�(KK��h�CH   d   \     (  B  �   &      d  �  $   N       �        �t�bhhK ��h��R�(KK��h�C@      J   �      �  �   &      M   �   �      �        �t�bhhK ��h��R�(KK��h�C   v     �t�bhhK ��h��R�(KK��h�Cd<  &   �   f           x         �         g     �      �         >     �        �t�bhhK ��h��R�(KK��h�C�  �      �     �t�bhhK ��h��R�(KK��h�C@   1  �  
   `   �      .      �          A        �t�bhhK ��h��R�(KK��h�C|   +   
   	  �      �  �   [  �          "     S              �     o   j   �  �     �  �        �t�bhhK ��h��R�(KK��h�C\!        (      
   X            g              "   �                     �t�bhhK ��h��R�(KK��h�C�	  �      �     i     �t�bhhK ��h��R�(KK��h�C>     �        �t�bhhK ��h��R�(KK��h�CH   e   '   )   9
  �  �           V   `     z   ,   �         �t�bhhK ��h��R�(KK��h�C8      =      +  4   
        �   �           �t�bhhK ��h��R�(KK	��h�C$,    
   ,      
            �t�bhhK ��h��R�(KK��h�CH                  �  �      
        &      U   �        �t�bhhK ��h��R�(KK��h�CZ      �               �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�CP        �       �      �     �     �  �      �     �        �t�bhhK ��h��R�(KK��h�Cp�  :
  �	  }     @   
         �     �           �             A        4     @         �t�bhhK ��h��R�(KK��h�C,#   !      v  '   
   3   6            �t�bhhK ��h��R�(KK��h�CD                 �  �        V   �                �t�bhhK ��h��R�(KK��h�C �     �   "   �  	         �t�bhhK ��h��R�(KK��h�C<      ~         �    n  B     %   �           �t�bhhK ��h��R�(KK��h�Ct         F     �  L      $   �      
  �   +     9   �        P   �   �  *   U     
  �        �t�bhhK ��h��R�(KK��h�C         ,         �t�bhhK ��h��R�(KK��h�C         �  �  r      �t�bhhK ��h��R�(KK��h�C<\        ?         <         �	                 �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK	��h�C$#   !   ?      
      F         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CD   
  +  5                                        �t�bhhK ��h��R�(KK
��h�C(!         Y     	      	         �t�bhhK ��h��R�(KK	��h�C$   '   
   B   �     4        �t�bhhK ��h��R�(KK��h�C4*      /   \  =  x         	      	         �t�bhhK ��h��R�(KK��h�C�     �  
   �      �t�bhhK ��h��R�(KK��h�CH   �   �   '   �
  e     �  M     �     �         h        �t�bhhK ��h��R�(KK��h�C@"   �     �     C      a   
   C   �         2        �t�bhhK ��h��R�(KK��h�C,      -   U      �     h          �t�bhhK ��h��R�(KK��h�C8E   &   r  �   �  h   �   �   :                  �t�bhhK ��h��R�(KK��h�C`"   �  '
     R         P   <      !      �              \      �      �        �t�bhhK ��h��R�(KK��h�C    �  �     B   �        �t�bhhK ��h��R�(KK
��h�C(-   �   ]   ,   O   -              �t�bhhK ��h��R�(KK��h�C@#   !   (      
   3   6         
   @     �  F         �t�bhhK ��h��R�(KK
��h�C(   '   �      (     �   S        �t�bhhK ��h��R�(KK��h�C0#   !      �  �  '   
   3   6   �         �t�bhhK ��h��R�(KK��h�C <  �  -      �   5        �t�bhhK ��h��R�(KK!��h�C�]   �     �        /   9   9  7               '  :   ]         �  �  0  s   p     r  C   
   �               �t�bhhK ��h��R�(KK��h�C,f     g  )                      �t�bhhK ��h��R�(KK	��h�C$;
  <
              �        �t�bhhK ��h��R�(KK��h�C,g   �   �  �   ;  �   =
              �t�bhhK ��h��R�(KK��h�C<G   �        0   <      �   �  �                �t�bhhK ��h��R�(KK��h�C �      (     +      �     �t�bhhK ��h��R�(KK��h�C8      u     !        �  $   0              �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK!��h�C�   �  ?   D  �  !   
   �   �   }                 {      �      �      p      �           G  w     x        �t�bhhK ��h��R�(KK��h�C
  v  	      	         �t�bhhK ��h��R�(KK��h�C         m  W           �t�bhhK ��h��R�(KK��h�C Z      �         �        �t�bhhK ��h��R�(KK��h�CP{   9   �     3           �  j      �           d   �           �t�bhhK ��h��R�(KK��h�C      �  W  7      �t�bhhK ��h��R�(KK��h�C0
   %   �  �        J	     D  ,         �t�bhhK ��h��R�(KK��h�C          �     �t�bhhK ��h��R�(KK��h�CX      0   �   �     �	  &      a   ;      �            N   �     W         �t�bhhK ��h��R�(KK��h�CZ                     �t�bhhK ��h��R�(KK��h�C,   '           +                  �t�bhhK ��h��R�(KK��h�C0   �  �     
   �           �         �t�bhhK ��h��R�(KK��h�C4            �  A      �   �  9         �t�bhhK ��h��R�(KK��h�C 1   #       4              �t�bhhK ��h��R�(KK��h�Cd
   3   6         p   ?      !      \      �            �          �              �t�bhhK ��h��R�(KK��h�CX     �      ;     �      ^     J   z   "   9  �   �  �  �     �        �t�bhhK ��h��R�(KK��h�Cu      O     �t�bhhK ��h��R�(KK��h�CL      �                i     >        G   �  �           �t�bhhK ��h��R�(KK��h�CL�      �      -   ;      A     K     �      �      ~            �t�bhhK ��h��R�(KK��h�C �     c  X  �  �         �t�bhhK ��h��R�(KK��h�CT      M   +         �        
   _      �              G  '        �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C,      �      �         �            �t�bhhK ��h��R�(KK��h�C1   #       �  �         �t�bhhK ��h��R�(KK��h�C8      \  �  "  )            5   �  ^        �t�bhhK ��h��R�(KK��h�Ch
   3   6      ?      !      �         0   <               V     +      m               �t�bhhK ��h��R�(KK��h�C�      L   "           �t�bhhK ��h��R�(KK��h�C`1   
   3   6         �  R   #     v           &   D  �  �  G   �      (        �t�bhhK ��h��R�(KK��h�Ch*      /   �     �      �   ;      M            J   �  H  '        M   �      D         �t�bhhK ��h��R�(KK��h�Cp            y      W           �  F                +         0                        �t�bhhK ��h��R�(KK	��h�C$�  �         N              �t�bhhK ��h��R�(KK��h�C*  �      �t�bhhK ��h��R�(KK��h�C4�  ;  &   3	  4     s   	  &               �t�bhhK ��h��R�(KK
��h�C(4            5   4               �t�bhhK ��h��R�(KK��h�C82      =         �  h      �  5  y  �        �t�bhhK ��h��R�(KK
��h�C(2      )   �   �   >
  
   �        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK	��h�C$	   �  	   �  	   �  	   �     �t�bhhK ��h��R�(KK��h�C4   w  (            �   *        �        �t�bhhK ��h��R�(KK��h�C,1           �  ,   	      	         �t�bhhK ��h��R�(KK��h�CD�  �       B       �             �               �t�bhhK ��h��R�(KK��h�Cj     �t�bhhK ��h��R�(KK��h�C <         	      	         �t�bhhK ��h��R�(KK��h�CX�      �   q     �      �   o   w   �   5  �     E   �   ^   �   �           �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C+  5  	      	         �t�bhhK ��h��R�(KK��h�C4      -  /      �      �  	      	         �t�bhhK ��h��R�(KK��h�C<�   �     �      I   p        q     N  7         �t�bhhK ��h��R�(KK��h�Cx      �      +      G        >      F        v                     y         �         k        �t�bhhK ��h��R�(KK	��h�C$�  �      �     9  j   �     �t�bhhK ��h��R�(KK��h�C�  4      �t�bhhK ��h��R�(KK��h�C,D   (   g                          �t�bhhK ��h��R�(KK��h�C`Z        �  V         R  �     �  �     �         z      2     B   a        �t�bhhK ��h��R�(KK��h�C;	  M     �t�bhhK ��h��R�(KK
��h�C(�     ,     .      �   q         �t�bhhK ��h��R�(KK��h�Ct�   �   )   x      �     l      �   :   M              �            �      �   �     R           �t�bhhK ��h��R�(KK��h�C�     	      	         �t�bhhK ��h��R�(KK��h�C@      5   �  <      �        �     �  j  /        �t�bhhK ��h��R�(KK
��h�C(      -   i     ?
     �        �t�bhhK ��h��R�(KK��h�C@:    c      e     �     l        �              �t�bhhK ��h��R�(KK��h�CD   `             �        .        q     k        �t�bhhK ��h��R�(KK
��h�C(     a     a  	      	         �t�bhhK ��h��R�(KK��h�C8�  �   x            �   "          �        �t�bhhK ��h��R�(KK��h�Cp                     �   ]  �         7      
     &      -   F  +      t   
   $   �        �t�bhhK ��h��R�(KK��h�C,f   [  o	  )   �  
   A   N  }         �t�bhhK ��h��R�(KK��h�C,9   �   _     �     N   <          �t�bhhK ��h��R�(KK��h�CL      5   <      [      $   �  �         �      n	  "           �t�bhhK ��h��R�(KK��h�C`            �   ]   �   O            8   ,   �   �      �      u	                 �t�bhhK ��h��R�(KK��h�C0�     j                 �  �        �t�bhhK ��h��R�(KK��h�C@#   !      �     C  3  ?      
   3   6      [        �t�bhhK ��h��R�(KK
��h�C(      A  M   c      �           �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�CT      �           �  h     &      �     c   #  "   $   �            �t�bhhK ��h��R�(KK��h�C@\   �        �  >   �    
   \   �  `   �   Y        �t�bhhK ��h��R�(KK��h�C4      z   �  i   �  _        j   4         �t�bhhK ��h��R�(KK��h�C06  �    
   �  �           @         �t�bhhK ��h��R�(KK��h�Ch            i  
            k               M     
   $   |  "   t      �           �t�bhhK ��h��R�(KK
��h�C(E              J     	         �t�bhhK ��h��R�(KK��h�C      ~        �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�C"   >  �      +         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C	     �        �t�bhhK ��h��R�(KK��h�C8      �              1     �     A        �t�bhhK ��h��R�(KK��h�C4,  R        |      �  V         �        �t�bhhK ��h��R�(KK��h�CI      ;      8        �t�bhhK ��h��R�(KK��h�C8   	      	      	   K   	     	   �   	   �     �t�bhhK ��h��R�(KK��h�CU   C  �      �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK
��h�C(2   �      �         G  E         �t�bhhK ��h��R�(KK��h�C1   #       �        �t�bhhK ��h��R�(KK
��h�C(.  G   �	     �   �     �        �t�bhhK ��h��R�(KK��h�C �     �                 �t�bhhK ��h��R�(KK	��h�C$m  -  
   �     �  y        �t�bhhK ��h��R�(KK��h�C@      �         �       �   
        l  w        �t�bhhK ��h��R�(KK��h�C4     C        �t�bhhK ��h��R�(KK��h�C\   �              .         %     �           )   U         $   /        �t�bhhK ��h��R�(KK
��h�C(      '      C  �              �t�bhhK ��h��R�(KK��h�CL      )   "   >                                         �t�bhhK ��h��R�(KK��h�C@�   0  s   l      �          3        �           �t�bhhK ��h��R�(KK��h�CX      �   �	       5         �   %   �         �     E  "   �           �t�bhhK ��h��R�(KK��h�C`      J      8   /   &   0                       &      
  L         Z        �t�bhhK ��h��R�(KK��h�Cu  �      �t�bhhK ��h��R�(KK��h�C�  �            �t�bhhK ��h��R�(KK	��h�C$�   &      w   �     @
        �t�bhhK ��h��R�(KK��h�C0      P   �   =     e   ^      _         �t�bhhK ��h��R�(KK��h�CDb  �
     b   #      (  s     "              <        �t�bhhK ��h��R�(KK��h�CD   ]   �         �      8   A
  �     �      q            �t�bhhK ��h��R�(KK��h�Cd/      O  X        ,            :  ,            �        �   �  �	     �        �t�bhhK ��h��R�(KK��h�C8
     �t�bhhK ��h��R�(KK��h�C,     �    �        !  n         �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C H      �   �     u         �t�bhhK ��h��R�(KK��h�C4     �     �           B
              �t�bhhK ��h��R�(KK��h�CD      �   .  "        $
              k               �t�bhhK ��h��R�(KK
��h�C(   f   3  '   -   A   �	  "        �t�bhhK ��h��R�(KK��h�C`   �     X   '   �         @   J  �     C
  l              �     �   B	        �t�bhhK ��h��R�(KK��h�C8�  o  �   7      '  c   �     I               �t�bhhK ��h��R�(KK��h�C4   (   8  :   2            g   �        �t�bhhK ��h��R�(KK��h�Cp�   &   �                             �   �   %               
   �     \   2      �         �t�bhhK ��h��R�(KK
��h�C(        �   '   B   �           �t�bhhK ��h��R�(KK��h�C=  �   Y  	         �t�bhhK ��h��R�(KK��h�C,"           e  +         �        �t�bhhK ��h��R�(KK��h�C      �             �t�bhhK ��h��R�(KK��h�C<   �      �           �      �      �   �	        �t�bhhK ��h��R�(KK��h�C0   �      B   �     d   �   
   #        �t�bhhK ��h��R�(KK��h�Cn     %     �t�bhhK ��h��R�(KK��h�C4I      ~      G        >   5  q   7        �t�bhhK ��h��R�(KK��h�CD   �  �     Q        (     �     <  �  9            �t�bhhK ��h��R�(KK��h�C0   e   '   �     0	        �  `        �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C �  	      	      	   K      �t�bhhK ��h��R�(KK��h�C      �        �t�bhhK ��h��R�(KK	��h�C$�	        F     0	  u         �t�bhhK ��h��R�(KK��h�C<!      �      �      @  ?      
   3   6   �        �t�bhhK ��h��R�(KK��h�C
   ,             �t�bhhK ��h��R�(KK��h�C0     �t�bhhK ��h��R�(KK��h�C �     c  X  �  �         �t�bhhK ��h��R�(KK��h�Ca     n     �     �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�CP*               &      \  t      �     
   D
  V         l        �t�bhhK ��h��R�(KK��h�CH      �  	      	      	   K   	   �   	   U  	   /  	   �     �t�bhhK ��h��R�(KK��h�C41   #      �     3   �  �        �         �t�bhhK ��h��R�(KK��h�C0       
   \   �  �       Z        �t�bhhK ��h��R�(KK��h�C0�      �                  D  �        �t�bhhK ��h��R�(KK	��h�C$�  �   
        
   �        �t�bhhK ��h��R�(KK
��h�C(   =            	      	         �t�bhhK ��h��R�(KK��h�C8*      �      �      �     g  �   `   �        �t�bhhK ��h��R�(KK��h�ChY      O         �   k            �     �     ?	           %      E
  C              �t�bhhK ��h��R�(KK��h�C<)   T   >   �          �        ]      +         �t�bhhK ��h��R�(KK��h�C0
            Z     �     �           �t�bhhK ��h��R�(KK��h�CL      �            �     "  �      �            �   �         �t�bhhK ��h��R�(KK��h�C\      N   �      6  C   ,                       �      �  L      u        �t�bhhK ��h��R�(KK��h�C�     T  	         �t�bhhK ��h��R�(KK��h�C<p      F
                 �     �               �t�bhhK ��h��R�(KK��h�C0�     �  \  �       %      m         �t�bhhK ��h��R�(KK��h�Ca   �  �    �         �t�bhhK ��h��R�(KK��h�C!         	         �t�bhhK ��h��R�(KK��h�CD      ;      �   �        
        �   
   $           �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C T      �  Q     +         �t�bhhK ��h��R�(KK��h�C4Z   Z     ,                              �t�bhhK ��h��R�(KK
��h�C(2   �      w        �          �t�bhhK ��h��R�(KK&��h�C�         `                  +                  O         
  Q         �   �   �   d  4         �	  �   �     Y      O         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C �   L        G   t         �t�bhhK ��h��R�(KK��h�C8     �     ;     �     �  /      �        �t�bhhK ��h��R�(KK��h�C|      <  R      �t�bhhK ��h��R�(KK��h�C    �      �  G   W         �t�bhhK ��h��R�(KK��h�CZ      �               �t�bhhK ��h��R�(KK��h�C4*   D      r     C  =  G         �        �t�bhhK ��h��R�(KK��h�Ch            �        \        $         9   �      7         0                    �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�CT         a        �  �     �           
   &  F         2        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C\   &   )  +      �	           �           �            c	     v            �t�bhhK ��h��R�(KK��h�C0!        �           Z              �t�bhhK ��h��R�(KK��h�C         	         �t�bhhK ��h��R�(KK��h�C@      ,        
  i   �   �   >      =      4         �t�bhhK ��h��R�(KK��h�C,      
   _         	      	         �t�bhhK ��h��R�(KK��h�C8   2     C         p   
        �   �  p      �t�bhhK ��h��R�(KK��h�CH      w   s        �   c   �  o     �     �               �t�bhhK ��h��R�(KK��h�C�        	         �t�bhhK ��h��R�(KK��h�CO             �t�bhhK ��h��R�(KK
��h�C(N        	      	      	   K      �t�bhhK ��h��R�(KK
��h�C("   I     '      �     �        �t�bhhK ��h��R�(KK��h�Ch  ?     �t�bhhK ��h��R�(KK��h�C�   �  2   �           �t�bhhK ��h��R�(KK
��h�C(   =      c  �  	      	         �t�bhhK ��h��R�(KK��h�CL      =      4      �      4      �  
     ^   �   �           �t�bhhK ��h��R�(KK	��h�C$�        �  i   h          �t�bhhK ��h��R�(KK	��h�C$      �  �	     .   �         �t�bhhK ��h��R�(KK��h�C8   .                  "                    �t�bhhK ��h��R�(KK��h�C!            �t�bhhK ��h��R�(KK��h�CL      5      &        r  '     �     >   D  
     &        �t�bhhK ��h��R�(KK��h�Cp               �   +      �  ;   [           ?      !        q	     &   M      
   �        �t�bhhK ��h��R�(KK��h�C
         Z         �t�bhhK ��h��R�(KK��h�C@!      c  	   K   	   �   	   I  	   U  	   /  	   s     �t�bhhK ��h��R�(KK��h�C8�     �  �   �             �  H   �         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK	��h�C$   �  �	  �  
   �            �t�bhhK ��h��R�(KK��h�C    R            |        �t�bhhK ��h��R�(KK��h�C0            i      .   %      �        �t�bhhK ��h��R�(KK��h�C<      �   +                  {         �        �t�bhhK ��h��R�(KK��h�C4�   I              P       �   $        �t�bhhK ��h��R�(KK���      h�C,.  M     �   �     �     ^        �t�bhhK ��h��R�(KK��h�C4   <  '      �     �     .     	        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�CD      )        x   �  A   �        .   �      G
        �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C         	         �t�bhhK ��h��R�(KK��h�C<         �         0      +  ^   =  b  *        �t�bhhK ��h��R�(KK
��h�C(     �        j   �            �t�bhhK ��h��R�(KK��h�C0	    
   T     �        h   �        �t�bhhK ��h��R�(KK��h�C �  �   (   �   7  �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C4�  �            �  h         R     7     �t�bhhK ��h��R�(KK��h�C,   �  �   (      <         1        �t�bhhK ��h��R�(KK��h�C!            �t�bhhK ��h��R�(KK��h�C�   -     �t�bhhK ��h��R�(KK��h�C4I  (      
   �	  F      :   �              �t�bhhK ��h��R�(KK��h�C8   X   '   P  �     i        h  �   �        �t�bhhK ��h��R�(KK��h�C{     �     �t�bhhK ��h��R�(KK��h�C�        a        �t�bhhK ��h��R�(KK
��h�C(|      �   �  q        �        �t�bhhK ��h��R�(KK
��h�C(   5      v      .  "           �t�bhhK ��h��R�(KK��h�C�  	      	         �t�bhhK ��h��R�(KK��h�C`     �t�bhhK ��h��R�(KK��h�Cp      u      �t�bhhK ��h��R�(KK��h�CX*         �         �     +            u        +      �              �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C1   #       �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CT   �   E     u      .      �      -       �             �        �t�bhhK ��h��R�(KK��h�C8�   =        �  �  �     �  �  �           �t�bhhK ��h��R�(KK��h�C<   X   '   �               A   s     B   �        �t�bhhK ��h��R�(KK
��h�C(-            0   4               �t�bhhK ��h��R�(KK��h�CL      5       
            &      �   D  �   +     �        �t�bhhK ��h��R�(KK��h�C4      	        �         G              �t�bhhK ��h��R�(KK��h�C<b                    Y         	      	         �t�bhhK ��h��R�(KK��h�C�     �         �t�bhhK ��h��R�(KK��h�C0�   >      �      L   G   �             �t�bhhK ��h��R�(KK��h�C4     T  C   :   m         �             �t�bhhK ��h��R�(KK��h�C0-         %     8           �        �t�bhhK ��h��R�(KK��h�CP�   (      b      $        %  d                                �t�bhhK ��h��R�(KK��h�C<y   �     s   l      �        �     �           �t�bhhK ��h��R�(KK��h�C   1         �t�bhhK ��h��R�(KK��h�CD      )        �                                   �t�bhhK ��h��R�(KK��h�C   $   n      �	     �t�bhhK ��h��R�(KK��h�Cv  	      	         �t�bhhK ��h��R�(KK��h�C�	       �  �   _     �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CD�    x  �          ^  @     �  �  �   �            �t�bhhK ��h��R�(KK��h�C�   �     �t�bhhK ��h��R�(KK��h�CTa  8   �   ~       "        =  �  p     +               "        �t�bhhK ��h��R�(KK��h�CD#   !         �          �   '   
   }  �  �  F         �t�bhhK ��h��R�(KK��h�C=      �      �t�bhhK ��h��R�(KK
��h�C(!      X        	      	         �t�bhhK ��h��R�(KK��h�C@   �   l         �              �     �  �         �t�bhhK ��h��R�(KK��h�C8D      ;      a   �      �  �   8  g           �t�bhhK ��h��R�(KK��h�C,$   �      v   c   U     8           �t�bhhK ��h��R�(KK��h�CD         �     *   D      �              �   �        �t�bhhK ��h��R�(KK��h�C1   #   
   �   F         �t�bhhK ��h��R�(KK��h�C 1        	      	         �t�bhhK ��h��R�(KK��h�C@
   3   6   �	  ?      !      %   $  .     3            �t�bhhK ��h��R�(KK��h�CD      �           S   Q   i         $           u     �t�bhhK ��h��R�(KK��h�C4      �  �  �   *         �     u        �t�bhhK ��h��R�(KK&��h�C�   8     0         �      �      .   �   {         A   �	        �   �              �  �  N            �  �  H
  
            �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C@%   �     �  *  �           V          b        �t�bhhK ��h��R�(KK��h�C{      	           �t�bhhK ��h��R�(KK��h�C
   K       4     �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C\y      7  +      �    &      F  +           �      �  h   z     �        �t�bhhK ��h��R�(KK��h�C,"   >  �        �                �t�bhhK ��h��R�(KK��h�CH
   k           �  2   �     d      �    �  9   �        �t�bhhK ��h��R�(KK��h�Ci     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CT      0   -  >      -   0                     .   :   W              �t�bhhK ��h��R�(KK��h�CX      J   �   h      �      5      �      g  �   `   �     ,               �t�bhhK ��h��R�(KK��h�C<   (   �  
   t      �        2     �           �t�bhhK ��h��R�(KK��h�C<   <      8           I   m  '      &           �t�bhhK ��h��R�(KK��h�C4!      1     n   ?      
   3   6           �t�bhhK ��h��R�(KK	��h�C$�   �         	      	         �t�bhhK ��h��R�(KK��h�C %         	      	         �t�bhhK ��h��R�(KK��h�C          	      	         �t�bhhK ��h��R�(KK��h�CM   .     �  I
        �t�bhhK ��h��R�(KK	��h�C$      �     �   J
     N     �t�bhhK ��h��R�(KK��h�C    0            W        �t�bhhK ��h��R�(KK��h�C,K
  "   �   �     
  	      	         �t�bhhK ��h��R�(KK��h�C<         -   s   �     s   `  �  C      �        �t�bhhK ��h��R�(KK
��h�C(      =         L
     ]         �t�bhhK ��h��R�(KK��h�C9     �t�bhhK ��h��R�(KK��h�C<   �   
   w  �     �        '         #        �t�bhhK ��h��R�(KK	��h�C$1   #   
   3   6      m         �t�bhhK ��h��R�(KK��h�C<   d     �           M
     D   �  �   �        �t�bhhK ��h��R�(KK��h�C</        W           @      %   N
     �        �t�bhhK ��h��R�(KK��h�C    $     	      	         �t�bhhK ��h��R�(KK��h�C     �     �t�bhhK ��h��R�(KK��h�C8;  &   �     �     �  �      {     J        �t�bhhK ��h��R�(KK��h�C`Y      O         �           �           %      E
  C                       �t�bhhK ��h��R�(KK��h�C    �     c  X  ;  r      �t�bhhK ��h��R�(KK��h�CD1   #      K     	  "            	  
      ]  T        �t�bhhK ��h��R�(KK	��h�C$P     �      (  ,   	         �t�bhhK ��h��R�(KK��h�C,"      (      x        j   �        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK
��h�C(/   (      (     �	  
            �t�bhhK ��h��R�(KK��h�CP2      =               K  �   �        I   /   9   -     V        �t�bhhK ��h��R�(KK��h�C 5         &     z	  r      �t�bhhK ��h��R�(KK��h�C8         �  �  (  q     q  �     �	        �t�bhhK ��h��R�(KK��h�C<         �  4      2        $   �     "	        �t�bhhK ��h��R�(KK��h�Cv  M          {     �t�bhhK ��h��R�(KK��h�C!         	         �t�bhhK ��h��R�(KK��h�CD   >   a      �     �t�bhhK ��h��R�(KK��h�C4%         
           �  �  �   �        �t�bhhK ��h��R�(KK��h�C4U        (      8   {         8   �        �t�bhhK ��h��R�(KK��h�C8   l         �        �	  �   3             �t�bhhK ��h��R�(KK��h�Cp      �   L         �  
   $   �   N     i        G      

     
      �                     �t�bhhK ��h��R�(KK��h�C �  -  C   �      
        �t�bhhK ��h��R�(KK��h�C<�   q   7        Y  /               a            �t�bhhK ��h��R�(KK	��h�C$        "                 �t�bhhK ��h��R�(KK��h�CT�     �     �   �          �     c  c  �        �              �t�bhhK ��h��R�(KK��h�C<         �   �   &      h  8        �   I         �t�bhhK ��h��R�(KK��h�CX        -   *               �         n         w   ~      �   n         �t�bhhK ��h��R�(KK��h�C8�   ]  �        �           	      	         �t�bhhK ��h��R�(KK��h�C2      )   z   }         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C`
   3  &      q  �  H   l      �       g       g       �         �        �t�bhhK ��h��R�(KK��h�Cp      �t�bhhK ��h��R�(KK��h�C@      J         �  �  �  
   �       
           �t�bhhK ��h��R�(KK��h�C@Z                  �      �     ?          �     �t�bhhK ��h��R�(KK��h�C          
   �  *        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C4   S         Q   O
           8   4         �t�bhhK ��h��R�(KK	��h�C$                 0        �t�bhhK ��h��R�(KK��h�C02      �      0   4   
   _      �        �t�bhhK ��h��R�(KK��h�CL�      )   �   5  �     o     �  &   �   �        J  V        �t�bhhK ��h��R�(KK��h�C�     	      	         �t�bhhK ��h��R�(KK	��h�C$�         x      v   �        �t�bhhK ��h��R�(KK��h�C,         �  3     $   E      �      �t�bhhK ��h��R�(KK��h�C<   8   S        .        �  5      s   �        �t�bhhK ��h��R�(KK��h�C8   �                  &   �  �    �        �t�bhhK ��h��R�(KK��h�CLq         ,            z  �  �     �           X           �t�bhhK ��h��R�(KK��h�C<!      !  �      E      >  '   
   �      F         �t�bhhK ��h��R�(KK��h�C8              #   !      R      �   �         �t�bhhK ��h��R�(KK��h�C`         F  +                 =      n     �  *            u              �t�bhhK ��h��R�(KK��h�C8"   �            2   �   �  �  p     P
        �t�bhhK ��h��R�(KK��h�CX*         i  
         J         i     n         �         
   �         �t�bhhK ��h��R�(KK
��h�C(_  #   
   3   6   �             �t�bhhK ��h��R�(KK��h�C,]     �   
     Q      �   [        �t�bhhK ��h��R�(KK
��h�C(!         	      	      	   K      �t�bhhK ��h��R�(KK��h�C4�      �   1     �   �      4  o  4         �t�bhhK ��h��R�(KK��h�C&  ,      �t�bhhK ��h��R�(KK*��h�C�!         	      	   K   	   �   	   �   	     	   I  	   U  	   �  	   �   	   �  	   �  	   �  	     	   s  	      	   )  	      	   �  	         �t�bhhK ��h��R�(KK ��h�C�   �  #              �  
            �      �            �  �     2         �   �     0   �   �        �t�bhhK ��h��R�(KK��h�C4@          _	                          �t�bhhK ��h��R�(KK��h�C\   (   2        r      �t�bhhK ��h��R�(KK��h�CD     X         �t�bhhK ��h��R�(KK��h�Ch      �      �           5   <         �   �     .     #   !      |      <  R         �t�bhhK ��h��R�(KK��h�C,-         �      \  �     �        �t�bhhK ��h��R�(KK��h�C     `      r      �t�bhhK ��h��R�(KK��h�C0�  1     �  1  ?      
   �  F         �t�bhhK ��h��R�(KK��h�C8   �  C      P   g      n   
      �  �        �t�bhhK ��h��R�(KK��h�CL   $   2     �  �      �  �   Q
  �   $   �   �	                �t�bhhK ��h��R�(KK��h�C<I      ;      �  �     )   %           N        �t�bhhK ��h��R�(KK
��h�C(*   D   �  >   2   F  �  X        �t�bhhK ��h��R�(KK��h�C,�      -   �     �   �  i   �        �t�bhhK ��h��R�(KK��h�C4      �             R
     �  \        �t�bhhK ��h��R�(KK��h�C<V  $  &   g              J  �     �  �        �t�bhhK ��h��R�(KK��h�C   {         �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�CPW      
   $   8  �  �   $   E            �  @     <     �        �t�bhhK ��h��R�(KK��h�CD
              ~   �                  0   �   �        �t�bhhK ��h��R�(KK��h�C     r         �t�bhhK ��h��R�(KK��h�CT      �  �   �      {  �     l  �       �        Y     �        �t�bhhK ��h��R�(KK��h�C8      F     �  5     $   E      
  $        �t�bhhK ��h��R�(KK��h�C             �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK
��h�C(   �  �      �        �        �t�bhhK ��h��R�(KK��h�C@   �      �t�bhhK ��h��R�(KK��h�C83   �  S
     s    #   !      m     �         �t�bhhK ��h��R�(KK��h�C    $   E   &      �         �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C      �        �t�bhhK ��h��R�(KK	��h�C$r  �        	      	         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C@�   >   %      ,        �     
   �                 �t�bhhK ��h��R�(KK��h�C2	          �t�bhhK ��h��R�(KK��h�CD
   �   F   '   !           �         0   �   S  �         �t�bhhK ��h��R�(KK��h�CH   /      �     �     �   �  O     �   �        7         �t�bhhK ��h��R�(KK��h�C0      -  �  %  |      �     @        �t�bhhK ��h��R�(KK��h�C<�       
      W  2     �   J     $   �         �t�bhhK ��h��R�(KK��h�C      g  �     	     �t�bhhK ��h��R�(KK��h�CX
      ]  T  ?      !      �         >   $  T      J   �  �               �t�bhhK ��h��R�(KK��h�CH�  L     %   ?  V      G     �               �  �        �t�bhhK ��h��R�(KK��h�C8      '            �           �            �t�bhhK ��h��R�(KK��h�C8P        L  �   m  {     �  �  �            �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK	��h�C$�   >   �   s   	  N   
        �t�bhhK ��h��R�(KK��h�C42      =      Q  "   �          <        �t�bhhK ��h��R�(KK��h�C,   �   R      u     /   9   -        �t�bhhK ��h��R�(KK��h�C0     �            �  {      �         �t�bhhK ��h��R�(KK��h�C0�      �     >  	      	      	   K      �t�bhhK ��h��R�(KK��h�CL   =  �     t     R	  
   l                  +      T
        �t�bhhK ��h��R�(KK��h�C8   @      W	     9                          �t�bhhK ��h��R�(KK��h�C@      J   a      �     �  �      U
  
   Q           �t�bhhK ��h��R�(KK
��h�C(�      h     B   [     �        �t�bhhK ��h��R�(KK��h�CL-   A   Y      �  O      �  C                 U  "   �	        �t�bhhK ��h��R�(KK��h�Ch*   �   _  o     �   
   c  �        \   �   D      A     K     ~   
      S   �        �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6            �t�bhhK ��h��R�(KK��h�CV
       �t�bhhK ��h��R�(KK��h�C1   #       9     �t�bhhK ��h��R�(KK��h�C      :         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�Cl"   �  (      )   �   
   �      ^   �     s  *      5   x      ~     /           �         �t�bhhK ��h��R�(KK��h�C   �     .     �        �t�bhhK ��h��R�(KK��h�C          M        W
     �t�bhhK ��h��R�(KK��h�C �     %   3     �  �     �t�bhhK ��h��R�(KK��h�CL   &   �   a      L  *      �            �   S   Q              �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C8*   �        c      �     �  +   
   "        �t�bhhK ��h��R�(KK��h�CD   �     �  -         
   �   �  =  h                 �t�bhhK ��h��R�(KK��h�CT�	  �   �     Y      O               Y      O      $   �  >   T        �t�bhhK ��h��R�(KK��h�C g     �  D   X
          �t�bhhK ��h��R�(KK$��h�C�         �           �     s           ;      0   [      �              :              [     �     8   E        �t�bhhK ��h��R�(KK��h�CL         <        n   &      U   �      %   o      h  u         �t�bhhK ��h��R�(KK��h�C`     ?  �   �      �  �       7   �  ;   R      [      p      {      o        �t�bhhK ��h��R�(KK��h�C D   _  C   )   �           �t�bhhK ��h��R�(KK��h�C<�     "   >  �     �          
      �        �t�bhhK ��h��R�(KK��h�CL�     �   -   �  +      �  �      �  �  g      n      +         �t�bhhK ��h��R�(KK��h�C/      A               �t�bhhK ��h��R�(KK��h�C             9      �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C,[         2      0   *   2      F     �t�bhhK ��h��R�(KK��h�C0�  <	  �           F  *      S        �t�bhhK ��h��R�(KK��h�C<*      	  �      [     W  �   �                 �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�CHD   _  C      S   �           �   �           B   �        �t�bhhK ��h��R�(KK��h�C <      �  	      	         �t�bhhK ��h��R�(KK��h�Cx#   !      \         0   4   '   
   3   �  �     �     �     �     /      K     �     h  6        �t�bhhK ��h��R�(KK
��h�C(�     j     #                �t�bhhK ��h��R�(KK��h�C4      n     �  r      �t�bhhK ��h��R�(KK��h�C   ,   	      	         �t�bhhK ��h��R�(KK��h�Cb   D  
   c        �t�bhhK ��h��R�(KK��h�C,A              t  %      o        �t�bhhK ��h��R�(KK��h�C�	     �t�bhhK ��h��R�(KK��h�CP  �   �     P	           �  �     ,         �  C      w        �t�bhhK ��h��R�(KK��h�C�  +     �t�bhhK ��h��R�(KK��h�C Z   �     K               �t�bhhK ��h��R�(KK��h�C4�   f     g  �     	      	      	   K      �t�bhhK ��h��R�(KK��h�CH         9     7            0   x        ^   �   &        �t�bhhK ��h��R�(KK��h�C     �   
   �         �t�bhhK ��h��R�(KK��h�C@Y           �  C  J       %         �   �         �t�bhhK ��h��R�(KK��h�CXk  "         �   Y
  !      �        �            �      _     �         �t�bhhK ��h��R�(KK��h�CH      5   :  <      [      &      U   $   N     i           �t�bhhK ��h��R�(KK��h�C
	     	         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CP           x   �  E      @  ^      �  �  Z      �               �t�bhhK ��h��R�(KK��h�CL*   D   �  s   7            
  �   `   Z
  )      v  '   �        �t�bhhK ��h��R�(KK��h�C<h        .   
   �        z         B   ^	         �t�bhhK ��h��R�(KK��h�C0
      �   D  >      v     �  w         �t�bhhK ��h��R�(KK��h�C@l  �  v     d   8          �         d   b        �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�CT            b         
  �            )   �   k  =  ^   F  F         �t�bhhK ��h��R�(KK��h�Cw     �t�bhhK ��h��R�(KK��h�C   @   '   H   W        �t�bhhK ��h��R�(KK��h�C`,   O         �  �      -   �           $  ,   �     �  3     t               �t�bhhK ��h��R�(KK��h�C2
              �t�bhhK ��h��R�(KK��h�CL
   �  F   '            ,   �   V         z   ,   
   �   �         �t�bhhK ��h��R�(KK	��h�C$1   #       �     �  m         �t�bhhK ��h��R�(KK��h�C@      w   s  *      \   �      J   N         `        �t�bhhK ��h��R�(KK��h�C,�   �             �  
            �t�bhhK ��h��R�(KK��h�C4   �               [                �t�bhhK ��h��R�(KK��h�CD*      �               z     �     4   
   8   �         �t�bhhK ��h��R�(KK��h�Cp           m         b      x   G      �     $   k      G      f   w        ;      @        �t�bhhK ��h��R�(KK��h�C �  T     
     U        �t�bhhK ��h��R�(KK
��h�C(               a      j        �t�bhhK ��h��R�(KK��h�C8   8   /   	  �   :     M   �      $   N        �t�bhhK ��h��R�(KK��h�C,b   #      �     &  �   
            �t�bhhK ��h��R�(KK��h�C�     /      �      �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C@R  �      u      �      -          ~     /         �t�bhhK ��h��R�(KK��h�C �      )                  �t�bhhK ��h��R�(KK��h�C'     g           �t�bhhK ��h��R�(KK��h�C                �t�bhhK ��h��R�(KK��h�C4*      �        &      }        �        �t�bhhK ��h��R�(KK��h�Ch@      �           V         b      Y
  !      @      �   R            {      �         �t�bhhK ��h��R�(KK��h�CH      5     �   �   �     &      �     �   T      �        �t�bhhK ��h��R�(KK��h�CT      -   �      6  �  �      �  �     �      �  ;        �        �t�bhhK ��h��R�(KK��h�Ch*      �  L      �        b      �
     �      &                       �   }         �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�CT   &   �   j        �  �   V   �          �             �        �t�bhhK ��h��R�(KK��h�C8O   :   h  ?  >   )  C   �  
   |      �         �t�bhhK ��h��R�(KK��h�ChR             n         .      �     �           �  �   z  �   O     �   �        �t�bhhK ��h��R�(KK��h�C1   #       �  �         �t�bhhK ��h��R�(KK
��h�C(   �  '        �      w        �t�bhhK ��h��R�(KK��h�CD[
    
   ,            w     %   e    )   
            �t�bhhK ��h��R�(KK��h�C,
   "  '            $   �  �        �t�bhhK ��h��R�(KK��h�C:   �   S   Q         �t�bhhK ��h��R�(KK��h�C<
   t   &      *  �               �              �t�bhhK ��h��R�(KK��h�C4      �     �t�bhhK ��h��R�(KK��h�C9     �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C�          �t�bhhK ��h��R�(KK��h�C,   <        o      �     \
        �t�bhhK ��h��R�(KK��h�C,            �     �     /         �t�bhhK ��h��R�(KK��h�CD5     �  &      T   n   x     �      )   r  �   3        �t�bhhK ��h��R�(KK��h�C0   �         0   4   
   _      �        �t�bhhK ��h��R�(KK��h�C,   �	        v      �     �        �t�bhhK ��h��R�(KK��h�C
            �t�bhhK ��h��R�(KK
��h�C(�   (   �   <      x         r      �t�bhhK ��h��R�(KK��h�CD!        �           n  �        �     ,   O         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C8     K    
   �   �   I   �      -  D         �t�bhhK ��h��R�(KK��h�CHD   >   N   9     7   �     �     �  T        4   V        �t�bhhK ��h��R�(KK��h�CT      �   *     �   N   �             �      %   !  (      n         �t�bhhK ��h��R�(KK��h�C<#   !      X     k   '   
   3   6   2              �t�bhhK ��h��R�(KK��h�CH?
     J                   �	     2   �     �            �t�bhhK ��h��R�(KK��h�CX
   �	  F      "      x    �   �        B        5      L             �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CD   f     g  )     #  6  (        �  /     X         �t�bhhK ��h��R�(KK	��h�C$�      y  �   &   T     t      �t�bhhK ��h��R�(KK��h�CP/      p        .   a   �
     �          �     �     �        �t�bhhK ��h��R�(KK��h�C4"   �   E  '           �  =  
           �t�bhhK ��h��R�(KK��h�CT            �     $   �        �        
   9    
   $           �t�bhhK ��h��R�(KK��h�C   �  �  9   �        �t�bhhK ��h��R�(KK
��h�C(+  �  �           �           �t�bhhK ��h��R�(KK��h�C,
      (      <      �	              �t�bhhK ��h��R�(KK	��h�C$      �     �      �        �t�bhhK ��h��R�(KK��h�C�      �      �t�bhhK ��h��R�(KK
��h�C(�   �   �   z    �   �   z         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C4      B
  H   �  q  
   B   �     @         �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK	��h�C$!            	      	         �t�bhhK ��h��R�(KK��h�C,�   ,   O      ]
  c         �  �      �t�bhhK ��h��R�(KK��h�C 
   j  �   -   �          �t�bhhK ��h��R�(KK��h�C1   Q  S     �t�bhhK ��h��R�(KK��h�C�     @      �t�bhhK ��h��R�(KK	��h�C$#   !      h                   �t�bhhK ��h��R�(KK��h�C0   B  �     3           �     �      �t�bhhK ��h��R�(KK��h�CL
         O  {     2      �        .                       �t�bhhK ��h��R�(KK��h�CH*      �  �      >
        d  -   A   q	     5     E         �t�bhhK ��h��R�(KK��h�CP*      ~         �      �  �     �       +   �   7      �        �t�bhhK ��h��R�(KK
��h�C(      �  �          �        �t�bhhK ��h��R�(KK��h�C`
   �  �   �      &  �  u      �               �      �      -  +     �  �     �t�bhhK ��h��R�(KK��h�C        �      4      �t�bhhK ��h��R�(KK��h�Ct*   �   1  �      5   <         �        �     �
        �   =            ^
                    �t�bhhK ��h��R�(KK��h�CX      �  �   �  Y  �  
      
       &      �   M   �                 �t�bhhK ��h��R�(KK
��h�C(                  �     `     �t�bhhK ��h��R�(KK��h�C*         F     �t�bhhK ��h��R�(KK��h�CD            �     -  �             �  G   �        �t�bhhK ��h��R�(KK��h�C4-   �     �     ;      0   �     �        �t�bhhK ��h��R�(KK��h�C       g  )               �t�bhhK ��h��R�(KK��h�C,      P   �   o   
      .           �t�bhhK ��h��R�(KK��h�C�  c            �t�bhhK ��h��R�(KK��h�C@   .        P   !      u  �        �      �        �t�bhhK ��h��R�(KK��h�CL
        a     �              P   W  
   B   [  
   ,         �t�bhhK ��h��R�(KK��h�C1   #       �      �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   6         �        �t�bhhK ��h��R�(KK	��h�C$  
   _                    �t�bhhK ��h��R�(KK��h�C0      P   �   =  
                    �t�bhhK ��h��R�(KK��h�C@"   �     Z  �              �      �   N  /        �t�bhhK ��h��R�(KK��h�C P        	      	         �t�bhhK ��h��R�(KK��h�CX*      J  +      �              )  +      )     �      $   �   d        �t�bhhK ��h��R�(KK��h�C               �t�bhhK ��h��R�(KK��h�CX1      �        
   3   6     g   d   t          �      /      V        �t�bhhK ��h��R�(KK��h�C�               a     �t�bhhK ��h��R�(KK��h�C      0   �        �t�bhhK ��h��R�(KK��h�C\y      m  )     B        5   �      `           >   )  `        �        �t�bhhK ��h��R�(KK��h�CDT   >   )   %   �         �        5  A     �   �         �t�bhhK ��h��R�(KK��h�C,      �   L   
     ^   $   N        �t�bhhK ��h��R�(KK��h�C1   #       A   d     �t�bhhK ��h��R�(KK��h�Cx         k               =      �  �  G   W      -     /   9   �   7      f     �  M     {        �t�bhhK ��h��R�(KK
��h�C(T      �           
   �        �t�bhhK ��h��R�(KK��h�CH   ?  V               �     �   S   Q                     �t�bhhK ��h��R�(KK��h�C      J   z      �     �t�bhhK ��h��R�(KK��h�C<      )   0   �  
   �  B   .
     q             �t�bhhK ��h��R�(KK��h�C�            �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�Cq   �     �t�bhhK ��h��R�(KK��h�C<      �   �              �   _
                �t�bhhK ��h��R�(KK��h�C42      H  �         7   .     g            �t�bhhK ��h��R�(KK	��h�C$9   �  (   D                 �t�bhhK ��h��R�(KK��h�CH      -   M   c   I     _     $   
  "   B   Z     �        �t�bhhK ��h��R�(KK��h�C,        �   �            9	        �t�bhhK ��h��R�(KK��h�C �     |     �             �t�bhhK ��h��R�(KK��h�C0|      �   h  R      �                �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�Cb           �      �t�bhhK ��h��R�(KK��h�C4
         �  �  H      :   �     e         �t�bhhK ��h��R�(KK��h�C,X            %   �  �     T        �t�bhhK ��h��R�(KK
��h�C(!      �        	      	         �t�bhhK ��h��R�(KK��h�CX)            �  }  (            �   
        S  ]      �             �t�bhhK ��h��R�(KK��h�C@�      ;      �     V        L   T         F        �t�bhhK ��h��R�(KK��h�C �     �  	      	         �t�bhhK ��h��R�(KK��h�C`   $   n      �	     .      H          �          f   �     %   I  �        �t�bhhK ��h��R�(KK��h�C�     �              �t�bhhK ��h��R�(KK	��h�C$�     �  �      �          �t�bhhK ��h��R�(KK��h�C         �     �t�bhhK ��h��R�(KK��h�C@            %     i	        =      �  :   P        �t�bhhK ��h��R�(KK��h�CT         m      @        P   <   "      .   C          $   k         �t�bhhK ��h��R�(KK��h�C0�     B  y   8   4      �   �	  c         �t�bhhK ��h��R�(KK��h�C�	           �t�bhhK ��h��R�(KK��h�CT      J   =         +     �        �     +  
   �  �  /  F         �t�bhhK ��h��R�(KK'��h�C�   $   �      �   +           L         �        �            ;      =      �                           �   �               �t�bhhK ��h��R�(KK
��h�C(   	      	      	   K   	   �      �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C 2      )   i             �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�CX      �      M   <         1  *      �  8   -           &   N   ~        �t�bhhK ��h��R�(KK��h�CP   �      y  �      �        �   *                            �t�bhhK ��h��R�(KK��h�C,  g     1  "      	      	         �t�bhhK ��h��R�(KK��h�C`
   �                 )   
   `
           S  [    D	  p	       �   �        �t�bhhK ��h��R�(KK
��h�C(M      +   �   *      @  t          �t�bhhK ��h��R�(KK��h�C0�   �   7     I   �    
   3           �t�bhhK ��h��R�(KK��h�CP      �     �   �        v               f          �        �t�bhhK ��h��R�(KK��h�C,�  �  (      �  C   �   q   7        �t�bhhK ��h��R�(KK	��h�C$!            	      	         �t�bhhK ��h��R�(KK��h�C%   �        �t�bhhK ��h��R�(KK��h�C8   >   �   �         
         %   �            �t�bhhK ��h��R�(KK��h�C                �t�bhhK ��h��R�(KK��h�Cl   �      o  �        +         J   a   �           =      
              �  �         �t�bhhK ��h��R�(KK��h�C|      �            m  �   e  [  i      Y      Q         Q     Q      x  �  $   �   �     �             �t�bhhK ��h��R�(KK��h�C@W   �  J  S  g      D      
     ~        <        �t�bhhK ��h��R�(KK��h�CL         k      l                 ;      ,  %   �           �t�bhhK ��h��R�(KK��h�C �  *      l  �            �t�bhhK ��h��R�(KK��h�C.          �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C!      ,         �t�bhhK ��h��R�(KK��h�C@      �         .   *      &   �                    �t�bhhK ��h��R�(KK��h�C8      0   4      �  >      a         �        �t�bhhK ��h��R�(KK��h�C    �  �  c   
            �t�bhhK ��h��R�(KK
��h�C(�        '   
   e   �   F         �t�bhhK ��h��R�(KK��h�C8      J         M      +   $   �     �
        �t�bhhK ��h��R�(KK"��h�C�               :      S   Y      Q   5      �      v         �  
   `   �       %   a
           �      +         �t�bhhK ��h��R�(KK��h�C,   X     �                       �t�bhhK ��h��R�(KK��h�C,      s   l  }      ,               �t�bhhK ��h��R�(KK
��h�C(%   H     *   2   m     o          �t�bhhK ��h��R�(KK��h�C89   �     �         )   �  `   �     ,         �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6            �t�bhhK ��h��R�(KK��h�C,	   �  	   �	  	   �  	   �  	   �     �t�bhhK ��h��R�(KK��h�C�      �   �     r      �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK	��h�C$                           �t�bhhK ��h��R�(KK	��h�C$         �          {     �t�bhhK ��h��R�(KK��h�C0
      �   D  >      v     �  w         �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK
��h�C(      ,  '   �  �     �        �t�bhhK ��h��R�(KK��h�Ch      �     4         �     �   _         .   �           a   ;      �               �t�bhhK ��h��R�(KK��h�Cp   5   7  4                     4      �        S   Y      Q            :  "      .        �t�bhhK ��h��R�(KK��h�CP         	      	      	   K   	     	   I  	   �  	   �   	   s     �t�bhhK ��h��R�(KK��h�C<   "   �      �t�bhhK ��h��R�(KK��h�C #   !   '   
   �  F         �t�bhhK ��h��R�(KK	��h�C$Z      �      Q              �t�bhhK ��h��R�(KK��h�CL^               %  2   (         X	     A   �     �           �t�bhhK ��h��R�(KK��h�CTg         �         
              /   0   �                       �t�bhhK ��h��R�(KK��h�C4         	     W   v   c         �        �t�bhhK ��h��R�(KK��h�CE         	         �t�bhhK ��h��R�(KK��h�C\�   �  >         �  �   �     %   �     �   �   �   �     y    	     �         �t�bhhK ��h��R�(KK
��h�C(�      r     t  %   e  �        �t�bhhK ��h��R�(KK��h�C!  �      /      �t�bhhK ��h��R�(KK��h�Cz  <     >     �t�bhhK ��h��R�(KK
��h�C(?  (      �           Z        �t�bhhK ��h��R�(KK��h�C4     R   h   m     	      	     	   �      �t�bhhK ��h��R�(KK��h�C�          �           �t�bhhK ��h��R�(KK��h�C�                   �t�bhhK ��h��R�(KK��h�CD        O  �                                  �t�bhhK ��h��R�(KK��h�C<:     )   N   �     C	     �   "        �        �t�bhhK ��h��R�(KK��h�C   g           �t�bhhK ��h��R�(KK
��h�C(      -   q     �     �         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C    �  �     �          �t�bhhK ��h��R�(KK��h�Ct      D  �   �        &      a      �      �      %   j	  �     �   �  �     $   �              �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK&��h�C�         O      �      %     z        Y      Q         Q     Q         x     �               z      >      F  $   �        �t�bhhK ��h��R�(KK��h�C�   �      �t�bhhK ��h��R�(KK��h�C      	         �t�bhhK ��h��R�(KK��h�C<�   =     �  i   *     �  c      o      n        �t�bhhK ��h��R�(KK��h�C0%   f     g  �	        �   )            �t�bhhK ��h��R�(KK��h�C s        �               �t�bhhK ��h��R�(KK��h�C1   #       �        �t�bhhK ��h��R�(KK	��h�C$        �                 �t�bhhK ��h��R�(KK	��h�C$   @      2   �     !        �t�bhhK ��h��R�(KK��h�CT      �            �       �      �      �  �      h     �         �t�bhhK ��h��R�(KK��h�C`W       *         6     �  
   �            �   �     I   $  
   �   :        �t�bhhK ��h��R�(KK��h�C    �   �        �  r      �t�bhhK ��h��R�(KK��h�CT%  +      %   $  .  
   }  S
     s     e      S
     s     @         �t�bhhK ��h��R�(KK
��h�C(:   �      �     �  b
  �        �t�bhhK ��h��R�(KK��h�C@      }     E   
   y     �     �   s     W         �t�bhhK ��h��R�(KK��h�C1   #               �t�bhhK ��h��R�(KK��h�C<      
        �   �        i      A   ?        �t�bhhK ��h��R�(KK
��h�C(P  &   �  �  �  _  g   c
        �t�bhhK ��h��R�(KK��h�C0g   �  ]     �         �   $   �         �t�bhhK ��h��R�(KK��h�C<         .  "     $  I      �      I   �        �t�bhhK ��h��R�(KK��h�C4K       �     �  �      �     �        �t�bhhK ��h��R�(KK��h�C#     �     �        �t�bhhK ��h��R�(KK��h�C\b     �   �          %  =	     �  �   �   *   2     �      �              �t�bhhK ��h��R�(KK��h�C\�        �  v                   �           I	  �        I  �        �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C,W      �     �   c   !  9   o        �t�bhhK ��h��R�(KK��h�C89   A            s   o  Y  f  
      6         �t�bhhK ��h��R�(KK��h�C,      
     �      �   �   �         �t�bhhK ��h��R�(KK��h�CL         E  Y  �        =      d
          3  "           �t�bhhK ��h��R�(KK��h�C8            m	  0  �   �           �        �t�bhhK ��h��R�(KK��h�C8
   }  '   L  �  x      1     \              �t�bhhK ��h��R�(KK��h�C,8     �     M   �      �   /         �t�bhhK ��h��R�(KK��h�C W  "      	      	         �t�bhhK ��h��R�(KK��h�CD      ,     �  �   �  �  s   �   y        
   		        �t�bhhK ��h��R�(KK��h�C@�            ;      �	     -   %        �   B	        �t�bhhK ��h��R�(KK��h�C    2   4  �   ,   �   r      �t�bhhK ��h��R�(KK��h�Cp
   3   6   �     �  '   !      �         0   <                    �  �          �         �t�bhhK ��h��R�(KK��h�C�   =  	      	         �t�bhhK ��h��R�(KK��h�C8#   !      �     �  �  (      
              �t�bhhK ��h��R�(KK'��h�C�      D  �  "      o      S          S   Y   �   Q     Q      &   �               �  �              8   {   �  A  �   �   �     �t�bhhK ��h��R�(KK	��h�C$t           	      	         �t�bhhK ��h��R�(KK��h�CP               4      �  
   _      �             
   �        �t�bhhK ��h��R�(KK��h�C@�      #  I           V           �     �        �t�bhhK ��h��R�(KK��h�C,   �  T  I   l      ~               �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�CH\   H     �   �     ,     \   �  $   2        �           �t�bhhK ��h��R�(KK��h�Co  e
     �t�bhhK ��h��R�(KK��h�CP         
   c        �  "     !        �           �         �t�bhhK ��h��R�(KK��h�CI   k  �     �t�bhhK ��h��R�(KK��h�C1   #       �          �t�bhhK ��h��R�(KK��h�C   $  �   �        �t�bhhK ��h��R�(KK��h�C<   �  �   7   
   �     �   %          �        �t�bhhK ��h��R�(KK��h�C@�  g  &   �   {	     �     e        ,               �t�bhhK ��h��R�(KK��h�CH�	     �     �  	      	   K   	     	   �  	   �   	   >     �t�bhhK ��h��R�(KK��h�C@      �                 �  &                    �t�bhhK ��h��R�(KK��h�C       �     �   s        �t�bhhK ��h��R�(KK��h�CD      P                    E  �  �      �   �         �t�bhhK ��h��R�(KK
��h�C(-   !  |     ;      �          �t�bhhK ��h��R�(KK��h�Ch      �        �     �         P   �           G   W                 �   f        �t�bhhK ��h��R�(KK��h�C44      2           5      4               �t�bhhK ��h��R�(KK	��h�C$�     |      �      �         �t�bhhK ��h��R�(KK	��h�C$Z       �  �     �        �t�bhhK ��h��R�(KK��h�C *           #   !         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C0�   �     9  �     �  i   %   �         �t�bhhK ��h��R�(KK��h�C@      5           &      �   �   L   G      o        �t�bhhK ��h��R�(KK��h�C�  	      	         �t�bhhK ��h��R�(KK��h�C@
   u  F   ?         �  �   %     V   �      �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CF            �t�bhhK ��h��R�(KK
��h�C(   e   '   �  �     �   5        �t�bhhK ��h��R�(KK��h�CD      $   f
  n      8   S  ]     �   �        G  ]     �t�bhhK ��h��R�(KK��h�CP   (   <         �      �  
         x      �   +         #        �t�bhhK ��h��R�(KK
��h�C(k        �    �  �   �         �t�bhhK ��h��R�(KK��h�C,#   !      �  (      :   @            �t�bhhK ��h��R�(KK��h�C\            L  �         .                     9   �  �   g
     '        �t�bhhK ��h��R�(KK��h�CP   ;        C      �   d  4       t      �           )        �t�bhhK ��h��R�(KK��h�C<   "      �     �t�bhhK ��h��R�(KK��h�C   �         .   �     �t�bhhK ��h��R�(KK��h�C 4         	      	         �t�bhhK ��h��R�(KK��h�C8   X      2   0   ,  
   ,                     �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C4>     %   W             �        7      �t�bhhK ��h��R�(KK��h�C4        -            �	     4   �         �t�bhhK ��h��R�(KK��h�CP      /           �         �         /  *     (     ]         �t�bhhK ��h��R�(KK
��h�C(   h
  �     :     $   �        �t�bhhK ��h��R�(KK��h�CP      U   �  *            �  m      @     ~     /      �         �t�bhhK ��h��R�(KK��h�C<*            �   >      F  +           <        �t�bhhK ��h��R�(KK��h�C<   �  C      �  B      �  y   2        �        �t�bhhK ��h��R�(KK��h�C�  )  	      	         �t�bhhK ��h��R�(KK
��h�C(      )   0      �   ~  "          �t�bhhK ��h��R�(KK��h�C\            ;      �   %   �        
           P   +         �   D        �t�bhhK ��h��R�(KK��h�Cl-      /      �           �   O         Y      Q      �     x  >   =      n     �        �t�bhhK ��h��R�(KK��h�CDB           �	     I   �   �           ;      0         �t�bhhK ��h��R�(KK��h�C<   �      �  x      �        �     �     �      �t�bhhK ��h��R�(KK��h�CH         &   D  0      �   ~  >   `   3  T     q   i
        �t�bhhK ��h��R�(KK��h�C`      .   �  �   +        n      )     	  5      a      �  �	     /  �        �t�bhhK ��h��R�(KK��h�C;	        �t�bhhK ��h��R�(KK��h�C4�   /        �      ;      6     �        �t�bhhK ��h��R�(KK��h�C'           �t�bhhK ��h��R�(KK��h�C0   }         .   �           /        �t�bhhK ��h��R�(KK
��h�C(
   *  +     �   G     ,        �t�bhhK ��h��R�(KK��h�C                �t�bhhK ��h��R�(KK��h�C       -  T     X          �t�bhhK ��h��R�(KK#��h�C�   �           �     �	  )     +            -   0   -      �  
               -         �              �        �t�bhhK ��h��R�(KK��h�C<1   #      ?        
   3   6   )  ?   �   �   r      �t�bhhK ��h��R�(KK��h�CL            �     C           C   
      S     i   �	        �t�bhhK ��h��R�(KK��h�C   0         �t�bhhK ��h��R�(KK��h�C 1   #       m      4         �t�bhhK ��h��R�(KK��h�C <  �   �        /         �t�bhhK ��h��R�(KK��h�Cx^      �        =         n   "   -     .  �     u  *        ?      )   
   -     .  /  F   *
     �t�bhhK ��h��R�(KK	��h�C$   l                        �t�bhhK ��h��R�(KK��h�C4�
     �	  �  �               A           �t�bhhK ��h��R�(KK��h�C 2
  R     �     >        �t�bhhK ��h��R�(KK��h�C@M     
   R  -         J   
  �        �   s        �t�bhhK ��h��R�(KK��h�C       z   ,               �t�bhhK ��h��R�(KK	��h�C$         Z  �     .        �t�bhhK ��h��R�(KK��h�CS  �  �         �t�bhhK ��h��R�(KK��h�CL   (        t    :   �  8   o         �     8   �           �t�bhhK ��h��R�(KK��h�C@�   &      	  <  N   $   k   �        �  �   n        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK
��h�C(_              �              �t�bhhK ��h��R�(KK��h�CLy         �        &      f     j
     ;      M              �t�bhhK ��h��R�(KK��h�C   P      �     �t�bhhK ��h��R�(KK��h�CL         E     +  �         =         �        G   �        �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C,1   �  
   3   6           �        �t�bhhK ��h��R�(KK	��h�C$U       �   �  �  �        �t�bhhK ��h��R�(KK��h�CT   >   �   �   �      �  E      W      %            5      $   �        �t�bhhK ��h��R�(KK��h�Cd      �  D      V        ;      M   c   /  k
  :   8   {   q  �  D   �  �   7         �t�bhhK ��h��R�(KK��h�CT*         
     U
           O  +         u  *  G   ;              �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C4           =               �  p        �t�bhhK ��h��R�(KK��h�C0     �t�bhhK ��h��R�(KK��h�C@}           �      B            .                  �t�bhhK ��h��R�(KK��h�C@   �            �   
   �   �      �   
               �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK	��h�C$�              
     &     �t�bhhK ��h��R�(KK��h�C8               G     6  �     Y            �t�bhhK ��h��R�(KK��h�CXl         �   k      e      0   '       e   �         .         �        �t�bhhK ��h��R�(KK��h�C|      �   �         �     F     �	  �  '  �      �  &   D  �   '           a   ;      [              �t�bhhK ��h��R�(KK��h�C 1   #       �     �  m      �t�bhhK ��h��R�(KK��h�C      a              �t�bhhK ��h��R�(KK��h�Cp�      2   0   �      2      �  �   �     8     }	  /      K     }	  /         l              �t�bhhK ��h��R�(KK	��h�C$%   ^  �                   �t�bhhK ��h��R�(KK��h�C\�        �        �  �  �                             .  a           �t�bhhK ��h��R�(KK��h�C  4  '  O  7         �t�bhhK ��h��R�(KK��h�C8   �   '   �     5     Q	     �  �   �        �t�bhhK ��h��R�(KK��h�C W         �     �        �t�bhhK ��h��R�(KK	��h�C$1   #       �  g  
   �        �t�bhhK ��h��R�(KK ��h�C�   �         �     1     �     T      �     �  b
  �           H   o         2     K  �    %        �t�bhhK ��h��R�(KK��h�C      m      �t�bhhK ��h��R�(KK��h�C4      �         J  C   B     j           �t�bhhK ��h��R�(KK��h�C8            -   �     2   �  D  "   Z        �t�bhhK ��h��R�(KK��h�C4               X         �              �t�bhhK ��h��R�(KK	��h�C$      -   t                 �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C;	           �      �t�bhhK ��h��R�(KK��h�C#       r      �t�bhhK ��h��R�(KK��h�CH            �             �     M   T   �               �t�bhhK ��h��R�(KK��h�C\l         �  �  �  #      V  9     "  7  J  C      !  "     �  �        �t�bhhK ��h��R�(KK��h�C4   >   �   z   
   �           `   �         �t�bhhK ��h��R�(KK	��h�C$      )   �  �     s        �t�bhhK ��h��R�(KK��h�C         �  h
        �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C�  <     �t�bhhK ��h��R�(KK��h�Chf     �      �  	      	      	   K   	   �   	   �   	     	   �  	   U  	   �   	   �     �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�CD   (               w      j   �   >   �                 �t�bhhK ��h��R�(KK��h�C�   p      ^  M     �t�bhhK ��h��R�(KK��h�C4   �   E  �  j      
        �  q	        �t�bhhK ��h��R�(KK��h�C0   5              $  $   �  G
        �t�bhhK ��h��R�(KK��h�C �     �  	      	         �t�bhhK ��h��R�(KK��h�C<   &   �   �            �  V     �  :   T        �t�bhhK ��h��R�(KK��h�CT�   -     %   f        ]  �        .      J  �            �	        �t�bhhK ��h��R�(KK��h�CDj   �        \  3  
   4     l
  �                     �t�bhhK ��h��R�(KK��h�C|     �t�bhhK ��h��R�(KK��h�CH`        "        f   �   0   R         �  �     �        �t�bhhK ��h��R�(KK��h�C         �      �t�bhhK ��h��R�(KK��h�C@�  "   &  �   +               �   {         �        �t�bhhK ��h��R�(KK��h�CH   �     A   �   �     j
  �  c   �  �         �   �         �t�bhhK ��h��R�(KK��h�C`
   ,      N           �  �      �     �     
   �     �  �      �     �     �t�bhhK ��h��R�(KK��h�C01   #   
   3   6              �        �t�bhhK ��h��R�(KK��h�C|         ?         n   V      J   �      d              +      �         �  n      
  g
  :   E        �t�bhhK ��h��R�(KK��h�C		     �t�bhhK ��h��R�(KK��h�C�   
          �	     �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C,#   !      �
  (      
   �   F         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C0)   �     e	     H   n  �  c   *        �t�bhhK ��h��R�(KK��h�C,      b   $   5     �     x         �t�bhhK ��h��R�(KK��h�C �     /         	         �t�bhhK ��h��R�(KK��h�C@   D            @     :  &         �     5        �t�bhhK ��h��R�(KK��h�CX            i  
            ;      k               B  ]   "   t         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C8�	  2  �  *   �   �      A     �  Y  �         �t�bhhK ��h��R�(KK��h�C4#  &   �   �      �         k         r      �t�bhhK ��h��R�(KK��h�CP�  �          �         /      �  �   �   �          �         �t�bhhK ��h��R�(KK��h�C�  a             �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�C8�     8           v     I   �  �  �        �t�bhhK ��h��R�(KK��h�C,   f   �   (         &  ^   D        �t�bhhK ��h��R�(KK��h�CD
   C  _        -     �     w  
   ,      
            �t�bhhK ��h��R�(KK��h�C<v     H   �  �     %      �         �  �         �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�C              �t�bhhK ��h��R�(KK��h�C�     	   K      �t�bhhK ��h��R�(KK��h�C4\   (   �      �  4            0  �   r      �t�bhhK ��h��R�(KK��h�Cm  �      �t�bhhK ��h��R�(KK��h�CH      �         $   k            k      l                 �t�bhhK ��h��R�(KK��h�C      
   ,         �t�bhhK ��h��R�(KK��h�C�  �      �t�bhhK ��h��R�(KK��h�CDd   �     )   ;      0   !      �     �  D      [        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C�         �     �t�bhhK ��h��R�(KK��h�C0d  -   
   \      �   �     �           �t�bhhK ��h��R�(KK��h�CL$   �           �                 #
  �            +         �t�bhhK ��h��R�(KK��h�C,1   #   
   3   6   �     �   f        �t�bhhK ��h��R�(KK	��h�C$m
     6  �   �     u         �t�bhhK ��h��R�(KK��h�C4:     (      #   !            B   3        �t�bhhK ��h��R�(KK
��h�C(�     
   ,            K         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C�  �      �t�bhhK ��h��R�(KK��h�Cd*                         �              n
     �     �   y  !      �         �t�bhhK ��h��R�(KK��h�C}      �t�bhhK ��h��R�(KK��h�C@g  _  �  �  �         �  �  �           �         �t�bhhK ��h��R�(KK��h�C      �            �t�bhhK ��h��R�(KK��h�C8U        �     *      �           %        �t�bhhK ��h��R�(KK��h�C8      �   �     I         I   &   �  �        �t�bhhK ��h��R�(KK��h�CD     o
     G    
   \   I                          �t�bhhK ��h��R�(KK��h�CLB           �                 �          
   $           �t�be(hhK ��h��R�(KK��h�C4   %  �        
      �  I               �t�bhhK ��h��R�(KK��h�CH�  
   8     #        �      �	  *   2   &   4              �t�bhhK ��h��R�(KK��h�C<	     p  9   �     �t�bhhK ��h��R�(KK	��h�C$      �	  +  �   
   y        �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C �    H  �      4         �t�bhhK ��h��R�(KK��h�C         	         �t�bhhK ��h��R�(KK��h�C�     	      	         �t�bhhK ��h��R�(KK��h�C�	     �	     �t�bhhK ��h��R�(KK��h�C0   �                  ,	  "   W         �t�bhhK ��h��R�(KK	��h�C$�      (  �   +      �        �t�bhhK ��h��R�(KK��h�C0#   !      �   �  '   9      ]          �t�bhhK ��h��R�(KK
��h�C("   �  �	  �     /      ^        �t�bhhK ��h��R�(KK��h�CT   A	  2   v           �t�bhhK ��h��R�(KK��h�C<      �   X  &      U   �           $   k         �t�bhhK ��h��R�(KK��h�C@   6           �     V   '      
   �  �  �        �t�bhhK ��h��R�(KK��h�C 2      �      \  2        �t�bhhK ��h��R�(KK��h�C@*   �  {  �  �  �   �      �  �  (   �   �   �        �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C!         	         �t�bhhK ��h��R�(KK��h�C              �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C8<      `             �  �  	      	         �t�bhhK ��h��R�(KK��h�C   X      �t�bhhK ��h��R�(KK��h�CH   (   #   !      �      G   �        Q   V      O
  &        �t�bhhK ��h��R�(KK��h�C4*   D   �   :  &      "   >  U     N        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CD!      R      �  "     �  (      
   3   6   Z          �t�bhhK ��h��R�(KK��h�C0     �     �     �  B   �          �t�bhhK ��h��R�(KK��h�C7        	         �t�bhhK ��h��R�(KK	��h�C$            �	     �        �t�bhhK ��h��R�(KK
��h�C(%   _  C   !  �        <         �t�bhhK ��h��R�(KK��h�Ct         O      �   Y      Q      �     x              +     &      F  +   "   H     t         �t�bhhK ��h��R�(KK��h�CT%     m  �            �  c           �     u      ~              �t�bhhK ��h��R�(KK��h�C4   �  
   b    T   %   A  y               �t�bhhK ��h��R�(KK��h�C�	     �t�bhhK ��h��R�(KK��h�C\               ;      �   %   �        
           6        �   �        �t�bhhK ��h��R�(KK��h�C,�   �   �  
   ,                     �t�bhhK ��h��R�(KK��h�C0w          h   p
        E           �t�bhhK ��h��R�(KK
��h�C(      E      5  	      	         �t�bhhK ��h��R�(KK��h�Cl   �   '   �     U  B   �      E                    �                                 �t�bhhK ��h��R�(KK��h�C4X  7     8        '   
      y           �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�CH      "     n      �   F     =            @   �   =        �t�bhhK ��h��R�(KK	��h�C$�      ,   �   
   4  	         �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�CT            �   !      @              A   �             m         �t�bhhK ��h��R�(KK��h�CD   e   '   �   �     �   9     �
  �     /      �         �t�bhhK ��h��R�(KK	��h�C$     9   �     K  A        �t�bhhK ��h��R�(KK��h�C�  �        	         �t�bhhK ��h��R�(KK��h�C!      �      	         �t�bhhK ��h��R�(KK��h�Cd�	     �     @      �        �     ,   	      	   K   	     	   �  	   �   	   >     �t�bhhK ��h��R�(KK��h�C      C      �t�bhhK ��h��R�(KK
��h�C(^            2   -   �           �t�bhhK ��h��R�(KK��h�CH
   $   �   N  (      #   !      \               $   k         �t�bhhK ��h��R�(KK��h�C�            �t�bhhK ��h��R�(KK
��h�C(�     j     �        �        �t�bhhK ��h��R�(KK��h�CH         E     �               0      �  4      �        �t�bhhK ��h��R�(KK	��h�C$[      V           	         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CD      �   V     v   :     (      �      �              �t�bhhK ��h��R�(KK��h�C4�  (     �   �   �        0   *  �         �t�bhhK ��h��R�(KK��h�Cd�         .   N         (   <         �  g      n      �        Q   �              �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C<   8   /            &      I           g        �t�bhhK ��h��R�(KK��h�C@[      �  q
     �     �  
     �   X     �         �t�bhhK ��h��R�(KK��h�C8�  �  �   �           "   B                  �t�bhhK ��h��R�(KK��h�C0D         �      )   2       �         �t�bhhK ��h��R�(KK��h�C\   .               B  /   �  �     A   �  Z  '        M   �      D         �t�bhhK ��h��R�(KK��h�C<�  !  �  
   ,                  �               �t�bhhK ��h��R�(KK��h�C4   �  �                          r
     �t�bhhK ��h��R�(KK��h�C .  M     �  ~            �t�bhhK ��h��R�(KK
��h�C(�     /         	      	         �t�bhhK ��h��R�(KK��h�CP%     �  �                      8        �   �              �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C              *	     �t�bhhK ��h��R�(KK��h�C8   ]   �              �     �     #        �t�bhhK ��h��R�(KK��h�C@              >     �      �  6  �   
   �        �t�bhhK ��h��R�(KK��h�CT      )   �  �   E      <    �   s              ^   �     s        �t�bhhK ��h��R�(KK��h�CT^   |      �         )   �           $   �        �     8   o         �t�bhhK ��h��R�(KK��h�Cl2      -   �     ;    j   3     ;    (      !   G      s
           s
                 �t�bhhK ��h��R�(KK��h�C�         �     �t�bhhK ��h��R�(KK��h�C p  �      5              �t�bhhK ��h��R�(KK��h�C E      �        	         �t�bhhK ��h��R�(KK��h�C	     Y      O      �t�bhhK ��h��R�(KK��h�Ce     n      �t�bhhK ��h��R�(KK��h�CT         /      &   �  +   �      �      |     <     "   X   �         �t�bhhK ��h��R�(KK��h�CH   X         z   
   �     �	     
   ,                     �t�bhhK ��h��R�(KK��h�C8               �     =        �   /         �t�bhhK ��h��R�(KK��h�C<
   �     ?      �     "         �     T        �t�bhhK ��h��R�(KK��h�Cx%               �   �       /      �  �     �     �      �  �     N  7      B        �         �t�bhhK ��h��R�(KK ��h�C�o         �	     >       �               %            (        0      �     �        �  "           �t�bhhK ��h��R�(KK��h�CH      ,  +        )   =      4         
   _      {         �t�bhhK ��h��R�(KK��h�C<      �   �   �                                �t�bhhK ��h��R�(KK��h�C<�
  �   �  �   "   @      X      e                �t�bhhK ��h��R�(KK��h�C<
            5     n     0   #   !      �        �t�bhhK ��h��R�(KK
��h�C(?     (     f   �  �            �t�bhhK ��h��R�(KK��h�C5         1  r      �t�bhhK ��h��R�(KK��h�Cx      ~         �     T  �  k      +                     �        %   l      ~         �         �t�bhhK ��h��R�(KK��h�CX      �  -   \         �  �           \      �  �         `            �t�bhhK ��h��R�(KK��h�CD�   >   -   �  0     �  �     x  �  �   g
              �t�bhhK ��h��R�(KK
��h�C(H  �   �     �   -   �   �         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C?     �     �t�bhhK ��h��R�(KK��h�CH         b         
  �         �              M        �t�bhhK ��h��R�(KK��h�Cs     �t�bhhK ��h��R�(KK��h�C   �         �t�bhhK ��h��R�(KK��h�CT                  �t�bhhK ��h��R�(KK��h�CH�        �  &   �     �   g   �  L             E         �t�bhhK ��h��R�(KK	��h�C$�  �         �   r	  r        �t�bhhK ��h��R�(KK��h�C8^   �         -   b      1     �      K        �t�bhhK ��h��R�(KK��h�C       +     -	     �t�bhhK ��h��R�(KK��h�C|   5   u     �   �      �      b     �         J   �   h      "
  �        >     (  p  
   ]  �        �t�bhhK ��h��R�(KK��h�C<T   (         �   ~  
   �   :        (   �        �t�bhhK ��h��R�(KK��h�Ct
           g     �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�CH�          �        ?           C  D     ,           �t�bhhK ��h��R�(KK��h�C,     �  �        �  
           �t�bhhK ��h��R�(KK*��h�C�            �     L  +      �  �     R            J   +
  `   �   �   �         0   !      �      D     [      �       :      ^  �        �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C4
   k     @     �	  �         �  �        �t�bhhK ��h��R�(KK���      h�C?           �t�bhhK ��h��R�(KK��h�C,  �      �   =	        �  �        �t�bhhK ��h��R�(KK��h�C                         �t�bhhK ��h��R�(KK	��h�C$�   �     �   �   �  �         �t�bhhK ��h��R�(KK��h�C0   �     �      (  �        B        �t�bhhK ��h��R�(KK	��h�C$         �  	      	         �t�bhhK ��h��R�(KK��h�CD*   D     
            �  \        �   �     �        �t�bhhK ��h��R�(KK��h�CH�     �  �  
   H   B   }   �   �         Y        =        �t�bhhK ��h��R�(KK��h�CR      �               �t�bhhK ��h��R�(KK��h�CT                              �  |     &      U   8   A
  �        �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�CD*      �      4              )   =         �   ~        �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C�              �t�bhhK ��h��R�(KK��h�C,"      �     �   (   D     g        �t�bhhK ��h��R�(KK��h�C�  
              �t�bhhK ��h��R�(KK��h�C@      �      B          �      V     v   :        �t�bhhK ��h��R�(KK��h�C4%         /  "   W      0      9   �         �t�bhhK ��h��R�(KK��h�C4I      J   6  C   I  ,      �              �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CH      F           �   &      *           �      �        �t�bhhK ��h��R�(KK��h�C      �	         �t�bhhK ��h��R�(KK��h�CP*               &      \  t      �     
   D
  V         l        �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�CY     �t�bhhK ��h��R�(KK
��h�C(   P    d   �
                 �t�bhhK ��h��R�(KK��h�C     r         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�Ct   $   2  �  �      �  �   Q
  (      U             �      �  T            �  �  �   _        �t�bhhK ��h��R�(KK��h�C�  
      �      �t�bhhK ��h��R�(KK
��h�C(�   �        I      �   �        �t�bhhK ��h��R�(KK��h�C1   #       m      4      �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CD      \  R  �
          5   !         }     o         �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�CD
        f     g  )        ?      !      @  R         �t�bhhK ��h��R�(KK��h�Ct
   3   6   I     +               ?      y  !      �        &   M   �      *                     �t�bhhK ��h��R�(KK��h�C`
               (      !      �     R           B   �     o      4  �         �t�bhhK ��h��R�(KK	��h�C$#  �   �   �  8	     �        �t�bhhK ��h��R�(KK*��h�C�         N     ]	  7   v     
   _      $   �        E
  +      f  �     �  
   �   �      �      r  �     "   >  )      L  �      +         �t�bhhK ��h��R�(KK��h�Cl   A     2   (       	     �     R      �  i      �  �   7      5   �  �    
            �t�bhhK ��h��R�(KK��h�CH�  �         ;      �     2     
   �   /      �  C         �t�bhhK ��h��R�(KK��h�CP|      �         �     �                              }        �t�bhhK ��h��R�(KK��h�CB          �t�bhhK ��h��R�(KK��h�C!      '        �t�bhhK ��h��R�(KK��h�C8�            �  ;            2  �   d        �t�bhhK ��h��R�(KK��h�Cl        /   P     �t�bhhK ��h��R�(KK
��h�C(%   /
     5                     �t�bhhK ��h��R�(KK	��h�C$   @   x  �     �   o         �t�bhhK ��h��R�(KK��h�C,      )   "           �            �t�bhhK ��h��R�(KK��h�C    (   #   !      �         �t�bhhK ��h��R�(KK��h�CB   e     �t�bhhK ��h��R�(KK��h�C4      �        )   w   u
  Q  $   �        �t�bhhK ��h��R�(KK��h�Cd�  &   *                                           �           �  �        �t�bhhK ��h��R�(KK��h�CH   �  '      H         3  C   
      �     ]     b         �t�bhhK ��h��R�(KK��h�CX      �   �      �	     6  
   �   �      �            2   j             �t�bhhK ��h��R�(KK��h�CD         v
     �
  �     %   l      v
  C              �t�bhhK ��h��R�(KK
��h�C(�        '  a        �        �t�bhhK ��h��R�(KK��h�C1   #       �  �         �t�bhhK ��h��R�(KK
��h�C(�        z  N                  �t�bhhK ��h��R�(KK��h�C\   �   %   B   }        �t�bhhK ��h��R�(KK
��h�C("     (      #   !               �t�bhhK ��h��R�(KK
��h�C(   ?   %   d	     ^   �   �        �t�bhhK ��h��R�(KK��h�C       �        T        �t�bhhK ��h��R�(KK��h�C �               r        �t�bhhK ��h��R�(KK��h�C@                  
       �         �   D        �t�bhhK ��h��R�(KK��h�C\         �     $  $   G
           `        0   x         O              �t�bhhK ��h��R�(KK��h�C   �  �     �t�bhhK ��h��R�(KK��h�CLf      �  "   >     
   �                 )                 �t�bhhK ��h��R�(KK��h�C<"               z   ,         
                  �t�bhhK ��h��R�(KK��h�CL7  (      N   �              Y       L  �     �  �        �t�bhhK ��h��R�(KK��h�CX      +         �  �      �                  k  �      %   �   .        �t�bhhK ��h��R�(KK��h�C �  $  �     $  �        �t�bhhK ��h��R�(KK��h�C@      P   !      �  
     
   ,                     �t�bhhK ��h��R�(KK��h�C�   >   `   �          �t�bhhK ��h��R�(KK��h�Cw
       �t�bhhK ��h��R�(KK��h�C8   �   �        �           Y      Q         �t�bhhK ��h��R�(KK��h�C0d   �   /     4     (   [               �t�bhhK ��h��R�(KK��h�Cr  �     L     �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C4�  
                 �       A        �t�bhhK ��h��R�(KK��h�C1   #       �        �t�bhhK ��h��R�(KK
��h�C(E  �               g            �t�bhhK ��h��R�(KK
��h�C(E  �               g            �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C ,     �  	      	         �t�bhhK ��h��R�(KK��h�C!   
         �t�bhhK ��h��R�(KK��h�C<1     �     �  !      .  '   
   �    _        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C�  p     �t�bhhK ��h��R�(KK��h�CL   �   �      5   `   3           �  8   �           �         �t�bhhK ��h��R�(KK��h�C%   �     6        �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C`S  G   H        �   �     S     $                    "   t      �           �t�bhhK ��h��R�(KK��h�C@   ?   !      �  
   F                    _        �t�bhhK ��h��R�(KK��h�C\   (      ~     H  *      R  4            *   $   �     Y      O   T        �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C8�        5   F  [      <      ;      �        �t�bhhK ��h��R�(KK��h�C@      �      L   �      �             \          �t�bhhK ��h��R�(KK��h�C@   (   #   !   
   3   6               Z  Y  �         �t�bhhK ��h��R�(KK��h�C8T   (         �   ~          (   8   4         �t�bhhK ��h��R�(KK��h�C �        	      	         �t�bhhK ��h��R�(KK��h�CA     �  Y  �      �t�bhhK ��h��R�(KK��h�C0�              	      	   K   	   �      �t�bhhK ��h��R�(KK��h�CDW      �  �   !      �  �   
   �  x
  y
        @         �t�bhhK ��h��R�(KK��h�C�      (     e      �t�bhhK ��h��R�(KK
��h�C(�   �        Z        i        �t�bhhK ��h��R�(KK��h�CH   %                    �   �  j      [    �            �t�bhhK ��h��R�(KK
��h�C(   (   �  3        �   �         �t�bhhK ��h��R�(KK��h�CL!           �   (      "   k     �  "   L     ~     p         �t�bhhK ��h��R�(KK��h�C�  �	  
   �        �t�bhhK ��h��R�(KK��h�C8      5   �  <            U   j  g  k        �t�bhhK ��h��R�(KK��h�C        �t�bhhK ��h��R�(KK��h�C@          _	     �t�bhhK ��h��R�(KK��h�C !      �
  	      	         �t�bhhK ��h��R�(KK
��h�C(*      �   �         �     V     �t�bhhK ��h��R�(KK��h�C,   �   �  *      �  �   $   E         �t�bhhK ��h��R�(KK	��h�C$   �         �   �           �t�bhhK ��h��R�(KK��h�C8   r  '  �   +      �  ;   R      $            �t�bhhK ��h��R�(KK��h�Cz
  �      �t�bhhK ��h��R�(KK��h�C�  k  �	         �t�bhhK ��h��R�(KK��h�CP      a  g      ]              -        <      �  
   Z        �t�bhhK ��h��R�(KK��h�C`#   !      )        �        �   d  ?      
   �   F      G                     �t�bhhK ��h��R�(KK��h�C8      J   �  �   &      =      G  G   t         �t�bhhK ��h��R�(KK��h�CD!      �   $   W                ?      
              �t�bhhK ��h��R�(KK��h�Cr  �     L     �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C8!         	      	      	   K   	   �   	        �t�bhhK ��h��R�(KK��h�C@   w  �      J  E      {     [     H              �t�bhhK ��h��R�(KK
��h�C(   A   {
  �      ,               �t�bhhK ��h��R�(KK��h�C8   (   !  )            ~   �      d           �t�bhhK ��h��R�(KK��h�C1        �         �t�bhhK ��h��R�(KK��h�C`      �  J   �   
   G   $   t        ?      #   !   
   3   6      �              �t�bhhK ��h��R�(KK��h�C4�  �   �   �     �	  �      �     q        �t�bhhK ��h��R�(KK��h�C   �	     �t�bhhK ��h��R�(KK��h�CL      �   F           �   &      j      �  ]      $           �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK
��h�C(   ]  �                       �t�bhhK ��h��R�(KK
��h�C(      �   �   �      ,   �         �t�bhhK ��h��R�(KK��h�C08     �       
      	      	         �t�bhhK ��h��R�(KK	��h�C$�   R   
      	      	         �t�bhhK ��h��R�(KK��h�C8*      ]              (         o  �        �t�bhhK ��h��R�(KK��h�C,   e   M  w     I        J        �t�bhhK ��h��R�(KK��h�C,�     f   W  V   �    
            �t�bhhK ��h��R�(KK��h�C |  �           �         �t�bhhK ��h��R�(KK��h�C        �t�bhhK ��h��R�(KK	��h�C$            r     �        �t�bhhK ��h��R�(KK��h�CD�   �  >      A     �  Y  �         K        �        �t�bhhK ��h��R�(KK��h�CT      -   t     �  �                 .      �     �	     �         �t�bhhK ��h��R�(KK	��h�C$L     }       `   �        �t�bhhK ��h��R�(KK��h�Ch   �  �     R   
   y        �  �  `   3     �     B        �     �	     
        �t�bhhK ��h��R�(KK��h�C�                �t�bhhK ��h��R�(KK��h�C0      =      4   
   �      �   �         �t�bhhK ��h��R�(KK��h�C\   �  �   Y     �t�bhhK ��h��R�(KK��h�C4     o     e      �        :   @         �t�bhhK ��h��R�(KK!��h�C�
   H   �  J   2      %   e              B         L  
   �     �      -   �
  �   �   B      "   T     �         �t�bhhK ��h��R�(KK��h�CLA     �  �  �  e                                         �t�bhhK ��h��R�(KK��h�C0      �         j   4      .             �t�bhhK ��h��R�(KK��h�C0
   �  �     �        Z     +         �t�bhhK ��h��R�(KK��h�C8   �   �  �  �   I      �   ~      �   n         �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�CL      �  w   �        `           ;             L         �t�bhhK ��h��R�(KK��h�CK     �t�bhhK ��h��R�(KK��h�C,�  �     L         �     n         �t�bhhK ��h��R�(KK	��h�C$%   �   p   h   H   B   3        �t�bhhK ��h��R�(KK��h�C        �t�bhhK ��h��R�(KK	��h�C$�        �  i   h          �t�bhhK ��h��R�(KK��h�CdW         S   �            :        �   �	     �           |
     @     �         �t�bhhK ��h��R�(KK��h�CH           I      2   5      M      C            �         �t�bhhK ��h��R�(KK��h�C,   6     x               }
        �t�bhhK ��h��R�(KK��h�C41   #      �   �  
   3   6        u        �t�bhhK ��h��R�(KK��h�CP�   �   z  �   l   �   :	  7               �     �  q              �t�bhhK ��h��R�(KK��h�CH         M        �t�bhhK ��h��R�(KK��h�C�   c     �t�bhhK ��h��R�(KK��h�C8      �   f        #   i      H   A   �        �t�bhhK ��h��R�(KK��h�C81   #      X     k   
   3   6   2              �t�bhhK ��h��R�(KK��h�CT/      ;         C  �  �        *   2     �      �     -  �         �t�bhhK ��h��R�(KK��h�C        e      @         �t�bhhK ��h��R�(KK��h�C0   '   
   f   �     
         y        �t�bhhK ��h��R�(KK	��h�C$e            6  �  ?        �t�bhhK ��h��R�(KK��h�C`�   5     7  �        �     /   9   -     %   8           �   �      �         �t�bhhK ��h��R�(KK��h�C,         =      �  4               �t�bhhK ��h��R�(KK��h�C0      #   !      j  
   3   6            �t�bhhK ��h��R�(KK��h�Cl      �    �   e  i   
   N                   j        M   �                       �t�bhhK ��h��R�(KK��h�C<u  *        ?      )   
   -     .  /  F   *
     �t�bhhK ��h��R�(KK$��h�C�@     �  "   ~  y     e   �   �  �           $     5   <           �        .   "   �      m      �     Q  m         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CP�  b     �   �     I   /      �     �    }          >        �t�bhhK ��h��R�(KK��h�C0O     `  �   x      D     �   �        �t�bhhK ��h��R�(KK��h�C0   f
  �                 B  *        �t�bhhK ��h��R�(KK��h�C      �   ^     �t�bhhK ��h��R�(KK��h�C8/      -    
      9     "   7     �        �t�bhhK ��h��R�(KK��h�Cl            �  �                      �      P      p      :          �           �t�bhhK ��h��R�(KK��h�C,z  +      �     |      <  �        �t�bhhK ��h��R�(KK��h�C E         	      	         �t�bhhK ��h��R�(KK��h�C<      �  �     �     x	     P     %   w	        �t�bhhK ��h��R�(KK��h�CH      5      ~     {            0      ~  )   
   2        �t�bhhK ��h��R�(KK��h�CD        Q  
     �     �                 �        �t�bhhK ��h��R�(KK��h�Cd   H      '         V   2   (   Y
  !                  \   2   &   J  C      �        �t�bhhK ��h��R�(KK��h�C@      5      &     &      �  ]   *      �  �        �t�bhhK ��h��R�(KK��h�C@   D              �     �  �        A   }         �t�bhhK ��h��R�(KK
��h�C(�  �                Z        �t�bhhK ��h��R�(KK��h�C4X  7     8        '   
      y           �t�bhhK ��h��R�(KK
��h�C(
   H   [  '   -   A      �	        �t�bhhK ��h��R�(KK��h�CH   r       �   \   �                   �     �         �t�bhhK ��h��R�(KK��h�CX�     /   9   �  7      "   m      �      �  0   <   "   C     �           �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C0      -   �   �      E   "      �        �t�bhhK ��h��R�(KK��h�Cm
  �               �t�bhhK ��h��R�(KK
��h�C(   &   N   M     �     �	        �t�bhhK ��h��R�(KK��h�CP
   u  F   '      H     %        B  �      *         �   �         �t�bhhK ��h��R�(KK��h�Cu     �t�bhhK ��h��R�(KK��h�C<
   H   �  [  '      H   u  *     &     0        �t�bhhK ��h��R�(KK��h�CD�     �  �   �     *   �              �     �        �t�bhhK ��h��R�(KK
��h�C(6  �   �   -   
         K         �t�bhhK ��h��R�(KK��h�C�  :   ?  �  Y      �t�bhhK ��h��R�(KK��h�C,b   
   �  
     y     &   R        �t�bhhK ��h��R�(KK��h�C \        	      	         �t�bhhK ��h��R�(KK	��h�C$      -   U   $   �   N        �t�bhhK ��h��R�(KK��h�C	  �               �t�bhhK ��h��R�(KK
��h�C(�     2                �      �t�bhhK ��h��R�(KK��h�CD   (   !         "   k     �  "   L     ~     p         �t�bhhK ��h��R�(KK��h�C4d  �     �     8     �     `          �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�C �     *        �        �t�bhhK ��h��R�(KK��h�C,   W  �  '   "   ~  y     e         �t�bhhK ��h��R�(KK��h�C  �   X     �t�bhhK ��h��R�(KK��h�C0   2   �   �         [     d   �        �t�bhhK ��h��R�(KK��h�C8       �t�bhhK ��h��R�(KK��h�C]     �t�bhhK ��h��R�(KK��h�C4      �     >   2   w   �   L               �t�bhhK ��h��R�(KK��h�Cx
   3   6   I     +               ?      y  !        A   �     �  M   �      y                     �t�bhhK ��h��R�(KK��h�CD      
      �    �  �      �      %   s               �t�bhhK ��h��R�(KK	��h�C$     9   �       A        �t�bhhK ��h��R�(KK��h�C�   �         	         �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK
��h�C(f   �  �   c  X  �     u         �t�bhhK ��h��R�(KK��h�C"     �t�bhhK ��h��R�(KK��h�C�  =  �  {     �t�bhhK ��h��R�(KK��h�C02      -   P   �   j   7	        �	        �t�bhhK ��h��R�(KK��h�CT�     �      �  *           g                    �   �           �t�bhhK ��h��R�(KK��h�CX   9
  �  �                     �   �               ,   �      G        �t�bhhK ��h��R�(KK
��h�C(      
     *  �   
   $        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK
��h�C(\   +  :  W    
   +   w         �t�bhhK ��h��R�(KK��h�C4�            S        .  M  �     T     �t�bhhK ��h��R�(KK	��h�C$
	     	      	      	   K      �t�bhhK ��h��R�(KK��h�C0@   �           �      �	     Z        �t�bhhK ��h��R�(KK��h�C       �      �  �        �t�bhhK ��h��R�(KK��h�C8"   m      �  /      -  �      .   /  i        �t�bhhK ��h��R�(KK��h�C    &   �        
        �t�bhhK ��h��R�(KK��h�CLg   z  U  w        
                 �  �  �               �t�bhhK ��h��R�(KK��h�C*         `   �      �t�bhhK ��h��R�(KK	��h�C$�  ?      
   X   �   F         �t�bhhK ��h��R�(KK
��h�C(   �  
   ,                     �t�bhhK ��h��R�(KK��h�CL      �               P   �         �      0     :            �t�bhhK ��h��R�(KK��h�Cth   Y            x     #     $     �     >   2   P   H        Q         O     2   �   �         �t�bhhK ��h��R�(KK��h�CT      0   �     �  >      u
  P   �      N         M   ~     �         �t�bhhK ��h��R�(KK��h�C\      �  �        E      �   �           %         �  u  �   �	           �t�bhhK ��h��R�(KK��h�C<�  �   �  <      �      �     E     A   !        �t�bhhK ��h��R�(KK	��h�C$  I   �     �     �        �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK
��h�C(�   �  �  "   �   �  0  ;        �t�bhhK ��h��R�(KK
��h�C(]   �           
   �   F         �t�bhhK ��h��R�(KK��h�CX              4         �  �   �   �   g            V  �   $     �     �t�bhhK ��h��R�(KK��h�C      �	         �t�bhhK ��h��R�(KK��h�CL      t     W     �     �      M   �      �   �     �        �t�bhhK ��h��R�(KK��h�CD`  �  =     X      H   �              -     .        �t�bhhK ��h��R�(KK��h�C0�   v     .            
  f   �        �t�bhhK ��h��R�(KK��h�C8      E      �     �  &     T   E   L        �t�bhhK ��h��R�(KK��h�C~
     �t�bhhK ��h��R�(KK��h�CX�     r  '  L     U           )      �      �   �      L     +         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C@     �     �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C8�  >        �        2   �  �   �   �        �t�bhhK ��h��R�(KK��h�Cp         $           �  b     6
        P  �  M
        P   �   @           G   W         �t�bhhK ��h��R�(KK��h�C|      <       �      �t�bhhK ��h��R�(KK��h�CH@   �      *  X     �   �   �     .   p      �     �         �t�bhhK ��h��R�(KK��h�C@   %
  �     �     !  o      o      �     E        �t�bhhK ��h��R�(KK	��h�C$Y     p                    �t�bhhK ��h��R�(KK��h�C4      5     &      �   U   $   �   N        �t�bhhK ��h��R�(KK��h�C+  2  {  h           �t�bhhK ��h��R�(KK��h�C,   �  
   `   �   
   ,               �t�bhhK ��h��R�(KK��h�C|           $   �         +   
   _      8             d     x      1  �   <           c           �t�bhhK ��h��R�(KK��h�C4�   a  2      .                          �t�bhhK ��h��R�(KK��h�C4      =                  :              �t�bhhK ��h��R�(KK��h�CZ  	         �t�bhhK ��h��R�(KK��h�C0)   %   6        [  �      0   <         �t�bhhK ��h��R�(KK��h�C<�     o           �	  �     !     u  *        �t�bhhK ��h��R�(KK��h�CXW  �     =      �  4      �      \  L   y              B    c         �t�bhhK ��h��R�(KK��h�C?     F     �t�bhhK ��h��R�(KK��h�C<*      �   �    7      �      �   �   �  b        �t�bhhK ��h��R�(KK
��h�C([      R     D  n               �t�bhhK ��h��R�(KK��h�C<   e   '              �         �              �t�bhhK ��h��R�(KK
��h�C(!      �        	      	         �t�bhhK ��h��R�(KK��h�C 3        (     ]  p      �t�bhhK ��h��R�(KK	��h�C$#           	      	         �t�bhhK ��h��R�(KK��h�C,      #   !   
   3   6      p         �t�bhhK ��h��R�(KK��h�C@         �  
   ,      "   >  )   
                  �t�bhhK ��h��R�(KK��h�C        O      �t�bhhK ��h��R�(KK
��h�C("   f        B   �   B   <        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�CX      �   u               :  �     �   p     �      -  p              �t�bhhK ��h��R�(KK��h�C4�         �  $   A     p                  �t�bhhK ��h��R�(KK��h�CX   5      =   �     Q     j   W   �   c                        �        �t�bhhK ��h��R�(KK��h�C,   f   ?     P  �  )   
           �t�bhhK ��h��R�(KK��h�C�     �  m      �t�bhhK ��h��R�(KK��h�C[      �      �t�bhhK ��h��R�(KK��h�C8      J         )        
     5           �t�bhhK ��h��R�(KK��h�CH   �   n     %   �   �                 �   -   
            �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�CR     	         �t�bhhK ��h��R�(KK��h�C<         	         �t�bhhK ��h��R�(KK��h�C   �   '   s   �         �t�bhhK ��h��R�(KK��h�C@W   \           ;      ,     
        $   E         �t�bhhK ��h��R�(KK��h�CP�  
   ,               �
  �     ,            X        A   }      �t�bhhK ��h��R�(KK��h�Cr  �     �t�bhhK ��h��R�(KK��h�Ch      '            �      &   I            �        a      �      M     �           �t�bhhK ��h��R�(KK��h�C&     �t�bhhK ��h��R�(KK	��h�C$   J    
   _              �t�bhhK ��h��R�(KK1��h�C�      z   "   �   B   �      �   n     7  �
        �        7  �	        ]              �        �
        �     �             #	        G	                 �t�bhhK ��h��R�(KK��h�Ct      �     �     �     S              '      .      7     !
     j        �   �   �        �t�bhhK ��h��R�(KK��h�C      �  	      	         �t�bhhK ��h��R�(KK��h�C            ^     �t�bhhK ��h��R�(KK��h�C@   ?   #   !      �  <   
   3   6   �
        1  r      �t�bhhK ��h��R�(KK��h�C8      �
        Y      @           @        �t�bhhK ��h��R�(KK��h�CL   f   �
     2   �   0   �   
            2                     �t�bhhK ��h��R�(KK��h�C,%   �   �  �
     �         �        �t�bhhK ��h��R�(KK��h�C     �      u      �t�bhhK ��h��R�(KK��h�C     �             �t�bhhK ��h��R�(KK��h�Cz  F     �     �t�bhhK ��h��R�(KK��h�C         !           �t�bhhK ��h��R�(KK��h�C   5  �     �        �t�bhhK ��h��R�(KK
��h�C(%   �  [   �   2         >        �t�bhhK ��h��R�(KK��h�C4$   �   5   J     �             �        �t�bhhK ��h��R�(KK
��h�C(1   #       �     /      �         �t�bhhK ��h��R�(KK��h�C8   �        .   �   �       _             �t�bhhK ��h��R�(KK��h�CH�  �        �  V      (      �      8   o        �
        �t�bhhK ��h��R�(KK
��h�C(!      �        	      	         �t�bhhK ��h��R�(KK	��h�C$      -   U   �     �        �t�bhhK ��h��R�(KK��h�C0      )   b      x   
   7
     u         �t�bhhK ��h��R�(KK��h�C`7      �              
      �  @         
   ,         "  q   �  "           �t�bhhK ��h��R�(KK��h�CD�  (         .   
   _           }     d     �        �t�bhhK ��h��R�(KK��h�C/      �     �t�bhhK ��h��R�(KK��h�C\   '   )   �              0            ~   �               �     3        �t�bhhK ��h��R�(KK��h�C4   &      w  -   v   %   �	  o
              �t�bhhK ��h��R�(KK��h�C�  
      �	     �t�bhhK ��h��R�(KK��h�C,�        �                        �t�bhhK ��h��R�(KK��h�C,            �
  \                 �t�bhhK ��h��R�(KK��h�Cd   7  S      o     8   �  -  �  �   7  :   .        �  9   %     �  �   �        �t�bhhK ��h��R�(KK��h�CX      J         )   R  D   
   �   S   y  h   @      g       �           �t�bhhK ��h��R�(KK	��h�C$            	      	         �t�bhhK ��h��R�(KK	��h�C$1   #       �  g     �        �t�bhhK ��h��R�(KK��h�CP      �        `        �      x     +   
   _                  �t�bhhK ��h��R�(KK��h�Cd�  �      v  	  l      
   _      �   �     �   \  5   <         �     �           �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C,      �  �        ;         �     �t�bhhK ��h��R�(KK	��h�C$�       �      �     9     �t�bhhK ��h��R�(KK��h�C<#   !      �          ?      
   3   6   �        �t�bhhK ��h��R�(KK��h�Cl         	  i     7            P   n   G         r                                   �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�C\   /     o  4   r      �t�bhhK ��h��R�(KK��h�CD$   �     T        :  "      �        �              �t�bhhK ��h��R�(KK��h�C0      �     4  �        �  )        �t�bhhK ��h��R�(KK��h�C[      �  	         �t�bhhK ��h��R�(KK��h�C`                     �
  �   O      j         -   a   
     ,      
   E         �t�bhhK ��h��R�(KK��h�C<   �     �  �        �  [         �  -        �t�bhhK ��h��R�(KK��h�C4#   !      �     �  ?      
   �   F         �t�bhhK ��h��R�(KK��h�C         	      	         �t�bhhK ��h��R�(KK��h�C 
        r  $  �        �t�bhhK ��h��R�(KK��h�C@      �                 &      �      �  E         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C8      -   �  +              <  =           �t�bhhK ��h��R�(KK��h�C8%   �     V  
            �      I   �        �t�bhhK ��h��R�(KK��h�C@
   C     d   |  �      D   (      <         5         �t�bhhK ��h��R�(KK��h�C<   ?   #   !            %   �     
   $  F         �t�bhhK ��h��R�(KK��h�C\
      (      -   !      \   �        :     *               �     �        �t�bhhK ��h��R�(KK��h�C        �  �        �t�bhhK ��h��R�(KK	��h�C$�	        >     X  �        �t�bhhK ��h��R�(KK��h�C0p           j              4        �t�bhhK ��h��R�(KK��h�C0q      [  \   H   E     �     u        �t�bhhK ��h��R�(KK��h�CD%            :      .          ,     H   �  q        �t�bhhK ��h��R�(KK��h�C,
   )        �                    �t�bhhK ��h��R�(KK��h�C<1   #       F     �     �     /   �              �t�bhhK ��h��R�(KK��h�C8O      A   ?  >   )  C   �  "   |      �         �t�bhhK ��h��R�(KK��h�C   	  	      	         �t�bhhK ��h��R�(KK��h�CX         �  �  
   _      �   �  q     �
  �   e     P   H              �t�bhhK ��h��R�(KK��h�C�  a            �t�bhhK ��h��R�(KK��h�Ck            �t�bhhK ��h��R�(KK��h�C0   P           +   b  �              �t�bhhK ��h��R�(KK
��h�C(      )   }     P     t         �t�bhhK ��h��R�(KK��h�C�     d   �  r      �t�bhhK ��h��R�(KK��h�C<#   !      /   "   �   '   
   3   6   �  "   �         �t�bhhK ��h��R�(KK
��h�C(c     |        q             �t�bhhK ��h��R�(KK��h�CT         J   $  �  w                       	  �        +         �t�bhhK ��h��R�(KK��h�C �    �  c   
   :        �t�bhhK ��h��R�(KK��h�CD   r  '           �   +      �     R      $            �t�bhhK ��h��R�(KK��h�C4)   �   f     g        �   �
  "   �        �t�bhhK ��h��R�(KK	��h�C$   �   9        �          �t�bhhK ��h��R�(KK��h�C0�     �      �  �        d  �        �t�bhhK ��h��R�(KK��h�C,?     �        �                  �t�bhhK ��h��R�(KK��h�C�     �         �t�bhhK ��h��R�(KK��h�C<   S        l           	     �              �t�bhhK ��h��R�(KK��h�C@      J   �      �         5         4      �         �t�bhhK ��h��R�(KK��h�C,K       a  �      �     �        �t�bhhK ��h��R�(KK��h�C4�      L   �   �   
   N     �               �t�bhhK ��h��R�(KK
��h�C(2           �  i   �  h        �t�bhhK ��h��R�(KK)��h�C��           �     	           V   l                  C  V  (   [      <      
   �        F   ?      �     �        d              �t�bhhK ��h��R�(KK��h�C4�  �   �      �     �  
   ,               �t�bhhK ��h��R�(KK��h�C
   ,         �t�bhhK ��h��R�(KK��h�C@   k     �t�bhhK ��h��R�(KK��h�C,k     �  �   �  �  T   �            �t�bhhK ��h��R�(KK	��h�C$Y        |  �  �     9     �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�CL      4  $   ;      e        ]  L         w         �
        �t�bhhK ��h��R�(KK��h�C,      �     f     $   E            �t�bhhK ��h��R�(KK��h�CDT   >         $   E           $   !   T     q   i
        �t�bhhK ��h��R�(KK��h�C<      >   i     �  
   w     �   �   k  L         �t�bhhK ��h��R�(KK��h�C4]   �     2      #     #                 �t�bhhK ��h��R�(KK��h�C 1   #       /   "   �         �t�bhhK ��h��R�(KK��h�CDd  -   
           `         �  �        %            �t�bhhK ��h��R�(KK��h�C8      ?      #   !   
        @   g           �t�bhhK ��h��R�(KK&��h�C�y      �      @  &      =      %   A               ;            .   
     �     �     �     �     �     �     (           �t�bhhK ��h��R�(KK��h�C�  
   ,   9     �t�bhhK ��h��R�(KK��h�C�              �t�bhhK ��h��R�(KK��h�C~     �t�bhhK ��h��R�(KK��h�C "   H   `  '   h  W        �t�bhhK ��h��R�(KK��h�C0   �     �	     �        0   4         �t�bhhK ��h��R�(KK��h�C0i           �               -         �t�bhhK ��h��R�(KK
��h�C(   D   ;      �     �  �        �t�bhhK ��h��R�(KK��h�C4K     �     :   �       �               �t�bhhK ��h��R�(KK��h�C0
   C        �    |     %   �         �t�bhhK ��h��R�(KK
��h�C(   &   �   �  $   �   |  �        �t�bhhK ��h��R�(KK��h�C4:    c   ^     �     D   �  N  7         �t�bhhK ��h��R�(KK��h�C<   Y      z  '   �     V   2      ~  i           �t�bhhK ��h��R�(KK��h�C<l  E   �   s   o  �   7      
   �     
           �t�bhhK ��h��R�(KK��h�CP           s        �  �      {   j        9   @     �        �t�bhhK ��h��R�(KK
��h�C(   (      ,
     �     �         �t�bhhK ��h��R�(KK��h�C#  &   �   �   r      �t�bhhK ��h��R�(KK��h�C,      �      n	  
   $   �   N        �t�bhhK ��h��R�(KK��h�CP   I   3     �                 �  3     5         �   ,        �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�CZ      �      �     �t�bhhK ��h��R�(KK��h�CH
   @   �   F   ?      !      l     @         �
     @         �t�bhhK ��h��R�(KK��h�C �  ?      
   j  F         �t�bhhK ��h��R�(KK��h�CT                     '     `           2     �   S   
   �         �t�bhhK ��h��R�(KK��h�C0�     
   �     �   f   _     �        �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C\4  �   �     .      �     	           �     �     %   �  !  j   <         �t�bhhK ��h��R�(KK��h�C@*      t       i        �       �   $   |        �t�bhhK ��h��R�(KK
��h�C(2   D          *   �  l        �t�bhhK ��h��R�(KK"��h�C�      J   H  �           F  +           &      a      �         u
  o         �           �     �  �        �t�bhhK ��h��R�(KK��h�CA   4            �t�bhhK ��h��R�(KK��h�C0      )   J  +      !                 �t�bhhK ��h��R�(KK��h�C,      �  �   .  M     k  #        �t�bhhK ��h��R�(KK��h�C0   �  m  �   7         m  s   7         �t�bhhK ��h��R�(KK��h�C01   #         �   
   3   6      �         �t�bhhK ��h��R�(KK��h�C<
   3   6      '   #   !      �                     �t�bhhK ��h��R�(KK��h�CH#   !      �     X   ?      
   X   �      g        F         �t�bhhK ��h��R�(KK��h�C�   x  "      .          �t�bhhK ��h��R�(KK��h�C4!      �     k  ?      
   3   6            �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�CL      J   a   #   !      R      �        U   0                 �t�bhhK ��h��R�(KK��h�C1   #       �      �t�bhhK ��h��R�(KK��h�C C     ;        �         �t�bhhK ��h��R�(KK��h�CX   2            O        2   �   Y  �  -   "      {        �
           �t�bhhK ��h��R�(KK��h�C4�         �  �   E      %  ^   �  F         �t�bhhK ��h��R�(KK��h�C4%      )   i  w     .         �   5        �t�bhhK ��h��R�(KK��h�CD-     b        S  u  �     �     l      �  b        �t�bhhK ��h��R�(KK��h�C      b         *      �t�bhhK ��h��R�(KK��h�C0      }     o           8   �         �t�bhhK ��h��R�(KK��h�C,      �     �         �           �t�bhhK ��h��R�(KK��h�C        9            �t�bhhK ��h��R�(KK
��h�C(  �         �   �              �t�bhhK ��h��R�(KK/��h�C�            O         Y      Q      Q     Q           t        O         �  Q         �               z      E  �
     �     >      v         :        �t�bhhK ��h��R�(KK��h�C$   k   �              �t�bhhK ��h��R�(KK��h�CL      �        5   <   �        U      W                   �t�bhhK ��h��R�(KK	��h�C$P     O  &   �  
   c        �t�bhhK ��h��R�(KK��h�C<#   !      �     e      @   ?      
      _        �t�bhhK ��h��R�(KK��h�C,     �     �  �
     ,   	         �t�bhhK ��h��R�(KK��h�C<      �  �     r  �     L     +   "   l        �t�bhhK ��h��R�(KK��h�C<
   �     m              2   &   D  *  !	        �t�bhhK ��h��R�(KK��h�C8*      �      �   �  `                        �t�bhhK ��h��R�(KK��h�Ch   �  n  5   �      3              �              �                     �         �t�bhhK ��h��R�(KK
��h�C(   �  E  &      �   j  /        �t�bhhK ��h��R�(KK"��h�C�   &   �
     �  �      h        7       l            7              �      %   l      S	           7        �t�bhhK ��h��R�(KK��h�Cd!      x      �         0   <      B   �  m      �  ?      
   3   6   �     �        �t�bhhK ��h��R�(KK	��h�C$�	  �     �  	      	         �t�bhhK ��h��R�(KK��h�C,1   #      o  
   T  Y      O         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C         	         �t�bhhK ��h��R�(KK��h�CHR  M  �   /      �   B   .
     _     �     �
             �t�bhhK ��h��R�(KK��h�CT   �  c                           �      �           :            �t�bhhK ��h��R�(KK��h�C4   "   �     �   �      ,   �   
            �t�bhhK ��h��R�(KK��h�C             �t�bhhK ��h��R�(KK	��h�C$   X   '   �                  �t�bhhK ��h��R�(KK��h�C0   �                        =         �t�bhhK ��h��R�(KK��h�C            �        �t�bhhK ��h��R�(KK	��h�C$I   m  &   �  ~	     �        �t�bhhK ��h��R�(KK��h�C�            �t�bhhK ��h��R�(KK��h�C   �   �   �     �t�bhhK ��h��R�(KK��h�C0d         �            j   d   �         �t�bhhK ��h��R�(KK	��h�C$�     �  =  Z     8   E     �t�bhhK ��h��R�(KK��h�C,*           t   &      M      +      �t�bhhK ��h��R�(KK��h�C   �   �     �t�bhhK ��h��R�(KK'��h�C�   (   �                 a  �   �   �     �	  �   $                 �  �     �   �                     D  *         H        �t�bhhK ��h��R�(KK��h�C8      �  v    �   M     p                 �t�bhhK ��h��R�(KK��h�C0q     �     �  	      	      	   K      �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C,   �           A        9	        �t�bhhK ��h��R�(KK��h�C     G           �t�bhhK ��h��R�(KK��h�CI  �     �           �t�bhhK ��h��R�(KK��h�CD      5      !  �  S           U      O	     �        �t�bhhK ��h��R�(KK��h�C #   !   ?      
           �t�bhhK ��h��R�(KK��h�C,%      �  �     I        4        �t�bhhK ��h��R�(KK��h�C@      �      d  
     }      J   F     8   /         �t�bhhK ��h��R�(KK��h�C0r                �  y   A           �t�bhhK ��h��R�(KK
��h�C(!      �	     >  	      	         �t�bhhK ��h��R�(KK��h�C�   p      �t�bhhK ��h��R�(KK��h�C=           �t�bhhK ��h��R�(KK��h�C g              �        �t�bhhK ��h��R�(KK��h�C)  	      	         �t�bhhK ��h��R�(KK��h�C4      2     �
  ^        M  *           �t�bhhK ��h��R�(KK��h�C�      �           �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C   i     �t�bhhK ��h��R�(KK��h�C   M  �     �t�bhhK ��h��R�(KK��h�Ct�  �  �   �      <         �  �   o   
   ,                  K      �      �      /     �        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK
��h�C()                    �         �t�bhhK ��h��R�(KK��h�C4.  h   (  �     �     /      �   ^        �t�bhhK ��h��R�(KK��h�C4=
                �      �      7         �t�bhhK ��h��R�(KK��h�C0   �  �   �   l         }     <        �t�bhhK ��h��R�(KK��h�CL   @   '   �  "     V   l      G        j   �      0            �t�bhhK ��h��R�(KK��h�CX   b  �  5         �
           (      .   :              �   

        �t�bhhK ��h��R�(KK��h�C@   �  �        �  v  �     �      �  �           �t�bhhK ��h��R�(KK��h�C@         @	  
   h              �      I  �         �t�bhhK ��h��R�(KK��h�CL   K        ~      D   �   J        K  G   %  D   ~   �        �t�bhhK ��h��R�(KK	��h�C$,      A   }         �         �t�bhhK ��h��R�(KK��h�CH   ?   !         �   f  
   3   �  
  �       �   �        �t�bhhK ��h��R�(KK��h�C   +   
   	     �t�bhhK ��h��R�(KK��h�C`   8   �  ,  �   �                              �  +      �  �  8   s        �t�bhhK ��h��R�(KK��h�C�  �         �t�bhhK ��h��R�(KK��h�C8%      ,     �     0	     h   p
     �        �t�bhhK ��h��R�(KK��h�C@         �         �   �         )   U   �            �t�bhhK ��h��R�(KK��h�C<         �   Z
     �         /   9   s   7         �t�bhhK ��h��R�(KK��h�C,l        W     �  D   ~            �t�bhhK ��h��R�(KK��h�C0   n  I   �  x  �   )   �   
            �t�bhhK ��h��R�(KK��h�Cq          �t�bhhK ��h��R�(KK	��h�C$     r  �                  �t�bhhK ��h��R�(KK��h�C4   S   "         
   �        �            �t�bhhK ��h��R�(KK��h�C,4         �     �      7   �        �t�bhhK ��h��R�(KK��h�C[   "     m      �t�bhhK ��h��R�(KK��h�C8�   �  !      �        '   
   3   6   �
        �t�bhhK ��h��R�(KK��h�C\)           +      H   �  w  
      (  %   �  �            ,               �t�bhhK ��h��R�(KK��h�CPr        %  t  (            �   (        
   _      �   F        �t�bhhK ��h��R�(KK��h�C3     	      	         �t�bhhK ��h��R�(KK��h�CX�  �                  8     Y            �         l  �     /         �t�bhhK ��h��R�(KK��h�C,   �    
   \   �  8   �           �t�bhhK ��h��R�(KK
��h�C(b   #         "   8   �   9        �t�bhhK ��h��R�(KK��h�C,        �  �     f   A   �         �t�bhhK ��h��R�(KK��h�CP      O      S   Q   i   %     z     Y      z     �     x        �t�bhhK ��h��R�(KK
��h�C(�  +      f  �  "   �      (     �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�Cb     	     �t�bhhK ��h��R�(KK��h�CDu   (   <      �  "   �   �           |      �            �t�bhhK ��h��R�(KK��h�C@;      �     �     \	        T   2   �    7         �t�bhhK ��h��R�(KK��h�CZ                  �t�bhhK ��h��R�(KK	��h�C$�   S  *      �     E         �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK��h�C8         P         c  c        J  E         �t�bhhK ��h��R�(KK ��h�C�   �         �        \   �   &   f  �   �        �     �     ;  �           J   �                    �t�bhhK ��h��R�(KK��h�CDV      �  �
  �   �     d  
        %      $           �t�bhhK ��h��R�(KK��h�CO
  B  �        �t�bhhK ��h��R�(KK��h�C   9       	         �t�bhhK ��h��R�(KK��h�C8   �  V   8   4   t	     �t�bhhK ��h��R�(KK	��h�C$   J    
   _              �t�bhhK ��h��R�(KK	��h�C$1   #       m      �      �     �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C0�                 �                 �t�bhhK ��h��R�(KK��h�C8�        u  F     l         �    7         �t�bhhK ��h��R�(KK��h�C�  b     �t�bhhK ��h��R�(KK��h�C4�  �   H  �      .   "            y        �t�bhhK ��h��R�(KK	��h�C$p  L     t      �           �t�bhhK ��h��R�(KK��h�C<W            �   +     G  �   #   i   �   �         �t�bhhK ��h��R�(KK��h�C<{         P        ,     �      j   D  2        �t�bhhK ��h��R�(KK��h�C,B  
     F     �         �        �t�bhhK ��h��R�(KK��h�C �     �      �   <         �t�bhhK ��h��R�(KK��h�C:     �        �t�bhhK ��h��R�(KK��h�C     �      9        �t�bhhK ��h��R�(KK��h�C_     �         �t�bhhK ��h��R�(KK��h�C0�   /      ;         \     �           �t�bhhK ��h��R�(KK��h�CD                          �  &      9      v        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK
��h�C(h      �   �      p     �        �t�bhhK ��h��R�(KK��h�C`      '   �   �   |        :         C  8  (  ]      �   �      �
  �   d        �t�bhhK ��h��R�(KK
��h�C(^     !     �  	      	         �t�bhhK ��h��R�(KK	��h�C$           j	  �  �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C`w  3        �        �   y  �      u            S   a             ?        �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C �         0   %           �t�bhhK ��h��R�(KK��h�C@      &   4           �   >      M   �      �          �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C �
     H   �     �        �t�bhhK ��h��R�(KK��h�Cd�          .   N   B   
        �   �           �     V                        �t�bhhK ��h��R�(KK��h�C,�     |  ?      
   X   �   F         �t�bhhK ��h��R�(KK��h�Cd   .   �      4   
   _      �  #   =  ;      �   i      �      �  
   _      �         �t�bhhK ��h��R�(KK	��h�C$�  �  '  O  7   �           �t�bhhK ��h��R�(KK��h�Cx      -   �   j   �        c     $   |     �       �      �     ?     l
  �      9     W        �t�bhhK ��h��R�(KK��h�C0%   �  @  :         �                 �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�CX      �   H      �      �   *             �      %   !  (      n         �t�bhhK ��h��R�(KK��h�C@      B
  �     
   �   �   *        x  +   f	        �t�bhhK ��h��R�(KK��h�C4{   �   +   w  {  ;         �   �            �t�bhhK ��h��R�(KK��h�C	     �t�bhhK ��h��R�(KK��h�C ]      �      �   "        �t�bhhK ��h��R�(KK��h�C   �        �        �t�bhhK ��h��R�(KK
��h�C(�   �   2      �     
   3        �t�bhhK ��h��R�(KK��h�CL      =         "   y        5      L
        v   `   `        �t�bhhK ��h��R�(KK��h�C	         �t�bhhK ��h��R�(KK��h�C      f  �        �t�bhhK ��h��R�(KK��h�C@   /   9   9  7         l        b  �   j      �      �t�bhhK ��h��R�(KK��h�C H   z  	
  (  �   �        �t�bhhK ��h��R�(KK ��h�C�      �        w         V  (   �  �
     �   �  �           U        8   �     �      L   G   �        �t�bhhK ��h��R�(KK
��h�C(1   #       m      �      �        �t�bhhK ��h��R�(KK��h�C@*         %     W   v   c   m              +         �t�bhhK ��h��R�(KK��h�C,�        �                        �t�bhhK ��h��R�(KK��h�C41   #      �  
   3   6   �
        &  r      �t�bhhK ��h��R�(KK��h�C0   f   W  �
          �               �t�bhhK ��h��R�(KK��h�CH%   �     9   {     9  _     �        
                  �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C@�  J  �            /   9     7      �               �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�CT   >   )        3     ,                  %      
   �   S   }         �t�bhhK ��h��R�(KK
��h�C(�   >   �  �  �     �   �         �t�bhhK ��h��R�(KK	��h�C$            �      �        �t�bhhK ��h��R�(KK��h�C,      )   �   L   G      �   

        �t�bhhK ��h��R�(KK��h�C0            "    �  �      �        �t�bhhK ��h��R�(KK��h�C4   �              %                     �t�bhhK ��h��R�(KK��h�C4      )  +   ^   &           �   X	        �t�bhhK ��h��R�(KK��h�C1         �t�bhhK ��h��R�(KK��h�CD      �   �
     �      �      �         �              �t�bhhK ��h��R�(KK��h�C@*      �       5         �     �   �   	  �        �t�bhhK ��h��R�(KK��h�C4!      �     /      �   '   
   �   F         �t�bhhK ��h��R�(KK��h�C4      �        @        �     X         �t�bhhK ��h��R�(KK��h�CE      �  	         �t�bhhK ��h��R�(KK��h�C4D      "   >  )   0                        �t�bhhK ��h��R�(KK��h�CE      0     m     �t�bhhK ��h��R�(KK
��h�C(Y      z     Q     z     x     �t�bhhK ��h��R�(KK	��h�C$<           	      	         �t�bhhK ��h��R�(KK
��h�C(-   !  |     ;      �          �t�bhhK ��h��R�(KK��h�C9     �t�bhhK ��h��R�(KK��h�C 1        	      	         �t�bhhK ��h��R�(KK��h�C,`  '                  8  3        �t�bhhK ��h��R�(KK��h�C8
      o  �  �        %   e  {   �  �        �t�bhhK ��h��R�(KK��h�C1   #       A   d        �t�bhhK ��h��R�(KK��h�C41   #           �   
   3   6      �        �t�bhhK ��h��R�(KK��h�C4|        ,      X  _  C         �         �t�bhhK ��h��R�(KK��h�C,*        $   n        �  �        �t�bhhK ��h��R�(KK��h�C01   #   
   3   6     �   �               �t�bhhK ��h��R�(KK��h�CQ  �     �t�bhhK ��h��R�(KK��h�C<      �     0     �   �     �  9   s   7         �t�bhhK ��h��R�(KK��h�CX*      /   �     �      �     �  �   7  H  '        M   �      D         �t�bhhK ��h��R�(KK��h�CD     �   �  2   �      �     D   ~   �      �           �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C<     p     �     <         �   	     A         �t�bhhK ��h��R�(KK��h�CD      �     j
  �  c      �      �         �   �         �t�bhhK ��h��R�(KK��h�C�             �t�bhhK ��h��R�(KK��h�C,   g  
           z     �        �t�bhhK ��h��R�(KK��h�CD
      R              2                 
   ,         �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C   ^     �t�bhhK ��h��R�(KK��h�C<4        C      �	           
     �            �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C ,   �     	      	   K      �t�bhhK ��h��R�(KK��h�C8�         )   �  �        E   ^   �  F         �t�bhhK ��h��R�(KK��h�CD      �  c      G  w  
   �  &      �   U   $           �t�bhhK ��h��R�(KK��h�C,G           �   �   �  i   �         �t�bhhK ��h��R�(KK��h�CP   �  -         	  �   �     %      �  )   �  S      -  {        �t�bhhK ��h��R�(KK��h�C<   �  �  �      '   
        R  9              �t�bhhK ��h��R�(KK	��h�C$         M     @            �t�bhhK ��h��R�(KK��h�C      �  �            �t�bhhK ��h��R�(KK
��h�C(�      '	  h     .   �   R          �t�bhhK ��h��R�(KK��h�C1        	         �t�bhhK ��h��R�(KK��h�CH         .   0   <      Q  m      �  �   <        �
        �t�bhhK ��h��R�(KK
��h�C(U   �   �   ,     !               �t�bhhK ��h��R�(KK��h�Ct      
   _      8   �  5      .      >  ,                0   U     ]   "   �     $   k         �t�bhhK ��h��R�(KK��h�C�
        �t�bhhK ��h��R�(KK5��h�C�      R  �     �      �                 |     �   E  
   _            d     �     �
        ]        
   _      �   �        T   }  
   _      ]         �     �   E        �t�bhhK ��h��R�(KK��h�C<                     (         W              �t�bhhK ��h��R�(KK��h�Cl   /      �           ,   	      	      	   K   	   �   	   I  	   U  	   �  	   �   	   �     �t�bhhK ��h��R�(KK��h�C8�         )   }        �  I  
   Q  �        �t�bhhK ��h��R�(KK��h�C	         �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C@      &   �  2     ,  9      �  L   y   �  l        �t�bhhK ��h��R�(KK��h�C<j   �         �   �     M   C   �   �              �t�bhhK ��h��R�(KK��h�C@   E  (      �   )                  k               �t�bhhK ��h��R�(KK��h�C0     �  r  
   ,                     �t�bhhK ��h��R�(KK��h�CDG   �   �        0   x      <      .   "   E      R         �t�bhhK ��h��R�(KK	��h�C$   Z        -   �   ,        �t�bhhK ��h��R�(KK��h�C   )  C      �     �t�bhhK ��h��R�(KK��h�C!            �t�bhhK ��h��R�(KK��h�CLt   �        '   �  Y  �  �  %   3     '   �     q   i
        �t�bhhK ��h��R�(KK��h�CP   v     �     �    �  G   �   �   �   #  �   9      �  y        �t�bhhK ��h��R�(KK
��h�C(2                J  E         �t�bhhK ��h��R�(KK��h�C`             �t�bhhK ��h��R�(KK��h�C8�     �     �  �   *      �  �             �t�bhhK ��h��R�(KK��h�C�     6     �        �t�bhhK ��h��R�(KK��h�Ck  
   B   }          �t�bhhK ��h��R�(KK��h�CP   �         �     D   0   e  �     l  �         C     �        �t�bhhK ��h��R�(KK��h�C,      '   U  �                    �t�bhhK ��h��R�(KK��h�C8
   X      �      �           �  �  �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�Ct      j        �t�bhhK ��h��R�(KK	��h�C$      �      ^   B   @        �t�bhhK ��h��R�(KK��h�CD�        R  �     �  0   4         
   �   �   _         �t�bhhK ��h��R�(KK��h�CT      D        �      �        �   &      I           $           �t�bhhK ��h��R�(KK��h�CX      
   _      8   �        �   �	        a   ;      �                 �t�bhhK ��h��R�(KK��h�CX   �      �     ~  �  �     �      ,         �      ^   �      (        �t�bhhK ��h��R�(KK��h�C@1   #      A     �  
   3   6         �  Y  �         �t�bhhK ��h��R�(KK��h�C0   *        �          �  �        �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�CT
   3   6         �  (      #   !      �        ;      �     �        �t�bhhK ��h��R�(KK	��h�C$�     �   '
        	         �t�bhhK ��h��R�(KK��h�CH   .      �           l  �      �  $   ;      �   �        �t�bhhK ��h��R�(KK��h�C<   �  �   �   
   _      l  ,   �      C           �t�bhhK ��h��R�(KK
��h�C(f	           Y    
   �         �t�bhhK ��h��R�(KK��h�C<
   �        2   �     U  �     �     +         �t�bhhK ��h��R�(KK��h�C`�   v     )         l        &   a   �  �        �     t                    �t�bhhK ��h��R�(KK��h�C    '   �  f
  ^  ^        �t�bhhK ��h��R�(KK��h�C8      -   �  +            u      $   x        �t�bhhK ��h��R�(KK��h�C               �t�bhhK ��h��R�(KK��h�CL   +                     +              �   �  
   �        �t�bhhK ��h��R�(KK��h�C�	  	      	         �t�bhhK ��h��R�(KK��h�C0
     �     i  8   h        �         �t�bhhK ��h��R�(KK��h�C0^   �        �   +
     .   �   �          �t�bhhK ��h��R�(KK	��h�C$   
      �    �  �   0     �t�bhhK ��h��R�(KK��h�C                       �t�bhhK ��h��R�(KK��h�C@      z   "        �  )               �   �         �t�bhhK ��h��R�(KK��h�C`      D   &   D  0   4   >   P  �   �  �        N   �        .   �     �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C4�     �      C  �     �                �t�bhhK ��h��R�(KK��h�C �     �      {   9   �
     �t�bhhK ��h��R�(KK��h�C1         �t�bhhK ��h��R�(KK��h�CL   =  �     t     R	  
   l                  +      T
        �t�bhhK ��h��R�(KK��h�Cl�      -           e  /         �                 �                                 �t�bhhK ��h��R�(KK��h�C �  �     k	  G   >        �t�bhhK ��h��R�(KK��h�C@         4           $     ;         �  �        �t�bhhK ��h��R�(KK
��h�C(        	      	      	   K      �t�bhhK ��h��R�(KK��h�C4      *     	      	      	   K   	   �      �t�bhhK ��h��R�(KK��h�C      $   x           �t�bhhK ��h��R�(KK��h�C    .   �      �  �        �t�bhhK ��h��R�(KK��h�CH      J   a      �  �  �           ]         �  �        �t�bhhK ��h��R�(KK��h�C�      �           �t�bhhK ��h��R�(KK��h�C<
   $        �   �             �  :   �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C4�      �  �  �  *   W     �      �        �t�bhhK ��h��R�(KK��h�C|*      �  
            ,                  6  +   &      R    }      p  
   $   �        $            �t�bhhK ��h��R�(KK��h�CD      �         �  [        .   W      |      �         �t�bhhK ��h��R�(KK��h�CT  �  �   �   7         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C2     �t�bhhK ��h��R�(KK��h�CH            �        c
     $   �   >   �                 �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK	��h�C$      F  +      f  �  =     �t�bhhK ��h��R�(KK	��h�C$-   �     �   .  "   �        �t�bhhK ��h��R�(KK	��h�C$�                 ,  r      �t�bhhK ��h��R�(KK��h�C 1   #       n             �t�bhhK ��h��R�(KK��h�C@I      w   �  �   %   J   �      -  J  C               �t�bhhK ��h��R�(KK��h�C9     �t�bhhK ��h��R�(KK��h�C #   !   '   
   3   6         �t�bhhK ��h��R�(KK��h�C �        �
     Z        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�CH�  �      $   Z  h        $   �      �
     P   �  �        �t�bhhK ��h��R�(KK��h�Cy     �t�bhhK ��h��R�(KK��h�C8         �   	     �  9      L   �	  Y        �t�bhhK ��h��R�(KK��h�C       �   -   H            �t�bhhK ��h��R�(KK��h�CT   �
     `   /      �              /   9     7                     �t�bhhK ��h��R�(KK
��h�C(A             �               �t�bhhK ��h��R�(KK��h�C<      �      p      �t�bhhK ��h��R�(KK	��h�C$   (   �   
   ,               �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK
��h�C(�  �	     8   ?     �           �t�bhhK ��h��R�(KK	��h�C$:  "   �   �        h
        �t�bhhK ��h��R�(KK��h�C4   &   �  �   �   $   E           <        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C@W   �  A           y     A  �  $  9   �   7         �t�bhhK ��h��R�(KK��h�C<�   &         �  '  y      a  +                  �t�bhhK ��h��R�(KK��h�C8   �  �   ,        D   ;      �  
   �        �t�bhhK ��h��R�(KK��h�C,      K  �  
   %  .	     �        �t�bhhK ��h��R�(KK��h�CH      �  q     $   �        �     q     
   �  �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CP   �      z     �  #     ?  �     �   S   X  i   ,               �t�bhhK ��h��R�(KK��h�C8*   D        $                             �t�bhhK ��h��R�(KK	��h�C$�   *  ?      
      F         �t�bhhK ��h��R�(KK��h�Cl   &     �        �        Y      Q              Y   
  �         5   &     �        �t�bhhK ��h��R�(KK��h�CJ     �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C�     =  	         �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C&  �  �      �     �t�bhhK ��h��R�(KK	��h�C$�   �   �            �        �t�bhhK ��h��R�(KK	��h�C$�     -                    �t�bhhK ��h��R�(KK��h�C@      �        J  E      A   F     {     [        �t�bhhK ��h��R�(KK��h�C8`           �                             �t�bhhK ��h��R�(KK��h�C 2      -   P   �   �        �t�bhhK ��h��R�(KK��h�Cj     �t�bhhK ��h��R�(KK��h�C,M   �      $   Z           W         �t�bhhK ��h��R�(KK��h�CD      �   �   $   E      u  
   %     F        �        �t�bhhK ��h��R�(KK��h�C@�  5                J                          �t�bhhK ��h��R�(KK��h�CPW  �     �   K     g  *      �     �      E     �     �        �t�bhhK ��h��R�(KK��h�CT      J   =      o  �   5         �  g  �   `   �     ,               �t�bhhK ��h��R�(KK��h�CH�     @   s   o  
         �  *   �     �  �      �        �t�bhhK ��h��R�(KK��h�CL      �
     Y       �            
     0   �  :            �t�bhhK ��h��R�(KK#��h�C�      U     �           ]
  c           �                   S  
   _      8   u  �                          �t�bhhK ��h��R�(KK��h�C  �   �         �t�bhhK ��h��R�(KK��h�C1   #       �      �t�bhhK ��h��R�(KK	��h�C$         `   b     �  y     �t�bhhK ��h��R�(KK��h�C       �
  	      	         �t�bhhK ��h��R�(KK��h�C4�     j              b         �        �t�bhhK ��h��R�(KK��h�C,�	       �              �        �t�bhhK ��h��R�(KK��h�CX-   �     0   <         �        �     �
        .   �         ^
        �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�C0%   5      .           �      �        �t�bhhK ��h��R�(KK��h�C,         I   �     0   Q  [
        �t�bhhK ��h��R�(KK��h�C�   �  �         �      �t�bhhK ��h��R�(KK��h�CD#   !      p        S      -  �   (      
   �  F         �t�bhhK ��h��R�(KK��h�C=     	      	         �t�bhhK ��h��R�(KK��h�CH   (   w   s        �   c   I   Z
     �     �      �         �t�bhhK ��h��R�(KK��h�C   M  �     �t�bhhK ��h��R�(KK	��h�C$      =
     A   �     �     �t�b�      hhK ��h��R�(KK	��h�C$�    
   ,      
            �t�bhhK ��h��R�(KK��h�C8
   |      <     '      �  �                 �t�bhhK ��h��R�(KK��h�CT      =               �     �   �         /   9   -     V        �t�bhhK ��h��R�(KK��h�C8      U     �   �      ^   �     \  x        �t�bhhK ��h��R�(KK
��h�C(V     I   �     �   �   R         �t�bhhK ��h��R�(KK"��h�C�"   t         0      �   ~              �     �     �           o  4      $   �     Y      O      "   H        �t�bhhK ��h��R�(KK	��h�C$K
     Y     ;     G        �t�bhhK ��h��R�(KK��h�Ck     �t�bhhK ��h��R�(KK	��h�C$1   #   
   3   6   (  O         �t�bhhK ��h��R�(KK��h�CD}  +   �        w  V         �     I  ,               �t�bhhK ��h��R�(KK��h�C8      a     �
     6  C         !  �        �t�bhhK ��h��R�(KK��h�C8      �     �     
       8   �            �t�bhhK ��h��R�(KK��h�C0
   �  F   '   #   !      S     !        �t�bhhK ��h��R�(KK
��h�C(q     �     �  	      	         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C8�   �  &   �   �   �  K  �     K              �t�bhhK ��h��R�(KK��h�C4�   �  �  "   �     �	     +     y        �t�bhhK ��h��R�(KK��h�Cd      G        #   i   �   �      5         �	     Y      O                        �t�bhhK ��h��R�(KK��h�C,I      ~         >   5  q   7        �t�bhhK ��h��R�(KK��h�C4   X   '   �  
      y        �           �t�bhhK ��h��R�(KK��h�C   �     7   v     �t�bhhK ��h��R�(KK��h�Cd      :  /   5            i  &      U        i           �   D     $   k         �t�bhhK ��h��R�(KK��h�C      �   $   �        �t�bhhK ��h��R�(KK��h�CH   �     $     "         �         9   �  "  P  �
        �t�bhhK ��h��R�(KK
��h�C(�      -   �  �     �   �         �t�bhhK ��h��R�(KK��h�C<q      	      	      	   K   	   �   	   I  	   /     �t�bhhK ��h��R�(KK��h�CT   '   �  H   }     �   *     �       �      I   }  (      n         �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK	��h�C$�        >   \  t   �        �t�bhhK ��h��R�(KK
��h�C(!               	      	         �t�bhhK ��h��R�(KK��h�C@   �     �t�bhhK ��h��R�(KK��h�C8�    �        /      �           �        �t�bhhK ��h��R�(KK��h�C@   @   '   �	     6        F     �     �  �         �t�bhhK ��h��R�(KK��h�C\     	      	         �t�bhhK ��h��R�(KK��h�C`   &   N   m  �  I     �       �  N      �      �   �  �     {      �        �t�bhhK ��h��R�(KK��h�CL   =                   �  
   b	     I         )            �t�bhhK ��h��R�(KK��h�CX   .      8  0   �        %              �      _  �   d   "           �t�bhhK ��h��R�(KK��h�C<   �   b     �   �        p  N   R     �         �t�be(hhK ��h��R�(KK��h�C 1   #   
   3   6            �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C    5   7  4               �t�bhhK ��h��R�(KK��h�C@�  "   &  �   +               �   {         �        �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�CZ          �            �t�bhhK ��h��R�(KK��h�C   q             �t�bhhK ��h��R�(KK��h�C�
           �t�bhhK ��h��R�(KK��h�C4   �           �         �              �t�bhhK ��h��R�(KK��h�C8     �       �              �           �t�bhhK ��h��R�(KK��h�C_     �  R          �t�bhhK ��h��R�(KK	��h�C$     �      �     �        �t�bhhK ��h��R�(KK��h�C<!         �         '   
   3   6                  �t�bhhK ��h��R�(KK��h�CL9   �     �   (      �          �   +      `   �    �         �t�bhhK ��h��R�(KK��h�CH      �         :   M        �      5         �   ~        �t�bhhK ��h��R�(KK��h�CH              F  �      U     
   $      
      6         �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C{      �      �t�bhhK ��h��R�(KK��h�CH1   #      r  
   3   �  7  �        L     �     r        �t�bhhK ��h��R�(KK
��h�C(b   #   G   �   �     R  �         �t�bhhK ��h��R�(KK��h�CX     :  {        �t�bhhK ��h��R�(KK��h�C,V             �  �      w        �t�bhhK ��h��R�(KK��h�Cx
   H   �     2   �  �     2      �      �      .   0  �  �     �     6  S  0  �  �     N        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK
��h�C(1   #       m      �      �        �t�bhhK ��h��R�(KK��h�C<         "     �  �      s  �  9   �           �t�bhhK ��h��R�(KK��h�C,�  {    ?              e        �t�bhhK ��h��R�(KK
��h�C(&  �   p        Z  �  �         �t�bhhK ��h��R�(KK��h�CD      =  
   �   �   �     �  �                        �t�bhhK ��h��R�(KK	��h�C$�  !      9  	      	         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C0               i      H   A   ?        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CD�  l     w  �   "   #  �  }     O  "   P  �  }        �t�bhhK ��h��R�(KK��h�C<   �   -   V     v      
      g      ]  L         �t�bhhK ��h��R�(KK��h�C,9     )   K     �     Q  �        �t�bhhK ��h��R�(KK��h�C�  "     �t�bhhK ��h��R�(KK��h�C      �         �t�bhhK ��h��R�(KK��h�C4   �  {  *   �     
  ~   
   �           �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�C�  	      	         �t�bhhK ��h��R�(KK
��h�C(            �  
   B           �t�bhhK ��h��R�(KK��h�C,�   
      �        �     @         �t�bhhK ��h��R�(KK��h�C/      �t�bhhK ��h��R�(KK��h�C01   #      �        
   3   6   N	        �t�bhhK ��h��R�(KK��h�C0�                 =         �
        �t�bhhK ��h��R�(KK ��h�C�           m              x   G     ^  @     �   
             @     Z               Z            �t�bhhK ��h��R�(KK��h�CP"         2      .   �  �     �   |     F	  �     }              �t�bhhK ��h��R�(KK
��h�C(�        �  �         S   Q      �t�bhhK ��h��R�(KK��h�C	  l      �t�bhhK ��h��R�(KK��h�C*   C     �     �t�bhhK ��h��R�(KK��h�C3      �t�bhhK ��h��R�(KK��h�CP   .   �  �  
  >                    �  �  >                 �t�bhhK ��h��R�(KK��h�C{     �   ,   	         �t�bhhK ��h��R�(KK��h�C@     �     �t�bhhK ��h��R�(KK��h�C<�                 C   
      S     i   �	        �t�bhhK ��h��R�(KK��h�CH
   @   �   F   ?         �  �   %   5     e     �   ,        �t�bhhK ��h��R�(KK��h�C<1     +      &   }                ,   	         �t�bhhK ��h��R�(KK��h�C4�	          �        �     ,   	         �t�bhhK ��h��R�(KK��h�C<            G             U      .   �        �t�bhhK ��h��R�(KK��h�C,       a  �      �     �        �t�bhhK ��h��R�(KK��h�C  �     �t�bhhK ��h��R�(KK��h�C`2            
  {                  %  }     �  �   �   \  2               �t�bhhK ��h��R�(KK��h�CP?
     �     a     .            3
        �         
   &        �t�bhhK ��h��R�(KK��h�CL      B  G         
      F         5      �      8   o         �t�bhhK ��h��R�(KK��h�CL         
            &        $   �      �     c
        �t�bhhK ��h��R�(KK��h�CH        �     /   9   -  (   2   <         i     Z        �t�bhhK ��h��R�(KK
��h�C(�     �      �	     d   �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�Cd         $           �  b     6
        P  �  M
        P   �   @  G   W         �t�bhhK ��h��R�(KK��h�C         J     	         �t�bhhK ��h��R�(KK��h�C       /      �             �t�bhhK ��h��R�(KK	��h�C$#   !   ?      
      F         �t�bhhK ��h��R�(KK��h�C0�           �
  �     .     :        �t�bhhK ��h��R�(KK��h�C@      4  �         *         �          i	        �t�bhhK ��h��R�(KK��h�C       �     ^           �t�bhhK ��h��R�(KK
��h�C(   d
  p   Y     z  �   7         �t�bhhK ��h��R�(KK
��h�C(   W        @      X   �        �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   6                  �t�bhhK ��h��R�(KK��h�CHe   �   �      	     %   �     �     9      /      V        �t�bhhK ��h��R�(KK��h�Ch     �t�bhhK ��h��R�(KK��h�CY         �            �t�bhhK ��h��R�(KK��h�CL
   �  '            o  �  :         �  �           
        �t�bhhK ��h��R�(KK��h�C�	     �     �t�bhhK ��h��R�(KK	��h�C$Z      �            z        �t�bhhK ��h��R�(KK��h�C      �  �         �t�bhhK ��h��R�(KK#��h�C�   �  "   �      (     ~  �  �     �     r  �                 L           �      +   *      �  +      �        �t�bhhK ��h��R�(KK��h�C0�   L   �   �   
   �     �               �t�bhhK ��h��R�(KK��h�C !      5  	      	         �t�bhhK ��h��R�(KK��h�Cd     �t�bhhK ��h��R�(KK	��h�C$1   #   
   3   6      �        �t�bhhK ��h��R�(KK��h�CD      P   �        �  �     p   �   �   ^   �   *        �t�bhhK ��h��R�(KK��h�C@     &  �  %   [     	  �  �         ]           �t�bhhK ��h��R�(KK��h�C,�  (     �   �   "  )              �t�bhhK ��h��R�(KK��h�C47  �     2     p      k     H	  �         �t�bhhK ��h��R�(KK��h�Cd�  5  C   �           S  �        �                  �  ~                    �t�bhhK ��h��R�(KK
��h�C(H   z  #  �        
            �t�bhhK ��h��R�(KK��h�C  �                 �t�bhhK ��h��R�(KK��h�C<   f   �   �  �       �      �     �           �t�bhhK ��h��R�(KK��h�C`f   ?  �     �   �      �   �      |     �        �  �   �        �  �        �t�bhhK ��h��R�(KK��h�Cd
   �  �   �      &  �  u      �               �      �      -  +     �  �        �t�bhhK ��h��R�(KK��h�CZ          �            �t�bhhK ��h��R�(KK��h�C<�   �   +   s  
   B   
  :      �        S         �t�bhhK ��h��R�(KK��h�CD�       
   4     l
  �  �     ?          �        �t�bhhK ��h��R�(KK	��h�C$      �   �  R      �        �t�bhhK ��h��R�(KK��h�C8   `   q     %           x  +      �         �t�bhhK ��h��R�(KK��h�CT              �   �   �   6	  
        �         
        {         �t�bhhK ��h��R�(KK��h�C1   #               �t�bhhK ��h��R�(KK��h�C0               	      	      	   K      �t�bhhK ��h��R�(KK��h�CD"        �	     �   -   A   �  O      ~         U        �t�bhhK ��h��R�(KK��h�CD   �  V        �
  �
  �  +  _  �  
      �  �        �t�bhhK ��h��R�(KK
��h�C(�   '      �
     �   B           �t�bhhK ��h��R�(KK��h�C08   ,
           $   A     �           �t�bhhK ��h��R�(KK��h�CH   &   \  �       h   �   �   g      a   �  E   
           �t�bhhK ��h��R�(KK
��h�C(      �  )                     �t�bhhK ��h��R�(KK��h�Cb   #   
   $   �        �t�bhhK ��h��R�(KK��h�C�  �   ,        �t�bhhK ��h��R�(KK��h�C8O       f              �                 �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C!      @  	  	         �t�bhhK ��h��R�(KK��h�CP      �      �        �   )      /      �        �  �  7         �t�bhhK ��h��R�(KK��h�CH         +  :         G  �   s   7   j   �  �  8   4         �t�bhhK ��h��R�(KK��h�CX
  $   |  �      �      \   �         v      "              0            �t�bhhK ��h��R�(KK��h�C [         	      	         �t�bhhK ��h��R�(KK��h�C�   �     �t�bhhK ��h��R�(KK��h�CS  �          �t�bhhK ��h��R�(KK��h�C	     �      �      �t�bhhK ��h��R�(KK��h�Ch*               >      �      �     6     F  +   "   t      �     
   $   �   �        �t�bhhK ��h��R�(KK	��h�C$�  (      N      �           �t�bhhK ��h��R�(KK��h�CH�      �  �           �      Q          u               �t�bhhK ��h��R�(KK��h�CD         D  2     �  �        {         �
           �t�bhhK ��h��R�(KK��h�C`      =      �                (   :            E   v  �     �     Z        �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C<1   #      ,   �       �  
   3   6   	  �         �t�bhhK ��h��R�(KK��h�Ct�	     �   7  4              ,  "   t      �                       ,     �     �           �t�bhhK ��h��R�(KK��h�CT]      �  �        �        J           
      *        �        �t�bhhK ��h��R�(KK��h�C   @        �t�bhhK ��h��R�(KK��h�C�     �  r      �t�bhhK ��h��R�(KK��h�CL*      �     �     �         �   �   
   +      �  $   0        �t�bhhK ��h��R�(KK��h�C�          �      �t�bhhK ��h��R�(KK��h�CH   .   �   "      �        �	           .        �        �t�bhhK ��h��R�(KK��h�Ch      6  +      �
                       6  
                                    �t�bhhK ��h��R�(KK��h�C2  	  	      	         �t�bhhK ��h��R�(KK��h�C01   #       n          2              �t�bhhK ��h��R�(KK
��h�C(9  �       2   �      �         �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C,              �     ,   K        �t�bhhK ��h��R�(KK��h�C[      �  	         �t�bhhK ��h��R�(KK��h�C9     �t�bhhK ��h��R�(KK
��h�C(p  9   �  7            �         �t�bhhK ��h��R�(KK��h�C   �   �      =           �t�bhhK ��h��R�(KK��h�C8�   x  �     e     R         .   '  R         �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�CX   D   �   5   �       q
  �  
   �   �     w     �      '              �t�bhhK ��h��R�(KK	��h�C$�  �           �           �t�bhhK ��h��R�(KK��h�C@         ,   _
        )   i  �  �  
      F         �t�bhhK ��h��R�(KK��h�C   
  
  �           �t�bhhK ��h��R�(KK��h�CH)         h     '   �     �        �           �        �t�bhhK ��h��R�(KK ��h�C�`            S              S                �  �                                      �   �     �t�bhhK ��h��R�(KK��h�CX         �   �     �           x           6     �	                 �t�bhhK ��h��R�(KK��h�C0   �   �     !  o      �    o         �t�bhhK ��h��R�(KK	��h�C$"   >  b  D      �   N        �t�bhhK ��h��R�(KK��h�C8g        y  �  2      T  �  �   #  o        �t�bhhK ��h��R�(KK��h�C   '   
   H   [        �t�bhhK ��h��R�(KK#��h�C�   D   (   �         Y      Q      &      =      n     Y      �  �     D      �  �     �  �        "   �  �        �t�bhhK ��h��R�(KK��h�C�     �  	         �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C<   �  �            �  �     $   �              �t�bhhK ��h��R�(KK��h�CH   �        �             �  ;     �  *   �  {        �t�bhhK ��h��R�(KK��h�C4      =      �	  G   B   �
                 �t�bhhK ��h��R�(KK	��h�C$         �     s           �t�bhhK ��h��R�(KK��h�C    >   �   w   �          �t�bhhK ��h��R�(KK��h�CL   �                           P   !      �  �     T        �t�bhhK ��h��R�(KK��h�CT   �        9                 $  �   �  j   %   L	                 �t�bhhK ��h��R�(KK��h�C4|      �      <  �  +   "   >     j        �t�bhhK ��h��R�(KK��h�C0  �     .   �
  
   �
     A            �t�bhhK ��h��R�(KK
��h�C(�        	      	      	   ^     �t�bhhK ��h��R�(KK��h�C�     �  �     �t�bhhK ��h��R�(KK��h�CH   ?   #   !         �        �  
   3   6   �              �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C8   	     %   �  #  �     `   b     �        �t�bhhK ��h��R�(KK��h�CDh   s   �  g      d   t    �  t        S     �        �t�bhhK ��h��R�(KK��h�C0   �     �        �                 �t�bhhK ��h��R�(KK	��h�C$�     �  u                 �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6            �t�bhhK ��h��R�(KK��h�C�  '     t         �t�bhhK ��h��R�(KK	��h�C$            �   l           �t�bhhK ��h��R�(KK��h�C         �	  �     �t�bhhK ��h��R�(KK��h�C0H   e  �  �      �      <               �t�bhhK ��h��R�(KK��h�C4           �      |      �   C     +      �t�bhhK ��h��R�(KK��h�C,      �   ~     �      x     +      �t�bhhK ��h��R�(KK��h�C,
   H   [  '   �        �  n
        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C   �   �            �t�bhhK ��h��R�(KK��h�CE      4      �        �t�bhhK ��h��R�(KK��h�CL      )   \  �  x
  y
              @         b      �        �t�bhhK ��h��R�(KK��h�C4#  &   �   R  *   �   �  }     +  n   r      �t�bhhK ��h��R�(KK
��h�C(�                     z
  �      �t�bhhK ��h��R�(KK��h�CT#   !      F     �  ?      
   X   �   �        
   &                 �t�bhhK ��h��R�(KK��h�C,1   #   
   3   6     �              �t�bhhK ��h��R�(KK��h�C    ?   �  "   $   /        �t�bhhK ��h��R�(KK��h�C0�   5      �  +      �  
   �            �t�bhhK ��h��R�(KK��h�C      �     �t�bhhK ��h��R�(KK��h�Cl�
     �     �
     X             �     �
     �        �     v        *          �t�bhhK ��h��R�(KK��h�CX   s  �              P     �     j
  :   �  �        *   A  {        �t�bhhK ��h��R�(KK��h�C   ,   	         �t�bhhK ��h��R�(KK��h�C*      �  /      �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK	��h�C$   '   u     %   .  �        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C[                 �t�bhhK ��h��R�(KK��h�C0      �  �           �               �t�bhhK ��h��R�(KK��h�C -       4  
   t         �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6            �t�bhhK ��h��R�(KK��h�C      $        �t�bhhK ��h��R�(KK��h�C8        	  C      2   �        2   �        �t�bhhK ��h��R�(KK
��h�C(   q   p  �   B         ^        �t�bhhK ��h��R�(KK��h�C,+  �   -   l        �     s        �t�bhhK ��h��R�(KK��h�CXT      /   C   c              �              f  c         %            �t�bhhK ��h��R�(KK��h�CZ     �t�bhhK ��h��R�(KK��h�C�  	      	         �t�bhhK ��h��R�(KK
��h�C(   M        q  �             �t�bhhK ��h��R�(KK
��h�C(�     �     v        7        �t�bhhK ��h��R�(KK��h�C`      6        �   D  )               ;      �      �        �              �t�bhhK ��h��R�(KK��h�C    �   '      �
  &        �t�bhhK ��h��R�(KK��h�C0         ;  �  �   *   %   �
  C         �t�bhhK ��h��R�(KK
��h�C(�            S         !        �t�bhhK ��h��R�(KK��h�C�     	      	         �t�bhhK ��h��R�(KK��h�CH"   _        0   !      �        .   >  "   m
              �t�bhhK ��h��R�(KK
��h�C(  �     �  (   �         r      �t�bhhK ��h��R�(KK��h�CH�     �  �      �     �        �    >      �   L         �t�bhhK ��h��R�(KK	��h�C$%            �               �t�bhhK ��h��R�(KK��h�Cd�         h  !      �     b  :   M     �     {   �   �   \      �  �   /  �        �t�bhhK ��h��R�(KK��h�C@�      c     �   m      �  
        �      �        �t�bhhK ��h��R�(KK��h�C0      0   �   >      a                  �t�bhhK ��h��R�(KK��h�CH      J   P         �   =  &      }        �     =        �t�bhhK ��h��R�(KK��h�C4g   :  
   A   F        6  �     �        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�CD      �      �    
         M      �      A   W
        �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C1   #       �  �         �t�bhhK ��h��R�(KK��h�CL   f   ?     D   ;      �  
   �  )   T      �  �     '        �t�bhhK ��h��R�(KK��h�CP   @   '   )   �   5  O              K      /     �      I        �t�bhhK ��h��R�(KK��h�C0�     �  �   �      ^   �     s         �t�bhhK ��h��R�(KK��h�C<              �   �   �         =               �t�bhhK ��h��R�(KK
��h�C(  	      	      	   K   	   U     �t�bhhK ��h��R�(KK��h�Cl  E      �  	         �t�bhhK ��h��R�(KK��h�CH*      �      +      G                 >                  �t�bhhK ��h��R�(KK��h�C@/    
   ,         �      �     �  )   
            �t�bhhK ��h��R�(KK��h�C                �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6            �t�bhhK ��h��R�(KK
��h�C(�       ?      
   X   F         �t�bhhK ��h��R�(KK��h�C0      b         
   $   �  "   k        �t�bhhK ��h��R�(KK	��h�C$H   7  C                     �t�bhhK ��h��R�(KK
��h�C(   O        )   �   j   4         �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK��h�CX   8   �     �  �  p     _     $   �     2           �  3  �        �t�bhhK ��h��R�(KK��h�CD         �   �        �     U   e   �   �              �t�bhhK ��h��R�(KK��h�C%   �  k     6        �t�bhhK ��h��R�(KK��h�C   �     z
  �      �t�bhhK ��h��R�(KK��h�C4T            .  �   �  i      �  p        �t�bhhK ��h��R�(KK��h�C 1   #       m      4         �t�bhhK ��h��R�(KK
��h�C(�  �   Q  �      �              �t�bhhK ��h��R�(KK��h�Cl"   @   {  '         ;     u   �   N  7      V         �   �        �         �   �         �t�bhhK ��h��R�(KK��h�C 2      -   P   �   �        �t�bhhK ��h��R�(KK��h�C8   >   �  I   ^  
   A  �   g   �  �            �t�bhhK ��h��R�(KK��h�C      L                �t�bhhK ��h��R�(KK
��h�C(      -   =      ~  :   t         �t�bhhK ��h��R�(KK��h�CD�  q     N      .                     �     �        �t�bhhK ��h��R�(KK��h�C,   w  7  C   D       �  O        �t�bhhK ��h��R�(KK��h�C0   :           `   �      �   s   7      �t�bhhK ��h��R�(KK��h�C\   5   a   �      �  /  �     �        D  v      �      �     A   �        �t�bhhK ��h��R�(KK��h�CX         <        }     �   o      6  �   
   3   6   7  }     o         �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�C0#   !      k  ?      
   3   6            �t�bhhK ��h��R�(KK��h�CPY      O               ,        -   �  �      (	     q   �	        �t�bhhK ��h��R�(KK��h�C\
   �  �  '   )                  V      %   C
  �                 B	        �t�bhhK ��h��R�(KK��h�CH   >   �   *      '   �   �   /            ]  d     <        �t�bhhK ��h��R�(KK��h�C@  &   N   b     �       /         J     &        �t�bhhK ��h��R�(KK��h�C0W  �           �	  `   �     L         �t�bhhK ��h��R�(KK
��h�C(         9   �                  �t�bhhK ��h��R�(KK
��h�C(O  �    �      i     �        �t�bhhK ��h��R�(KK��h�C<   t   �  $   �     T  `   U  �  )              �t�bhhK ��h��R�(KK��h�CD   �  �         �   �     O        Q   V      E  �      �t�bhhK ��h��R�(KK��h�C   �    7         �t�bhhK ��h��R�(KK��h�C@�  )
        )
     �   p     �           [        �t�bhhK ��h��R�(KK��h�C    �                   �t�bhhK ��h��R�(KK��h�Cm                 �t�bhhK ��h��R�(KK��h�CD      5   B              -   M   �      @     �        �t�bhhK ��h��R�(KK��h�CL   �      $     �     
  :   �   3  �         �	     �         �t�bhhK ��h��R�(KK��h�C   �   '   E           �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�C0               �     	      	         �t�bhhK ��h��R�(KK��h�Cl        C                  0  %   c        }
        %   N
        }
                 �t�bhhK ��h��R�(KK��h�CX#   !      R      	  (      :     ^  @     �   
     �   �                �t�bhhK ��h��R�(KK��h�C�   �     �t�bhhK ��h��R�(KK��h�CT
   3   6   Y      O   ?      !      �           A     i      �        �t�bhhK ��h��R�(KK��h�C  �           �t�bhhK ��h��R�(KK��h�C          f   �  �        �t�bhhK ��h��R�(KK��h�C@/   9   N  7   �     7     �     z  s   �  �        �t�bhhK ��h��R�(KK��h�C|S        X  �              g      u  �  �  B        9         �           L   T   q               �t�bhhK ��h��R�(KK��h�C       )   �     �        �t�bhhK ��h��R�(KK��h�Cl              �         T      E  {      
   �  &      �   M   �   ]   
   $   �        �t�bhhK ��h��R�(KK��h�C     r  �         �t�bhhK ��h��R�(KK��h�C4n     �     Y      O   (     �            �t�bhhK ��h��R�(KK��h�CH!      B        	      	      	   K   	     	   �   	   �     �t�bhhK ��h��R�(KK��h�C,         �t�bhhK ��h��R�(KK��h�C9  	         �t�bhhK ��h��R�(KK��h�C82   �  �   (     m   �  y   %   �     �        �t�bhhK ��h��R�(KK	��h�C$�     E      2     �        �t�bhhK ��h��R�(KK	��h�C$0     �  p  "        .     �t�bhhK ��h��R�(KK��h�C:     -        �t�bhhK ��h��R�(KK��h�C,   �   ,  )      ~                 �t�bhhK ��h��R�(KK	��h�C$�
        ]  �     �        �t�bhhK ��h��R�(KK��h�C\     �     �t�bhhK ��h��R�(KK��h�C   �  g	     �t�bhhK ��h��R�(KK��h�C@      z     N         M   .        �  
   A         �t�bhhK ��h��R�(KK��h�C
  =  �  M     �t�bhhK ��h��R�(KK��h�C�           �     �t�bhhK ��h��R�(KK
��h�C(   �      �  �  �      ]         �t�bhhK ��h��R�(KK��h�C8�   &   �     !        %   b        �        �t�bhhK ��h��R�(KK��h�C8
         2      
         �     
            �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C      �   �   F     �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C@   s  �  {  �  j   e  
      �     �     A        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK	��h�C$
   3   6              r      �t�bhhK ��h��R�(KK	��h�C$      ~   H        =        �t�bhhK ��h��R�(KK��h�CP   @	  
      �        .   N      o          �  �               �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�CL            �  G   �      (  L     r  '     �  
   �        �t�bhhK ��h��R�(KK��h�CH      0        :      �  T      �  P  "   |      �         �t�bhhK ��h��R�(KK��h�C8#   !      �  ?      
   3   6   �             �t�bhhK ��h��R�(KK��h�C �       A  ,  a        �t�bhhK ��h��R�(KK��h�C       l         ]  \     �t�bhhK ��h��R�(KK��h�C%     �t�bhhK ��h��R�(KK��h�C8      �  �      V
        �     �  &         �t�bhhK ��h��R�(KK��h�CPA     .        �     	     N         �        �              �t�bhhK ��h��R�(KK��h�C 1        	      	         �t�bhhK ��h��R�(KK��h�CH   �  �      +         J  +      |      �      f  �        �t�bhhK ��h��R�(KK
��h�C(�	     �  �   �        �   O      �t�bhhK ��h��R�(KK��h�C%   '   d     T        �t�bhhK ��h��R�(KK��h�C8!      b     �      �  h      	      	         �t�bhhK ��h��R�(KK��h�C@         V     .   �     �     J                 �t�bhhK ��h��R�(KK��h�C,9   �        =      �     >        �t�bhhK ��h��R�(KK��h�C0      ;  +      G     $   �   �        �t�bhhK ��h��R�(KK��h�C@     �  B        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�CX�  q     )   N      .                       �                        �t�bhhK ��h��R�(KK��h�C   f     g            �t�bhhK ��h��R�(KK	��h�C$�  �         �               �t�bhhK ��h��R�(KK��h�C@            �     `  ,     )      %      /         �t�bhhK ��h��R�(KK��h�C0     ^       9     ]	     �        �t�bhhK ��h��R�(KK��h�CP      -   P   !      �   
  
      .   q   R     �        F         �t�bhhK ��h��R�(KK��h�CT@      z             �     k     ,      �  �           X        �t�bhhK ��h��R�(KK��h�Cl               �            �   f     z  +   
   �      (  �  
   $     �     f        �t�bhhK ��h��R�(KK.��h�C��  �   �       �         %   �      v        �   7                          �       7        C  D     ,           �      �           �        �t�bhhK ��h��R�(KK��h�C8         2   �   `  �  "   `     "           �t�bhhK ��h��R�(KK	��h�C$f   �	     )   �  A   �        �t�bhhK ��h��R�(KK��h�C(     �t�bhhK ��h��R�(KK��h�CW   v  	      	         �t�bhhK ��h��R�(KK	��h�C$   &   -   �     :            �t�bhhK ��h��R�(KK��h�CX   �     �  0  +      $   �            9      ]  L   &   �   
   �        �t�bhhK ��h��R�(KK��h�CHb   #   "   7
     u            $   k         "   $  �        �t�bhhK ��h��R�(KK��h�C\�   *           �      �        �     8   %     �  $   �        �         �t�bhhK ��h��R�(KK��h�C,�  q  �      .      ?     �        �t�bhhK ��h��R�(KK
��h�C(f   ?     -   �     A           �t�bhhK ��h��R�(KK��h�C0  �   d   :  6  �   *   �     �         �t�bhhK ��h��R�(KK#��h�C�   ;     �     �  �  �  "   �      *      �  �  �	     ;              ;     �     �  �  �     ;              �t�bhhK ��h��R�(KK
��h�C(            o      B   3        �t�bhhK ��h��R�(KK��h�C T   �   P  e   �           �t�bhhK ��h��R�(KK��h�CP         F  9      
  L   (      �   �   9   m     �  L   �        �t�bhhK ��h��R�(KK	��h�C$      )         �            �t�bhhK ��h��R�(KK��h�C 4      r  	      	         �t�bhhK ��h��R�(KK��h�C0        J   �        :     �        �t�bhhK ��h��R�(KK��h�C 1   #   
   X   �   F         �t�bhhK ��h��R�(KK
��h�C(   �  q     �  
   �   �	        �t�bhhK ��h��R�(KK��h�C,*      5   �   5      �               �t�bhhK ��h��R�(KK��h�C8!         =        ?      
   3   6   �        �t�bhhK ��h��R�(KK��h�C8�   R      �                k               �t�bhhK ��h��R�(KK)��h�C�      -   =      8     L              $   t     �   O         w      O            Q         J   �        5   L        �               �t�bhhK ��h��R�(KK��h�C0�        4  :            S   Q   r      �t�bhhK ��h��R�(KK��h�CT            �        �  �     &      w   �  q          �        �t�bhhK ��h��R�(KK��h�C<1   #   
   3   6        u       g   d   t        �t�bhhK ��h��R�(KK��h�C1   #          �t�bhhK ��h��R�(KK��h�C�	     �     	         �t�bhhK ��h��R�(KK��h�C`�  �     +                  �        �
     ,   	      	      	   K   	   �      �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�CS  (         �t�bhhK ��h��R�(KK��h�Cm     	         �t�bhhK ��h��R�(KK��h�C4�   q   7     I   /   �
    �     }        �t�bhhK ��h��R�(KK��h�CX      �         �     �   �   S        �  U   q   �  �    �  O        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C4n     )   c         *     %   �  c         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C8�        �      �     *   �      g   n         �t�bhhK ��h��R�(KK��h�C�	    {   !           �t�bhhK ��h��R�(KK��h�CT-   �               J  
   C      S  q  n
     �	                �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8   $  )   m     �     �      �   ,   �         �t�bhhK ��h��R�(KK��h�C �  {  �          �     �t�bhhK ��h��R�(KK��h�C-   �  �   �        �t�bhhK ��h��R�(KK��h�C�     m     �t�bhhK ��h��R�(KK��h�CH*      �  t  (      /   T     �  �     d   �     �        �t�bhhK ��h��R�(KK��h�C4!      �         ?      
   3   6   �        �t�bhhK ��h��R�(KK��h�C@      0   4   
   _      �     8   /   ~               �t�bhhK ��h��R�(KK��h�C4�   &   �     �              �   �         �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�C    L  �     +   w        �t�bhhK ��h��R�(KK��h�C �      K	  �   
           �t�bhhK ��h��R�(KK��h�Cm      �      �     �t�bhhK ��h��R�(KK��h�C\   �     �     p  "   �   ,   9     �      9     �      ^  "   �   {        �t�bhhK ��h��R�(KK��h�CT�   �     ;         ~	             �  *   %     �      
   �        �t�bhhK ��h��R�(KK��h�C 
   )     H   �           �t�bhhK ��h��R�(KK��h�C,   d  w   \   �   ,	     J   M         �t�bhhK ��h��R�(KK��h�C,�     -   �  
   s      �  7         �t�bhhK ��h��R�(KK��h�C�  
   ,         �t�bhhK ��h��R�(KK��h�C,      �      9   I   Z  
   �        �t�bhhK ��h��R�(KK��h�C8�  �      �                �  �   �        �t�bhhK ��h��R�(KK��h�C@�   =     �      i   *     2   �     o      n        �t�bhhK ��h��R�(KK��h�C   �            �t�bhhK ��h��R�(KK��h�C<e   @     �  "   ~  y  �  l      ~              �t�bhhK ��h��R�(KK%��h�C�!         �      �     o         N     	      	      	   �   	   �   	   I  	   /  	   s  	   )  	   �  	   �  	   �  	   �     �t�bhhK ��h��R�(KK��h�CX         <        }     �   o      6  �   
   3   6   7  }     o         �t�bhhK ��h��R�(KK��h�C0      5      �         U   $            �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�CP              �   �               =      �     �  G   W         �t�bhhK ��h��R�(KK	��h�C$   �     H   �              �t�bhhK ��h��R�(KK��h�CD               J   �   8  5         �      `   8        �t�bhhK ��h��R�(KK��h�C,           �      	      	         �t�bhhK ��h��R�(KK:��h�C��     B     8   E           S   Q   V      G  ~           -   =      8     4            $   �     �     �   O         w      O            Q         J   �        5   L        �               �t�bhhK ��h��R�(KK��h�C<�      -   r     �	     v  �     �      �         �t�bhhK ��h��R�(KK��h�C{     �     �t�bhhK ��h��R�(KK��h�C`      �     �  
         �     �        �     ,      K                     �t�bhhK ��h��R�(KK	��h�C$5         r   �     �  m      �t�bhhK ��h��R�(KK��h�Cr     	         �t�bhhK ��h��R�(KK��h�C%   �      h           �t�bhhK ��h��R�(KK��h�C   �      �t�bhhK ��h��R�(KK��h�C,O     P  (   N   A    (  I        �t�bhhK ��h��R�(KK��h�C�  �              �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�Cl      5   x      �     -  ~     /      �              �      L   G   C     �           �t�bhhK ��h��R�(KK��h�C   }     o      �t�bhhK ��h��R�(KK��h�C4   (   !      �        
   3   6   n        �t�bhhK ��h��R�(KK��h�CX   $           �            �           ;      %   �     �   �        �t�bhhK ��h��R�(KK��h�C<        �      N     q        �  �  �        �t�bhhK ��h��R�(KK��h�C0      �   "     z   "      �           �t�bhhK ��h��R�(KK��h�Cb   �     W         �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK	��h�C$�  	     �      -           �t�bhhK ��h��R�(KK��h�C,M      +      3     �     �        �t�bhhK ��h��R�(KK��h�CT   P           5   v      %           5         �  +      "        �t�bhhK ��h��R�(KK��h�C0      �  A      &      a      }        �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C  &     �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�CD*         1
           j  �      �   +   "               �t�bhhK ��h��R�(KK��h�C<�  �     �     �  �      �     {     J        �t�bhhK ��h��R�(KK��h�C                        �t�bhhK ��h��R�(KK��h�C<           (      �        `   �     A         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C0�  4      �   �    [   �      0         �t�bhhK ��h��R�(KK	��h�C$:     Q                     �t�bhhK ��h��R�(KK��h�C<      i              
         3
     �
        �t�bhhK ��h��R�(KK��h�CD      �      6  
   �       �   �        O  �        �t�bhhK ��h��R�(KK
��h�C(            v     .             �t�bhhK ��h��R�(KK��h�C8      V
  X                �        "     �t�bhhK ��h��R�(KK��h�C�     T  
   &        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C,�  7     �     ;      P   �         �t�bhhK ��h��R�(KK��h�Cd   �      >     �     l      &   �  �   o         �      �      �     �   o         �t�bhhK ��h��R�(KK��h�C �  "   �  	      	         �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�CHR      	        .   y        �     �           �         �t�bhhK ��h��R�(KK��h�C<   5  �            *      j        ^            �t�bhhK ��h��R�(KK	��h�C$        Z     8   �        �t�bhhK ��h��R�(KK��h�C@
   �   �             �	  [   �     0               �t�bhhK ��h��R�(KK��h�C0%   �         �     �      d   �         �t�bhhK ��h��R�(KK��h�C0�  �      �      �      )      �         �t�bhhK ��h��R�(KK��h�C             �t�bhhK ��h��R�(KK��h�C<H     e     �
        �     H     d  �        �t�bhhK ��h��R�(KK��h�C`I   /         �   �   �            �       P     %   >   2        �   �         �t�bhhK ��h��R�(KK��h�C4
   3   6      ?      #   !   ;     E        �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6            �t�bhhK ��h��R�(KK��h�CDD   _  C   -   B        �   �     6  C   �  !  �        �t�bhhK ��h��R�(KK��h�C	         �t�bhhK ��h��R�(KK��h�C<      �     �   G  &      �   �  a               �t�bhhK ��h��R�(KK��h�CS  {           �t�bhhK ��h��R�(KK	��h�C$%   B         3      �        �t�bhhK ��h��R�(KK��h�C^     �t�bhhK ��h��R�(KK��h�CD         
  8     /         �   )      m  
   �        �t�bhhK ��h��R�(KK��h�Cp�  !        �     �	           �            %   �      2  �   Y  �   �     �   �   t        �t�bhhK ��h��R�(KK	��h�C$�  �     �                 �t�bhhK ��h��R�(KK��h�CP   �  :   7      7      �      �  C      B  �  �   
     F         �t�bhhK ��h��R�(KK
��h�C(9   �  L            �  �         �t�bhhK ��h��R�(KK	��h�C$�     �     %   �            �t�bhhK ��h��R�(KK��h�C,�                 p     �        �t�bhhK ��h��R�(KK��h�Ca  �  �   �        �t�bhhK ��h��R�(KK��h�C !      �  	      	         �t�bhhK ��h��R�(KK��h�C0                  �  R              �t�bhhK ��h��R�(KK	��h�C$[      �      /      V        �t�bhhK ��h��R�(KK	��h�C$W        A  0        f     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C4      �t�bhhK ��h��R�(KK��h�C4      P         �  
   }                 �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�CD�   �  �  �
  w     |     $                         �t�bhhK ��h��R�(KK��h�C0      )   =      4   
   �   �   _         �t�bhhK ��h��R�(KK��h�C,      �        -        &        �t�bhhK ��h��R�(KK��h�CL%   �  �   �        �   J   �  C      �   {      �
  !  �        �t�bhhK ��h��R�(KK��h�C ^     �   �  
   �        �t�bhhK ��h��R�(KK��h�C8B  -            .      ;      �     @        �t�bhhK ��h��R�(KK��h�CX         &   D  0      �  >      a   �  b        v   (    j   m         �t�bhhK ��h��R�(KK��h�C5  %            �t�bhhK ��h��R�(KK��h�C8   5      �   �   L         \  |      �         �t�bhhK ��h��R�(KK
��h�C(1   #   
   T      Q              �t�bhhK ��h��R�(KK��h�C8         0   �     D           �  5        �t�bhhK ��h��R�(KK
��h�C(         i      H   A   }         �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6   �        �t�bhhK ��h��R�(KK��h�C{  b     �  �     �t�bhhK ��h��R�(KK��h�C4�
     ,            	   �   	   /  	   >     �t�bhhK ��h��R�(KK��h�C@   L  e  
     �   d   t     G   |  g   d   t        �t�bhhK ��h��R�(KK��h�C`*         E   &      \  q   �  x  +         �  $   0     *  �   �     �        �t�bhhK ��h��R�(KK��h�Cr  �     �t�bhhK ��h��R�(KK��h�C           
   �        �t�bhhK ��h��R�(KK	��h�C$5     �   �  	      	         �t�bhhK ��h��R�(KK��h�C@         .   a      �      @     �  m      �         �t�bhhK ��h��R�(KK��h�CH"         �  B   w     :      �  #       �              �t�bhhK ��h��R�(KK��h�Cd�  
   �  �  �  �      
   �     D   �  y   �              �     �              �t�bhhK ��h��R�(KK
��h�C(
        2   z   H   B   �        �t�bhhK ��h��R�(KK��h�C4      =      B  
     ^   �   �           �t�bhhK ��h��R�(KK��h�CD         m      s     �           M   �      b        �t�bhhK ��h��R�(KK��h�C<�   �  !      �  '   
   �     T  �              �t�bhhK ��h��R�(KK��h�C,2      -   �   �
  Z                 �t�bhhK ��h��R�(KK��h�Ch               �     y      W           $                        �     �        �t�bhhK ��h��R�(KK	��h�C$   (     )      �   ~        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK
��h�C(      �  �        I  	         �t�bhhK ��h��R�(KK��h�C,            �  
   �   �  �        �t�bhhK ��h��R�(KK��h�C@      	      	         �t�bhhK ��h��R�(KK��h�C       -   N      U        �t�bhhK ��h��R�(KK��h�C�            �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CT                                �       h           �         �t�bhhK ��h��R�(KK��h�C�   p      �t�bhhK ��h��R�(KK
��h�C(!      �
        	      	         �t�bhhK ��h��R�(KK��h�C             �t�bhhK ��h��R�(KK��h�C8d   8     �        �  �      D   5            �t�bhhK ��h��R�(KK��h�C1   #       �         �t�bhhK ��h��R�(KK��h�C<B  #  �  �     .      �     %        �        �t�bhhK ��h��R�(KK��h�CH      �  #            �        �   �  
   T  
  �        �t�bhhK ��h��R�(KK��h�C@   .      �     �         �  2         	           �t�bhhK ��h��R�(KK��h�C      -     �         �t�bhhK ��h��R�(KK��h�C0M      +      �  �          �        �t�bhhK ��h��R�(KK��h�C<Q  $        9                                �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C4
   Z        )   q        	     /         �t�bhhK ��h��R�(KK��h�CP'  �   [      x      G     �       �      V	  9   h     �         �t�bhhK ��h��R�(KK��h�C0V         �                 4         �t�bhhK ��h��R�(KK)��h�C�      >   $  �      �   [     �         ,                    '   �   S   }      �        D                f   �   a   ;      �        �t�bhhK ��h��R�(KK��h�C�   �   T     �t�bhhK ��h��R�(KK��h�C4U        $   �  (   N   �     �   �         �t�bhhK ��h��R�(KK��h�C   	      	      	   K      �t�bhhK ��h��R�(KK��h�C|   �      @      �     t      ~     �     �   �  x
  y
        $           ~     �     =           �t�bhhK ��h��R�(KK��h�CT#   !      �  �  %   B   u  �     %  (      
   u          F         �t�bhhK ��h��R�(KK��h�C4   �     �        �  �         +        �t�bhhK ��h��R�(KK��h�C@         O         S   Q   >      \  �      (        �t�bhhK ��h��R�(KK��h�CZ            �t�bhhK ��h��R�(KK��h�CH
   3   6   �     /         '   !      \   /                  �t�bhhK ��h��R�(KK��h�C1   #               �t�bhhK ��h��R�(KK��h�CX      (   �  
   $   E      4               8         >      �            �t�bhhK ��h��R�(KK
��h�C(              �  �           �t�bhhK ��h��R�(KK��h�C.     |        �t�bhhK ��h��R�(KK��h�C@y         =      4   >      �  +      �              �t�bhhK ��h��R�(KK��h�CD�         �  )         u         /  "   �      (        �t�bhhK ��h��R�(KK��h�C,   �  �  �   ]            �        �t�bhhK ��h��R�(KK��h�C�  R     �
  �        �t�bhhK ��h��R�(KK	��h�C$�      d        �  �        �t�bhhK ��h��R�(KK��h�C,      )   �      �  
   �  �        �t�bhhK ��h��R�(KK
��h�C({     ;     �  `     �        �t�bhhK ��h��R�(KK��h�C8      @      �   �      
   �  �     X         �t�bhhK ��h��R�(KK��h�CdD      0   4   
   _      �     P  �   �  8     4               K  ~               �t�bhhK ��h��R�(KK��h�C4   .   �   (      �  �   /      �  C         �t�bhhK ��h��R�(KK��h�Cx      M   �         `  h   t                   +   �              �   U    
        Z            �t�bhhK ��h��R�(KK��h�C     �     �t�bhhK ��h��R�(KK��h�C4   �        ;      �      �  9   �        �t�bhhK ��h��R�(KK	��h�C$f   w    �  �      �	        �t�bhhK ��h��R�(KK��h�CW   �          �t�bhhK ��h��R�(KK��h�Cp   
   A   F     �t�bhhK ��h��R�(KK��h�C 1        	      	         �t�bhhK ��h��R�(KK	��h�C$E      
     	      	         �t�bhhK ��h��R�(KK��h�C,�         
      �                 �t�bhhK ��h��R�(KK��h�CD            M      C      *        �         S        �t�bhhK ��h��R�(KK��h�C_     �t�bhhK ��h��R�(KK��h�C|�
     b     �      �        �     ,   	      	      	   K   	   �   	   �   	   I  	   U  	   �  	   �      �t�bhhK ��h��R�(KK��h�CU     �     U     �t�bhhK ��h��R�(KK��h�C   9     �t�bhhK ��h��R�(KK��h�C 1   #            �        �t�bhhK ��h��R�(KK��h�C4      =      Q  "   �     $   �   x        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C<   "     m      �t�bhhK ��h��R�(KK��h�C�   p         �t�bhhK ��h��R�(KK
��h�C(   (   I  G         8   E        �t�bhhK ��h��R�(KK��h�Ct   �  (      �   h      �        �  �              k            ;      �   
   _      {         �t�bhhK ��h��R�(KK��h�C                     �t�bhhK ��h��R�(KK��h�CP            ,                    &  *      	  �      [        �t�bhhK ��h��R�(KK��h�C0�   �     �   �   S     
   +  �        �t�bhhK ��h��R�(KK��h�Cp�   (      d  %   �   *   �      �     �            q           �     M           x        �t�bhhK ��h��R�(KK��h�C@
      ,   �	  F   '      �  �   A   �  �              �t�bhhK ��h��R�(KK��h�CdP     O  (  "      �             �     �   d     (   S     �   �      �         �t�bhhK ��h��R�(KK��h�C       	  x     k         �t�bhhK ��h��R�(KK��h�C Z      �         �        �t�bhhK ��h��R�(KK��h�CL9   �  �
     �      �  �               l      �   
   �        �t�bhhK ��h��R�(KK��h�C              �t�bhhK ��h��R�(KK��h�CH   �  L        �  #   
        f     g  )              �t�bhhK ��h��R�(KK��h�C t        �   l           �t�bhhK ��h��R�(KK��h�C0
   f   �  >   2   D  �  ,               �t�bhhK ��h��R�(KK��h�C,     �  �  d        �           �t�bhhK ��h��R�(KK	��h�C$      	     �  
   �        �t�bhhK ��h��R�(KK��h�C<|
        b        5                         �t�bhhK ��h��R�(KK#��h�C�               k                          f                 �  a   ;      �         :   W   
   �   �   _         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK
��h�C(   �  �   �         �           �t�bhhK ��h��R�(KK��h�C �  �   �        �  O      �t�bhhK ��h��R�(KK��h�C4�        �  �   �	     (  �              �t�bhhK ��h��R�(KK��h�C4     i  7                    �   7      �t�bhhK ��h��R�(KK
��h�C(      �   j    :   I            �t�bhhK ��h��R�(KK��h�C<2      -   �  C      �     .      �      �        �t�bhhK ��h��R�(KK��h�C�        {        �t�bhhK ��h��R�(KK��h�C   �                �t�bhhK ��h��R�(KK��h�C<         _  C   �   :   �     B        u        �t�bhhK ��h��R�(KK	��h�C$1   #       �     /      �      �t�bhhK ��h��R�(KK��h�C8   (      N      �     �           B        �t�bhhK ��h��R�(KK��h�CD*      a  g      +        �  g   �     .   
           �t�bhhK ��h��R�(KK��h�C l            7     �      �t�bhhK ��h��R�(KK)��h�C�            �     �        Q                                         G     ]     9      �  L   g      a        �              �t�bhhK ��h��R�(KK��h�Cq      �         �t�bhhK ��h��R�(KK��h�C�        ,   	         �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�C8#   !   '   
                        _        �t�bhhK ��h��R�(KK��h�C4q     d   t    :   �                    �t�bhhK ��h��R�(KK��h�CK     �   �     �t�bhhK ��h��R�(KK��h�C,    
   5              �        �t�bhhK ��h��R�(KK��h�C/      q     �t�bhhK ��h��R�(KK	��h�C$!      �     	      	         �t�bhhK ��h��R�(KK��h�C,   �     u  Y        �  R         �t�bhhK ��h��R�(KK
��h�C(�     
   ,            K         �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C4   @   '   H   `     �
     s              �t�bhhK ��h��R�(KK��h�C<      �     �t�bhhK ��h��R�(KK��h�C`T      D   )   6  C   ,            A   }         �	     }      �	                 �t�bhhK ��h��R�(KK��h�CHW  �        $   E   *            Z     @  �	     c         �t�bhhK ��h��R�(KK��h�CD�  �  $   �     �        0             H  �         �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   6         �        �t�bhhK ��h��R�(KK��h�C4
     '   H   �     *           �
        �t�bhhK ��h��R�(KK��h�C    
   I            �t�bhhK ��h��R�(KK��h�C<   ?   #   !   
   w
  F   
   ,                     �t�bhhK ��h��R�(KK��h�CL      �  o   �	  K  w           9  A     	  �              �t�bhhK ��h��R�(KK��h�C   {     �t�bhhK ��h��R�(KK��h�C0P     )   ;      B                    �t�bhhK ��h��R�(KK��h�Cd   2               �  �  &   �   j   �  8  �     G       %   H  �     �         �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�CL         0      �                       �   �               �t�bhhK ��h��R�(KK��h�C4   >   v   �  *      �  �   E      4         �t�bhhK ��h��R�(KK��h�C<
        �       �      |	     /   9   -        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C8        �   �  �     ,   �      Y  �        �t�bhhK ��h��R�(KK��h�C<            �        -   �       
           �t�bhhK ��h��R�(KK	��h�C$e     a      .   �             �t�bhhK ��h��R�(KK��h�C8#   !      .     	  ?      
   e   �   �
        �t�bhhK ��h��R�(KK��h�CD]  '   �          �     q  �      
   �   B   }         �t�bhhK ��h��R�(KK��h�Cl  E      E  	         �t�bhhK ��h��R�(KK��h�CX      5   �     8                   �           U                  �t�bhhK ��h��R�(KK��h�C<e   �   �   B   R      	        .   
              �t�bhhK ��h��R�(KK
��h�C(t  �  D   -   '  �   g   �        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C8�   �  &      �  K  �        K              �t�bhhK ��h��R�(KK��h�CX*      �      n     �           
   �     -   K     0      �   ~        �t�bhhK ��h��R�(KK��h�C0      =      R         G   �   �        �t�bhhK ��h��R�(KK��h�C%   �        6        �t�bhhK ��h��R�(KK��h�Cx   8   �            z  �            �  a   ;              �   �         
   _            ,        �t�bhhK ��h��R�(KK
��h�C(�  �     �  "                 �t�bhhK ��h��R�(KK��h�C   �      �t�bhhK ��h��R�(KK��h�C	     �t�bhhK ��h��R�(KK��h�C�             �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6            �t�bhhK ��h��R�(KK��h�C�       �t�bhhK ��h��R�(KK
��h�C(�      �            �  �        �t�bhhK ��h��R�(KK��h�CL'  �  c   �
     A     �     -  �     �          �        �t�bhhK ��h��R�(KK	��h�C$      �     0  �      �      �t�bhhK ��h��R�(KK��h�C,      -   �         G   �  z        �t�bhhK ��h��R�(KK��h�C>           �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C�	       �  �   _     �t�bhhK ��h��R�(KK��h�C<      J   �  �	     �         �  P  "      .     �t�bhhK ��h��R�(KK��h�C0
     �   F         �  ?              �t�bhhK ��h��R�(KK��h�C�       �t�bhhK ��h��R�(KK	��h�C$   @   '   �   |      �        �t�bhhK ��h��R�(KK��h�C@      =      n     �     $   �           �        �t�bhhK ��h��R�(KK	��h�C$�      w           <         �t�bhhK ��h��R�(KK
��h�C(#  �  �   R  y   �   r	  �  r      �t�bhhK ��h��R�(KK
��h�C(#  a  �         l  �  '  r      �t�bhhK ��h��R�(KK��h�C0      �      >
  
   @  �  /  F         �t�bhhK ��h��R�(KK
��h�C(   >   )   �  +         ,        �t�bhhK ��h��R�(KK��h�C1   #       �         �t�bhhK ��h��R�(KK��h�C,   �   �  �     m     7   �        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�CD   ?      !            8   �              
           �t�bhhK ��h��R�(KK��h�C�   R         S          �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C0   >   K        �  �     $   Z        �t�bhhK ��h��R�(KK��h�C0   �   �              Y      O         �t�bhhK ��h��R�(KK��h�CH$      >   N   �   q     �        >        �  �   �        �t�bhhK ��h��R�(KK��h�CD         5   �  �           d  �   �   
      L         �t�bhhK ��h��R�(KK	��h�C$2      -         H           �t�bhhK ��h��R�(KK��h�C�	        �t�bhhK ��h��R�(KK��h�Ch      �               �   9   �  �            a   ;      �     /         �   t        �t�bhhK ��h��R�(KK��h�C�
     ,            �t�bhhK ��h��R�(KK��h�Ce   @     �     �t�bhhK ��h��R�(KK��h�CP         O         
  Q               &      F  +   "   t         �t�bhhK ��h��R�(KK��h�CP�
  �      R     �     I   �                 �  :   C           �t�bhhK ��h��R�(KK��h�C             �t�bhhK ��h��R�(KK
��h�C(*      �   �         �     V     �t�bhhK ��h��R�(KK��h�C01   #   
   3   6              �        �t�bhhK ��h��R�(KK��h�C00        �   �      �  	      	         �t�bhhK ��h��R�(KK��h�C\      �   ;   r      �t�bhhK ��h��R�(KK��h�CT   .   W      �        H     �     �     f   w     &     �        �t�bhhK ��h��R�(KK��h�Cd                     �   ]  �      �      7   &      -   F  +           t         �t�bhhK ��h��R�(KK��h�C      z   "   �   �     �t�bhhK ��h��R�(KK��h�CL         .         o               �     &   �  �           �t�bhhK ��h��R�(KK��h�C*      j  j  /         �t�bhhK ��h��R�(KK��h�C<   �           v      �     �                 �t�bhhK ��h��R�(KK��h�C81   #      �     r  
   3   6   �     r        �t�bhhK ��h��R�(KK
��h�C(C  �   p        g  
   �        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK
��h�C(b   $     \   �                 �t�bhhK ��h��R�(KK��h�C8*      �      ;  >      a         �           �t�bhhK ��h��R�(KK
��h�C(b   �  3     �  "   W           �t�bhhK ��h��R�(KK��h�Cx      �             +      �  j   <         �   
            6  +   \      �   �      D   V         �t�bhhK ��h��R�(KK��h�C   '      �   E        �t�bhhK ��h��R�(KK��h�C8&  �   +   x      p      {      "     �        �t�bhhK ��h��R�(KK��h�C    	      	      	   K      �t�bhhK ��h��R�(KK��h�CD      5     �         �  :   s   �  
   ,               �t�bhhK ��h��R�(KK��h�Cp   �  �              ;  �     �  �  �  �  0           C
  �        �     �  V	        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C ;         	      	         �t�bhhK ��h��R�(KK	��h�C$   %   �   �  �   �  �        �t�bhhK ��h��R�(KK��h�Cq   �  �      �t�bhhK ��h��R�(KK��h�CD{  *   Y  �                   q  7   �  �  w        �t�bhhK ��h��R�(KK��h�C8   X   '   H   B   j        .         �        �t�bhhK ��h��R�(KK	��h�C$      >   >        T        �t�bhhK ��h��R�(KK��h�C@
   k  �  2      �     d      �    �  9   �        �t�bhhK ��h��R�(KK��h�C`�  �  �   -   �      �     �           \      &   6           =      �        �t�bhhK ��h��R�(KK��h�CL      G        �   �   j   �  5         =      n     �        �t�bhhK ��h��R�(KK��h�C1   #       q        �t�bhhK ��h��R�(KK��h�Cu      �   p      �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�Cr  
   ,      �t�bhhK ��h��R�(KK��h�CD   ,  '      �  �  �           �         
  |        �t�bhhK ��h��R�(KK��h�C�     X     �t�bhhK ��h��R�(KK��h�C0T   5           v                     �t�bhhK ��h��R�(KK��h�C@   ?   *     �  c      o      n  ^      
           �t�bhhK ��h��R�(KK��h�C�            �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�CL   �  �  
   �   �   _   i   X  �        A   6     0   4         �t�bhhK ��h��R�(KK��h�CB           �         �t�bhhK ��h��R�(KK��h�C  �        �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6            �t�bhhK ��h��R�(KK��h�C8   '   �  �           �  D  }             �t�bhhK ��h��R�(KK��h�CT      �   w     D  
     &     v      �     ]         �   "        �t�bhhK ��h��R�(KK
��h�C(   @   '      -   H   �   �        �t�bhhK ��h��R�(KK��h�Cd*         �   >      �  ]      W            (   �   �                 N  �        �t�bhhK ��h��R�(KK��h�CX
      F   '   �              V         P      b           b           �t�bhhK ��h��R�(KK��h�C4      D  �      5   �           +         �t�bhhK ��h��R�(KK��h�C1     
  	         �t�bhhK ��h��R�(KK��h�Cj     �t�bhhK ��h��R�(KK��h�C8M      +   3           *      �      J        �t�bhhK ��h��R�(KK��h�C   �  /         �t�bhhK ��h��R�(KK��h�CD   f     g  )     �  6  (        �  /     �         �t�bhhK ��h��R�(KK��h�CT
   H            I  $   �     �     %     �      �      �  �         �t�bhhK ��h��R�(KK��h�C8�      �
  9              j  :   �            �t�bhhK ��h��R�(KK��h�C      ;      �  r      �t�bhhK ��h��R�(KK
��h�C(         �      U   Y	  Z	        �t�bhhK ��h��R�(KK��h�C4q      �   x        �     �              �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�CX      )  W        ^   �        �  )  :   +           �  �  �        �t�bhhK ��h��R�(KK��h�C       )         �        �t�bhhK ��h��R�(KK��h�CH   '   -   A   |  �     .   >      D  *  \         +         �t�bhhK ��h��R�(KK��h�C	         �t�bhhK ��h��R�(KK	��h�C$      �	  %   �              �t�bhhK ��h��R�(KK��h�CH   .   &   2   a           �     ]  L   �   2   �   f        �t�bhhK ��h��R�(KK��h�C<�      r     �  �     I   �   �      v   o
        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C\   9   �        Z     u  �   �   j   �     5         =      n     �        �t�b�      hhK ��h��R�(KK
��h�C(@      X   R  �       X         �t�bhhK ��h��R�(KK��h�C8      �  �        �   �         b
  ?        �t�bhhK ��h��R�(KK��h�C\!      @      �        �     ,   	      	      	   K   	   �   	   U  	   /     �t�bhhK ��h��R�(KK	��h�C$         '   
   H   [        �t�bhhK ��h��R�(KK��h�C<[              �            �                 �t�bhhK ��h��R�(KK��h�C K  �   Y  	      	         �t�bhhK ��h��R�(KK��h�C0   V        H     �  �      4         �t�bhhK ��h��R�(KK��h�CP"     �        z      .   }      	     �     2     �  q        �t�bhhK ��h��R�(KK��h�C�      M     �t�bhhK ��h��R�(KK��h�C,                  �               �t�bhhK ��h��R�(KK��h�C�     �      �      �t�bhhK ��h��R�(KK��h�C        �t�bhhK ��h��R�(KK��h�C   �   �         �t�bhhK ��h��R�(KK��h�C�  
              �t�bhhK ��h��R�(KK	��h�C$9   �     �     K           �t�bhhK ��h��R�(KK��h�C          	      	         �t�bhhK ��h��R�(KK��h�C]     �t�bhhK ��h��R�(KK��h�C@*   E         5     �  
   8   [      �     �
        �t�bhhK ��h��R�(KK��h�C   �   �      �t�bhhK ��h��R�(KK��h�C      M  w     J        �t�bhhK ��h��R�(KK��h�C<y         0      4   >      �     �               �t�bhhK ��h��R�(KK��h�C<   f     g        �  )                       �t�bhhK ��h��R�(KK��h�C0!      <         	      	      	   K      �t�bhhK ��h��R�(KK��h�C       ;     �           �t�bhhK ��h��R�(KK	��h�C$�  1  '   
   e   �   F         �t�bhhK ��h��R�(KK��h�C      �     �t�bhhK ��h��R�(KK��h�CX   �
     �  a   ;                  �   �   �                         �t�bhhK ��h��R�(KK��h�C0   &   �   �   =      �   @  G   W         �t�bhhK ��h��R�(KK��h�C�   l     �           �t�bhhK ��h��R�(KK��h�CS  �
         �t�bhhK ��h��R�(KK��h�C<�  �     e  '      �   e     �  e     @         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�Ch                    �        �     �   n               i  +      �   n   �         �t�bhhK ��h��R�(KK��h�C9          �t�bhhK ��h��R�(KK��h�C!      �     �     �t�bhhK ��h��R�(KK��h�C   @   �   �     �t�bhhK ��h��R�(KK��h�C                    �t�bhhK ��h��R�(KK��h�C8      (
        i     �      G              �t�bhhK ��h��R�(KK��h�C4T   �
     �  q     c  w  
      �        �t�bhhK ��h��R�(KK��h�C@   (   )   [   *      �  
         &   �     o         �t�bhhK ��h��R�(KK��h�C !      �  	      	         �t�bhhK ��h��R�(KK��h�C\      �  2   �     :      s    �   �      v  �                 �	        �t�bhhK ��h��R�(KK��h�C   D      (   o  �      �t�bhhK ��h��R�(KK��h�CLX     "   �   ,   9     �   {     ,         "   �      9        �t�bhhK ��h��R�(KK��h�C    �  �     �  �        �t�bhhK ��h��R�(KK	��h�C$f	     �   �  8	     �        �t�bhhK ��h��R�(KK��h�C47   U  �     G     6  �     Y            �t�bhhK ��h��R�(KK��h�C@�  '   
   �   B   �              [        �        �t�bhhK ��h��R�(KK��h�C [      �         �	  �     �t�bhhK ��h��R�(KK��h�C4�  
   $   �    
   \      b              �t�bhhK ��h��R�(KK��h�CT"   �      *   �     ]  >   �   5     d   �     �     �      {        �t�bhhK ��h��R�(KK��h�Ct      ~     e   �     �t�bhhK ��h��R�(KK��h�CT      5   <      x      �     `   a
  �      M   T   �   �      �        �t�bhhK ��h��R�(KK��h�C            �  �      �t�bhhK ��h��R�(KK��h�C      �     �t�bhhK ��h��R�(KK��h�C0                       C      �     �t�bhhK ��h��R�(KK	��h�C$6  �           �           �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   6   3              �t�bhhK ��h��R�(KK��h�C         �            �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C8U     ;        O  \  (  �  U     �         �t�bhhK ��h��R�(KK��h�C,   �              �     U        �t�bhhK ��h��R�(KK��h�CHH   ~   -   �	  :   E              x        �	     N        �t�bhhK ��h��R�(KK��h�CT�   B   j  �   �  M  �   �   �     z   �
       �   �  }      �
        �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK	��h�C$A     &          *        �t�bhhK ��h��R�(KK��h�C,�     /   9   9     	      	         �t�bhhK ��h��R�(KK��h�C,#     8   �  �   $   �        r      �t�bhhK ��h��R�(KK��h�C|     �t�bhhK ��h��R�(KK��h�C   >   z   
   �        �t�bhhK ��h��R�(KK	��h�C$#   !   ?      ^   �            �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C4      -   �     �     �                  �t�bhhK ��h��R�(KK��h�C!      �     	         �t�bhhK ��h��R�(KK��h�CW   	                 �t�bhhK ��h��R�(KK��h�C m  
         �            �t�bhhK ��h��R�(KK	��h�C$#   !   ?      
   j  F         �t�bhhK ��h��R�(KK��h�C<�             H   x     0     �   >   5        �t�bhhK ��h��R�(KK��h�CL      �     �   	  �
              �   �      )      ^        �t�bhhK ��h��R�(KK��h�C�      �   �   �     �t�bhhK ��h��R�(KK
��h�C(v     H
  
   |     R           �t�bhhK ��h��R�(KK	��h�C$N     �   %     �   �        �t�bhhK ��h��R�(KK
��h�C(!      q   B     	      	         �t�bhhK ��h��R�(KK��h�C4         B          F        �        �t�bhhK ��h��R�(KK��h�C,   �   '   �     B        4        �t�bhhK ��h��R�(KK��h�C4      5   �  <      �     �  j  /        �t�bhhK ��h��R�(KK��h�CD$   �     T              t        �   l              �t�bhhK ��h��R�(KK��h�C1   #       �     �t�bhhK ��h��R�(KK	��h�C$   9     �	  9     �        �t�bhhK ��h��R�(KK��h�C@=     �   x     =  b  *           g              �t�bhhK ��h��R�(KK��h�C      �     �t�bhhK ��h��R�(KK��h�C0�     )   �             �   �        �t�bhhK ��h��R�(KK��h�C4�   C  8                     $           �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�Ct   h	       p      u      2   z      ,   �         ,   f           �  C   �        �   �        �t�bhhK ��h��R�(KK��h�C8:     -           �  
         �	  �        �t�bhhK ��h��R�(KK��h�CX                 �              +      .      l                    �t�bhhK ��h��R�(KK��h�C�  	      	         �t�bhhK ��h��R�(KK	��h�C$C     =  "      9   �        �t�bhhK ��h��R�(KK��h�C8   �  N   d   �  e  �      d        �        �t�bhhK ��h��R�(KK	��h�C$   �      _
                �t�bhhK ��h��R�(KK ��h�C�   �     p  �   2   9     ^   l  �     �     2      �  �	     2         :   O     �  F
                 �t�bhhK ��h��R�(KK	��h�C$�      �     �  �     N     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C9     �     �t�bhhK ��h��R�(KK��h�C0!         ?      
   �
  F      �        �t�bhhK ��h��R�(KK��h�CL      ;     l         �   (
       C  �     �     �        �t�bhhK ��h��R�(KK��h�C,�   7  &   �   v   �                �t�bhhK ��h��R�(KK��h�CH�  0  �     D   >   T	        .         �     �  <        �t�bhhK ��h��R�(KK��h�CL  L  "   t            �   �   E      A  "   %  .	     �        �t�bhhK ��h��R�(KK��h�C,�   �        �     	      	         �t�bhhK ��h��R�(KK	��h�C$1   #       m      �      �     �t�bhhK ��h��R�(KK	��h�C$�  �     ,  g   H  8        �t�bhhK ��h��R�(KK��h�C      �     @         �t�bhhK ��h��R�(KK��h�CX�   v           �  
   _         �          .         2   �  E        �t�bhhK ��h��R�(KK��h�C�      l  :	     �      �t�bhhK ��h��R�(KK��h�C *              "        �t�bhhK ��h��R�(KK
��h�C(   f   �   (        ^   D        �t�bhhK ��h��R�(KK��h�CL%   �  �   �        �   J   �  C      �   {      �
  !  �        �t�bhhK ��h��R�(KK��h�CD     g     �                 �        5   {	        �t�bhhK ��h��R�(KK��h�C 7      �                 �t�bhhK ��h��R�(KK��h�C�   j   �     �t�bhhK ��h��R�(KK��h�Cd                        �           �           0   �   :                     �t�bhhK ��h��R�(KK��h�C   g  k         �t�bhhK ��h��R�(KK��h�C)
     �t�bhhK ��h��R�(KK��h�CL   v  w     �   �      �      �  �  g              �        �t�bhhK ��h��R�(KK��h�C       �      �  �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C0!         �   �      �  	      	         �t�bhhK ��h��R�(KK��h�C _     �        	         �t�bhhK ��h��R�(KK��h�CdX   �   �   �      	     �     /      %   �     �     9   M        /      V        �t�bhhK ��h��R�(KK��h�C   "   �   /     �t�bhhK ��h��R�(KK��h�C1   #       q        �t�bhhK ��h��R�(KK��h�C0   /   9        C  �     ~            �t�bhhK ��h��R�(KK��h�C8q   a     �  I   �   3     o      I            �t�bhhK ��h��R�(KK��h�Cu        �t�bhhK ��h��R�(KK��h�C<I      �         �	  &   �   �      E      ,        �t�bhhK ��h��R�(KK��h�Cd   f   �   �     �      �   :   [        �  �        -   >   2   )  `     [        �t�bhhK ��h��R�(KK��h�C8�  �      �                �  �   �        �t�bhhK ��h��R�(KK��h�C,X        u  p   ;     �  �        �t�bhhK ��h��R�(KK��h�C4   @   '   H   B            �   B            �t�bhhK ��h��R�(KK*��h�C�      0   �	  �        9           �  9   z  �   k  L      �
     ]  j  �     (   �     �      �                �     Q  $           �t�bhhK ��h��R�(KK��h�C                �t�bhhK ��h��R�(KK��h�CL6  �  `   �     $   A     d  
          x  +      �         �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�Cp   5      ~  *      	  �   G   [        �   �           �         .   e	        $   �         �t�bhhK ��h��R�(KK��h�CL
   3   6      '   #   !      �               
   _      
        �t�bhhK ��h��R�(KK��h�CT*         
     �  �  :   q           =      4      �  G   H        �t�bhhK ��h��R�(KK��h�C�  	         �t�bhhK ��h��R�(KK��h�C �      e   '               �t�bhhK ��h��R�(KK��h�C     	         �t�bhhK ��h��R�(KK��h�C      �
  
         �t�bhhK ��h��R�(KK��h�Cx:            M  �  �     �   :   ?  �  Y      Q  a   ;      f   �        .   �          f        �t�bhhK ��h��R�(KK��h�C 1   �  
   3   6   �        �t�bhhK ��h��R�(KK��h�CX   �                   |  V   �  �     �      �                   �t�bhhK ��h��R�(KK��h�Cd   �   �     �t�bhhK ��h��R�(KK��h�C,�  �   |           �     �         �t�bhhK ��h��R�(KK��h�CP�   �   �  ~
     �  
   ,               �     �  )   
            �t�bhhK ��h��R�(KK��h�C<'  �  �        �      �  �        �  �         �t�bhhK ��h��R�(KK��h�C@�     �  �  *         a  #  �   �        )        �t�bhhK ��h��R�(KK��h�C{      s     �t�bhhK ��h��R�(KK��h�C<         :      r  �            �  /  �        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�CH/      O  8     �  C         ;      �  A  �      �         �t�bhhK ��h��R�(KK��h�CP      0   �  �  '   �  |     >      y         "     0   �        �t�bhhK ��h��R�(KK��h�CT*   2      E  �        2   =      ;      �  �      �         P
        �t�bhhK ��h��R�(KK��h�C�      u      �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C!      �      	         �t�bhhK ��h��R�(KK��h�C0.  �  
   ,                  /        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C         o  e
     �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�C<            +    n  �               �
        �t�bhhK ��h��R�(KK��h�CP�         &                    �         "                     �t�bhhK ��h��R�(KK��h�CF            �t�bhhK ��h��R�(KK��h�CH@         �        �   <      �     �
     �  �            �t�bhhK ��h��R�(KK��h�C8   �
  _  C   �     �	  �   }      �           �t�bhhK ��h��R�(KK��h�C,
    �      .      (     �        �t�bhhK ��h��R�(KK��h�C   }     o      �t�bhhK ��h��R�(KK��h�C[      �   M     �t�bhhK ��h��R�(KK��h�C �        	      	         �t�bhhK ��h��R�(KK��h�C4   %   e        2   �     �   
  k        �t�bhhK ��h��R�(KK��h�C4           x   �   �      �              �t�bhhK ��h��R�(KK��h�C �  �     �   ,   <        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C�  �      �     O     �t�bhhK ��h��R�(KK��h�C�   =     �t�bhhK ��h��R�(KK��h�C                �t�bhhK ��h��R�(KK��h�CP      �         t     W  �     
   c          5      &        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK	��h�C$=     l   9        	         �t�bhhK ��h��R�(KK��h�C<        �   �     �         �
     �  ?        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CH   �  c                  �   
	     �         B   �        �t�bhhK ��h��R�(KK
��h�C(U   8   �  �   *                  �t�bhhK ��h��R�(KK��h�C,�   f     g  �  {      �  	         �t�bhhK ��h��R�(KK��h�C:  q     �t�bhhK ��h��R�(KK��h�C,p      ,         I  	      	         �t�bhhK ��h��R�(KK��h�CD*      �   ~     �           +      �  z      �        �t�bhhK ��h��R�(KK��h�C,%   �        `   �     A   [        �t�be(hhK ��h��R�(KK��h�C   �        a        �t�bhhK ��h��R�(KK��h�C,   �   W           A               �t�bhhK ��h��R�(KK��h�CD   �	  }  �  :
  �   �        �  :           �        �t�bhhK ��h��R�(KK��h�C   (      �           �t�bhhK ��h��R�(KK��h�C`      -         �  �                2                 
   _      �         �t�bhhK ��h��R�(KK��h�C[      �     �t�bhhK ��h��R�(KK
��h�C(�      �  4	  9       7         �t�bhhK ��h��R�(KK��h�C8
   �   F   ?      -   1     \        +        �t�bhhK ��h��R�(KK	��h�C$q      �  �            ,     �t�bhhK ��h��R�(KK��h�C~   �            �t�bhhK ��h��R�(KK��h�C    �  �  �               �t�bhhK ��h��R�(KK
��h�C(     /      a  	      	         �t�bhhK ��h��R�(KK��h�C�  �         �   �      �t�bhhK ��h��R�(KK��h�C0m           q  G   7     G   �        �t�bhhK ��h��R�(KK��h�CPE      r     <         �  �   s     4     ^   �     s        �t�bhhK ��h��R�(KK��h�Cu     !     �t�bhhK ��h��R�(KK��h�C*      �        �t�bhhK ��h��R�(KK��h�C         �     �t�bhhK ��h��R�(KK��h�C,-   j     �  �   �        p        �t�bhhK ��h��R�(KK
��h�C(   ?   �  
   �  R     F         �t�bhhK ��h��R�(KK
��h�C(2        t        Y      O      �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�CD   D         �   9         �      �   �  �     �         �t�bhhK ��h��R�(KK��h�Cx      P   	                   
  D     *                 �   �   7   g            9  7         �t�bhhK ��h��R�(KK��h�C#     �t�bhhK ��h��R�(KK��h�C4     K     2   w   �     ~     D         �t�bhhK ��h��R�(KK	��h�C$�     �        K  �	         �t�bhhK ��h��R�(KK
��h�C(n          �                 �t�bhhK ��h��R�(KK
��h�C(      �      L   
   �           �t�bhhK ��h��R�(KK��h�Ch      ~                          �  g      �     ,   �        +   �   �            �t�bhhK ��h��R�(KK��h�C  
         �t�bhhK ��h��R�(KK��h�C   '   s   �  �        �t�bhhK ��h��R�(KK��h�Cl   ;  �  o  T   )  {  
   _            }        �   �  6        g      K              �t�bhhK ��h��R�(KK��h�C4            <	     p  &      U   �        �t�bhhK ��h��R�(KK��h�C8      =   :   �     �	  [      -     /         �t�bhhK ��h��R�(KK��h�Ct      �  8   /   '  )   g   ]         ;      N      :   8   {      �      /   �  D   �  �   7         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�CP   D         �  �   �        �  O     �      �   0     �         �t�bhhK ��h��R�(KK��h�CP                 �     d                                   �t�bhhK ��h��R�(KK��h�CL      w   �       �   �                &  *      �        �t�bhhK ��h��R�(KK��h�CP*   D   �  s   7            
  M   c   
             _  �        �t�bhhK ��h��R�(KK��h�CH   q   '   m        �     L  z  ,     �  �      �        �t�bhhK ��h��R�(KK��h�C@      =      B  =  ^   �   �        
   �  �        �t�bhhK ��h��R�(KK��h�Ch�  �   I   w  8  N  9
  �  /        c      �     �      �        �                 �t�bhhK ��h��R�(KK��h�C �        	      	   K      �t�bhhK ��h��R�(KK
��h�C(         	      	      	   K      �t�bhhK ��h��R�(KK��h�Cpq   �  �    �  O     �        �  �     �   [      <      B          �     �  p        �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�CX!         	      	      	   K   	   �   	   �   	     	   �  	   �   	   �     �t�bhhK ��h��R�(KK��h�C     �           �t�bhhK ��h��R�(KK��h�C   g  k         �t�bhhK ��h��R�(KK��h�Cl            �      �   }      &      b            "       &  *      �  L      �        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�CK
  "   �   �     �     �t�bhhK ��h��R�(KK��h�Cdu           �  �        (         �  
   �   �     I   A         �              �t�bhhK ��h��R�(KK	��h�C$   �           
           �t�bhhK ��h��R�(KK	��h�C$�      ,   �   
   4  	         �t�bhhK ��h��R�(KK��h�C<         �     7         U   0  "     N        �t�bhhK ��h��R�(KK��h�C,      V     z  9  �     �        �t�bhhK ��h��R�(KK
��h�C(�   �     �  
   s   k  "        �t�bhhK ��h��R�(KK��h�CH            �
        =  5     �   z  q  7               �t�bhhK ��h��R�(KK��h�C       }     $   0        �t�bhhK ��h��R�(KK��h�C 6  �  I                �t�bhhK ��h��R�(KK��h�C<      -   P   �   �     j   $   �     /	  �	        �t�bhhK ��h��R�(KK��h�C@   �   
   B   �           �          
   �        �t�bhhK ��h��R�(KK
��h�C(   ]   �  �         :            �t�bhhK ��h��R�(KK��h�C0/      �     0   �           V        �t�bhhK ��h��R�(KK��h�Cl"   �   -        z      �  +   c  ;     c     I   ^	  �  h   _	     �     <     =        �t�bhhK ��h��R�(KK��h�C@!      \      �      B  '   9     7  =      4         �t�bhhK ��h��R�(KK��h�C       '      B           �t�bhhK ��h��R�(KK��h�C,     �t�bhhK ��h��R�(KK��h�C0      0   �     C	     $   �   �        �t�bhhK ��h��R�(KK��h�Cp   H                      
         �        C   
   �              
   1     �        �t�bhhK ��h��R�(KK��h�C8#   !      P  (      
   u          F         �t�bhhK ��h��R�(KK��h�C1     �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�CX%	  $  o  )         �      �      o  g      $   �  �   �  W              �t�bhhK ��h��R�(KK��h�CD      �   �      D      V     h  �  C      d            �t�bhhK ��h��R�(KK��h�C@   %     )                     M        ]         �t�bhhK ��h��R�(KK��h�CD9   �     �  '         8  �     "   Q  �     @         �t�bhhK ��h��R�(KK
��h�C(-      J  /      �      �         �t�bhhK ��h��R�(KK��h�C%           �t�bhhK ��h��R�(KK��h�C<   "   �     �  -      *     �  c      �         �t�bhhK ��h��R�(KK��h�Ck              �t�bhhK ��h��R�(KK��h�C4b   #      �  "   $   �   N     i           �t�bhhK ��h��R�(KK��h�Ct%   J   �      3   �  �     �            "     !  ?     A   �     ;  C      �   -               �t�bhhK ��h��R�(KK��h�C   �        �   n      �t�bhhK ��h��R�(KK��h�Cg   �     �t�bhhK ��h��R�(KK��h�C8�         )   "     �        "               �t�bhhK ��h��R�(KK��h�C4*           |      �   &      M      +      �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK,��h�C��
     �     �
              @   �         ;      �  *    �        ,                 �           
   &        A   �  �  �   R  a        �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK&��h�C�<      �        	      	      	   K   	   �   	   �   	     	   U  	   �  	   �   	   �  	   �  	   �  	     	   )  	   �  	   >     �t�bhhK ��h��R�(KK��h�C8�   x  �     e     R         .   '  R         �t�bhhK ��h��R�(KK��h�CL�         .         �            J  +                        �t�bhhK ��h��R�(KK
��h�C(   �   �     G   I   `   �         �t�bhhK ��h��R�(KK
��h�C(   �
     �                    �t�bhhK ��h��R�(KK��h�C       /      �  	         �t�bhhK ��h��R�(KK��h�C 1  �    
   Q           �t�bhhK ��h��R�(KK��h�Cc       �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK
��h�C(      �     B         k        �t�bhhK ��h��R�(KK��h�C@
   Z        R  �  
               
      ,         �t�bhhK ��h��R�(KK��h�C�                  �t�bhhK ��h��R�(KK��h�Chp      :     �                 "       �     ;     �      J   �      �           �t�bhhK ��h��R�(KK��h�C`      _  +   
   _         $   �  �   �    W  Y  +      8   4   �            �t�bhhK ��h��R�(KK
��h�C(      0   �     A  �  �         �t�bhhK ��h��R�(KK��h�C�        (   �         �t�bhhK ��h��R�(KK'��h�C�      �      �  4   �   g      8   3  4   a  c      (         +         9   �  T   E   �  �         ;      �   y      S  �  4         �t�bhhK ��h��R�(KK��h�C4Z   �               �     K               �t�bhhK ��h��R�(KK��h�CH        �     �     �  �  +      {         �   �         �t�bhhK ��h��R�(KK	��h�C$�	     �  �      N          �t�bhhK ��h��R�(KK��h�C8   �      L        x    �   �              �t�bhhK ��h��R�(KK��h�C\I         �  
   3   F   
   I   }      -  �     ;                          �t�bhhK ��h��R�(KK��h�CP                  �     +   j   �   :   $   �   ]   �     �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C   {  �     �t�bhhK ��h��R�(KK��h�C4          *   D        Y  �  P        �t�bhhK ��h��R�(KK��h�C �      c  	   K   	   �      �t�bhhK ��h��R�(KK��h�CL      �   �     Z     �     �  �      �     q     Z         �t�bhhK ��h��R�(KK��h�CHH   o         2       �     H     H        �   �         �t�bhhK ��h��R�(KK��h�CX      5   #   %              .         &      �   �   L   G      �        �t�bhhK ��h��R�(KK��h�C@      =      �                                 �t�bhhK ��h��R�(KK��h�C8   '   )   H   �  V         0   !      [         �t�bhhK ��h��R�(KK��h�CD      E
  +      �  "   �      (     $   ?        Z     �t�bhhK ��h��R�(KK��h�C   I  ,      �t�bhhK ��h��R�(KK��h�C�     �     M     �t�bhhK ��h��R�(KK	��h�C$!      �      	      	         �t�bhhK ��h��R�(KK��h�CD   5   �  �     �     �     j      w   �      L         �t�bhhK ��h��R�(KK��h�C4�
                      %   A            �t�bhhK ��h��R�(KK��h�CW     L      N        �t�bhhK ��h��R�(KK
��h�C(b      �  �      G     ]         �t�bhhK ��h��R�(KK��h�C    @   '   )   H   �        �t�bhhK ��h��R�(KK��h�C0      �   �   
   ,            K         �t�bhhK ��h��R�(KK��h�C�      �
        �t�bhhK ��h��R�(KK��h�CP         �  j   �   �   �      w              S  %               �t�bhhK ��h��R�(KK��h�CP�                      n  I   �      �  �           �         �t�bhhK ��h��R�(KK��h�C<      �      �     �  �     i        �        �t�bhhK ��h��R�(KK��h�C<9        �   �   g         A   E      �  �         �t�bhhK ��h��R�(KK��h�C�            �t�bhhK ��h��R�(KK��h�C4      P      H   B   �        J  E         �t�bhhK ��h��R�(KK��h�C\O      Y      z     $     �     x     )  C      �  ^   |      <           �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C8   �         �  :   s   �  
   ,               �t�bhhK ��h��R�(KK��h�C�  T   �         �t�bhhK ��h��R�(KK��h�CT�  7  �     S   
     
   _      L  �  h   �      �   @     �        �t�bhhK ��h��R�(KK��h�CL            �     %                  �         C  �        �t�bhhK ��h��R�(KK��h�CL,     I     �      �  �     �   5  �            �  �        �t�bhhK ��h��R�(KK��h�C0?     `        	      	     	   �      �t�bhhK ��h��R�(KK��h�Cz  F     �     �t�bhhK ��h��R�(KK��h�C�        �      u      �t�bhhK ��h��R�(KK��h�C4#   !            ^
  (      
   �  F         �t�bhhK ��h��R�(KK	��h�C$   �  �   5      �  �        �t�bhhK ��h��R�(KK0��h�C�              �         �     �   �   1        +   
   _      8           Y  �       0  `     �             d     x      1  �   <         �  �        �t�bhhK ��h��R�(KK��h�C@�   �   $   E   
        �   �        "   �  �        �t�bhhK ��h��R�(KK
��h�C(n     �           Y      O      �t�bhhK ��h��R�(KK��h�C<*           t   &      M      +   w  �   �         �t�bhhK ��h��R�(KK��h�C<      d  &  -   *           �         �        �t�bhhK ��h��R�(KK��h�CD      5   �           �        U   �   �   �	  �	        �t�bhhK ��h��R�(KK��h�CD      5   <         �   \  &        �                  �t�bhhK ��h��R�(KK��h�C8         �  4   
   _      �        �  u     �t�bhhK ��h��R�(KK��h�C@   (   H              R  H     4   
   A   �        �t�bhhK ��h��R�(KK��h�C8]     
   4     A   u  o	  �  �      D         �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C8�  
   4      �              Y      O         �t�bhhK ��h��R�(KK��h�CD*   D   l     5  �  2   �      �      I        P	        �t�bhhK ��h��R�(KK��h�C,)   �            0                 �t�bhhK ��h��R�(KK��h�C N  �      "  +  "        �t�bhhK ��h��R�(KK��h�C�  N        �     �t�bhhK ��h��R�(KK��h�C@^   �   i  j        P   !   g      3        D
        �t�bhhK ��h��R�(KK��h�Cd   �   
   B   n                           M           
   
  n                 �t�bhhK ��h��R�(KK��h�Cp�	        t        Y      O   R     �  7         �  L      �        Y  �  i   �  7         �t�bhhK ��h��R�(KK��h�C0   "   �     �  +      }     �        �t�bhhK ��h��R�(KK��h�C4            y     &     y               �t�bhhK ��h��R�(KK��h�CL"   X   E	     g          N     B     �     �   Y  �        �t�bhhK ��h��R�(KK��h�C|�   ?     %     z     �           #     $        &
                                            �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C l  �   �        �         �t�bhhK ��h��R�(KK ��h�C�      0   <              e     �   1           k        
        �  �                 �           �t�bhhK ��h��R�(KK��h�C�         	         �t�bhhK ��h��R�(KK��h�CX   �   -   V     v                     N        Q   V      ~   �         �t�bhhK ��h��R�(KK��h�CB     R            �t�bhhK ��h��R�(KK��h�C\      �     �t�bhhK ��h��R�(KK��h�C"     �t�bhhK ��h��R�(KK��h�Cd      ;  +           �      M   �      �  
   $   �   �     �      U   G  �         �t�bhhK ��h��R�(KK��h�C?     �	     �t�bhhK ��h��R�(KK
��h�C(   	      	      	   K   	   U     �t�bhhK ��h��R�(KK��h�C@�     �  �      �     9     $  G            �     �t�bhhK ��h��R�(KK��h�C�      �        �t�bhhK ��h��R�(KK��h�C j  &   a   �      �        �t�bhhK ��h��R�(KK��h�C<      0   4   
   _      �  >      N   d   �        �t�bhhK ��h��R�(KK��h�C �  R        �
  �        �t�bhhK ��h��R�(KK��h�CH�     c        �     +   �  :   \   �         y  y         �t�bhhK ��h��R�(KK��h�C<     G     �     �      �  y      �  f        �t�bhhK ��h��R�(KK��h�C�      N      .      �t�bhhK ��h��R�(KK��h�CZ            �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK
��h�C(1   #          J  C      !        �t�bhhK ��h��R�(KK��h�C@�   �     d   8     �        d   �                 �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C:  &            �t�bhhK ��h��R�(KK&��h�C�   $   �  �   �  �   8  �   �     
  �     M    
     g   ]   &   E      4   r  �   h   �   �   g      �  
  �   
   �   E         �t�bhhK ��h��R�(KK��h�Ck  5	  	      	         �t�bhhK ��h��R�(KK��h�C8G   y        0   <      x            `        �t�bhhK ��h��R�(KK��h�C1     �       �t�bhhK ��h��R�(KK��h�C<�  '   
   �   B   �                  >  c        �t�bhhK ��h��R�(KK	��h�C$      �      [     �        �t�bhhK ��h��R�(KK��h�C1   #       j        �t�bhhK ��h��R�(KK��h�C<
   f   �        .   y     ,  2   )   9            �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�CD"   �          �   =     %   !             5
        �t�bhhK ��h��R�(KK��h�C,   &   -   a      �     �           �t�bhhK ��h��R�(KK��h�CH*            n         �      -   M      ]                 �t�bhhK ��h��R�(KK��h�CD      0   4      �   >      w   �      8   o               �t�bhhK ��h��R�(KK��h�C,         i  �  �   "   �   K        �t�bhhK ��h��R�(KK��h�C8�  �  
        
   �     �     @            �t�bhhK ��h��R�(KK��h�C E      +     �  	         �t�bhhK ��h��R�(KK��h�C�  �        8   �     �t�bhhK ��h��R�(KK��h�C,�     0   B   �  U     �            �t�bhhK ��h��R�(KK��h�C,              7	  /      �        �t�bhhK ��h��R�(KK��h�C,�  L     &   M     N              �t�bhhK ��h��R�(KK
��h�C(�   q   7  &   I     �  �        �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C^  |         	         �t�bhhK ��h��R�(KK��h�CD         �         P      +        ;  �     �         �t�bhhK ��h��R�(KK��h�C<   Q          G     J  �   0   1     x         �t�bhhK ��h��R�(KK��h�Cq      	      	         �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK	��h�C$      F        !  <         �t�bhhK ��h��R�(KK
��h�C(   �   O  �  �         �        �t�bhhK ��h��R�(KK��h�C       -   �  `   �        �t�bhhK ��h��R�(KK��h�C4      �     �        �	        c         �t�bhhK ��h��R�(KK	��h�C$�  �  )           �        �t�bhhK ��h��R�(KK	��h�C$�     `  	
  (  B   Z        �t�bhhK ��h��R�(KK��h�C X   �       �  �        �t�bhhK ��h��R�(KK��h�C�   �
  d   d        �t�bhhK ��h��R�(KK��h�C�             �t�bhhK ��h��R�(KK��h�Cd      G        �           0      �   ~        �     .   
   _      8   {         �t�bhhK ��h��R�(KK��h�CD�      �	     �     �   �   �                          �t�bhhK ��h��R�(KK��h�C@�   B   9
  �  �      �     E  
   B   �     X         �t�bhhK ��h��R�(KK	��h�C$�  �  -   �   �              �t�bhhK ��h��R�(KK��h�C,        
   �  0  +      D        �t�bhhK ��h��R�(KK
��h�C(�  (      
   _      �   R
        �t�bhhK ��h��R�(KK��h�C 2  =  <      a  	         �t�bhhK ��h��R�(KK��h�CH#   !      �               �  �  ?      
   3   �  �	        �t�bhhK ��h��R�(KK��h�Cp      9      �  L   �   �         :     e  /   9   9  7         P               :   W         �t�bhhK ��h��R�(KK��h�Cl      ,                 a   ;         �        �  )                  k               �t�bhhK ��h��R�(KK��h�C�      D      �t�bhhK ��h��R�(KK	��h�C$1   #   
   X   �  ?  F         �t�bhhK ��h��R�(KK��h�CT   &        �                �   �         )         ,  �         �t�bhhK ��h��R�(KK��h�C4j     �      I   p        �     N        �t�bhhK ��h��R�(KK��h�Cd%   M       a     o           M   c        d        �  �      A  �  z        �t�bhhK ��h��R�(KK��h�C   �   9     7      �t�bhhK ��h��R�(KK��h�C�     �  	         �t�bhhK ��h��R�(KK��h�C�   p         �t�bhhK ��h��R�(KK��h�CX         �      @                    0      �              I        �t�bhhK ��h��R�(KK��h�C4           �t�bhhK ��h��R�(KK	��h�C$Z     
   ,      
            �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�       9     �t�bhhK ��h��R�(KK��h�C   �     �     �t�bhhK ��h��R�(KK��h�C1   #       x        �t�bhhK ��h��R�(KK��h�CH
   f   [  '      5        �  
   A   }   i   ,               �t�bhhK ��h��R�(KK��h�C 	        	      	         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C1   #       �        �t�bhhK ��h��R�(KK	��h�C$      �	  %   �  +           �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CL         �     �  �   +     "     �        �   ~           �t�bhhK ��h��R�(KK��h�C@      -   M   c   I     Z
  �        .   g   b        �t�bhhK ��h��R�(KK��h�C	   >     �t�bhhK ��h��R�(KK
��h�C(   >   w   t  $   �              �t�bhhK ��h��R�(KK#��h�C�I   �   �        �         %   �      �   :   ?  �  Y   �   Q     �           �        �            �  
            �t�bhhK ��h��R�(KK��h�C�        	         �t�bhhK ��h��R�(KK��h�C*         �     �t�bhhK ��h��R�(KK��h�CH2   (      �  v                    P     �     �         �t�bhhK ��h��R�(KK
��h�C(!         =      	      	         �t�bhhK ��h��R�(KK��h�C*   D      �     �t�bhhK ��h��R�(KK��h�CL         �         m      $   2           U   �     u         �t�bhhK ��h��R�(KK��h�Cx         9      7   v     ~      X               �         �           0   x           3        �t�bhhK ��h��R�(KK
��h�C(      )   b      x   G   W         �t�bhhK ��h��R�(KK��h�CDH     �  :   �          �    `  w  �   �  V        �t�bhhK ��h��R�(KK��h�C j  &   a   �   �  �        �t�bhhK ��h��R�(KK��h�C1   #       +        �t�bhhK ��h��R�(KK��h�C,            ;  �                �t�bhhK ��h��R�(KK��h�C!            �t�bhhK ��h��R�(KK	��h�C$!         �   �      �   �     �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C4�   (            h   %     >   �            �t�bhhK ��h��R�(KK��h�C,   :   8
  
     �  	      	         �t�bhhK ��h��R�(KK	��h�C$   )  C      f     	         �t�bhhK ��h��R�(KK��h�C<      2     �   9   �	     
   �     
   �        �t�bhhK ��h��R�(KK��h�C0   5      ~        $   �      �        �t�bhhK ��h��R�(KK��h�CD�  �      �   �     �  �	     J   �  �                 �t�bhhK ��h��R�(KK��h�C�   ?   �   �   r      �t�bhhK ��h��R�(KK��h�C   '     �t�bhhK ��h��R�(KK��h�CD   �  "   |      �   �   �      +         �  �  3        �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�C,   
      �        �     �        �t�bhhK ��h��R�(KK��h�CT      0      �      8   �          �      �
     �      �  �         �t�bhhK ��h��R�(KK��h�C   �  
   H   B   }         �t�bhhK ��h��R�(KK��h�C44                 !  �   �   7            �t�bhhK ��h��R�(KK��h�C0*   z  �           �     /
           �t�bhhK ��h��R�(KK
��h�C(   (   T   $   Q     ;           �t�bhhK ��h��R�(KK��h�C0�        %   B   i  '   
   u  F         �t�bhhK ��h��R�(KK��h�C �  h              �     �t�bhhK ��h��R�(KK��h�C4   �   �  �        �      %               �t�bhhK ��h��R�(KK(��h�C��     �      �        �        �     ,   	      	      	   K   	   �   	   �   	     	   I  	   �  	   U  	   �   	   �  	   �  	        �t�bhhK ��h��R�(KK��h�C_  +   ,            �t�bhhK ��h��R�(KK	��h�C$!      �     	      	         �t�bhhK ��h��R�(KK��h�C    (   �      �
  �         �t�bhhK ��h��R�(KK��h�C8m           �           �         �        �t�bhhK ��h��R�(KK��h�CL      F     l  h      7   g      2      �   �                �t�bhhK ��h��R�(KK
��h�C(;
     )   �        0  �        �t�bhhK ��h��R�(KK��h�C�   �     .             �t�bhhK ��h��R�(KK��h�CH*               >      =      4   G   H     F  $   �        �t�bhhK ��h��R�(KK��h�C0      n  �  c   *  )      �
  z        �t�bhhK ��h��R�(KK��h�C }  �     	      	   K      �t�bhhK ��h��R�(KK��h�C?     �t�bhhK ��h��R�(KK��h�C8   @   �   ,     I        H   5     e        �t�bhhK ��h��R�(KK"��h�C�     �     �  �              &   �      
        $   n         �                                        �t�bhhK ��h��R�(KK��h�C1   #       	  l         �t�bhhK ��h��R�(KK��h�C,1   #   
   3   6   �  g  �   �        �t�bhhK ��h��R�(KK��h�Cm      �     �t�bhhK ��h��R�(KK��h�C �      :  	      	         �t�bhhK ��h��R�(KK��h�Cc  X     R        �t�bhhK ��h��R�(KK��h�C0                                   �t�bhhK ��h��R�(KK��h�CX      �         �        �   5     U   �      5                       �t�bhhK ��h��R�(KK��h�CpD      0   4   
   _      �     P  �   �  K     �   O      �        �   O      ~               �t�bhhK ��h��R�(KK��h�C8!         =        ?      
   3   6   �        �t�bhhK ��h��R�(KK��h�C       '   )   �            �t�bhhK ��h��R�(KK��h�C8   ?   #   !      .   
               _        �t�bhhK ��h��R�(KK��h�C,w  l     E     �        �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C<      /   �   :  9     r  �      �      �         �t�bhhK ��h��R�(KK��h�CT�        f   �   )              G        S   �     Q     Q         �t�bhhK ��h��R�(KK��h�C\   ;        �     �     -  �     �              �  �  �  0  ;        �t�bhhK ��h��R�(KK��h�C0O        �        ;     �   ^        �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�CL      5     <      �  
   `
           �  U  
   Z            �t�bhhK ��h��R�(KK��h�C,T              
   �
  �  �        �t�bhhK ��h��R�(KK
��h�C(/      a   -  5     f   �        �t�bhhK ��h��R�(KK��h�C4$   |  \  \            `   �               �t�bhhK ��h��R�(KK��h�C0*     5  q     )   e  i               �t�bhhK ��h��R�(KK��h�C0b   #      ]   "   �     8   �   Q         �t�bhhK ��h��R�(KK��h�C   {     �t�bhhK ��h��R�(KK
��h�C(               n             �t�bhhK ��h��R�(KK��h�C�      	      	         �t�bhhK ��h��R�(KK��h�C8%      0      +  4   *   �     �  �  7         �t�bhhK ��h��R�(KK��h�C,   �     B   3  V   �     v         �t�bhhK ��h��R�(KK��h�C�  $   E      �         �t�bhhK ��h��R�(KK��h�C`   `   �            .   Y  �  i   s   7      &   �  �  �  �      �      �        �t�bhhK ��h��R�(KK��h�C\     �      �t�bhhK ��h��R�(KK��h�C8   �   �   )     y  �     �                 �t�bhhK ��h��R�(KK��h�CZ  '   )   
   y        �t�bhhK ��h��R�(KK
��h�C(W  �     �           L         �t�bhhK ��h��R�(KK��h�C  N     �t�bhhK ��h��R�(KK	��h�C$      �  �                 �t�bhhK ��h��R�(KK��h�C,)   D   >   N   
  *   �  r  �         �t�bhhK ��h��R�(KK��h�C@�      P                          	      	         �t�bhhK ��h��R�(KK��h�C@g         �  (         �     �  5        �        �t�bhhK ��h��R�(KK��h�CH�  �  
   ,               �   
   A   }      <      &        �t�bhhK ��h��R�(KK��h�C  p   �       �t�bhhK ��h��R�(KK��h�C 1   #       4              �t�bhhK ��h��R�(KK��h�CL   (   �  7  �              �     *      :  "   �   �
        �t�bhhK ��h��R�(KK��h�C         �  
        �t�bhhK ��h��R�(KK��h�C                    �t�bhhK ��h��R�(KK��h�Clq   �  �    �  O     �        �  �     �   [      <      B          �     �        �t�bhhK ��h��R�(KK
��h�C()     �  '   
   @   �   F         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CLT      (      n   &      �      �                   ;        �t�bhhK ��h��R�(KK��h�C8�   �  2      �      J  N                    �t�bhhK ��h��R�(KK��h�C
                �t�bhhK ��h��R�(KK��h�C<�      R     8     K     �      $   �            �t�bhhK ��h��R�(KK��h�C0@   �                    �	          �t�bhhK ��h��R�(KK��h�CP*      �  
      4           (      �  !         �              �t�bhhK ��h��R�(KK��h�C03         R                          �t�bhhK ��h��R�(KK	��h�C$�  �  	      	      	   K      �t�bhhK ��h��R�(KK��h�Ct      �  �                     �           0        {     �  <   "     k     
           �t�bhhK ��h��R�(KK��h�CX   t     M     �     �  /   (   2   <            �     i     Z        �t�bhhK ��h��R�(KK��h�C4   �  M     �           8   �   o         �t�bhhK ��h��R�(KK��h�CL      '   �   @   �  �     @      �     @      �              �t�bhhK ��h��R�(KK��h�C�            �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   6   �
     �         �t�bhhK ��h��R�(KK��h�CH   @   '   )   �  v     V   X     �   S   i   ,               �t�bhhK ��h��R�(KK��h�C !              	         �t�bhhK ��h��R�(KK��h�C   �        �t�bhhK ��h��R�(KK��h�C                   �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C       #        �        �t�bhhK ��h��R�(KK��h�C86  J     	      	      	     	   �  	   �      �t�bhhK ��h��R�(KK��h�CP            ,                    &  *      	  �      [        �t�bhhK ��h��R�(KK��h�CX   S   �   �                     
        
   U        5               �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C<            $  �        .                     �t�bhhK ��h��R�(KK��h�C4      )   �          *  �      H        �t�bhhK ��h��R�(KK	��h�C$      \    �
     �        �t�bhhK ��h��R�(KK��h�CDB                       &     �     �     <        �t�bhhK ��h��R�(KK��h�C4      �
     �     �      c     \         �t�bhhK ��h��R�(KK��h�CX�   �
             
   %            H   !     
      �                 �t�bhhK ��h��R�(KK��h�C           Q      �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C      :   �      �t�bhhK ��h��R�(KK��h�C,�  �     �  �     
     -
        �t�bhhK ��h��R�(KK��h�CP   �  �        �  _  C         B     �   �   �     �   �        �t�bhhK ��h��R�(KK"��h�C��   '   
   ,                  K      �      �           I     �     U     �     �      %   B         �        �t�bhhK ��h��R�(KK��h�C0�        �  $  )   !  �              �t�bhhK ��h��R�(KK��h�C0�            
       �  �        �t�bhhK ��h��R�(KK��h�CPQ       �      ;      �   �         <     �      $  �          �t�bhhK ��h��R�(KK��h�CX         �           �        k            ;      ,  %   �           �t�bhhK ��h��R�(KK��h�C�      ,      ^     �t�bhhK ��h��R�(KK��h�C,�   R   �   	     �  C   �  '        �t�bhhK ��h��R�(KK��h�C1          �t�bhhK ��h��R�(KK��h�C�   �      �   �        �t�bhhK ��h��R�(KK��h�CL*      #     �  &      M      +   �  �	  2     D               �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C`   $   �
  Y       a     �     &      �           $   �      �  
   c        �t�bhhK ��h��R�(KK��h�CD*              c  c     &      a      �  �  A        �t�bhhK ��h��R�(KK��h�C      0   -
           �t�bhhK ��h��R�(KK��h�C0
      �   N  >   �  w   v     �        �t�bhhK ��h��R�(KK��h�CX      /                  '        ]  &      �   j          /        �t�bhhK ��h��R�(KK��h�C@   �  (              ]     >      �     
        �t�bhhK ��h��R�(KK��h�C#       %  r      �t�bhhK ��h��R�(KK��h�CZ            �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK
��h�C(n        �     	      	         �t�bhhK ��h��R�(KK��h�Cl      C   B     �  *  �             0
     �           �              *  �        �t�bhhK ��h��R�(KK��h�C1   #       �         �t�bhhK ��h��R�(KK��h�C4   e   '   �        
   B   �     4        �t�bhhK ��h��R�(KK��h�C\   �        �  
   �     &      U                  8   �     8           �t�bhhK ��h��R�(KK��h�CD   ?   !      |      <  R   
   3   6   �     �   f        �t�bhhK ��h��R�(KK��h�C<         �         0      +  ^   =  b  *        �t�bhhK ��h��R�(KK��h�C {   j   5  	      	         �t�bhhK ��h��R�(KK��h�C %   �     	      	         �t�bhhK ��h��R�(KK��h�C \   �   �      c  X  r      �t�bhhK ��h��R�(KK��h�CDx  &   N   �   �  �   �     $   �       &   N   �        �t�bhhK ��h��R�(KK��h�C8-   /   9        ;      �  �      f   �         �t�bhhK ��h��R�(KK��h�C`      �   ~              �              �      5   [         D  �   B        �t�bhhK ��h��R�(KK��h�C8       �t�bhhK ��h��R�(KK��h�C@�   3        .   <     �     �                  �t�bhhK ��h��R�(KK��h�C0      �   P     8   �   <              �t�bhhK ��h��R�(KK��h�C &     �     �  �         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�CH#   !   (      
        �     �           
      F         �t�bhhK ��h��R�(KK��h�C �         h   0        �t�bhhK ��h��R�(KK��h�C8   8   o                  ?     j            �t�bhhK ��h��R�(KK��h�CP     �   d  �     S               �
  d     W  
   1  |        �t�bhhK ��h��R�(KK��h�CD            i  
      �  �     6     c   
   �        �t�bhhK ��h��R�(KK	��h�C$         �   -      e        �t�bhhK ��h��R�(KK��h�C\      -      �      �              S   Q              v	     ?  V         �t�bhhK ��h��R�(KK��h�C1   #             �t�bhhK ��h��R�(KK��h�C,#   !      %  H  �        W         �t�bhhK ��h��R�(KK��h�C,   �      �  &   �  �   3	  I        �t�bhhK ��h��R�(KK%��h�C��      �  P   ;      �  
   �     D   5   �  [      .         6  C      ,   �      
   _         �   r  C         �  |        �t�bhhK ��h��R�(KK	��h�C$�  �           �           �t�bhhK ��h��R�(KK��h�CP*      �         �   �  (   �      �   �   �  0  �                 �t�bhhK ��h��R�(KK��h�C W   �         �   &        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK
��h�C(n        
   4  	      	         �t�bhhK ��h��R�(KK��h�C4   R      �  �     [     ,     u         �t�bhhK ��h��R�(KK��h�CD      �      ,                        �      �        �t�bhhK ��h��R�(KK	��h�C$      (   �        e        �t�bhhK ��h��R�(KK��h�C8d  
   #  �   �  �	     `        8   �        �t�bhhK ��h��R�(KK��h�C0                       �   �        �t�bhhK ��h��R�(KK��h�C      �  	      	         �t�bhhK ��h��R�(KK��h�C    �        �   �         �t�bhhK ��h��R�(KK��h�C�  �                 �t�bhhK ��h��R�(KK��h�C\      J         )   R  D   
   �   S   y  h   y  @      g       �           �t�bhhK ��h��R�(KK��h�C,T      ]     C  ]        
        �t�bhhK ��h��R�(KK��h�C   R      �        S      �t�bhhK ��h��R�(KK��h�C@      i     
   �  F      
            
            �t�bhhK ��h��R�(KK��h�C\         �            Q     �  5                  �         }  �        �t�bhhK ��h��R�(KK��h�C@      �                �     %                 �t�bhhK ��h��R�(KK��h�CX"      '      �  6     �   h  W     �     B     �  W     �     �     �t�bhhK ��h��R�(KK��h�CL      t        O         Y      Q         Q     Q      x     �t�bhhK ��h��R�(KK��h�CD   �      '   )      
         "   >     2   �   �        �t�bhhK ��h��R�(KK$��h�C�"   y        )   =         B  �           5   %                    �           �
                 >              �t�bhhK ��h��R�(KK��h�C+     �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK
��h�C(      w           r  �        �t�bhhK ��h��R�(KK��h�C      �     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C4      w   U   C     �                   �t�bhhK ��h��R�(KK��h�C8   �   �   �   �         ,   �      �   �         �t�bhhK ��h��R�(KK��h�Ch      �     9   �        Z     u  �   �   j   �     5         =      n     �        �t�bhhK ��h��R�(KK��h�C,�     �      -   �  $     8        �t�bhhK ��h��R�(KK��h�C4   5   �     v   8
     I   �   |  �	         �t�bhhK ��h��R�(KK��h�CX      J   }                    =      4      �        F              �t�bhhK ��h��R�(KK��h�CH�      =      @             m                 @        �t�bhhK ��h��R�(KK��h�C\           �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�CTG   C  (   /      �      �  <      m      -  ~     /      �           �t�bhhK ��h��R�(KK��h�C`   �      ;      �      �        �  %   �     �      �         �   �   {         �t�bhhK ��h��R�(KK��h�Cp         1
  L      �         �            	  �           �     L      �   �  �  y         �t�bhhK ��h��R�(KK��h�C<g      >      �	  $   E         �  a  g   n         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK	��h�C$f   �   �        �   m        �t�bhhK ��h��R�(KK��h�C<   f   ?     2            �  
      S           �t�bhhK ��h��R�(KK��h�C4e	       %
  �     �      m     o         �t�bhhK ��h��R�(KK��h�C0v   �  �  
            �     �        �t�bhhK ��h��R�(KK��h�CP   5      y                    ,  
                           �t�bhhK ��h��R�(KK
��h�C(      �	     ?                 �t�bhhK ��h��R�(KK��h�C=        �t�bhhK ��h��R�(KK��h�C4K       �     �  �      �     �        �t�bhhK ��h��R�(KK��h�C0      �  �  �   #   i   
   �  [        �t�bhhK ��h��R�(KK��h�C8        	      	      	     	   �  	   �      �t�bhhK ��h��R�(KK��h�C<      -   )  +         r  '  "   |      �         �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C@      ;  �  v  ;      O                         �t�bhhK ��h��R�(KK��h�CE      |
     �t�bhhK ��h��R�(KK��h�C+        �t�bhhK ��h��R�(KK��h�C@
      (      <      �      m      �         @        �t�bhhK ��h��R�(KK��h�C 
      A	  2   v  �        �t�bhhK ��h��R�(KK��h�C8g   �     2   P           �                �t�bhhK ��h��R�(KK��h�C7      �              �t�bhhK ��h��R�(KK��h�Cd%   [  -   4  `   �  �      $   h                �         �      c              �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6            �t�bhhK ��h��R�(KK��h�C,%   h          n
  �              �t�bhhK ��h��R�(KK	��h�C$      i  Q  
              �t�bhhK ��h��R�(KK��h�C�   !            �t�bhhK ��h��R�(KK��h�C8v  	      	   K   	   �   	   �   	   �  	   >     �t�bhhK ��h��R�(KK��h�C ,            q            �t�bhhK ��h��R�(KK��h�C �     �  	      	         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C p        	      	         �t�bhhK ��h��R�(KK��h�C    e     �              �t�bhhK ��h��R�(KK��h�C,�  �  �  �   %                     �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C�      9     �t�bhhK ��h��R�(KK��h�C,�                 i      �        �t�bhhK ��h��R�(KK��h�CH   d  �   (      �  
   i  �  
      9   %   �    	        �t�bhhK ��h��R�(KK��h�C,�     $   E   I  �
     {   �         �t�bhhK ��h��R�(KK��h�C      �     �      �t�bhhK ��h��R�(KK��h�CH   A       Z     �  L   i      7         �  �   �         �t�bhhK ��h��R�(KK��h�C �      l  :	     z
  �      �t�bhhK ��h��R�(KK��h�C`#   !         �   �         ?      
   �   F      
   3   6     �   �               �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C0   e   '   �   +  
   B   �     4        �t�bhhK ��h��R�(KK
��h�C(�   !        '   
   �  F         �t�bhhK ��h��R�(KK��h�C4*      �   �  [  d   8  \   l  &   �         �t�bhhK ��h��R�(KK��h�C8\   �  2   ~      �    
      �     >        �t�bhhK ��h��R�(KK��h�C�  	      	         �t�bhhK ��h��R�(KK	��h�C$%   �	     �  �              �t�bhhK ��h��R�(KK��h�C4�         �         
   z        �        �t�bhhK ��h��R�(KK��h�CL   ]   �         (        Q   V      �   y      W              �t�bhhK ��h��R�(KK��h�Ch         f     �      &   6  �      	  
   �     .   :   �     �      {      V        �t�bhhK ��h��R�(KK��h�C1       �  O         �t�bhhK ��h��R�(KK	��h�C$z                        �t�bhhK ��h��R�(KK��h�C,
        �  #      i   
   n        �t�bhhK ��h��R�(KK��h�C4        �     �   �   �   d     X         �t�bhhK ��h��R�(KK��h�CP   �     p       .   !
     A     �       9         �        �t�bhhK ��h��R�(KK��h�C@         `     �  �  5  �  %   &   �  C            �t�bhhK ��h��R�(KK��h�C    \            +         �t�bhhK ��h��R�(KK��h�CLI  (      e  "   �  
           
   �     
     �   F         �t�bhhK ��h��R�(KK��h�C�        	            �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�C<�              0      
      &  �  i   �         �t�bhhK ��h��R�(KK��h�C�     �  	         �t�bhhK ��h��R�(KK��h�CP<     )   �  +                 i  �               <  �
        �t�bhhK ��h��R�(KK��h�C,     �     `        r  /         �t�bhhK ��h��R�(KK��h�CPA              �        u      �        r  �  �   g   �        �t�bhhK ��h��R�(KK��h�CL{       '   
   H   [        %   e    '   )     
            �t�bhhK ��h��R�(KK��h�C@1   #           /         
   3   6      e  /         �t�bhhK ��h��R�(KK��h�CX^            0            �  +   *        {      �     |     o         �t�bhhK ��h��R�(KK��h�C8   �        .               >      �        �t�bhhK ��h��R�(KK��h�CP   .   �     H   
     R   �     �  #         i      h  �        �t�bhhK ��h��R�(KK��h�C8      P   �   �     �      $   �  �   �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CT                        �  c      �      |     U   8   A
  �        �t�bhhK ��h��R�(KK��h�C8           l        9   �      �  L         �t�bhhK ��h��R�(KK"��h�C�B               �  �           �    &     7        �  �           �  �              <                 �t�bhhK ��h��R�(KK��h�Cl   �    *   0     �   �        �        {      U             �   h  �     |        �t�bhhK ��h��R�(KK��h�C,   �   �	           �              �t�bhhK ��h��R�(KK��h�CL      �      M     
   \   �                              �t�bhhK ��h��R�(KK��h�C  h   t     �t�bhhK ��h��R�(KK��h�CH      
     �     �   8   4   �	  c         �     c         �t�bhhK ��h��R�(KK��h�C      �             �t�bhhK ��h��R�(KK��h�C1   #       j        �t�bhhK ��h��R�(KK��h�C      '   #           �t�bhhK ��h��R�(KK��h�C@      �        �      �     x     /      �         �t�bhhK ��h��R�(KK��h�Cl               x  V   8   �     $     >      �  +      �  �  "   Z  
   $   !  �        �t�bhhK ��h��R�(KK��h�C �                        �t�bhhK ��h��R�(KK��h�Cx      5   f  <      �            4      E      o  �      �         U   �        
     
   w        �t�bhhK ��h��R�(KK��h�C8  S     �t�bhhK ��h��R�(KK��h�CL1   #         �       �  
   3   6           �              �t�bhhK ��h��R�(KK
��h�C(P     )  L  �   7      [        �t�bhhK ��h��R�(KK��h�C       �     9            �t�bhhK ��h��R�(KK��h�C	     �     �t�bhhK ��h��R�(KK
��h�C(q   �  9      �  7   �            �t�bhhK ��h��R�(KK��h�C4      -   z   "              9          �t�bhhK ��h��R�(KK��h�CP   #     v           �  �   �  &   �         �         [        �t�bhhK ��h��R�(KK��h�CH      �      &  *      J         �    w      �   �        �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�CP   �        �     �   �  �      %  =         G         X        �t�bhhK ��h��R�(KK��h�C    '   H                  �t�bhhK ��h��R�(KK��h�C      <     `        �t�bhhK ��h��R�(KK��h�C E      E  	      	         �t�bhhK ��h��R�(KK��h�C,#   !   '   
   3   6   2              �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C4
     �  O        0   �
     !           �t�bhhK ��h��R�(KK
��h�C(   �   e     X  ,               �t�bhhK ��h��R�(KK��h�CL�
              �        &             K                  �t�bhhK ��h��R�(KK��h�C %      �         }         �t�bhhK ��h��R�(KK��h�CX~
           �        9   �                >     <         �        �t�bhhK ��h��R�(KK��h�C,           %   �  �     T        �t�bhhK ��h��R�(KK��h�C4   �   �  U  �  �	        �              �t�bhhK ��h��R�(KK��h�C<      ]     
        �  �     �     P        �t�bhhK ��h��R�(KK��h�C`%     �        K              �	     �   !      �   �     �        K        �t�bhhK ��h��R�(KK��h�C8W   �   c  �      �   l      ^        ,        �t�bhhK ��h��R�(KK��h�C�   T     �t�bhhK ��h��R�(KK��h�C�  	         �t�bhhK ��h��R�(KK
��h�C(�    �     g     7            �t�bhhK ��h��R�(KK
��h�C(  �   �  �      N     q        �t�bhhK ��h��R�(KK��h�C`!         	      	      	   �   	   �   	   I  	   �  	   /  	   s  	   )  	   �     �t�bhhK ��h��R�(KK��h�C4      N   �     �     n        "        �t�bhhK ��h��R�(KK
��h�C(�  ;  >   N   
   �  "            �t�bhhK ��h��R�(KK)��h�C�                     �   :   Y      �        Q     Q      x          �         �   �         9   $   2     )   *   $   2     X
        �t�bhhK ��h��R�(KK��h�C8      }     E   
   &     #        W         �t�bhhK ��h��R�(KK
��h�C(E      �   �      	      	         �t�bhhK ��h��R�(KK��h�Cg  �   �      �  �     �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK	��h�C$q         z                �t�bhhK ���      h��R�(KK��h�C        �     �t�bhhK ��h��R�(KK
��h�C(S        	      	   K   	   �      �t�bhhK ��h��R�(KK��h�CP      -   =      /  �
     $   |  (                 
  L         �t�bhhK ��h��R�(KK��h�C!         	         �t�bhhK ��h��R�(KK��h�C                    �t�bhhK ��h��R�(KK��h�C0   e   '   �   +  
   B   �     4        �t�bhhK ��h��R�(KK	��h�C$   �     �        6         �t�bhhK ��h��R�(KK��h�C0`   �     A   C     /  -              �t�bhhK ��h��R�(KK��h�C@      J   A     �  Z       ]   *      �  �        �t�bhhK ��h��R�(KK��h�C      �
  `   �         �t�bhhK ��h��R�(KK��h�C,   d  �      )  C      &           �t�bhhK ��h��R�(KK
��h�C(   �  �     �                 �t�bhhK ��h��R�(KK��h�C0   �  C      �  �        �   g        �t�bhhK ��h��R�(KK��h�CH�        {      �         N   y  *              {         �t�bhhK ��h��R�(KK��h�C0   n  �  )   �   .  M        '         �t�bhhK ��h��R�(KK��h�C<      �           �      a     k  G   �        �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�Ch   �  �      �        �      s   7         l  �        /                     �     �t�bhhK ��h��R�(KK��h�C    ?   �  !      �        �t�bhhK ��h��R�(KK��h�Cp*      �   F  &      �   U   $   �   N     i        V         �   L   G      o        i        �t�bhhK ��h��R�(KK��h�CpN  �     �  c         l   h        �     ,        �     Q     Q      x                 �t�bhhK ��h��R�(KK��h�CXI           F   V         P   !      �	  �     �	  `   �  �   �          �t�bhhK ��h��R�(KK��h�C0   s  �           �   o              �t�bhhK ��h��R�(KK��h�C2   (            �t�bhhK ��h��R�(KK��h�CT9   �     �  '   �     /   9   9  7   "   ~  y     
   d     @         �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C`�    $     .   �        :       �           �  �  �               �     �t�bhhK ��h��R�(KK��h�C       �  	      	         �t�bhhK ��h��R�(KK��h�CH9   �  T   $   E   �        0   �      �  "      �   \        �t�bhhK ��h��R�(KK��h�C     y     �t�bhhK ��h��R�(KK��h�C@                �t�bhhK ��h��R�(KK��h�CHW      v   c   U           �      >   w   �                �t�bhhK ��h��R�(KK��h�C,   �  �      :     
  
   �        �t�bhhK ��h��R�(KK��h�C0%   h           �   �                �t�bhhK ��h��R�(KK��h�C      p           �t�bhhK ��h��R�(KK��h�CPW   �  �      K     �      �             �      P              �t�bhhK ��h��R�(KK��h�C,�   W     l      }     �  �        �t�bhhK ��h��R�(KK��h�C0      �        �      
   N  /        �t�bhhK ��h��R�(KK��h�C,1   #       [      �      /      V     �t�bhhK ��h��R�(KK��h�C�  �         �t�bhhK ��h��R�(KK��h�C,
   )     %   �                   �t�bhhK ��h��R�(KK��h�C�        	         �t�bhhK ��h��R�(KK��h�C		     �t�bhhK ��h��R�(KK��h�C8      �   �     2   �  
      �              �t�bhhK ��h��R�(KK��h�CP      @  U       9   �  &      �   �      K     �              �t�bhhK ��h��R�(KK��h�C*      �
  +            �t�bhhK ��h��R�(KK��h�CL   <         �	  (      ^  !         x           <           �t�bhhK ��h��R�(KK��h�C@      	  u      �         �      	  u               �t�bhhK ��h��R�(KK
��h�C(G     �     �   s   d	  �        �t�bhhK ��h��R�(KK��h�CD*      �  �     �  ;  �   (     %   &   �     �         �t�bhhK ��h��R�(KK��h�C,   .     �      @      X   �        �t�bhhK ��h��R�(KK��h�C0%   �   )   �   y  !      R      �        �t�bhhK ��h��R�(KK	��h�C$      N   �     s           �t�bhhK ��h��R�(KK��h�C�          �           �t�bhhK ��h��R�(KK��h�C %  H  �  	      	         �t�bhhK ��h��R�(KK��h�CL         .   N   
  p     {      �      w     �               �t�bhhK ��h��R�(KK��h�C4�   �     �     �  �                   �t�bhhK ��h��R�(KK��h�CD   '   )      �              .      a      �            �t�bhhK ��h��R�(KK��h�C|   d   K     4   
   _         �     �      �     v     �        �  �        D   &   D  0   4         �t�bhhK ��h��R�(KK��h�C               �t�bhhK ��h��R�(KK��h�CLb   #   "   $   �   N  9   �  �     �  �   �  
   $   \  F         �t�bhhK ��h��R�(KK	��h�C$1   #       5         1  r      �t�bhhK ��h��R�(KK
��h�C(�  �        W
     �
           �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C4
              (   
         G   t         �t�bhhK ��h��R�(KK��h�C�   h                 �t�bhhK ��h��R�(KK��h�C8"   �    �           �    h  9   �        �t�bhhK ��h��R�(KK��h�C0H	  l  g      t  �      :     �        �t�bhhK ��h��R�(KK"��h�C�      =      	              �           $        	              
   \   �             Y              �t�bhhK ��h��R�(KK
��h�C(]   �           �     �         �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK	��h�C$�  �   �  �      f   W        �t�bhhK ��h��R�(KK��h�CL�     ~     �      }                       S     �        �t�bhhK ��h��R�(KK��h�CD  �  =              �                 .            �t�bhhK ��h��R�(KK��h�C	     �          �t�bhhK ��h��R�(KK��h�C   �   �
  �  %        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C        9         �t�bhhK ��h��R�(KK��h�CL"   m      @        P   <      .   "   C          $   k         �t�bhhK ��h��R�(KK��h�C@                 @  �  
   #  (                  �t�bhhK ��h��R�(KK��h�C      0   B            �t�bhhK ��h��R�(KK	��h�C$�              �           �t�bhhK ��h��R�(KK
��h�C(      -   0   I     �   s        �t�bhhK ��h��R�(KK��h�C�  	      	         �t�bhhK ��h��R�(KK��h�C r     �     �  �        �t�bhhK ��h��R�(KK��h�CP�      0     �     r  �        |        �  i   �     �        �t�bhhK ��h��R�(KK
��h�C(d     �  0  �   �   C           �t�bhhK ��h��R�(KK��h�C<�
  -  �  �   B  �
                C  V        �t�bhhK ��h��R�(KK��h�C\      e                       D             d    #     J   a         �t�bhhK ��h��R�(KK��h�C  &   N   ^        �t�bhhK ��h��R�(KK��h�C@�   q   7  (              
   _      �   �  q        �t�bhhK ��h��R�(KK��h�C|          �t�bhhK ��h��R�(KK��h�C�
     `   /      �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C      ;      �t�bhhK ��h��R�(KK��h�C,         Y  
           2
        �t�bhhK ��h��R�(KK��h�CL      -   �        �        $      �     �     9   �        �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C\   7  �      +  r      �t�bhhK ��h��R�(KK	��h�C$      -   b   �   "            �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C$  =  �  �     �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�Ch   &         �           �   }                    }     S  ]      �             �t�bhhK ��h��R�(KK
��h�C(!      t     �  	      	         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C<         P   �      �t�bhhK ��h��R�(KK*��h�C�               h   Q        O      �   S   Q   i               6  �        Q     Q      x     5         4         �     o               �t�bhhK ��h��R�(KK��h�C0     e  �   �                       �t�bhhK ��h��R�(KK��h�CH1   #      �  �     �   /   
   3   6   �     /               �t�bhhK ��h��R�(KK
��h�C(�     a   B   <     B   ?        �t�bhhK ��h��R�(KK��h�C<              �	     -      %   N   �  M        �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6            �t�bhhK ��h��R�(KK��h�C4   �   +   !      �     �        R         �t�bhhK ��h��R�(KK��h�C4V      2   I     m      0   <      [         �t�bhhK ��h��R�(KK��h�CT     �   `           �            %   �      2  �   Y     t        �t�bhhK ��h��R�(KK��h�C4�   �  �  "   �     �	     +     y        �t�bhhK ��h��R�(KK��h�C4*   �  �  A        �  �        U	        �t�bhhK ��h��R�(KK
��h�C(      )   U   K
  �  ^   �        �t�bhhK ��h��R�(KK��h�Ct
   �     
   f      �         &   �  �     �         C            �        M   �      �        �t�bhhK ��h��R�(KK��h�C,T   >      d  
   '     �
  �         �t�bhhK ��h��R�(KK��h�C\     �     �t�bhhK ��h��R�(KK��h�CL   D      �  �  7   >   2   0   d   8  �         �  d   �         �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK	��h�C$      G  �  �      �        �t�bhhK ��h��R�(KK��h�C87  &   N      ;     q   7     5  \           �t�bhhK ��h��R�(KK��h�C<�      ;     �     �           }     �        �t�bhhK ��h��R�(KK	��h�C$   Y  �        B            �t�bhhK ��h��R�(KK��h�C,   .   
   L  �
     n  �            �t�bhhK ��h��R�(KK��h�C@k     X      �  �     �     �   
   H   B           �t�bhhK ��h��R�(KK��h�CX  �
  �  �         �   �     �             �       x    S        �t�bhhK ��h��R�(KK��h�C0     �t�bhhK ��h��R�(KK��h�C�  j     u      �t�bhhK ��h��R�(KK
��h�C(   ,     0   �     �           �t�bhhK ��h��R�(KK��h�CPb      �         G         $   k         "   �     7
     u         �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK	��h�C$�          �     �  r      �t�bhhK ��h��R�(KK	��h�C$e      �  T     [  
        �t�bhhK ��h��R�(KK��h�C8�  $   E         �     �  �      
           �t�bhhK ��h��R�(KK��h�C   �         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C,   �   (         �
  9  a  
        �t�bhhK ��h��R�(KK��h�C@V     p     M   �   �        (  g  :   A   ?        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C�  �     z  �  �      �t�bhhK ��h��R�(KK	��h�C$   �      �  �   "   �        �t�bhhK ��h��R�(KK��h�Cq     �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C,0  �  �              �  �         �t�bhhK ��h��R�(KK��h�CX      '      B   R      Q  $   �     �   +      �       6  +   �         �t�bhhK ��h��R�(KK��h�C,   w  &   �   �    �               �t�bhhK ��h��R�(KK��h�CL
   �  #  2               	              S                  �t�bhhK ��h��R�(KK��h�Ch�     v  &   q  
   8        -   &      a      g  �      r
     �        	  1        �t�bhhK ��h��R�(KK��h�CLd  �  &   \           h           X        �              �t�bhhK ��h��R�(KK��h�CHf   %     �  �     9        T   5   2      2     �        �t�bhhK ��h��R�(KK��h�CH   z  �	           �t�bhhK ��h��R�(KK��h�CP      �   i     �   �  �        5      �  8   <  *      j        �t�bhhK ��h��R�(KK��h�C               �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�CP      J   a   �   
         &      �  �   $   b   ^      h  F         �t�bhhK ��h��R�(KK��h�C,"   >  �  �     �     �  5        �t�bhhK ��h��R�(KK��h�CH�   �  f     $     E      4   �           ;      �         �t�bhhK ��h��R�(KK��h�Ch     %              v   �     �      �        �     �   =      !  �  "   >        �t�bhhK ��h��R�(KK	��h�C$         
                 �t�bhhK ��h��R�(KK��h�C8     
   $   �      �  %        >   �         �t�bhhK ��h��R�(KK��h�CP#   !               ?      
   3   6   �     �                     �t�bhhK ��h��R�(KK&��h�C�V        �                �              .        ?             �
     a     
      C     ,              �        �t�bhhK ��h��R�(KK��h�C@   /         �         �  (        "               �t�bhhK ��h��R�(KK��h�C,�         �     �                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�CDB     �           $   �  j      �         $            �t�bhhK ��h��R�(KK��h�Cl         �      .  "     �         U   �   �  ^   �     s  
   �        .              �t�bhhK ��h��R�(KK��h�C�  �              �t�bhhK ��h��R�(KK	��h�C$     '   -         5        �t�bhhK ��h��R�(KK��h�C               7   v     �t�bhhK ��h��R�(KK��h�C      
     �         �t�bhhK ��h��R�(KK��h�CH      =      !  )               .   �      f     �         �t�bhhK ��h��R�(KK
��h�C(�   
         �            �     �t�bhhK ��h��R�(KK��h�C           �	  	         �t�bhhK ��h��R�(KK��h�C	     u      �     �t�bhhK ��h��R�(KK��h�C Z       �     @         �t�bhhK ��h��R�(KK��h�C@*      (   4      �  $   �     (        G  !         �t�bhhK ��h��R�(KK��h�CH   �
  _  C   �     S                  �   �             �t�bhhK ��h��R�(KK��h�C8�   -  �     p      u      J   P              �t�bhhK ��h��R�(KK��h�C0   e   '   6     #  �
     �           �t�bhhK ��h��R�(KK��h�C,v   �  �   *            �  �        �t�bhhK ��h��R�(KK��h�C4�  �      N            �   -               �t�bhhK ��h��R�(KK��h�Cd   &   �
  8  �            7                      l      S	           7        �t�bhhK ��h��R�(KK��h�C�	           �t�bhhK ��h��R�(KK
��h�C(         �  U     )      `     �t�bhhK ��h��R�(KK��h�C8      
  |        �     2   7  C   <         �t�bhhK ��h��R�(KK��h�C0      �        J  E      A   F        �t�bhhK ��h��R�(KK��h�Ct      @      �t�bhhK ��h��R�(KK��h�C8
     '   H         u     e                 �t�bhhK ��h��R�(KK��h�CT   �      A      ,     C   w      �  �     C   w      %   �   $        �t�bhhK ��h��R�(KK��h�C <   "      	      	         �t�bhhK ��h��R�(KK��h�CLN     d  E         8   %  �   :  *      �         �  �         �t�bhhK ��h��R�(KK	��h�C$   �   '   �   B   3  �        �t�bhhK ��h��R�(KK��h�C *      �     V     V     �t�bhhK ��h��R�(KK��h�CL'  �   �  ~  ?  
                  3                       �t�bhhK ��h��R�(KK��h�C<               %            
      �          �t�bhhK ��h��R�(KK��h�Cp   /         �  \        �     )   0   �        /   9   9  7         9                    �t�bhhK ��h��R�(KK��h�Cp�  !     �  !           �     �   �             �         �      �      ;     �	        �t�bhhK ��h��R�(KK��h�C4   &   �           $   E      �  4         �t�bhhK ��h��R�(KK��h�C09   �        "        �  "   ]        �t�bhhK ��h��R�(KK��h�C@%   d	        �   9   B               [  :   �        �t�bhhK ��h��R�(KK��h�Cl�     	                �   B        �      g              
                        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK	��h�C$u                         �t�bhhK ��h��R�(KK	��h�C$   =      �  	      	         �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C4      =      �            )   �   �         �t�bhhK ��h��R�(KK��h�CL*      J   }     o   &      S  d  
               �            �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�CPv  �  �   )   T      /              .   �  �         �
  �         �t�bhhK ��h��R�(KK	��h�C$   @  �     �              �t�bhhK ��h��R�(KK��h�C      y     �t�bhhK ��h��R�(KK
��h�C(   �  �     %   H  �     �      �t�bhhK ��h��R�(KK��h�Ct      
  4      $   k   '               �   .  h      �   t  
   �        %   h  k     <        �t�bhhK ��h��R�(KK��h�C,      )   �  D         �   D        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CT   �      f  *   �      �         �  �   �        �   z     �        �t�bhhK ��h��R�(KK��h�CT   8   /               .  |        U   C     �        $   k         �t�bhhK ��h��R�(KK��h�C<      J         ;  +      G     $   �   �        �t�bhhK ��h��R�(KK��h�Cd      )  +      �  "   |      �   e  "      $  |      �      
   |      <  F         �t�bhhK ��h��R�(KK��h�C4N  E      %  
   �   }                    �t�bhhK ��h��R�(KK��h�CC     �t�bhhK ��h��R�(KK��h�CL         �   J   $  D   '  g   �
        �      �   0   �        �t�bhhK ��h��R�(KK��h�CD�   l     E     �     .              �     �        �t�bhhK ��h��R�(KK��h�CL   .   �        �                V      �  �   G   [        �t�bhhK ��h��R�(KK��h�C@      )   �  c      
   y     �   �         �        �t�bhhK ��h��R�(KK��h�C	  	         �t�bhhK ��h��R�(KK��h�C0�               �      *              �t�bhhK ��h��R�(KK��h�C	  O     	         �t�bhhK ��h��R�(KK��h�C,   .           {  
      �        �t�bhhK ��h��R�(KK��h�CD              �           (      v     �           �t�bhhK ��h��R�(KK��h�CL   �   ~   �        @      e            -   P   T              �t�bhhK ��h��R�(KK��h�C        
           �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C   b     ;      y     �t�bhhK ��h��R�(KK��h�C*   &   �   P   <   r      �t�bhhK ��h��R�(KK��h�CD         .   
     �          a   _
                �t�bhhK ��h��R�(KK
��h�C(-   �  �   �     /      �         �t�bhhK ��h��R�(KK
��h�C(   ?   �     k  
      F         �t�bhhK ��h��R�(KK��h�C4�     �        �  �     $             �t�bhhK ��h��R�(KK��h�C   ]                 �t�bhhK ��h��R�(KK��h�Cd   �  �     
               8   �        G            N      �        �         �t�bhhK ��h��R�(KK��h�C   �  M  �     �t�bhhK ��h��R�(KK��h�C O     �  	      	         �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�CT�  8  �  �      �      %     o   �   �   �     
  
   �   B   }         �t�bhhK ��h��R�(KK��h�C,[      �     9        �  "   &     �t�bhhK ��h��R�(KK��h�CH   a              .                                    �t�bhhK ��h��R�(KK��h�C`                     �   ]  �   &      -   F  +           t      �           �t�bhhK ��h��R�(KK
��h�C(#   !         (      :           �t�bhhK ��h��R�(KK��h�CL-   %   l            ;         �   t           \  �   �        �t�bhhK ��h��R�(KK��h�C<�	  �   +   �      �	     2     "
  �              �t�bhhK ��h��R�(KK��h�Cd9   A            s   �  Y  f      �      	              �     	                 �t�bhhK ��h��R�(KK	��h�C$     �    D   �  O        �t�bhhK ��h��R�(KK	��h�C$   ?     e  8	     �        �t�bhhK ��h��R�(KK��h�C<   "   �  �      �t�bhhK ��h��R�(KK��h�Cx
   *  +     �   G     ,     \
  �     *           .   `                   %                  �t�bhhK ��h��R�(KK��h�CP   .   %                          �     �   B                  �t�bhhK ��h��R�(KK��h�C@      �          T   �
  `  �	  �   �   W  a        �t�bhhK ��h��R�(KK��h�C,�     �     z   "   %   �   �        �t�bhhK ��h��R�(KK��h�Cd      �      �t�bhhK ��h��R�(KK��h�C\      �	           h        �     %      �           �  f     	        �t�bhhK ��h��R�(KK��h�Cd�     $        8   L                               �      *   8   L  �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C@      R  Y      4      m     Y                      �t�bhhK ��h��R�(KK��h�CT         Y      O         =      ~          �      n     �        �t�bhhK ��h��R�(KK��h�C       �        �        �t�bhhK ��h��R�(KK��h�C<n     2     �     7  J   M   .     P  �        �t�bhhK ��h��R�(KK��h�C4�   �   �     ,     I   �  7      /         �t�bhhK ��h��R�(KK��h�CD      �   "           �   �     �                     �t�bhhK ��h��R�(KK��h�C  	      	         �t�bhhK ��h��R�(KK��h�C4
      ]  T  '   #   !         �   �        �t�bhhK ��h��R�(KK��h�C@         $   k      X            ,  %   �           �t�bhhK ��h��R�(KK��h�C      �   s   q        �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C,   >   -   )  +                    �t�bhhK ��h��R�(KK��h�CE            �t�bhhK ��h��R�(KK��h�Cl   �     
  �           �     &   2   =      4      D   h   �   �   :      �  
  �        �t�bhhK ��h��R�(KK��h�C4  �   d   :  6  �   *   �   [     �        �t�bhhK ��h��R�(KK��h�C,         �     �     �  w        �t�bhhK ��h��R�(KK��h�C0   �  C      =      n   
   �   �        �t�bhhK ��h��R�(KK��h�CDy      �      �  &      K           $   5     �        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C   e   '   �   �
        �t�bhhK ��h��R�(KK��h�C<�      �  �     {      0   <           ?        �t�bhhK ��h��R�(KK!��h�C�!            	      	   K   	   �   	     	   �  	   �  	   �   	   �  	   �  	     	      	      	      	         �t�bhhK ��h��R�(KK��h�C      �     �t�bhhK ��h��R�(KK��h�C`      b         �   �         �     @   "   k     �  "   L     ~     p         �t�bhhK ��h��R�(KK��h�C0      �   �     I   $  
   �   :        �t�bhhK ��h��R�(KK��h�CX�      2           
               o  
   �              
            �t�bhhK ��h��R�(KK
��h�C(�   g   ]   T  8   /              �t�bhhK ��h��R�(KK��h�CX   D         S   X  i   ,            (   �  [            ,               �t�bhhK ��h��R�(KK��h�C4�
  �        	      	      	   K   	   �      �t�bhhK ��h��R�(KK��h�CD   �          c           }
        0
              �t�bhhK ��h��R�(KK��h�C      �   '   "   2        �t�bhhK ��h��R�(KK��h�CX      -   U   �      K  #   !               �   �         �     Q        �t�bhhK ��h��R�(KK��h�C`!            �     �     ,   	      	   K   	     	   U  	   �  	   �   	   �     �t�bhhK ��h��R�(KK��h�C,�   �            .   �   �   R
         �t�bhhK ��h��R�(KK��h�CD      �      �   �      �       E   ^   �     s        �t�bhhK ��h��R�(KK��h�C�      /      �t�bhhK ��h��R�(KK��h�C<      -   �  
      S   �     �  "              �t�bhhK ��h��R�(KK��h�C@      �     d        �     c                     �t�bhhK ��h��R�(KK��h�C4�  )      E      4   $   �         #        �t�bhhK ��h��R�(KK��h�C               �t�bhhK ��h��R�(KK��h�CD      =      �   "   �           Y  �  7      
        �t�bhhK ��h��R�(KK��h�C q     G                 �t�bhhK ��h��R�(KK��h�C`      
   c  D        5   �   �        ]  L            s  �     �   #        �t�bhhK ��h��R�(KK��h�CDg   b     D   �     �     �     �         D   '        �t�bhhK ��h��R�(KK��h�C,}        �  �         �   f        �t�bhhK ��h��R�(KK��h�CD�     B     8   E           S   Q   V      G  ~        �t�bhhK ��h��R�(KK*��h�C�         O      �      %     z        Y      Q         Q     Q         x     �               �      �     o      >      F  $   �        �t�bhhK ��h��R�(KK��h�Cm                 �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�CPH   �        )         z      �            %   �  �     ]        �t�bhhK ��h��R�(KK��h�C0j          �        p              �t�bhhK ��h��R�(KK��h�C0%      )         �         ,   �         �t�bhhK ��h��R�(KK��h�C4      P   !      l                       �t�bhhK ��h��R�(KK��h�C!                  �t�bhhK ��h��R�(KK��h�C0#     ;      �     6     
   [        �t�bhhK ��h��R�(KK��h�C             �t�bhhK ��h��R�(KK��h�C   �	     �t�bhhK ��h��R�(KK	��h�C$�  �  "           �        �t�bhhK ��h��R�(KK��h�C`   6	  8  �        f     g  )     �  )     �   -   K  �                   �t�bhhK ��h��R�(KK��h�C0   -   
     �              5         �t�bhhK ��h��R�(KK��h�CP�         x  z  :   U     �         �   �   z     o
              �t�bhhK ��h��R�(KK��h�C,   5   �   �      ]        ;        �t�bhhK ��h��R�(KK��h�Cd%         .   �  +            ]
  c         ]     �  F       �        �         �t�bhhK ��h��R�(KK��h�Ce     �t�bhhK ��h��R�(KK��h�C0               �               �     �t�bhhK ��h��R�(KK��h�CH�          �        ?           C  D     ,           �t�bhhK ��h��R�(KK��h�C�      y  �      �t�bhhK ��h��R�(KK��h�CL      �   X  
   _                  ]     &      U   �        �t�bhhK ��h��R�(KK��h�CD         /        �     �   &      M   �      |        �t�bhhK ��h��R�(KK��h�C %   5      a   �  �         �t�bhhK ��h��R�(KK��h�C|      �         �   �     �     �      $        W           
   _      h     �         H  '        �t�bhhK ��h��R�(KK��h�C1   #       	  l         �t�bhhK ��h��R�(KK��h�C             �t�bhhK ��h��R�(KK
��h�C(H   z     �  �      �  3        �t�bhhK ��h��R�(KK
��h�C(   �     j      	      	         �t�bhhK ��h��R�(KK��h�C�       �t�bhhK ��h��R�(KK��h�CE           �t�bhhK ��h��R�(KK��h�C4V   (      <   *        n      !           �t�bhhK ��h��R�(KK��h�C H      -                  �t�bhhK ��h��R�(KK��h�CH   "	       =      ;     �  �         A   j     [        �t�bhhK ��h��R�(KK��h�C0�  ~   2            �  �
     �        �t�bhhK ��h��R�(KK��h�C,*           t   &      M      +      �t�bhhK ��h��R�(KK"��h�C�h                 �           ,   	      	      	   K   	   �   	   �   	     	   I  	   U  	   �  	   �  	   ^     �t�bhhK ��h��R�(KK��h�CL
   �  m       -   4  �   e        .   '                    �t�bhhK ��h��R�(KK��h�CD      )   b      A   �           .   �        �         �t�bhhK ��h��R�(KK��h�Cl      �     �            �   �   �      &      =      �     �     Y      O   G   H        �t�bhhK ��h��R�(KK��h�CD   5   7              �  �  7   �      M  �           �t�bhhK ��h��R�(KK��h�C0      �      L        
      F         �t�bhhK ��h��R�(KK��h�CD           !      �      ,            u   G   l        �t�bhhK ��h��R�(KK
��h�C(!               	      	         �t�bhhK ��h��R�(KK��h�CLl   9     7      u     ;      0   I   %   �     h     (         �t�bhhK ��h��R�(KK��h�C      E     �t�bhhK ��h��R�(KK��h�Cl
   .  �            x      \         �       �        �  �  �	        �    �        �t�bhhK ��h��R�(KK��h�C@      �  �                      �      �         �t�bhhK ��h��R�(KK��h�CT
   j     �
  �  7                       �   �     �     �        �t�bhhK ��h��R�(KK��h�CD�  0  �     D   >   T	     .         �     �  <        �t�bhhK ��h��R�(KK��h�C�   p      �   u      �t�bhhK ��h��R�(KK��h�C�   [         .      �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C,#   !   '   
   3   6        u        �t�bhhK ��h��R�(KK��h�C    	      	      	   K      �t�be(hhK ��h��R�(KK��h�C      �         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK
��h�C(      �        $  �           �t�bhhK ��h��R�(KK��h�CP      (   U        �     &      �  $   �      �  g     c
        �t�bhhK ��h��R�(KK��h�CT_           �   h          �           �     �  !              �t�bhhK ��h��R�(KK��h�C,      -   P   �  :   W              �t�bhhK ��h��R�(KK&��h�C�      &   �         �  �   Q     Q              �   �         9      L   T      ,     u     )      �   �  �  i   #  �         �t�bhhK ��h��R�(KK��h�CD4     R  4     
   \         �                       �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6            �t�bhhK ��h��R�(KK��h�C,�        �   �     {      �        �t�bhhK ��h��R�(KK��h�C`7         4        K  ;               �  �                              �t�bhhK ��h��R�(KK��h�C8      P                  >  ^   �   n        �t�bhhK ��h��R�(KK��h�C\      >   �           �       $   n         0   �     ]      $   k         �t�bhhK ��h��R�(KK��h�C#  �  �   �   r      �t�bhhK ��h��R�(KK��h�C@�      )   �     M      0  �  �         J  <        �t�bhhK ��h��R�(KK��h�Cm      �      �     �t�bhhK ��h��R�(KK��h�C8�     �                       �  �         �t�bhhK ��h��R�(KK��h�Cl      5   �  [      %     :  �  
   _      �        &      =      �   ^   E      g        �t�bhhK ��h��R�(KK��h�C �     �  [     �        �t�bhhK ��h��R�(KK��h�C\f   l         .   �     l      �        �     �     %   �  !  j   <         �t�bhhK ��h��R�(KK��h�C[                 �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C             �t�bhhK ��h��R�(KK��h�CX         �  "   �   n          n  �      ^   �  E                     �t�bhhK ��h��R�(KK��h�CX         /   9   �  7      1     �  +      M   �      C     �           �t�bhhK ��h��R�(KK��h�CH@   �   �   R      l      �        .        �     
        �t�bhhK ��h��R�(KK��h�CL�      L   "        M      +      �  �     �	        �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK	��h�C$�     ;     /   9   -        �t�bhhK ��h��R�(KK	��h�C$�   �      �   :   $           �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C4�      k	        �        �  ;  �         �t�bhhK ��h��R�(KK��h�C4                     J     �   l         �t�bhhK ��h��R�(KK	��h�C$�    2   �     �   h        �t�bhhK ��h��R�(KK��h�C\   �         �t�bhhK ��h��R�(KK
��h�C(            &   �  
   �         �t�bhhK ��h��R�(KK��h�CX         ;  �  �      �      l  �  :      �  T   E         A   �        �t�bhhK ��h��R�(KK��h�CL         O         Q   �  Y      >      =      4               �t�bhhK ��h��R�(KK��h�C \   �  m  r   ,   	         �t�bhhK ��h��R�(KK��h�C             �t�bhhK ��h��R�(KK��h�C�	          �t�bhhK ��h��R�(KK��h�C8H  [  H
  
   $            R  H              �t�bhhK ��h��R�(KK��h�C%   !  �   �  
        �t�bhhK ��h��R�(KK
��h�C(-   H   �   o   �         /         �t�bhhK ��h��R�(KK��h�C =
  ;           �        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C1        �   �        �t�bhhK ��h��R�(KK��h�C<'  
   q      �      M              �           �t�bhhK ��h��R�(KK��h�CP   �          �   �   (               �   �     (               �t�bhhK ��h��R�(KK��h�CX   D         �      �        �        �  0     �   �      �   �         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK-��h�C�   J    
   _      }     �     �     }      d     �     �                   �     h     �     �  q     �   �         $           �         �t�bhhK ��h��R�(KK��h�C\   B        .   N         ]           V  �	           �   �     �         �t�bhhK ��h��R�(KK��h�C4�	     �  �   �  �   8  �   �        �     �t�bhhK ��h��R�(KK��h�C I            0   4         �t�bhhK ��h��R�(KK��h�ChO      �     Q     z     )  C      �  
   y     |      <  "  �  �     R   "        �t�bhhK ��h��R�(KK��h�CX
   3   6   �
  ?      #   !      \        n      A   �      Q     �         �t�bhhK ��h��R�(KK��h�CHW  �     )  +   -   �   g   �      X        �              �t�bhhK ��h��R�(KK��h�C0�
  �     %   l      v
  C              �t�bhhK ��h��R�(KK��h�Cm     �      �t�bhhK ��h��R�(KK��h�C �     �  	      	         �t�bhhK ��h��R�(KK��h�Cn          �t�bhhK ��h��R�(KK��h�C [      -     �  	         �t�bhhK ��h��R�(KK��h�C
   ,      Z         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   6   �              �t�bhhK ��h��R�(KK��h�C8       �   :   U                          �t�bhhK ��h��R�(KK��h�C    5   -      o  ~        �t�bhhK ��h��R�(KK��h�C4-   D        2     (  &   �               �t�bhhK ��h��R�(KK��h�C@   �      ,  ~  l         �  �            v
        �t�bhhK ��h��R�(KK��h�CH�  :   �        �
  �     ,            X        A   }      �t�bhhK ��h��R�(KK��h�C\%     m  �            �  c           �     �   �
             �        �t�bhhK ��h��R�(KK��h�C8[  L  
   y       �   �   M     {  _        �t�bhhK ��h��R�(KK��h�CH   r  �     L  �     +      �      (           �        �t�bhhK ��h��R�(KK��h�C�   R      �     �t�bhhK ��h��R�(KK��h�C 1        	      	         �t�bhhK ��h��R�(KK	��h�C$�	                �        �t�bhhK ��h��R�(KK��h�C02   5           �   :      .   �        �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C�      y  �      �t�bhhK ��h��R�(KK��h�CT      :  �      J   �            n  5         4   
   _      �        �t�bhhK ��h��R�(KK��h�C,�      �     �  �      �
     �     �t�bhhK ��h��R�(KK��h�C8      �     W     *      �     �          �t�bhhK ��h��R�(KK��h�CP           �  
   �  &      U      "   �	     j      
           �t�bhhK ��h��R�(KK��h�C      |        �t�bhhK ��h��R�(KK��h�C  I   _  �  �        �t�bhhK ��h��R�(KK��h�C0?  V      �      �  �  	      	         �t�bhhK ��h��R�(KK��h�C,Z      �     �  �      �     �     �t�bhhK ��h��R�(KK��h�C@
   �     G     %   �         �           �        �t�bhhK ��h��R�(KK
��h�C(      -   i     ?
     �        �t�bhhK ��h��R�(KK��h�CC  �   $
     �t�bhhK ��h��R�(KK��h�C 4       t      n        �t�bhhK ��h��R�(KK
��h�C(      �   �     �	  ;           �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�CDf   5     �       �  �          �  {      �         �t�bhhK ��h��R�(KK��h�CZ          �            �t�bhhK ��h��R�(KK��h�Cf   �              �t�bhhK ��h��R�(KK��h�C�  �           �t�bhhK ��h��R�(KK	��h�C$   ?   �       
           �t�bhhK ��h��R�(KK��h�C@      b   #      '     �  "   l     |      �         �t�bhhK ��h��R�(KK��h�C8"      l  >  �      E     H        �        �t�bhhK ��h��R�(KK��h�CP         '     %      N         ,   )               �   S         �t�bhhK ��h��R�(KK6��h�C�         
  L   i                 &      -   )  ]      W      �     �             �   �               �      A     7         $   ;         �   �         �   9   $   �  �         �t�bhhK ��h��R�(KK��h�CX
        q           '      H     %        P      &        z	        �t�bhhK ��h��R�(KK��h�CP       h  �   h   H         �         �      J   �  
           �t�bhhK ��h��R�(KK��h�C0�    �     /         	      	         �t�bhhK ��h��R�(KK��h�CT      ;            .   T            �     �              �
        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�Cy  <      
     �t�bhhK ��h��R�(KK��h�CX            �  �      u  *     *     �      �  u  ;  �               �t�bhhK ��h��R�(KK��h�C8g   (  )     .  M        ,   �     �        �t�bhhK ��h��R�(KK��h�C8B   P          �     �     �     �        �t�bhhK ��h��R�(KK1��h�C�           �     I        3  }          }              e
     �     }      d     �     �     �     h     �  q     �   �   �     $  P     �  �         �t�bhhK ��h��R�(KK��h�CD   &   �  +      N  �        Q   V         $   Z        �t�bhhK ��h��R�(KK��h�C,�      �     �  �      �
     �     �t�bhhK ��h��R�(KK��h�C4�     e   �     :               �        �t�bhhK ��h��R�(KK��h�C     �   
        �t�bhhK ��h��R�(KK��h�C,!         �         	      	         �t�bhhK ��h��R�(KK��h�C<           m         b      x   G   Q  �        �t�bhhK ��h��R�(KK��h�Cd        �t�bhhK ��h��R�(KK��h�C�  	      	         �t�bhhK ��h��R�(KK��h�C8�     @   �   =     0  i   %      �   =        �t�bhhK ��h��R�(KK��h�C(   @        �t�bhhK ��h��R�(KK��h�C\      �              �     �   x      �      -  �  �      |	              �t�bhhK ��h��R�(KK��h�CX  �	     �t�bhhK ��h��R�(KK��h�C   X         �t�bhhK ��h��R�(KK��h�C,   &   �     �   �     s   �        �t�bhhK ��h��R�(KK��h�C-     �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK	��h�C$   �   
   C   �   N
           �t�bhhK ��h��R�(KK��h�CR      �     �t�bhhK ��h��R�(KK��h�CH   S   
              '      �     *           �
        �t�bhhK ��h��R�(KK��h�C@o        �      b        ;     �  c      �        �t�bhhK ��h��R�(KK	��h�C$p  L  
   t      �           �t�bhhK ��h��R�(KK��h�C8�        �  
     }   V   I         �        �t�bhhK ��h��R�(KK��h�CL         
   n           �     
      �       
   J        �t�bhhK ��h��R�(KK��h�C3     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C �  �   T     d   �        �t�bhhK ��h��R�(KK��h�CD1   #      �  
   3   �       u       g   d   t        �t�bhhK ��h��R�(KK��h�CT   /            S   X  i   ,         _  C   ,            �  }         �t�bhhK ��h��R�(KK	��h�C$1   #       ,         �         �t�bhhK ��h��R�(KK��h�CP
             R  �     �          �     	     �   S         �t�bhhK ��h��R�(KK��h�C<�   &      	  <  N   $   k         �  �   n        �t�bhhK ��h��R�(KK��h�C8E   &   r  �   �  �   y      5   �  h   p        �t�bhhK ��h��R�(KK��h�C01   
   �   I  *   \    c      M        �t�bhhK ��h��R�(KK��h�CD*      5   <      �        �     �     k  j  /        �t�bhhK ��h��R�(KK��h�C�      4      �t�bhhK ��h��R�(KK��h�C       Z  (   �  [        �t�bhhK ��h��R�(KK��h�C               �t�bhhK ��h��R�(KK��h�CD�             �     %   �     5     �      <        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK0��h�C�
        1     S      }        �  ~      �   �   S     G      K        �     �        �       /      B    
   $      
   �   F      "      W      �        �t�bhhK ��h��R�(KK��h�C<      �      �t�bhhK ��h��R�(KK��h�C<�         0     *           �   7               �t�bhhK ��h��R�(KK��h�C<      �                �  0                 �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�Ch
   3   6   �     �      �  '   3     '        �  +         0   <   "   m      @        �t�bhhK ��h��R�(KK��h�C�     ,     �t�bhhK ��h��R�(KK��h�C          A  �  �         �t�bhhK ��h��R�(KK��h�C,*      /   �     (   D   o  �         �t�bhhK ��h��R�(KK��h�C@   P        >   4  c   �  �      v   %      �        �t�bhhK ��h��R�(KK��h�C@      B  Q         �  *  �  i         q            �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK
��h�C(      0        	     
        �t�bhhK ��h��R�(KK��h�C,   �  '   !      .     H   ?        �t�bhhK ��h��R�(KK��h�C4      �     �t�bhhK ��h��R�(KK��h�C	  	         �t�bhhK ��h��R�(KK��h�C|         '   �   >     8         q   i
     &      �   �                  :   D     8   E     t         �t�bhhK ��h��R�(KK��h�Cl   �      >     �     l      J   }     o            �      �      �        �   o         �t�bhhK ��h��R�(KK��h�C@*      ]  &   2   �  \   �   �     `  V  �           �t�bhhK ��h��R�(KK��h�C�
     ,            �t�bhhK ��h��R�(KK��h�C,                 	      	         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CP
         �  �   H               	                 h  �        �t�bhhK ��h��R�(KK��h�C�  �  �        r      �t�bhhK ��h��R�(KK��h�C4      �     �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   6   2              �t�bhhK ��h��R�(KK��h�C4H   �  �   �	           l      I           �t�bhhK ��h��R�(KK��h�CH   �     �     %   J   #  �         �           �         �t�bhhK ��h��R�(KK��h�C1   #       �        �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C�     %     �t�bhhK ��h��R�(KK��h�CT   (   �   j        �  �  V   �     �      �     
        �        �t�bhhK ��h��R�(KK��h�C4   P                 F     �  �        �t�bhhK ��h��R�(KK
��h�C(     �  �  �         7         �t�bhhK ��h��R�(KK��h�CL   f   �   (         &  �   D        	  �     �             �t�bhhK ��h��R�(KK��h�CH            �   �     �  {      2         ,               �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK'��h�C�   8   o      o        >    �            �  �   %              0      L
     &      b            0      �     �  G           �t�bhhK ��h��R�(KK��h�Cx�      Y        	      	      	   �   	   �   	   I  	   /  	   s  	   )  	   �  	   �  	   �  	   �     �t�bhhK ��h��R�(KK
��h�C(      �     L     G          �t�bhhK ��h��R�(KK��h�CL0   o  �           i     �                �              �t�bhhK ��h��R�(KK
��h�C(�   &      v            �         �t�bhhK ��h��R�(KK
��h�C(   �              r  s        �t�bhhK ��h��R�(KK��h�C4�     j              b         �        �t�bhhK ��h��R�(KK��h�C+  5  	      	         �t�bhhK ��h��R�(KK��h�C0"   m         b   x   G   �     �        �t�bhhK ��h��R�(KK��h�C         �        �t�bhhK ��h��R�(KK��h�C8   /   9   -  L              �  �  �        �t�bhhK ��h��R�(KK��h�CL*      #     �  &      M      +   �  �	  2     D               �t�bhhK ��h��R�(KK��h�C �     ^     �   �        �t�bhhK ��h��R�(KK��h�CD      z      .      S   }         �     	     �        �t�bhhK ��h��R�(KK
��h�C(   '      �   �  
   V  F         �t�bhhK ��h��R�(KK��h�C4m     ]                  �	     �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C4      F  +   "   @   �  "   t      ~        �t�bhhK ��h��R�(KK��h�C8         Y      O         �     �            �t�bhhK ��h��R�(KK
��h�C(!      k     '   
   �           �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK$��h�C�-   A   6     ,   O   i      �  �   �        8     8       /        /         f   �   0   4         
   _      �        �t�bhhK ��h��R�(KK��h�CD+  "   @   �   @     �  �   u   �     4        C         �t�bhhK ��h��R�(KK��h�C   	  �          �t�bhhK ��h��R�(KK��h�C1               �t�bhhK ��h��R�(KK��h�C,T   �  H   a  
   B   �     @         �t�bhhK ��h��R�(KK��h�CL!         P   {         ?      
   3   6       �   ?   �   �   r      �t�bhhK ��h��R�(KK	��h�C$     @   �                 �t�bhhK ��h��R�(KK��h�C       �   �   c   U        �t�bhhK ��h��R�(KK��h�CZ   �     �t�bhhK ��h��R�(KK��h�C`      �     s   �     �              ,   	      	   K   	   �   	   I  	   �     �t�bhhK ��h��R�(KK��h�CL   �  (      �  )                  k         4               �t�bhhK ��h��R�(KK��h�C,      �  �  �
     �      7         �t�bhhK ��h��R�(KK��h�C       f     F  �         �t�bhhK ��h��R�(KK��h�C      f  �     �t�bhhK ��h��R�(KK��h�C+  �             �t�bhhK ��h��R�(KK��h�C0               �     �              �t�bhhK ��h��R�(KK��h�C8	          I        "   T                 �t�bhhK ��h��R�(KK��h�C   
   j  �        �t�bhhK ��h��R�(KK��h�CD  w  2     @               O           �           �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK	��h�C$�    
   ,      
            �t�bhhK ��h��R�(KK��h�C@`     �      �     %   �      �  �  �     `        �t�bhhK ��h��R�(KK��h�C8   (   �  1     \      �     �  "            �t�bhhK ��h��R�(KK��h�C4   e   '   �      V   2            !        �t�bhhK ��h��R�(KK��h�C )                        �t�bhhK ��h��R�(KK��h�ClX   �   R      u      g        �   +   !      �     @     �        �      B      R         �t�bhhK ��h��R�(KK��h�CH      &   �                    )   �         j   4         �t�bhhK ��h��R�(KK��h�C`   H       *  �   
   $              ;      �   9   �  T            �        �t�bhhK ��h��R�(KK��h�C�     �     �     �t�bhhK ��h��R�(KK��h�C8      �   �      �      L        
           �t�bhhK ��h��R�(KK��h�C8   �     w     �      (                    �t�bhhK ��h��R�(KK��h�Cu     	         �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�C�	     �     
        �t�bhhK ��h��R�(KK��h�C�        	         �t�bhhK ��h��R�(KK��h�C �      M        �         �t�bhhK ��h��R�(KK��h�C�       �     �t�bhhK ��h��R�(KK��h�CLM   �            �     s        �        �  �              �t�bhhK ��h��R�(KK��h�C<�     X     2        >  ^   �   |      �        �t�bhhK ��h��R�(KK��h�CX      5   x      [         �       p      ,   �      U   @   �            �t�bhhK ��h��R�(KK��h�C\      0   R  B           �  D  J  
   +         .                        �t�bhhK ��h��R�(KK��h�C@0     ;      
   8  0      �     �   *   x  {        �t�bhhK ��h��R�(KK��h�C         !           �t�bhhK ��h��R�(KK��h�CX�  �  "   >     �        �        �           �         :  �         �t�bhhK ��h��R�(KK��h�C<         	         �t�bhhK ��h��R�(KK��h�C�   ~     �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C<T      H   z  
           @        
            �t�bhhK ��h��R�(KK��h�C|         
     �     �	     �      �	  9   �   L   
   y     M   �            �  �   �   
   N           �t�bhhK ��h��R�(KK��h�C<  �     �   p        �t�bhhK ��h��R�(KK
��h�C(!         	      	      	   K      �t�bhhK ��h��R�(KK��h�C	  l      �t�bhhK ��h��R�(KK
��h�C(         H   �	                 �t�bhhK ��h��R�(KK��h�C�  F      �t�bhhK ��h��R�(KK��h�C      u      �t�bhhK ��h��R�(KK��h�C,            �          E        �t�bhhK ��h��R�(KK��h�CP      b      x   "   �     �        \     
        $   k         �t�bhhK ��h��R�(KK��h�C0h        .               �           �t�bhhK ��h��R�(KK��h�C0      r       %   �
     �  �
        �t�bhhK ��h��R�(KK��h�CD�       L  
   `     �       9  7   '     7         �t�bhhK ��h��R�(KK��h�C     e      �t�bhhK ��h��R�(KK��h�Cl   f   w     :  -     c      M              $   �  �   �          �   �               �t�bhhK ��h��R�(KK��h�C@   e          q  �
             p	  
   `
        �t�bhhK ��h��R�(KK
��h�C(  '   �           #            �t�bhhK ��h��R�(KK��h�C,      �  �     A   �  :            �t�bhhK ��h��R�(KK��h�CD�   �     �  �	     �   
              �   "   �        �t�bhhK ��h��R�(KK��h�CP   >   =         �  4   
   _      {   y   8   4      �    c         �t�bhhK ��h��R�(KK��h�C1         �t�bhhK ��h��R�(KK��h�C*     p     �      �t�bhhK ��h��R�(KK��h�C4   ?      �  �   >     ,   
   �	  F         �t�bhhK ��h��R�(KK��h�C0�      �           �  V     H        �t�bhhK ��h��R�(KK��h�C<   @   '   )   A           .   "         �        �t�bhhK ��h��R�(KK��h�C       #      i            �t�bhhK ��h��R�(KK��h�C�              �t�bhhK ��h��R�(KK��h�C\�     �  +            ]
  c         ]     �  F     �          �         �t�bhhK ��h��R�(KK��h�C8`            0   4         
   _      �        �t�bhhK ��h��R�(KK��h�C<
   f   [     �     >     
         �   �        �t�bhhK ��h��R�(KK��h�C<I      0   �                          �         �t�bhhK ��h��R�(KK��h�C b   #      $   �  h        �t�bhhK ��h��R�(KK��h�CB          �t�bhhK ��h��R�(KK��h�C4   �   '   �   5     Q	     �  �   �        �t�bhhK ��h��R�(KK��h�CT^   
  �        �   L   
        b   �     x      F     �  �         �t�bhhK ��h��R�(KK	��h�C$   �                      �t�bhhK ��h��R�(KK��h�C8�
        	      	      	   K   	   U  	   /     �t�bhhK ��h��R�(KK��h�C>
     5     �t�bhhK ��h��R�(KK��h�C�  	      	         �t�bhhK ��h��R�(KK��h�C81   #   
   3   6         2   =      o  �   r      �t�bhhK ��h��R�(KK��h�C     /   9   9  7      �t�bhhK ��h��R�(KK��h�C,#   !      ]   '   
   3   6            �t�bhhK ��h��R�(KK
��h�C(!      4         	      	         �t�bhhK ��h��R�(KK��h�C1   #   
   3   6   �     �t�bhhK ��h��R�(KK��h�CP         '      Z	  
   �           G           U   8           �t�bhhK ��h��R�(KK��h�C�  �  �         �t�bhhK ��h��R�(KK��h�C E            �   �         �t�bhhK ��h��R�(KK��h�C8�         (   -     �   �                    �t�bhhK ��h��R�(KK��h�CX!      �        �           f     �  
   ,                  K         �t�bhhK ��h��R�(KK	��h�C$     �     �   u  C        �t�bhhK ��h��R�(KK��h�CH|  �  �     �   �  &   �      	     �     {     J        �t�bhhK ��h��R�(KK��h�C@      �  ?           r     .   ^      �           �t�bhhK ��h��R�(KK
��h�C(      ;      �   g               �t�bhhK ��h��R�(KK��h�CZ     �t�bhhK ��h��R�(KK��h�CP            ;      �   %   �   �        P   <   
      �   D        �t�bhhK ��h��R�(KK��h�C             �t�bhhK ��h��R�(KK��h�CT                    �     �      �        &      U   $   N        �t�bhhK ��h��R�(KK��h�CE      �t�bhhK ��h��R�(KK��h�CH#   !      �     �   (         W      $   5                �t�bhhK ��h��R�(KK��h�C      �  	         �t�bhhK ��h��R�(KK��h�C,   �
                            �t�bhhK ��h��R�(KK��h�Ch
         �  �     z     �     S     �  #   �         �  �     �  i               �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C   �  �      �         �t�bhhK ��h��R�(KK��h�C0   '   )   -  �  �	                    �t�bhhK ��h��R�(KK��h�C�	           �t�bhhK ��h��R�(KK��h�CD�       8   ~     `   1          �                 �t�bhhK ��h��R�(KK��h�CD#   !      �  '   
   @     �        �        F         �t�bhhK ��h��R�(KK��h�CD   �       �     �   �     �
     �         �
  r      �t�bhhK ��h��R�(KK��h�C�        	         �t�bhhK ��h��R�(KK��h�C	  E	         �t�bhhK ��h��R�(KK��h�C4      �t�bhhK ��h��R�(KK��h�C8�  E   �  )   ]  \   �          :  �         �t�bhhK ��h��R�(KK
��h�C(1   #      �  
   3   6   t        �t�bhhK ��h��R�(KK��h�C !         �   �            �t�bhhK ��h��R�(KK��h�C_     �         �t�bhhK ��h��R�(KK��h�C01   #      �        
   3   6   N	        �t�bhhK ��h��R�(KK��h�C       ?        *        �t�bhhK ��h��R�(KK
��h�C(�   &   2     �         �        �t�bhhK ��h��R�(KK��h�CX     �   -   �        i            [         �  �  �      D         �t�bhhK ��h��R�(KK��h�CH         0   4      �        j      �  �  :   q           �t�bhhK ��h��R�(KK��h�C0         �  J  �  #         M        �t�bhhK ��h��R�(KK��h�C<      5        �    &      �      �  D        �t�bhhK ��h��R�(KK��h�Cp   &   -   �           L     |      �      2     %   R      �	     |      �   �      +         �t�bhhK ��h��R�(KK��h�CD      (   A   �   �        9   �
        $   
  �        �t�bhhK ��h��R�(KK��h�C4
   %   �  3  �
  I   �  }     �   �        �t�bhhK ��h��R�(KK��h�CT      5   $     �     �     8   E  &      M   �      8   �  �        �t�bhhK ��h��R�(KK��h�C`         �               )   M   �      t     �	        �                 �t�bhhK ��h��R�(KK��h�C       -   z   
           �t�bhhK ��h��R�(KK��h�CL   d        �        �     C              D   �           �t�bhhK ��h��R�(KK��h�C0�               
   *                 �t�bhhK ��h��R�(KK��h�C\            W           �           &      M         *      @           �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CL      �   �     4           1   #   
   3   6   �              �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C�     =     �t�bhhK ��h��R�(KK��h�CL�     >        ?         
   �
  F   
   ,                     �t�bhhK ��h��R�(KK��h�C �        	      	         �t�bhhK ��h��R�(KK��h�C@   [  [     X     2     "
  �     �               �t�bhhK ��h��R�(KK��h�Ch�     �     0   �     �  �       �        �   �     �   �      D   9   B   Z        �t�bhhK ��h��R�(KK��h�C,m  �  �     �     ,      X        �t�bhhK ��h��R�(KK��h�C              �t�bhhK ��h��R�(KK��h�C81   #      .     �  
   3   6   1     	        �t�bhhK ��h��R�(KK��h�CX      J   �        o                  �        �        �   �        �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK
��h�C(!            �  	      	         �t�bhhK ��h��R�(KK	��h�C$   �  �   �       �        �t�bhhK ��h��R�(KK��h�C@               ;     �  T   �   �   �      D         �t�bhhK ��h��R�(KK	��h�C$X      i         �           �t�bhhK ��h��R�(KK��h�CL      �     �           �   O      �    7   �  
   n        �t�bhhK ��h��R�(KK��h�C<
     �  c   g   �
     �  �      A  s   z        �t�bhhK ��h��R�(KK
��h�C(M     
   �      W     '         �t�bhhK ��h��R�(KK��h�C   (   o  �         �t�bhhK ��h��R�(KK��h�C8      [        .      G           W	        �t�bhhK ��h��R�(KK��h�C<�   $   �        �        �        $   E         �t�bhhK ��h��R�(KK��h�CP   %   �       2   -   ;  C   �      }           
     F         �t�bhhK ��h��R�(KK��h�C�     �  m      �t�bhhK ��h��R�(KK��h�C@   �     �  I     I   �  �  �          b        �t�bhhK ��h��R�(KK��h�C      �  H   �        �t�bhhK ��h��R�(KK��h�C41   #      J  
   3   6   �        K        �t�bhhK ��h��R�(KK��h�CL      �                          �     �                  �t�bhhK ��h��R�(KK��h�CpD         �      0     �   �      �   �   9   %  �      �   :  ,                  f   �        �t�bhhK ��h��R�(KK��h�C8h   t        ;      �     
   ,               �t�bhhK ��h��R�(KK��h�C@"   n        �                  P
                 �t�bhhK ��h��R�(KK��h�CD      =      :  :   W   e  ^   �   I           �        �t�bhhK ��h��R�(KK��h�C        �t�bhhK ��h��R�(KK��h�Cd   '   f   |        0   �     %   �     |      �   C     �   |  �	     $   |        �t�bhhK ��h��R�(KK��h�Ct               �         J  E      �  
        �  �  H   �        "     P      
           �t�bhhK ��h��R�(KK��h�CH�            )      �                    :               �t�bhhK ��h��R�(KK��h�CD      �  c         �              <   "              �t�bhhK ��h��R�(KK��h�C@   �        �     7  %  p      v     �   �        �t�bhhK ��h��R�(KK��h�C8d  
           `           �  %            �t�bhhK ��h��R�(KK��h�CP*      �   �            0   �        t  M
  *   )        b        �t�bhhK ��h��R�(KK��h�C<            9      �  L      0  f              �t�bhhK ��h��R�(KK��h�C"         2            �t�bhhK ��h��R�(KK��h�CLd   �     �   O      �   �              �      �     �        �t�bhhK ��h��R�(KK��h�C�      ;             �t�bhhK ��h��R�(KK��h�C   �  �        W
     �t�bhhK ��h��R�(KK��h�C1   #               �t�bhhK ��h��R�(KK
��h�C(      '   s            �         �t�bhhK ��h��R�(KK��h�C   �   �              �t�bhhK ��h��R�(KK��h�C�     n         �t�bhhK ��h��R�(KK��h�C4      '      �         
   I   [        �t�bhhK ��h��R�(KK��h�CH�     �  �      �     �        �    >      �   L         �t�bhhK ��h��R�(KK��h�C         ,   O      �t�bhhK ��h��R�(KK��h�CT      $        �     2   0      �     e  0     {     �  �        �t�bhhK ��h��R�(KK��h�C,   Q  R   �     .   	     b        �t�bhhK ��h��R�(KK ��h�C�            �     �        Q                                         ]     A  s   7               �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK
��h�C(   �  
   _                     �t�bhhK ��h��R�(KK��h�C<      �  �   G   +         b   #                  �t�bhhK ��h��R�(KK��h�C 8   �   �  *         �      �t�bhhK ��h��R�(KK��h�C0         /       �  $      �         �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C8      "     �   `  "   �        �   `        �t�bhhK ��h��R�(KK	��h�C$      �  �   �     O  �     �t�bhhK ��h��R�(KK��h�C        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�CX  �     �t�bhhK ��h��R�(KK��h�CX   l  g      t  �      :          �  �          �   �     �        �t�bhhK ��h��R�(KK��h�C   5         $   �     �t�bhhK ��h��R�(KK	��h�C$#     �   z      c  X  r      �t�bhhK ��h��R�(KK��h�C,   
   �     �t�bhhK ��h��R�(KK��h�CH)      �  �
        q  �  h  V   �  (  
      �  }         �t�bhhK ��h��R�(KK��h�C�          �t�bhhK ��h��R�(KK��h�Ch*        <   G      1           �      f                    �  V      5   <         �t�bhhK ��h��R�(KK	��h�C$      �   p  m     �        �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�C1     �  	         �t�bhhK ��h��R�(KK��h�C�  �           �t�bhhK ��h��R�(KK��h�C0g   O        z   
   �                �t�bhhK ��h��R�(KK��h�C�          �           �t�bhhK ��h��R�(KK��h�C8%   �  �        �   G
     7   ^     �        �t�bhhK ��h��R�(KK
��h�C(B  �      �    �
             �t�bhhK ��h��R�(KK��h�CZ      �               �t�bhhK ��h��R�(KK��h�C@!         �   �      %        	      	      	   �     �t�bhhK ��h��R�(KK��h�CT4                                           �   n              �t�bhhK ��h��R�(KK��h�C,T   �
        �     -   �           �t�bhhK ��h��R�(KK	��h�C$K     A       9   �        �t�bhhK ��h��R�(KK��h�C�  	         �t�bhhK ��h��R�(KK��h�C4               �     *  �      �        �t�bhhK ��h��R�(KK��h�C4�                              
         �t�b�      hhK ��h��R�(KK��h�Cd     �t�bhhK ��h��R�(KK��h�C      c  
            �t�bhhK ��h��R�(KK��h�C,      �        �  �  �  3        �t�bhhK ��h��R�(KK��h�C\     $               $         \  L   �            �      �              �t�bhhK ��h��R�(KK��h�C<�        �   �        �  s   �  y   5  ]        �t�bhhK ��h��R�(KK��h�C   �            �t�bhhK ��h��R�(KK��h�CX      �     �     4            �   B     �       H  �               �t�bhhK ��h��R�(KK	��h�C$#   !   '   
   @      F         �t�bhhK ��h��R�(KK��h�C�   S  �      �t�bhhK ��h��R�(KK"��h�C�      �         �     L  %   �                             �   �         @                  �   
   �        �t�bhhK ��h��R�(KK��h�C [      �  	      	         �t�bhhK ��h��R�(KK��h�CH      J    �        �  3         �      &   �         �t�bhhK ��h��R�(KK��h�C^     �t�bhhK ��h��R�(KK��h�C�  �      �           �t�bhhK ��h��R�(KK��h�C �        	      	         �t�bhhK ��h��R�(KK��h�C                      �t�bhhK ��h��R�(KK��h�C\!  &   �   7  )        �   3     ,   O      C  �        Y  �      7         �t�bhhK ��h��R�(KK��h�Cp                     �   ]  �         7      
     &      -   F  +      t   
   $   �        �t�bhhK ��h��R�(KK��h�C`*      &   \       M      +   $   �  E      �	        
   5  �   �             �t�bhhK ��h��R�(KK��h�C    	      	      	   K      �t�bhhK ��h��R�(KK��h�C4      a   ;      0   [   :   8   �   E        �t�bhhK ��h��R�(KK��h�C`   ?   #   !         �   �         
   �   F      
   3   6     �   �               �t�bhhK ��h��R�(KK��h�CX2   (   �     �   +  �  i      �  +     �        �   n      �   �        �t�bhhK ��h��R�(KK��h�C   �	     	  �     �t�bhhK ��h��R�(KK��h�C/      8     �     �t�bhhK ��h��R�(KK��h�CD#   !         i     �   n   (      
   P     G            �t�bhhK ��h��R�(KK��h�C8         �t�bhhK ��h��R�(KK��h�C	  N        �     �t�bhhK ��h��R�(KK��h�C82      )  C      w  e  =           �        �t�bhhK ��h��R�(KK��h�C k    
   H   B   }         �t�bhhK ��h��R�(KK��h�C0�     3     d   �      �  
   J        �t�bhhK ��h��R�(KK��h�C@�      �  %         )   �  B   �  "     �   �         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�CT               k            -                x  V      G        �t�bhhK ��h��R�(KK��h�C4   R         .   D     �      r  �        �t�bhhK ��h��R�(KK��h�Cl      �  #      n     d   t           l     D   
   3   6       *      /   �              �t�bhhK ��h��R�(KK��h�C (            �   �        �t�bhhK ��h��R�(KK��h�CH�           �     p  '      �         �
        @         �t�bhhK ��h��R�(KK
��h�C(  �     �  �      �     �     �t�bhhK ��h��R�(KK��h�C\         ~   �            �   j   n      M   T   �      8   �  �              �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�CD�   )   �      �      |      �         $  �     �        �t�bhhK ��h��R�(KK��h�C    �     	      	         �t�bhhK ��h��R�(KK��h�C<      �           �t�bhhK ��h��R�(KK��h�Ch            V   �  �  P     �  �     �  �        T   �	  (   7     �   '            �t�bhhK ��h��R�(KK��h�C                     �t�bhhK ��h��R�(KK��h�C h        	      	         �t�bhhK ��h��R�(KK��h�C,1   #       A     �  Y  �            �t�bhhK ��h��R�(KK��h�CT   q        �                 �               �     �  �        �t�bhhK ��h��R�(KK��h�C`   �  �
        �t�bhhK ��h��R�(KK��h�CP�   s  (      :   Q     z  
     j  �     �  A  �   k  �
        �t�bhhK ��h��R�(KK��h�C�  	      	         �t�bhhK ��h��R�(KK��h�C,�	     j      
  �  	      	         �t�bhhK ��h��R�(KK��h�C@"            �   s  �      z   
   �                 �t�bhhK ��h��R�(KK��h�C4   ?   *        
   �        
           �t�bhhK ��h��R�(KK��h�C w  �  +   �              �t�bhhK ��h��R�(KK��h�C|�  !      \   2   �  C      A  �   3                                                   Z            �t�bhhK ��h��R�(KK��h�C@0     ;      0         V        #  U             �t�bhhK ��h��R�(KK
��h�C(      �     :                  �t�bhhK ��h��R�(KK��h�CT   p  �  �          .         q                               �t�bhhK ��h��R�(KK	��h�C$   �   �   �     �            �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C�        .          �t�bhhK ��h��R�(KK��h�CT*         
                       =      �   "   $         W         �t�bhhK ��h��R�(KK��h�CD/   _  C   !  }        )               �     �        �t�bhhK ��h��R�(KK��h�CL
   t   C  2   )            "     F     k            +         �t�bhhK ��h��R�(KK��h�Cp      M  	         �t�bhhK ��h��R�(KK��h�C      e      �t�bhhK ��h��R�(KK��h�C   �  �        �t�bhhK ��h��R�(KK��h�C  "  >   �   a   r      �t�bhhK ��h��R�(KK
��h�C(   W        ~  y     e         �t�bhhK ��h��R�(KK��h�C,9   �  L   x        X     �        �t�bhhK ��h��R�(KK��h�CP   D         S   X  i   ,            <  �  �      d   �   X        �t�bhhK ��h��R�(KK��h�C      �               �t�bhhK ��h��R�(KK��h�Cd        �t�bhhK ��h��R�(KK��h�CL
   3   6   �        �   ?      !      �     z   ,               �t�bhhK ��h��R�(KK��h�C   �      �t�bhhK ��h��R�(KK��h�C           �   r      �t�bhhK ��h��R�(KK��h�CT     �
        �  �       �     2   �  �  j      �     o         �t�bhhK ��h��R�(KK
��h�C(   <     a           �        �t�bhhK ��h��R�(KK��h�CP   D         k                  =      >     [      �   �         �t�bhhK ��h��R�(KK	��h�C$�  -      n      a  g         �t�bhhK ��h��R�(KK��h�C8      �   -   �  h  V      �     �  �        �t�bhhK ��h��R�(KK��h�C81   #   
   3   6   �           2              �t�bhhK ��h��R�(KK��h�C@      �    
   �  &      �   M   �      $            �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C<   �	     Z  �  )        e      X              �t�bhhK ��h��R�(KK	��h�C$�  /     .      �   w         �t�bhhK ��h��R�(KK��h�C ]      �     �   �        �t�bhhK ��h��R�(KK��h�C4�        �       �      �
     �        �t�bhhK ��h��R�(KK��h�C*     p     �      �t�bhhK ��h��R�(KK��h�CP            �     (         .     +        L
        �        �t�bhhK ��h��R�(KK��h�CL   5      k         D  �   �  R      �       �     5        �t�bhhK ��h��R�(KK
��h�C(        n  �   ;      �         �t�bhhK ��h��R�(KK��h�CL   �      $     �     
  :   �   3  �         �	     �         �t�bhhK ��h��R�(KK��h�C0      a  Z  h   %   �     �  z        �t�bhhK ��h��R�(KK��h�C !        	      	         �t�bhhK ��h��R�(KK��h�C`   D         :   �      .   
   _      \  &      �  �      ]   
   �  ^   \        �t�bhhK ��h��R�(KK��h�C             �t�bhhK ��h��R�(KK��h�C0/      �        .                     �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK	��h�C$[        �  	      	         �t�bhhK ��h��R�(KK��h�C�	     	      	         �t�bhhK ��h��R�(KK��h�C $   |       �   �        �t�bhhK ��h��R�(KK��h�Ct
   w        �  c      �     B  
      Y     S      �  �        E  �           �           �t�bhhK ��h��R�(KK
��h�C(�   �   �        �   �             �t�bhhK ��h��R�(KK��h�C        �         �t�bhhK ��h��R�(KK��h�C4W   �   #   !      �
  [           	        �t�bhhK ��h��R�(KK	��h�C$      L  �                 �t�bhhK ��h��R�(KK	��h�C$   (   �  3  :   �   �        �t�bhhK ��h��R�(KK��h�C@*      �   F  &      U        i     
   $   �        �t�bhhK ��h��R�(KK��h�CH   R   �   �      "   �   �        �           d   I
        �t�bhhK ��h��R�(KK��h�C      
  �  �     �t�bhhK ��h��R�(KK��h�C@!         �   �            Y        	      	         �t�bhhK ��h��R�(KK
��h�C(         �  �          �     �t�bhhK ��h��R�(KK��h�CT      �  $        &         $        �        .   �     2        �t�bhhK ��h��R�(KK	��h�C$"   �  (      !               �t�bhhK ��h��R�(KK��h�CP�  �     p  -   7     H               .   �          �        �t�bhhK ��h��R�(KK��h�C1     t      @          �t�bhhK ��h��R�(KK��h�C0   \              �        F        �t�bhhK ��h��R�(KK��h�CD"   �          �   =     %   !             5
        �t�bhhK ��h��R�(KK��h�C8#   !         ?      
   X   �   F      �        �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C,   �   w      �      -   U   C        �t�bhhK ��h��R�(KK��h�CH   5      �      \  |      �                  �   ]         �t�bhhK ��h��R�(KK��h�C4#   !         P     ?      
   T  �        �t�bhhK ��h��R�(KK��h�C0�  "  J     8     �     A   [        �t�bhhK ��h��R�(KK��h�C�   n     �t�bhhK ��h��R�(KK��h�C0
   e   �   F   '   �           K        �t�bhhK ��h��R�(KK��h�CT
   2           .   0        �  $   �     b      �     -  �        �t�bhhK ��h��R�(KK��h�C2     �
  	         �t�bhhK ��h��R�(KK��h�C\   5      *      �      0              m           G   W      �           �t�bhhK ��h��R�(KK��h�CP   P  X
     {     �     �   :     �         R                 �t�bhhK ��h��R�(KK
��h�C(   =      H  �  	      	         �t�bhhK ��h��R�(KK��h�C   }     o         �t�bhhK ��h��R�(KK��h�C8�                   �                    �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C,�      �  
            j   v        �t�bhhK ��h��R�(KK��h�C0   �     X     )     �   B   }         �t�bhhK ��h��R�(KK��h�C8         2   
      _                       �t�bhhK ��h��R�(KK��h�C,�  (                  $   �        �t�bhhK ��h��R�(KK��h�C^    �        �t�bhhK ��h��R�(KK��h�C\      U   k     8   /      m         �      m      �         J   a   <         �t�bhhK ��h��R�(KK��h�C<b   G   W            ;      �     �   S   U        �t�bhhK ��h��R�(KK��h�Cdg   b     e  �     �  M   c      /  k
        M   �      D   �  D   �  �   7         �t�bhhK ��h��R�(KK��h�C�              �t�bhhK ��h��R�(KK��h�C,b   $   �   #    
   $   �  �        �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   6   Y      O         �t�bhhK ��h��R�(KK��h�CH9   �  ;  �      %   p     ?        +      �   8   E        �t�bhhK ��h��R�(KK��h�CX   �      /      [  o        �  &   �   �      L   G   |     <           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C      	         �t�bhhK ��h��R�(KK��h�C,   �     %           
   3        �t�bhhK ��h��R�(KK��h�CT�   v        w     8   4      �              r     a      4         �t�bhhK ��h��R�(KK��h�CL      �            
   c        �               "   �        �t�bhhK ��h��R�(KK��h�C R  �
     	      	         �t�bhhK ��h��R�(KK��h�C4!      1     �  ?      
   3   6   	        �t�bhhK ��h��R�(KK��h�C�
     �t�bhhK ��h��R�(KK��h�CL#   !      �     4      U    :      S   t      �     |        �t�bhhK ��h��R�(KK	��h�C$   5      =   �              �t�bhhK ��h��R�(KK��h�C8      P   �  G      �  h         $   k         �t�bhhK ��h��R�(KK��h�C0"   �  (      <      [         w        �t�bhhK ��h��R�(KK��h�C*      /   \     �t�bhhK ��h��R�(KK��h�C0<      �             �  �  	         �t�bhhK ��h��R�(KK��h�C         \  9   �        �t�bhhK ��h��R�(KK��h�C8      M   �        *         �    7         �t�bhhK ��h��R�(KK��h�C u     �  
   f   �         �t�bhhK ��h��R�(KK��h�C[   �     �        �t�bhhK ��h��R�(KK��h�CD3     T        S   <     �     �      �             �t�bhhK ��h��R�(KK	��h�C$
   3   6   )  ?   �   �   r      �t�bhhK ��h��R�(KK��h�C0
   �  F   '   �   !      �              �t�bhhK ��h��R�(KK��h�C      ;     u         �t�bhhK ��h��R�(KK��h�C�	     j      
        �t�bhhK ��h��R�(KK��h�C0      �   0   <   "   �     +  �  r      �t�bhhK ��h��R�(KK��h�CH           
   )  9           
   �  �     q          �t�bhhK ��h��R�(KK��h�C        �            �t�bhhK ��h��R�(KK��h�C   �  B   �          �t�bhhK ��h��R�(KK��h�CP
   3   6   )  ?   �   �   r   (      !      \        {               �t�bhhK ��h��R�(KK��h�Cm      �     �t�bhhK ��h��R�(KK��h�C\1   #   
   3   6      [      9     �     �     V     V  
   T  Z          �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C0�  j  /           b         �        �t�bhhK ��h��R�(KK��h�C,I      (   -  �     �              �t�bhhK ��h��R�(KK��h�C B  �        
            �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK
��h�C(B   �   �      �  /      ^        �t�bhhK ��h��R�(KK��h�C`�  h  �   	     ^   �     s  *      5         �      -             �         �t�bhhK ��h��R�(KK��h�CP      ;                           %     �     j     �        �t�bhhK ��h��R�(KK	��h�C$   �        �      �        �t�bhhK ��h��R�(KK��h�C8M   �   �         �	  V      J   �      �        �t�bhhK ��h��R�(KK��h�C0w     ;     u          "   5        �t�bhhK ��h��R�(KK��h�C<   �        �     (      !            W        �t�bhhK ��h��R�(KK��h�C�  	      	         �t�bhhK ��h��R�(KK��h�C,!      
     	      	      	   K      �t�bhhK ��h��R�(KK��h�C`      D  �         5      �   e     4      m     �   �   
     4               �t�bhhK ��h��R�(KK��h�Ck     �        �t�bhhK ��h��R�(KK��h�CD�   �     �  �	     �   
              �   "   �        �t�bhhK ��h��R�(KK��h�C �         	      	         �t�bhhK ��h��R�(KK��h�CH   �   '      ~       O  s      �              �	        �t�bhhK ��h��R�(KK��h�C4�  ,         p  )   A   {
  }               �t�bhhK ��h��R�(KK+��h�C�      �   :      Q               Y      Q         Q     Q      x              z   5      �   a         Z     8   E        0   4               �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C -        �     �        �t�bhhK ��h��R�(KK��h�CTX   �   �   )                       9     �  /      r     V        �t�bhhK ��h��R�(KK��h�C8I   l                       0      �        �t�bhhK ��h��R�(KK��h�C   9     �t�bhhK ��h��R�(KK��h�C,   %   �        X  ,               �t�bhhK ��h��R�(KK��h�CP)   O      Y      ?       ?     C        ;      �      z         �t�bhhK ��h��R�(KK��h�C,]   v     $   �       �           �t�bhhK ��h��R�(KK��h�C,   >   �     �      J   &	  +         �t�bhhK ��h��R�(KK
��h�C(   S   >  5         �  �         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C|      �   �      �t�bhhK ��h��R�(KK��h�C,O
        A  G   |     $   k         �t�bhhK ��h��R�(KK��h�C�            �t�bhhK ��h��R�(KK��h�C    X   '   -   �   �        �t�bhhK ��h��R�(KK��h�C_  
         �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C  n  
   4  	         �t�bhhK ��h��R�(KK��h�CX$        8   }      $   d     �  �	     �  �      8   �  -               �t�bhhK ��h��R�(KK��h�C �        	      	         �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6            �t�bhhK ��h��R�(KK��h�C(  	  	         �t�bhhK ��h��R�(KK��h�CD      �     2   	  s   �	  	     �     �
              �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK	��h�C$   �	  ,                     �t�bhhK ��h��R�(KK��h�C�   	  	         �t�bhhK ��h��R�(KK��h�CP      -   =      H   �  4      Y      n  
        �   �           �t�bhhK ��h��R�(KK��h�C[      :     =  �	     �t�bhhK ��h��R�(KK��h�C�     	      	         �t�bhhK ��h��R�(KK��h�C4�  �   {     �  7      W  
      �         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C 1        	      	         �t�bhhK ��h��R�(KK��h�C0�     �     �  �        �   [	        �t�bhhK ��h��R�(KK��h�C`      M   c   k
              +      �      �  9   �   �  �   9      �  y        �t�bhhK ��h��R�(KK��h�C4V   (      )            �     A            �t�bhhK ��h��R�(KK��h�CP      J   4  c   �  �   >      �                       ;        �t�bhhK ��h��R�(KK��h�C,   �  ?      !      �     @         �t�bhhK ��h��R�(KK��h�CI   `   �           �t�bhhK ��h��R�(KK��h�C0         3              j            �t�bhhK ��h��R�(KK��h�CE      4      �t�bhhK ��h��R�(KK��h�C�     v     �t�bhhK ��h��R�(KK��h�C�     �    ,         �t�bhhK ��h��R�(KK��h�C0   _  +   �   �           �            �t�bhhK ��h��R�(KK	��h�C$         0                  �t�bhhK ��h��R�(KK��h�CL1   #      .     	           =   �   
   3   6   1     	        �t�bhhK ��h��R�(KK��h�C<      -   N            i  �                    �t�bhhK ��h��R�(KK��h�C 1   #       �     _        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�Cz  �                 �t�bhhK ��h��R�(KK��h�C4�  �     `     /      N   �     s        �t�bhhK ��h��R�(KK	��h�C$Z      �                     �t�bhhK ��h��R�(KK��h�C  �      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK	��h�C$�                     r      �t�bhhK ��h��R�(KK��h�CP�     �     9   �  L         o     �     �  N      �            �t�bhhK ��h��R�(KK��h�C       -   \  �   c	        �t�bhhK ��h��R�(KK��h�Cl         E  �      �   S   Q         d  �      b     �         D  �      z               �t�bhhK ��h��R�(KK��h�Cd        �   O         �t�bhhK ��h��R�(KK��h�C0      
   �     %   9  �  y  y         �t�bhhK ��h��R�(KK��h�C@   .     M                @   (      �     �     �t�bhhK ��h��R�(KK��h�CX         �     7   y      �  f           0   
     �  i      _        �t�bhhK ��h��R�(KK%��h�C�         �     7      X      $   k         �  �   X   �   `     �
        �     �                                       �t�bhhK ��h��R�(KK
��h�C(         �     )  ^            �t�bhhK ��h��R�(KK��h�CDu   (   <      �  "   �   �           |      �            �t�bhhK ��h��R�(KK��h�C8   &   G  ~        Q   V      �      L        �t�bhhK ��h��R�(KK��h�C     �            �t�bhhK ��h��R�(KK��h�C8�                       0  �      �         �t�bhhK ��h��R�(KK��h�C~     �t�bhhK ��h��R�(KK��h�CL         <        n   &      U   �      %   o      h  u         �t�bhhK ��h��R�(KK
��h�C(�	     �  �   �        �  O      �t�bhhK ��h��R�(KK��h�C      u      �t�bhhK ��h��R�(KK��h�C<      L  �   t	  �           .                  �t�bhhK ��h��R�(KK��h�C!            �t�bhhK ��h��R�(KK��h�C�   L  �   �        �t�bhhK ��h��R�(KK��h�CL   (      @
  �      �   �         �  8   <     $   !          �t�bhhK ��h��R�(KK��h�C01   #   
             �     �         �t�bhhK ��h��R�(KK��h�Cl   2   J     :  �     �   �  B     >   2   �   �  C   �   7      A  :   �   �     �         �t�bhhK ��h��R�(KK��h�C�             �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C0T   (               �     :   k        �t�bhhK ��h��R�(KK��h�C<      )  +   e  ^         �  G   |      �         �t�bhhK ��h��R�(KK��h�C0      )   6     X   �     6  �        �t�bhhK ��h��R�(KK��h�C 4         	      	         �t�bhhK ��h��R�(KK��h�CP   �     �       .   !
     A     n                �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C<  �   5      r      �        �     ,   	         �t�bhhK ��h��R�(KK��h�C0            w     :   �             �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CH   ?   �   !         �     o         
   �   �     �        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C8   �      (         "   A   g  �     �	        �t�bhhK ��h��R�(KK��h�CT      �  �  =     $   E      �   ]      �  ^   8   �        t        �t�bhhK ��h��R�(KK��h�CP   X   '   H   �  j     �     A   j  ^        -      �  �        �t�bhhK ��h��R�(KK��h�Cx*   x  {     0  ;      0         %   _     �      �         
  �           "   �     '           �t�bhhK ��h��R�(KK��h�C<   �        �   W                 _  �        �t�bhhK ��h��R�(KK��h�C �          �              �t�bhhK ��h��R�(KK��h�C@
   u  F   '      �  �   %   �        %   R  �        �t�bhhK ��h��R�(KK��h�C,      5      &     7  H          �t�bhhK ��h��R�(KK��h�C8   �         �  �     Q
     �   �   a        �t�bhhK ��h��R�(KK��h�C0�  �  �  �      .     �	     �        �t�bhhK ��h��R�(KK��h�C1   #       �      D      �t�bhhK ��h��R�(KK��h�C\   u  �   
   m  
           �     
   �   �        .                     �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C<   c        p               �     $   �         �t�bhhK ��h��R�(KK��h�Cv  �     �     �t�bhhK ��h��R�(KK��h�C8`     �     �  5     �  %   �
  C            �t�bhhK ��h��R�(KK��h�C0W   �   �   
   �   )   
   K      �         �t�bhhK ��h��R�(KK��h�C=     �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C8r     N   �        '      �  �     ]         �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C�   (   �   <   r      �t�bhhK ��h��R�(KK��h�C8   /         	  �     -      �  8           �t�bhhK ��h��R�(KK��h�CX   8   /      k      l              �      �   ;      ,  %   �           �t�bhhK ��h��R�(KK(��h�C�   .   
                 (   /  
   _      8   u  �        2   "         (        &      ,   �                    J	     �         �t�bhhK ��h��R�(KK
��h�C(R	     )   �  ]     j            �t�bhhK ��h��R�(KK��h�CX      2   f  �   b  �      �     �  Z  '           M   �      D         �t�bhhK ��h��R�(KK
��h�C(!      [         	      	         �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   6   Y      O         �t�bhhK ��h��R�(KK��h�C{
        �t�bhhK ��h��R�(KK��h�C4b   #                  &  �   G            �t�bhhK ��h��R�(KK	��h�C$           	      	        �t�bhhK ��h��R�(KK��h�C@.     �     u      @      �  N  7         4         �t�bhhK ��h��R�(KK��h�C0   .                  H      �        �t�bhhK ��h��R�(KK��h�C4      5         �     M   �              �t�bhhK ��h��R�(KK��h�C�     	      	         �t�bhhK ��h��R�(KK��h�C{     �      �t�bhhK ��h��R�(KK��h�CT      �     �   �     2      (   �        �     /   9     7         �t�bhhK ��h��R�(KK��h�C<�         �   Y  k                         �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�CD   e   '   `     �               A   s     B   �        �t�bhhK ��h��R�(KK��h�C�  �        	         �t�bhhK ��h��R�(KK��h�C,
      �  2   �  
      B           �t�bhhK ��h��R�(KK ��h�C�      5   !      w     L	     �           \   �
        �         3  W  &      �   F    �  9            �t�bhhK ��h��R�(KK��h�C4g  
   c             E  
   ,            �t�bhhK ��h��R�(KK	��h�C$4     )  �      9   �        �t�bhhK ��h��R�(KK	��h�C$   =      )  	      	         �t�bhhK ��h��R�(KK
��h�C(=  �     )   �  ^  `   :        �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�C�  !      9  	         �t�bhhK ��h��R�(KK��h�C      �  �           �t�bhhK ��h��R�(KK��h�C   
         �t�bhhK ��h��R�(KK��h�CX   �   5   <         �        �     -  �     �   =                     �t�bhhK ��h��R�(KK��h�C8p   =  �  `   �                 �  �         �t�bhhK ��h��R�(KK��h�C   �     X          �t�bhhK ��h��R�(KK��h�C4   (   w   s    N  8   /   &   O           �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C`                 �     s     U         <      !  �                       �t�bhhK ��h��R�(KK��h�C@            z   
   ,            �  )   
            �t�bhhK ��h��R�(KK��h�C<         ;      �        =         "   W         �t�bhhK ��h��R�(KK��h�CL         �          �            0   <      x   "           �t�bhhK ��h��R�(KK��h�C4�      �  �  �   V     �                 �t�bhhK ��h��R�(KK��h�C@      -   0              
   f     �   ,            �t�bhhK ��h��R�(KK��h�C0>     �          u     �  O         �t�bhhK ��h��R�(KK��h�C�   "   G	     M     �t�bhhK ��h��R�(KK��h�Cd      0      4      �      &      D  *     $     |  �   +   �     #              �t�bhhK ��h��R�(KK��h�C0   5   �     .      $   �      �        �t�bhhK ��h��R�(KK��h�C\     �      ;     p     ^        $          J   �  �   �     ,         �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�C      T  	      	         �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK
��h�C(�	     �        	      	         �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C4�   �   (      /  
   ,                     �t�bhhK ��h��R�(KK��h�C<�  �              &   �   �                     �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�CX      N   �     �     n   S     
   *     e  i   �  �     e          �t�bhhK ��h��R�(KK��h�C,�      �  �   �   �     %   J         �t�bhhK ��h��R�(KK��h�C<�  h    "   �     i        �	                 �t�bhhK ��h��R�(KK��h�CZ             �t�bhhK ��h��R�(KK��h�C1   #   �          �t�bhhK ��h��R�(KK��h�C4      =      B  
        �   �           �t�bhhK ��h��R�(KK��h�C@      J   }     �   o            0   <   "            �t�bhhK ��h��R�(KK��h�C<   '   -              *	           �            �t�bhhK ��h��R�(KK��h�C01   #   
   3   6      �   4  o  4   r      �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C   �   �              �t�bhhK ��h��R�(KK
��h�C(�      �   �  �            �     �t�bhhK ��h��R�(KK
��h�C(      N   �     �   �   �        �t�bhhK ��h��R�(KK
��h�C(�  �      E      G     t         �t�bhhK ��h��R�(KK��h�CK        1        �t�bhhK ��h��R�(KK
��h�C(d   �           l        /      �t�bhhK ��h��R�(KK
��h�C(      A     �  Y     	         �t�bhhK ��h��R�(KK��h�C8   �   
   ,            K      �      �         �t�bhhK ��h��R�(KK��h�C<|      �      |      s	     �   +      P   {         �t�bhhK ��h��R�(KK	��h�C$      '   -      �   M        �t�bhhK ��h��R�(KK��h�C~     �t�bhhK ��h��R�(KK��h�C4*      @  t      M      +   �   �   �         �t�bhhK ��h��R�(KK	��h�C$-      �      N      �        �t�bhhK ��h��R�(KK��h�C    ?   �  
   �
  F         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CH2      =                 ,   D     W   T   4      �        �t�bhhK ��h��R�(KK��h�C!                    �t�bhhK ��h��R�(KK��h�C0         �   7  l   9     7   /         �t�bhhK ��h��R�(KK��h�C4   (   �  �   �   *         
     4         �t�bhhK ��h��R�(KK��h�C8@      �                 9   �     4        �t�bhhK ��h��R�(KK��h�CX�    
   %   b     K     �     �  *   I   �     )            	        �t�bhhK ��h��R�(KK��h�CD   �  �      {           2   �           �          �t�bhhK ��h��R�(KK��h�C8.     	    �           V                 �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CP
      �  (      !           �   �        �     %   �            �t�bhhK ��h��R�(KK��h�C      U     �        �t�bhhK ��h��R�(KK��h�C4�      I              �     ^           �t�bhhK ��h��R�(KK��h�C0   �  C   -      M      �
     U        �t�bhhK ��h��R�(KK��h�C               �      �t�bhhK ��h��R�(KK��h�Ck     Q        �t�bhhK ��h��R�(KK��h�C<�  �     �     �  �      �     {     J        �t�bhhK ��h��R�(KK��h�CD   �  �   �           �      �         G              �t�bhhK ��h��R�(KK��h�CH�           a	     �  -      
  V     a                 �t�bhhK ��h��R�(KK��h�C4�     j              b         �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CP*              #
           L     P           %     X        �t�bhhK ��h��R�(KK��h�C0G  8     r  �      %  .	     �        �t�bhhK ��h��R�(KK��h�C      	         �t�bhhK ��h��R�(KK��h�C   �        ^        �t�bhhK ��h��R�(KK��h�C<     �t�bhhK ��h��R�(KK��h�C,            �t�bhhK ��h��R�(KK
��h�C(1   #      �  
   3   6            �t�bhhK ��h��R�(KK	��h�C$   ?   �  ^   $   \  F         �t�bhhK ��h��R�(KK��h�C,      �     
   y                 �t�bhhK ��h��R�(KK"��h�C�%   �   h     �  �         �  �      �  �        �  �      �  $  G   B   [        �   y    �      �  �        �t�bhhK ��h��R�(KK��h�CP         k               �   L            �  
   $   �   N        �t�bhhK ��h��R�(KK��h�C%                 �t�bhhK ��h��R�(KK��h�C`"   W       X    p      Y  �  h   �     �          Z     [     \        �t�bhhK ��h��R�(KK	��h�C$i     a     .   
   w        �t�bhhK ��h��R�(KK��h�C,      0      �      A     7         �t�bhhK ��h��R�(KK��h�C�   =     �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C0�  �        �  ^     �   A   �         �t�bhhK ��h��R�(KK��h�C;     �t�bhhK ��h��R�(KK��h�C<�      �   d  
   %     [      �     �	  +         �t�bhhK ��h��R�(KK��h�C4      ?      �           �  �   �        �t�bhhK ��h��R�(KK��h�CH      O      Y      x     �           �  $   �           �t�bhhK ��h��R�(KK	��h�C$�              �  M        �t�bhhK ��h��R�(KK��h�C)   �     �  i        �t�bhhK ��h��R�(KK��h�C    �                    �t�bhhK ��h��R�(KK��h�CX      �   L     �         x     K     L        !  �                 �t�bhhK ��h��R�(KK��h�C<            �t�bhhK ��h��R�(KK��h�C<      5           y        \  j  q   �        �t�bhhK ��h��R�(KK��h�C`�   7  (   F     d  �      .   
   _      L  �     d     �   *   %   d  �        �t�bhhK ��h��R�(KK��h�C,2   �         �   
         �        �t�bhhK ��h��R�(KK��h�C4I      ~      G        >   5  q           �t�bhhK ��h��R�(KK��h�CH           &  *      �        �       �   �  w         �t�bhhK ��h��R�(KK��h�C"   K     �
  �        �t�bhhK ��h��R�(KK��h�C0   �       C     '                  �t�bhhK ��h��R�(KK	��h�C$$  �   
   4  	      	         �t�bhhK ��h��R�(KK��h�CX                              �  `   �              0   h  �        �t�bhhK ��h��R�(KK	��h�C$�        l   �              �t�bhhK ��h��R�(KK ��h�C��        	        q        �                       �        �   q     @      e      X              �t�bhhK ��h��R�(KK	��h�C$1   #          }     o         �t�bhhK ��h��R�(KK��h�CD   :  �     "   �      (  j   "      �     �   �	        �t�bhhK ��h��R�(KK��h�C,      %   �      �
    �            �t�bhhK ��h��R�(KK��h�C0   Y  '   -   H      :      .            �t�bhhK ��h��R�(KK��h�C   /            �t�bhhK ��h��R�(KK��h�C4�          t  
           �   �        �t�bhhK ��h��R�(KK��h�C4   ?      �  �   >     ,   
   �	  F         �t�bhhK ��h��R�(KK��h�C8V        �  �     
     Q      j           �t�bhhK ��h��R�(KK
��h�C(1   #       �     �	              �t�bhhK ��h��R�(KK��h�C,p   
   A   F     �  R     Y        �t�bhhK ��h��R�(KK��h�CL        @
  �      �            �  8   <     $   !          �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�C0           (     %     �   q         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�Ch  �     �     �t�bhhK ��h��R�(KK
��h�C(      �  �     ,   I  	         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C8      N           d              �        �t�bhhK ��h��R�(KK��h�CZ   .     �t�bhhK ��h��R�(KK��h�Cv     :     �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�CX           /   �      $   8     T      �  
     �   9   s   �  L         �t�bhhK ��h��R�(KK��h�C,�   �  �  P  �  �        �         �t�bhhK ��h��R�(KK��h�C8
               m  �         ?      !         �t�bhhK ��h��R�(KK��h�C,   >   -   w                        �t�bhhK ��h��R�(KK��h�C4v         �  )         �  �     �        �t�bhhK ��h��R�(KK��h�CHd   �     y   D         D   �  	  �            C          �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CD      )        <            D  %  �     &   U         �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�CP   �  l   �   �  -              �  <            ^     V        �t�bhhK ��h��R�(KK��h�C B        Z     7         �t�bhhK ��h��R�(KK��h�C 7       0  `     �     �t�bhhK ��h��R�(KK��h�CT         Y     �  �   7      �           0   
     A  ,  _        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C,[           l   9                 �t�bhhK ��h��R�(KK ��h�C�   q        �  �     �                >      �      g  :   �     �   �   Q      A     �     t         �t�bhhK ��h��R�(KK	��h�C$   K        /   9     7      �t�bhhK ��h��R�(KK��h�Ct      �
          Y  �      �  L   y                 %      )   a   ;      �  :      u        �t�bhhK ��h��R�(KK��h�C8   4  '   �                  C      �        �t�bhhK ��h��R�(KK��h�C8      0   �      .   "                        �t�bhhK ��h��R�(KK��h�C<*                     \        �   S            �t�bhhK ��h��R�(KK��h�CL   �     y  �   >   2         �	              t      n        �t�bhhK ��h��R�(KK��h�CP�  �   �  z  *   %   5   $  �      ,   [        .   =      �  �     �t�bhhK ��h��R�(KK��h�C\      &   G        #   i   �  _        Y      O      >      F  $   �        �t�bhhK ��h��R�(KK1��h�Cč   �     8           (   �    
   _      }     L        �     �     }      d     �     �     h           �  q        �   �   �     $  P     �  �         �t�bhhK ��h��R�(KK��h�C,%        g   O     9             �t�bhhK ��h��R�(KK��h�C4E      �  =  ^   �   F            �        �t�bhhK ��h��R�(KK��h�Cd      �     -                   G  �  �   �     &      $   �  g   $            �t�bhhK ��h��R�(KK��h�C|   H  �        �                        %   �         �  C        |	           C     �        �t�bhhK ��h��R�(KK��h�C<   �   *         "  �        �   �  y   '        �t�bhhK ��h��R�(KK��h�C =     K  	      	         �t�bhhK ��h��R�(KK
��h�C(�  p     ^     z   "   �        �t�bhhK ��h��R�(KK��h�C`                        �   �        i       s     t  
   w  j   �        �t�bhhK ��h��R�(KK��h�CH   �      ;  C         N        �     N     �  8  �      �t�bhhK ��h��R�(KK��h�C,�      ,         I  	      	         �t�bhhK ��h��R�(KK��h�C\	     �t�bhhK ��h��R�(KK��h�C    �          {        �t�bhhK ��h��R�(KK��h�CH            
   /      �                        7        �t�bhhK ��h��R�(KK��h�CP      �     @        �           �      �  ~   �               �t�bhhK ��h��R�(KK��h�C�  
      �	     �t�bhhK ��h��R�(KK	��h�C$_          �  !           �t�bhhK ��h��R�(KK��h�C4           �   �            0   �  r      �t�bhhK ��h��R�(KK��h�Cl:      (      )   �   
   �      ^   �     s  *      5   x      ~     /           �         �t�bhhK ��h��R�(KK��h�C`G   C     "   $
  (   /      �      �  <      m      -  ~     /      �           �t�bhhK ��h��R�(KK��h�C@*   2           �     �
        �  
   k  n        �t�bhhK ��h��R�(KK��h�Cm      �     �t�bhhK ��h��R�(KK��h�Ct     �t�bhhK ��h��R�(KK��h�CT   �      �   q       C         �   w     �                        �t�bhhK ��h��R�(KK��h�CL   ?   !      �      ,      .   G   �                        �t�bhhK ��h��R�(KK��h�C�   |      �     �t�bhhK ��h��R�(KK��h�C1   #          �t�bhhK ��h��R�(KK��h�CL   /   9   �   7      N      �  �  
   �  9   �     �  k
        �t�bhhK ��h��R�(KK��h�C<      U   6  )   *      t     �  +      �         �t�bhhK ��h��R�(KK��h�C@      ~               a   ;      0                 �t�bhhK ��h��R�(KK��h�C4
        �       �     �               �t�bhhK ��h��R�(KK��h�C,V   ?   2   �  
   �   9  B   }         �t�bhhK ��h��R�(KK	��h�C$+  4      �     R            �t�bhhK ��h��R�(KK��h�C�          �t�bhhK ��h��R�(KK��h�CD!         =      H  ?      
   3   6   �        �        �t�bhhK ��h��R�(KK
��h�C(   �   '   �  5     �   5        �t�bhhK ��h��R�(KK��h�CD         &   D  0   4   >      a   �  �     8   �        �t�bhhK ��h��R�(KK��h�C`G      �            6       0      n      �   �     N   �  i      �   =        �t�bhhK ��h��R�(KK��h�C-   H   o   �   �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�CL            �   ]   �   O         
   �  _   0   4               �t�bhhK ��h��R�(KK��h�C\�   �  !     �  !           �     �   �             �   �     �         �t�bhhK ��h��R�(KK��h�CX   5      �         �         �            J            �  �   �        �t�bhhK ��h��R�(KK	��h�C$�           	      	         �t�bhhK ��h��R�(KK��h�C8V           \  (  
   B        B           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CD         <     )	     b      x   "   �     $   k         �t�bhhK ��h��R�(KK
��h�C(         P   H     +   w         �t�bhhK ��h��R�(KK��h�CD      �   �  �     �
  �
        ,            e         �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C<g   ]   ~         �   
   "     �   "  �   �        �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   6   2              �t�bhhK ��h��R�(KK��h�C@         �  <  �        �  a  y      "  �        �t�bhhK ��h��R�(KK��h�C            �         �t�bhhK ��h��R�(KK��h�CpU            5   x      <      "     J   6  +   ,            2     k     a     2  �	        �t�bhhK ��h��R�(KK
��h�C(H     $   E           �         �t�bhhK ��h��R�(KK��h�C   '   )   
           �t�be(hhK ��h��R�(KK��h�C �     �         >	        �t�bhhK ��h��R�(KK��h�C8         �           �                     �t�bhhK ��h��R�(KK��h�C<�     n     �     Y      O      �   �            �t�bhhK ��h��R�(KK��h�C`  �   X   �            �t�bhhK ��h��R�(KK��h�C,�        (   �      	      	         �t�bhhK ��h��R�(KK��h�C4A                c   %  �
     5         �t�bhhK ��h��R�(KK��h�C8*            n         �      M      ]        �t�bhhK ��h��R�(KK��h�C �  W  �  '      @          �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C,
   y  ?      �  
   H   B   �        �t�bhhK ��h��R�(KK��h�C\�  "   Q  �       a  �      O                   �      �             �t�bhhK ��h��R�(KK��h�C        �              �t�bhhK ��h��R�(KK��h�C;     	      	         �t�bhhK ��h��R�(KK��h�C@W  �     �  $   �      �  �  s   �   y      l        �t�bhhK ��h��R�(KK��h�C�  (  �          �t�bhhK ��h��R�(KK��h�C �   p      ^  M  	         �t�bhhK ��h��R�(KK��h�CD;     =      �   �      -         �  $  �      �        �t�bhhK ��h��R�(KK��h�C1   #       m  �         �t�bhhK ��h��R�(KK��h�Cp         &   D  0   4      v        f   �      �	        �  �        �  �                  �t�bhhK ��h��R�(KK��h�C   O        
         �t�bhhK ��h��R�(KK��h�C�   p      M     �t�bhhK ��h��R�(KK��h�C,   5      o  ~        �          �t�bhhK ��h��R�(KK
��h�C(%     �           N   �        �t�bhhK ��h��R�(KK��h�C1   #       4     �      �t�bhhK ��h��R�(KK��h�CLq   �  �   �                    �   o     �     B   �        �t�bhhK ��h��R�(KK��h�C,'   !      �     �	        �        �t�bhhK ��h��R�(KK��h�CP�     t        �  +      `   V  �            �     u
  �        �t�bhhK ��h��R�(KK��h�C4   5   a      ~  *      	  �      [        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C<c  �   �                     W      �           �t�bhhK ��h��R�(KK��h�CpH  �              �         F        
      �     q
     q   �  �                       �t�bhhK ��h��R�(KK��h�C<         k      @            �   %   �   �        �t�bhhK ��h��R�(KK��h�C\      �  �        u     !        M     
   %  
     �  P              �t�bhhK ��h��R�(KK��h�C_     (         �t�bhhK ��h��R�(KK��h�C�  a         �t�bhhK ��h��R�(KK��h�C`            8        r  �     $   |  �     �      (     �     $   x        �t�bhhK ��h��R�(KK��h�CL      -   �   L   "               e  �     �      $   �        �t�bhhK ��h��R�(KK	��h�C$   \	     u  �	              �t�bhhK ��h��R�(KK��h�CP   m        G        <  �           �  *   �      �            �t�bhhK ��h��R�(KK��h�C@   �           V      �  V	  �   j      N   �        �t�bhhK ��h��R�(KK��h�C�  �     	         �t�bhhK ��h��R�(KK��h�C�          �t�bhhK ��h��R�(KK��h�C4*            9                �        �t�bhhK ��h��R�(KK��h�C\$   8             �         �   s   7         %        l  �        /      �t�bhhK ��h��R�(KK��h�C<   �   k     �  �      '   -   7       �        �t�bhhK ��h��R�(KK��h�C    R     �     >        �t�bhhK ��h��R�(KK��h�CX#   !      4      m     �   ?      
   T              �        �         �t�bhhK ��h��R�(KK��h�C`      �     �         
  i   �   �      >      F  $   �  G   H     �           �t�bhhK ��h��R�(KK��h�C4         4      �   +   ;      �            �t�bhhK ��h��R�(KK��h�C0   X   '   6     #  �
     �           �t�bhhK ��h��R�(KK��h�C8E  �                  *         �  �         �t�bhhK ��h��R�(KK��h�CP   J  C      !                            �  9   I   �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C1   #       �        �t�bhhK ��h��R�(KK��h�C8#   !      8  ?      
   3   6         8        �t�bhhK ��h��R�(KK	��h�C$      �                    �t�bhhK ��h��R�(KK��h�C;     :     �t�bhhK ��h��R�(KK��h�C@�       �     )   �   
   �  �            �        �t�bhhK ��h��R�(KK��h�C    �  '      �
  &        �t�bhhK ��h��R�(KK��h�CL      P      &     z	     <         
   q           F         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK
��h�C(      )   b   $   ]     ,         �t�bhhK ��h��R�(KK!��h�C�%   �     �   �     v           ;      �               8   �   �               $   2  Y     �   �  �         �t�bhhK ��h��R�(KK��h�C<�  �      S      �          �                 �t�bhhK ��h��R�(KK��h�C@        �     ,     �   p   �   
   ,               �t�bhhK ��h��R�(KK��h�CD!         #        �        ?      
   3   6            �t�bhhK ��h��R�(KK��h�C�      �      W      �t�bhhK ��h��R�(KK��h�C'  �         �t�bhhK ��h��R�(KK��h�C,#   !   (      "   �     $   k         �t�bhhK ��h��R�(KK��h�C8      a   ;      j     �   �   |      �         �t�bhhK ��h��R�(KK��h�C      �              �t�bhhK ��h��R�(KK��h�C8
   f   [     )   �     �        �	  �        �t�bhhK ��h��R�(KK��h�C8               �     =        �   /         �t�bhhK ��h��R�(KK��h�C4      -   �   L      Z  
      �   N        �t�bhhK ��h��R�(KK��h�C|   �      �     �     �     �      K     ~      D      �  A        K     ~   e  U   |     <        �t�bhhK ��h��R�(KK��h�C,           �        '  �        �t�bhhK ��h��R�(KK��h�C                   �t�bhhK ��h��R�(KK��h�C   	      	   K      �t�bhhK ��h��R�(KK��h�C�         	     �t�bhhK ��h��R�(KK��h�CH      �   (  *        �  V     v   �  �                 �t�bhhK ��h��R�(KK��h�C1   #       ,     �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK
��h�C("   >     �  �  �     Z        �t�bhhK ��h��R�(KK��h�Ci  n      �t�bhhK ��h��R�(KK
��h�C(2      -   �   �        C        �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   6   �             �t�bhhK ��h��R�(KK��h�C@     �t�bhhK ��h��R�(KK��h�CLi     i     �   +            �             �   h   �         �t�bhhK ��h��R�(KK��h�C_     �t�bhhK ��h��R�(KK��h�Cp2  R      �  
   I   �  V   �  �        .   
   �     y     �   	                 	        �t�bhhK ��h��R�(KK��h�C\�
  :  "                                 ^  :  �   "   �     �
           �t�bhhK ��h��R�(KK��h�C!      $  R      �t�bhhK ��h��R�(KK��h�C�   T     �t�bhhK ��h��R�(KK��h�C8#   !      .     �  ?      
   X   �   F         �t�bhhK ��h��R�(KK	��h�C$�   R         	      	         �t�bhhK ��h��R�(KK��h�C<      �  �     '       X     �  
   �        �t�bhhK ��h��R�(KK��h�C�            �t�bhhK ��h��R�(KK��h�C,1   #          }     o               �t�bhhK ��h��R�(KK��h�C8   >   =      8     4   y      �               �t�bhhK ��h��R�(KK��h�CX         Y     �  �   7      �           0   �  �     A  ,  _        �t�bhhK ��h��R�(KK��h�C`�  (         �      f   �
        .            W     �      *  �               �t�bhhK ��h��R�(KK��h�C   e   '   �   �         �t�bhhK ��h��R�(KK��h�C0!      �     o      r  	      	         �t�bhhK ��h��R�(KK��h�CD      �     L      A        Z  g            �         �t�bhhK ��h��R�(KK��h�C,   $     .        �     &
        �t�bhhK ��h��R�(KK��h�C8
         �  �  e      %        H            �t�bhhK ��h��R�(KK��h�C(   2   �   �   r      �t�bhhK ��h��R�(KK��h�C82           
   �   �        �     �        �t�bhhK ��h��R�(KK��h�C�   =  	      	         �t�bhhK ��h��R�(KK��h�C�      �      �t�bhhK ��h��R�(KK��h�C,$     .   $   �   N                 �t�bhhK ��h��R�(KK��h�CL   �   l      S	  &   2              �  �      �  �  7         �t�bhhK ��h��R�(KK��h�CZ             �t�bhhK ��h��R�(KK��h�C\   H              �t�bhhK ��h��R�(KK��h�C4                     2	        A         �t�bhhK ��h��R�(KK��h�C4         P         {        J  E         �t�bhhK ��h��R�(KK��h�C\�      .   8   �     $        |      �        \   �     N  G  
            �t�bhhK ��h��R�(KK
��h�C(      )   }     P  
   t         �t�bhhK ��h��R�(KK��h�C8      b      �  �     .   "   e   �            �t�bhhK ��h��R�(KK��h�CP!      P  	      	      	   K   	   �   	     	   �  	   �   	   �     �t�bhhK ��h��R�(KK��h�C   g     �t�bhhK ��h��R�(KK��h�CX
      +        �     B   �     �        �  �  �      �  
            �t�bhhK ��h��R�(KK��h�C   e   '   �   �        �t�bhhK ��h��R�(KK��h�C1   #       �         �t�bhhK ��h��R�(KK��h�C0      -   P   �  :   W   )              �t�bhhK ��h��R�(KK��h�C1   #       +     �t�bhhK ��h��R�(KK��h�C1   #               �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C4�            �   �
     �  ^  7            �t�bhhK ��h��R�(KK��h�C�     �	           �t�bhhK ��h��R�(KK��h�C  �   ^     �t�bhhK ��h��R�(KK��h�C      �   �         �t�bhhK ��h��R�(KK��h�C<      �   L   a  �      �     9  
   N  �        �t�bhhK ��h��R�(KK��h�C   6  n     �         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CD�  �  $   �     �        0             H  �         �t�bhhK ��h��R�(KK��h�C4      0   �  �            k               �t�bhhK ��h��R�(KK��h�C\      \       �  c         ]  (        ^  )      $   k         X         �t�bhhK ��h��R�(KK��h�Cl         �                   f   '        V        5      �  +      }     �         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C4|               E     �  a  r           �t�bhhK ��h��R�(KK%��h�C�      P                    E     o  �        �  �      �  �        c                         J  E      �        �t�bhhK ��h��R�(KK��h�C,!          	      	      	   �     �t�bhhK ��h��R�(KK��h�C\            �      �        �     ,   	      	      	   K   	   �   	        �t�bhhK ��h��R�(KK
��h�C(        	      	     	   �      �t�bhhK ��h��R�(KK��h�C<         m      8   �      �        U   C        �t�bhhK ��h��R�(KK��h�C0*      �     �  I  5      �            �t�bhhK ��h��R�(KK��h�C<   ?   !         �   �  
   3   6     �   �        �t�bhhK ��h��R�(KK��h�CP            2        I     �  Z     �     -     �          �t�bhhK ��h��R�(KK��h�C        �t�bhhK ��h��R�(KK��h�C<1  �       
         7      *   x     b        �t�bhhK ��h��R�(KK��h�C�  �  �     �t�bhhK ��h��R�(KK��h�C\   �  $        j      A   7	  �   J    J  n            �     �  �
        �t�bhhK ��h��R�(KK��h�C   D     �t�bhhK ��h��R�(KK��h�CD     $  �      �   �  �   �     .      �     	        �t�bhhK ��h��R�(KK	��h�C$#   !   (      
   u  F         �t�bhhK ��h��R�(KK��h�C4#   !      Q     (      "   $   �   N        �t�bhhK ��h��R�(KK��h�C8   �  �  
        %               �        �t�bhhK ��h��R�(KK��h�CP           m      �     �     �        �  0   <   "   �
        �t�bhhK ��h��R�(KK��h�Cd
   "       1     S   1        �                �           4
     �        �t�bhhK ��h��R�(KK��h�C  7      �t�bhhK ��h��R�(KK��h�C4      "        �  c      +      �        �t�bhhK ��h��R�(KK��h�C         9     �t�bhhK ��h��R�(KK��h�C,   >  H  %
        <
     �
        �t�bhhK ��h��R�(KK��h�CD   t  5      �   �     �               �      z         �t�bhhK ��h��R�(KK��h�CD*         1
  L                 �     �      L         �t�bhhK ��h��R�(KK	��h�C$W          �     �         �t�bhhK ��h��R�(KK��h�C4;
  <
   	     �                         �t�bhhK ��h��R�(KK��h�C              }        �t�bhhK ��h��R�(KK��h�C4�       �       �      �
     �        �t�bhhK ��h��R�(KK��h�C8[        "           �     �     �         �t�bhhK ��h��R�(KK��h�C@      �   =         r
          �         �        �t�bhhK ��h��R�(KK��h�C4      �   O      �    7   �  
   n        �t�bhhK ��h��R�(KK��h�C0M     p            �  m           �t�bhhK ��h��R�(KK��h�C �     N   A  �  _        �t�bhhK ��h��R�(KK��h�C\           8   /      $      5               <      &      U      �        �t�bhhK ��h��R�(KK��h�C�  G   p     �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6            �t�bhhK ��h��R�(KK��h�CL#   !      t
     �  (      G   t      G   8   �  �              �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�C       P     G   W         �t�bhhK ��h��R�(KK��h�C4f   �  �  (      �  w                     �t�bhhK ��h��R�(KK��h�C@      U   k                    �               �t�bhhK ��h��R�(KK��h�CD              �   �         �  W      �      �        �t�bhhK ��h��R�(KK��h�C,�     S      >   2   �   i  w         �t�bhhK ��h��R�(KK��h�CT   �        9  
   ,      �	  
         �	  
         4  
   K         �t�bhhK ��h��R�(KK��h�CD   �      �                 �  ;   �     �           �t�bhhK ��h��R�(KK��h�C0      (      �         �  �   �         �t�bhhK ��h��R�(KK��h�C0$   �  �   /	  b  1     
   $   �        �t�bhhK ��h��R�(KK��h�C0   �  �              �   �          �t�bhhK ��h��R�(KK��h�C4      P   �   o      .         
   &        �t�bhhK ��h��R�(KK��h�Cp   �
  �
              ;     9     �     �     �      �              �   �               �t�bhhK ��h��R�(KK��h�CP   H     �t�bhhK ��h��R�(KK��h�CP"   ^  |      �     �           (      <         �     �        �t�bhhK ��h��R�(KK��h�C,   .   &         �   �             �t�bhhK ��h��R�(KK��h�CP   ,   �              �        �	  H
  
   8   �     8           �t�bhhK ��h��R�(KK��h�C >        	      	         �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C4U        $   8  (   N   �     �   �         �t�bhhK ��h��R�(KK��h�C<�   &   �   s   	        �  �  7   N   
   �        �t�bhhK ��h��R�(KK��h�CDe     y  =  i  z                 �   �	     T        �t�bhhK ��h��R�(KK��h�CP              4         �  �   *      �     #  �      u        �t�bhhK ��h��R�(KK��h�C P        	      	         �t�bhhK ��h��R�(KK��h�C6        	  u      �t�bhhK ��h��R�(KK��h�C1   #       j        �t�bhhK ��h��R�(KK&��h�C�            k                 �   �   _   �   +   ;      ,  %   �           >      v      P     �  %      �     �   �        �t�bhhK ��h��R�(KK��h�CP     �      N      .   �                 h                    �t�bhhK ��h��R�(KK	��h�C$k  �   +      }     E         �t�bhhK ��h��R�(KK��h�C4      -   P   <         t        �        �t�bhhK ��h��R�(KK��h�C@   �  C      P   <               �      �             �t�bhhK ��h��R�(KK��h�C>     �        �t�bhhK ��h��R�(KK��h�CT      �           �        �                 Q   V   �           �t�bhhK ��h��R�(KK��h�C|g  |      �     |      s	     �   E  R      l      �  
      �  �      �         
   �     �  �         �t�bhhK ��h��R�(KK��h�C      c     �t�bhhK ��h��R�(KK��h�C<      b   #      .  "   `	          8   �        �t�bhhK ��h��R�(KK��h�Cp
   3   6   �        K  '   !        U     �     ~      �   /      0      �      ~   �         �t�bhhK ��h��R�(KK��h�CL      �        �     ,   	      	   K   	   �   	     	   �      �t�bhhK ��h��R�(KK
��h�C(  �     �                    �t�bhhK ��h��R�(KK��h�C   N     ]	  7   v     �t�bhhK ��h��R�(KK	��h�C$      �     	      	         �t�bhhK ��h��R�(KK��h�C41   #      �  �   
   3   �  t     �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C@      �   �   "   �   �
  �     (                    �t�bhhK ��h��R�(KK��h�C,   5      �  8   <  T      j        �t�bhhK ��h��R�(KK
��h�C(=  �     )   �  ^  `   :        �t�bhhK ��h��R�(KK��h�Cp      5   [               D         �        \  L        x      .   "        Q           �t�bhhK ��h��R�(KK��h�C  ^     	         �t�bhhK ��h��R�(KK��h�CD�        L  
   `     �  �       7   m  �
  7         �t�bhhK ��h��R�(KK��h�C 1   #       /   "   �         �t�bhhK ��h��R�(KK��h�C`   f   q  5            4      m     �      5   �      4      R     f   �        �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C"  4  '     7         �t�bhhK ��h��R�(KK��h�C4*           �  v     .  b     �         �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C0      �  V     d  �  
      n         �t�bhhK ��h��R�(KK��h�Cl      �   ;  �  H   �        �                          B   �                       �t�bhhK ��h��R�(KK��h�C,4      �     R     A     7         �t�bhhK ��h��R�(KK��h�CD|      �   �  
     ^   T        R                     �t�bhhK ��h��R�(KK��h�C4�          l   9     7     h            �t�bhhK ��h��R�(KK	��h�C$i     k  5	  	      	         �t�bhhK ��h��R�(KK��h�CP   $   �     �        P   �  
           9   %   �  #  �        �t�bhhK ��h��R�(KK��h�C,      �   �     I   �     g        �t�bhhK ��h��R�(KK	��h�C$U   �  �      �     �        �t�bhhK ��h��R�(KK��h�C,   (   I  :   t      
   �  F         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C W              �  �     �t�bhhK ��h��R�(KK	��h�C$      (         ,  �        �t�bhhK ��h��R�(KK��h�C,  {   �  /   9   -     C  �        �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�C   S   �      �        �t�bhhK ��h��R�(KK��h�CP   �  [	     	  �  �         4  8   �  �   *      (   o  �         �t�bhhK ��h��R�(KK	��h�C$#   !   ?      
   �  F         �t�bhhK ��h��R�(KK��h�C2  �     �t�bhhK ��h��R�(KK��h�Cj     �t�bhhK ��h��R�(KK��h�CP         9     7         0                  
   �   �            �t�bhhK ��h��R�(KK��h�C,   L  �               �  �         �t�bhhK ��h��R�(KK��h�CH5     e  a  �         �  q  �   ]         C     >        �t�bhhK ��h��R�(KK��h�CX                 �                  U      �         �          �t�bhhK ��h��R�(KK#��h�C��     $   �     �	     .         (      �           �
  +         �   O         �         0     �  �               �t�bhhK ��h��R�(KK��h�Cd7               %     Y      z  �  J  J
     �              �   �   �   J
        �t�bhhK ��h��R�(KK��h�C!	     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK	��h�C$W      {          t        �t�bhhK ��h��R�(KK��h�CL   �       �            .   �      2     /     B           �t�bhhK ��h��R�(KK��h�C,b     �      �     K	  G   �        �t�bhhK ��h��R�(KK��h�C0      \  >      w   v                  �t�bhhK ��h��R�(KK	��h�C$B               B            �t�bhhK ��h��R�(KK	��h�C$!      �  �  	      	         �t�bhhK ��h��R�(KK��h�C<      l     �   �      7   T   D   �  P  7         �t�bhhK ��h��R�(KK���      h�C`         �         =         +  ^   =  b  *     �  �  	     �  *           �t�bhhK ��h��R�(KK��h�C8
   3   6         b      x   ?      #   h        �t�bhhK ��h��R�(KK ��h�C��  G  
      V         3     J  C   �   j	              .      (
  -  �     �     �        �  *        �t�bhhK ��h��R�(KK��h�CD   5  �     8   ?        ~         ,        �
        �t�bhhK ��h��R�(KK��h�C1   #       k        �t�bhhK ��h��R�(KK��h�C<            �t�bhhK ��h��R�(KK��h�C@        �  O  >        �  8     (             �t�bhhK ��h��R�(KK��h�C�       �t�bhhK ��h��R�(KK��h�CL�     '      �      �     �              .                  �t�bhhK ��h��R�(KK��h�C     �     �         �t�bhhK ��h��R�(KK��h�CL
   �                    ;  �     �              �
        �t�bhhK ��h��R�(KK��h�C0b   #      ]   "   �     8   �   Q         �t�bhhK ��h��R�(KK��h�C@      0   ,	  -   *         +               ^        �t�bhhK ��h��R�(KK��h�C    '                    �t�bhhK ��h��R�(KK��h�C1   #       k        �t�bhhK ��h��R�(KK��h�C8   X   '   H   �   	     )   �   �      /         �t�bhhK ��h��R�(KK��h�C,              �          �     �t�bhhK ��h��R�(KK
��h�C(      �  N   �  :   �            �t�bhhK ��h��R�(KK��h�C@   (   !      \      ]     n   
   3   6      n         �t�bhhK ��h��R�(KK��h�C,�     �           q               �t�bhhK ��h��R�(KK��h�CT      6        �   �  )               ;      �      �      R         �t�bhhK ��h��R�(KK��h�C<   �     z     a     L  z     a     b        �t�bhhK ��h��R�(KK��h�CD�   �     �  �	     �   
              �   "   �        �t�bhhK ��h��R�(KK��h�C`   /        a   �  o  �      �         S   Q            A   u  o	  �  �         �t�bhhK ��h��R�(KK
��h�C(   ?   �     J  
   �   F         �t�bhhK ��h��R�(KK��h�Cd      �         :  �   7      g
     :                  .               "        �t�bhhK ��h��R�(KK��h�CP%   �   �  -  :      �  T   $   �  �   �  �   8  �   �             �t�bhhK ��h��R�(KK��h�CT      �   �  [        f        �      �        �
  -               �t�bhhK ��h��R�(KK��h�C,   .     @      X   �     X         �t�bhhK ��h��R�(KK��h�C<                     z            0   �        �t�bhhK ��h��R�(KK��h�CP   %   �     �  �      �     �
  %  =	       $   �  �   �         �t�bhhK ��h��R�(KK��h�C0   �  �     �  �      k               �t�bhhK ��h��R�(KK��h�C,�                  .
     _        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C1   #       �        �t�bhhK ��h��R�(KK��h�C0�     �        �     	      	         �t�bhhK ��h��R�(KK ��h�C��   |      �  �  8  �   �   V     l
           �      �     �  �   4        �      �     �  
   N        �t�bhhK ��h��R�(KK��h�CD�        +      �  �     8   �     a                 �t�bhhK ��h��R�(KK��h�Cm         �       �t�bhhK ��h��R�(KK��h�C 8            4   �        �t�bhhK ��h��R�(KK��h�C          G      �        �t�bhhK ��h��R�(KK��h�C8B   P          �     �     �              �t�bhhK ��h��R�(KK��h�C�      	         �t�bhhK ��h��R�(KK
��h�C(�  $  0     �  `  
            �t�bhhK ��h��R�(KK��h�C�  "   �   �     �t�bhhK ��h��R�(KK��h�C   %     �         �t�bhhK ��h��R�(KK��h�CT         &   D  P      +  G   4     &      a   4      �      7         �t�bhhK ��h��R�(KK
��h�C(   '   )   A         !  �         �t�bhhK ��h��R�(KK!��h�C�
   3   6      w     e   ?      3     '        �  +      e         0   <   "   �     �  m      m      �         �t�bhhK ��h��R�(KK��h�C8         
   _      $   �  5   <         &     �t�bhhK ��h��R�(KK��h�CX!      �        �   X     d  (               �     B   
               �t�bhhK ��h��R�(KK��h�C`�     �  �          �         /      �  �      �      �          �         �t�bhhK ��h��R�(KK��h�CL*         H       n   �       s  +         J   a            �t�bhhK ��h��R�(KK��h�C`   �      �           %   H  �     �         �      �      �   �     �        �t�bhhK ��h��R�(KK	��h�C$�         �  �  �  �        �t�bhhK ��h��R�(KK	��h�C$
   Z        -   �   ,        �t�bhhK ��h��R�(KK��h�C8                  
            -            �t�bhhK ��h��R�(KK
��h�C(         .        �           �t�bhhK ��h��R�(KK��h�C�      	      	         �t�bhhK ��h��R�(KK��h�C,H  [        &   R  4               �t�bhhK ��h��R�(KK��h�C�     �            �t�bhhK ��h��R�(KK��h�C4!      1     n   ?      
   3   6           �t�bhhK ��h��R�(KK��h�CH            ;      �   %   �           U      �            �t�bhhK ��h��R�(KK��h�C   z            �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�Cl#   !         (      
                              @     �        �        _        �t�bhhK ��h��R�(KK��h�C�  v     �t�bhhK ��h��R�(KK��h�Cd            o  e
           �  �               R  4         
   _      ]         �t�bhhK ��h��R�(KK��h�CH                        )              �              �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�C<         f  �     �t�bhhK ��h��R�(KK��h�C`*              +      �  �	     T
                         I
     N        �t�bhhK ��h��R�(KK��h�C      0   �        �t�bhhK ��h��R�(KK��h�C 2   >   v                 �t�bhhK ��h��R�(KK��h�C@   �
  �   O   �     �         
  o  �   "   �        �t�bhhK ��h��R�(KK��h�C@         O      �   S   Q   5         4      m        �t�bhhK ��h��R�(KK��h�C`w  3        �     �   u   y  �         �      S   �          Q     �        �t�bhhK ��h��R�(KK��h�C!            	         �t�bhhK ��h��R�(KK
��h�C(      �   K     �     .          �t�bhhK ��h��R�(KK	��h�C$�      �      �               �t�bhhK ��h��R�(KK��h�CX   J                �            �           �     .              �t�bhhK ��h��R�(KK
��h�C(T   �  D       �      �        �t�bhhK ��h��R�(KK��h�Cf     E      �        �t�bhhK ��h��R�(KK	��h�C$   X   '   H   �              �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK
��h�C(�        j   %   �      v        �t�bhhK ��h��R�(KK��h�CP2            �   �      �   2      J        �        �   n         �t�bhhK ��h��R�(KK��h�C l     �         �         �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�C        �t�bhhK ��h��R�(KK��h�C8�        �   )         A   8     C            �t�bhhK ��h��R�(KK��h�Cx         E  `  �      J     `   �               0   !        "   �  R      �      '
     .        �t�bhhK ��h��R�(KK	��h�C$            �  �  �        �t�bhhK ��h��R�(KK	��h�C$   (   !      �   "   0        �t�bhhK ��h��R�(KK��h�C<m        �   q   �  $  I   /      ~               �t�bhhK ��h��R�(KK��h�CD      �  �  =     $   E   �   ]      �  ^   8   t        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK	��h�C$         �     �   �         �t�bhhK ��h��R�(KK��h�C0M      +      �  3  *      �          �t�bhhK ��h��R�(KK��h�CL   .   �  �         �  w   4     �  �   �   �  �	     �        �t�bhhK ��h��R�(KK��h�C   p      M  	         �t�bhhK ��h��R�(KK��h�C  �     �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�Ch#   !      <      /      G  w  (      
   3   6   )  ?   �   <   *   /      �      m   r      �t�bhhK ��h��R�(KK��h�C       '   P              �t�bhhK ��h��R�(KK��h�CH�                �      �     9        �      q     �     �t�bhhK ��h��R�(KK��h�C,      i     
   �
  �     F         �t�bhhK ��h��R�(KK��h�C             �t�bhhK ��h��R�(KK��h�C       
   �        �t�bhhK ��h��R�(KK��h�Cl   �     ;              �  �  e  0     {     %   _  C            �     ;  �        �t�bhhK ��h��R�(KK	��h�C$   �  (        
   Z        �t�bhhK ��h��R�(KK��h�C[            �t�bhhK ��h��R�(KK��h�CH#   !      {      	        ?      
   3   6   S
     s        �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C   9          X     �t�bhhK ��h��R�(KK��h�C !     �   �     �        �t�bhhK ��h��R�(KK��h�C0   �   Z  h      �   t  a     5        �t�bhhK ��h��R�(KK��h�C4I      *        �        %   �   �        �t�bhhK ��h��R�(KK��h�C  �  r      �t�bhhK ��h��R�(KK��h�C\            ;      �   %   �        
           �   L   
      �   D        �t�bhhK ��h��R�(KK��h�C �     K  	      	         �t�bhhK ��h��R�(KK��h�C<   �        �  �     ^     s   �     /         �t�bhhK ��h��R�(KK��h�CD#   !      4      �   ?      
   3   6      �               �t�bhhK ��h��R�(KK	��h�C$        >        4        �t�bhhK ��h��R�(KK��h�C      �                  �t�bhhK ��h��R�(KK
��h�C(�     )  �   �     9            �t�bhhK ��h��R�(KK��h�C      �          �t�bhhK ��h��R�(KK��h�CL      5   �       &      �   D  �   +     �  �               �t�bhhK ��h��R�(KK��h�CD
   `     F   '   #   !         R      �  �   Y
          �t�bhhK ��h��R�(KK��h�CH�      �        V           �         �  �     W         �t�bhhK ��h��R�(KK��h�Ch      0   �  �  :   *  <              �       G     �  �  �  y      �  f        �t�bhhK ��h��R�(KK��h�C8
   l	  �  ?      �   !      .  
   B   [        �t�bhhK ��h��R�(KK
��h�C(#        	      	      	   K      �t�bhhK ��h��R�(KK��h�C<   ?   �      �  "         
                     �t�bhhK ��h��R�(KK��h�C,   R           f         �        �t�bhhK ��h��R�(KK��h�C#     �   �   r      �t�bhhK ��h��R�(KK��h�C    
   4  	      	         �t�bhhK ��h��R�(KK��h�CH      )  8   /      �   ^   &     �      \  �   
            �t�bhhK ��h��R�(KK��h�C,      P   n     
   H   B   �        �t�bhhK ��h��R�(KK��h�C�
  !      �t�bhhK ��h��R�(KK��h�CX   �   �         �           8   f
  S              -   G     u        �t�bhhK ��h��R�(KK��h�C<Q     z     6        �   #     $     �        �t�bhhK ��h��R�(KK��h�C,h            /   9     7         �t�bhhK ��h��R�(KK
��h�C(
        �       ]           �t�bhhK ��h��R�(KK��h�CdP     O  (  "      �             �     �   d     (   S     �   �      �         �t�bhhK ��h��R�(KK��h�C �   J  �   /      �         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CP�     ~           -   P   T     �   /      e      @      X         �t�bhhK ��h��R�(KK
��h�C(        �   &  V     �         �t�bhhK ��h��R�(KK��h�C4            [  /  $            �        �t�bhhK ��h��R�(KK��h�CH            o  ~        P   +  G   @   �   ^               �t�bhhK ��h��R�(KK��h�CDb   #      ?  
   k        �  
        l     W        �t�bhhK ��h��R�(KK ��h�C�                     �                 -   %   �   (   �   ,  �  T      V  �      �     /  C           �t�bhhK ��h��R�(KK��h�C,   5      �  8   <  *      j        �t�bhhK ��h��R�(KK��h�C@E      )        <    �   s     ^   �     s        �t�bhhK ��h��R�(KK��h�C�      N          �t�bhhK ��h��R�(KK��h�C,%   �  �      S  �  �   c  P
        �t�bhhK ��h��R�(KK��h�Cp      -  �      �t�bhhK ��h��R�(KK��h�C8     �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C
   �  1     �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C      	      	         �t�bhhK ��h��R�(KK��h�C8   5      �  :   q           `              �t�bhhK ��h��R�(KK��h�C4   e  /      0   g     d   �              �t�bhhK ��h��R�(KK��h�CV     �t�bhhK ��h��R�(KK��h�C �     '      �   E        �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK	��h�C$T     #      �  i           �t�bhhK ��h��R�(KK	��h�C$              �  �        �t�bhhK ��h��R�(KK��h�C<�              @           [                �t�bhhK ��h��R�(KK��h�Cu        �t�bhhK ��h��R�(KK
��h�C(   �     .                     �t�bhhK ��h��R�(KK
��h�C(   �        �   �   �  7         �t�bhhK ��h��R�(KK��h�Cl      5   �      L      |      �   &      U   |      �   �   �   �      �      L   
   �        �t�bhhK ��h��R�(KK.��h�C�X  �     R        �  �        |     
   _            d     �
        ]                          @             �     �   E     �               �t�bhhK ��h��R�(KK*��h�C�      =         �               J   �        =  M                    �  Y  �  �   7      y  y      �         
     �  
   A   F        �t�bhhK ��h��R�(KK��h�C4   D         -        U         W        �t�bhhK ��h��R�(KK��h�C   �  �     .          �t�bhhK ��h��R�(KK��h�C@         :      �    :      T           �        �t�bhhK ��h��R�(KK��h�CH      J   P         �   =  &      }        �     =        �t�bhhK ��h��R�(KK��h�C8      )   \  �  x
  y
              @         �t�bhhK ��h��R�(KK��h�C<      �  �        �
  `   �     ,               �t�bhhK ��h��R�(KK��h�C4�  �  >      �  ^     �   �   A   �        �t�bhhK ��h��R�(KK��h�C 1        	      	         �t�bhhK ��h��R�(KK	��h�C$      =      @  G   W         �t�bhhK ��h��R�(KK��h�C`         
  $   ~  �   e  i   "   t      J   a      k      >      )   \  t         �t�bhhK ��h��R�(KK��h�C<r     �           0   #   L   
   +      v         �t�bhhK ��h��R�(KK��h�Cx9   %   /
     (   2      N            .   �
  
         �  
     
   �        �   I	  �     3        �t�bhhK ��h��R�(KK��h�C    �        9           �t�bhhK ��h��R�(KK��h�C�  �     3          �t�bhhK ��h��R�(KK��h�C,�   q   7     �     `  �           �t�bhhK ��h��R�(KK��h�C 1   #            �        �t�bhhK ��h��R�(KK��h�C�	     /      �      �t�bhhK ��h��R�(KK��h�CX              �t�bhhK ��h��R�(KK��h�CP           .   N                                 �          �t�bhhK ��h��R�(KK��h�C<   �      �  ;     �                 �        �t�bhhK ��h��R�(KK��h�C    �   �  �      �  r      �t�bhhK ��h��R�(KK��h�Ch      �   �  R      �           C              %   &   D  �   '  �   �     "        �t�bhhK ��h��R�(KK��h�CX	  �
        �        �      �     �     �	           W      �        �t�bhhK ��h��R�(KK
��h�C(\   �  m  r   ,   	      	         �t�bhhK ��h��R�(KK��h�C@         W       4           �   �     �        �t�bhhK ��h��R�(KK
��h�C(*                    '        �t�bhhK ��h��R�(KK��h�C8         �  $   �  ^   �     s     4        �t�bhhK ��h��R�(KK��h�C|   7  �            O  ,           C  D     &   �
  f     �      �         �         �   b	        �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK	��h�C$      0   �  9   :           �t�bhhK ��h��R�(KK��h�C�     �  U     P     �t�bhhK ��h��R�(KK��h�CL           <         �     G   |     <        $   k         �t�bhhK ��h��R�(KK��h�C`*      '              8   �            �      z     �   �         �   �        �t�bhhK ��h��R�(KK��h�C9        �t�bhhK ��h��R�(KK��h�C            
         �t�bhhK ��h��R�(KK��h�C<M   -     
      "  �  %               `        �t�bhhK ��h��R�(KK��h�C   �      r  	         �t�bhhK ��h��R�(KK��h�C4�  j  /           b         �  �        �t�bhhK ��h��R�(KK
��h�C(      �   �     G   I   C        �t�bhhK ��h��R�(KK��h�Cc  �      $           �t�bhhK ��h��R�(KK��h�C            �  S     �t�bhhK ��h��R�(KK��h�C,      -      .   U                  �t�bhhK ��h��R�(KK��h�C5       �     �t�bhhK ��h��R�(KK��h�CX   @   '      �           V      �        /      8     	  �  '        �t�bhhK ��h��R�(KK��h�CS  �          �t�bhhK ��h��R�(KK��h�Cd     z          L  9  �     ,         �        �  �     S   }      X        �t�bhhK ��h��R�(KK
��h�C(   	      	      	   K   	   U     �t�bhhK ��h��R�(KK��h�CD   �   o      h     	  -   �  :      Q         S         �t�bhhK ��h��R�(KK��h�CP*      �      �  &      M                              L         �t�bhhK ��h��R�(KK��h�C	     �     �t�bhhK ��h��R�(KK��h�CT   u           �  �           0   �  
   _      �   }              �t�bhhK ��h��R�(KK��h�C�             �t�bhhK ��h��R�(KK��h�CD   �  :  2   ,            �   S                        �t�bhhK ��h��R�(KK��h�C -   �       
           �t�bhhK ��h��R�(KK��h�C8         �   �     �  �  �     �   �         �t�bhhK ��h��R�(KK��h�C       r  �   ^   &        �t�bhhK ��h��R�(KK��h�C�       r     �t�bhhK ��h��R�(KK��h�C81   #              
   3   6   1     	        �t�bhhK ��h��R�(KK��h�C   h
  -  �          �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK	��h�C$1   #       �  �      S        �t�bhhK ��h��R�(KK	��h�C$   %   �    '               �t�bhhK ��h��R�(KK��h�C@�     0   �     .   ^                              �t�bhhK ��h��R�(KK#��h�C�              Y     A   Y      ?  i            �   Q                             a   ;      �  :   �   ?        �t�bhhK ��h��R�(KK��h�C@"   e   �               (      #   !      �   R         �t�bhhK ��h��R�(KK	��h�C$�      p  "                  �t�bhhK ��h��R�(KK��h�C8�        0  B   �  �  m   0  �     �         �t�bhhK ��h��R�(KK	��h�C$�
  
      �     B            �t�bhhK ��h��R�(KK��h�CH�	     �   �  W        .   �           �   �               �t�bhhK ��h��R�(KK��h�C,�     @      C  6     U            �t�bhhK ��h��R�(KK��h�C0   @   '   H   d        �      I         �t�bhhK ��h��R�(KK��h�CG	     �t�bhhK ��h��R�(KK��h�CX
   �  _      4   R     .         K        b       7   v     �         �t�bhhK ��h��R�(KK
��h�C(   :  "           c          �t�bhhK ��h��R�(KK��h�CG           c     �t�bhhK ��h��R�(KK��h�CD      -   �   L   G               ~  "      �   D        �t�bhhK ��h��R�(KK��h�C01   #      o  �   
   3   6   	  �         �t�bhhK ��h��R�(KK��h�C,D  �       T   (                 �t�bhhK ��h��R�(KK��h�C                          �t�bhhK ��h��R�(KK��h�CL   �               i     %   0   <                 ^
        �t�bhhK ��h��R�(KK��h�CTj          �  V   %   �                  �        �     �         �t�bhhK ��h��R�(KK��h�C:  �     �     �      �t�bhhK ��h��R�(KK��h�C �
  Y     z  #  �         �t�bhhK ��h��R�(KK
��h�C(�      l      �  �     	         �t�bhhK ��h��R�(KK��h�C0Z         �     �  �      �     9     �t�bhhK ��h��R�(KK	��h�C$   ;         	      	         �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   6                  �t�bhhK ��h��R�(KK��h�C0I   /  h   t     ;      8  j           �t�bhhK ��h��R�(KK��h�CX      P   !                                 .   
            _        �t�bhhK ��h��R�(KK��h�Cq     �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C,   <         D  '     .   �          �t�bhhK ��h��R�(KK��h�CP      D  =         +  G   4     >      a   4      �      7         �t�bhhK ��h��R�(KK��h�C_     �         �t�bhhK ��h��R�(KK��h�CS  �         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C<   �	     �         &      �   �     B           �t�bhhK ��h��R�(KK��h�C0W   	  )   %              �   ^        �t�bhhK ��h��R�(KK��h�C          I   �            �t�bhhK ��h��R�(KK��h�C3         �t�bhhK ��h��R�(KK
��h�C(      �  �   j   �     s   7      �t�bhhK ��h��R�(KK��h�C�	  �   S   }         �t�bhhK ��h��R�(KK��h�C �      ,   �   "   �   n     �t�bhhK ��h��R�(KK��h�C 1     �        �         �t�bhhK ��h��R�(KK��h�C\            ;      �   %   �              ;      �  ~	  h      �   t        �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C4   o  �   5         g     w    �        �t�bhhK ��h��R�(KK��h�C\-   @   g  �        7  �
        �     X      V     �   
         �        �t�bhhK ��h��R�(KK��h�Cn             �t�bhhK ��h��R�(KK��h�Cpy      �      o  �         �      M     
      �  �   -      3        Q   V         O         �t�bhhK ��h��R�(KK��h�CD
       d   �      
        �      V     )   	        �t�bhhK ��h��R�(KK��h�C02      �                 '  �        �t�bhhK ��h��R�(KK��h�CL]   v        �  �      E      �  h      7   g   $   �  �         �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C\!           �   (      "   k     �  "   L     ~     p      "   �  �        �t�bhhK ��h��R�(KK��h�C<            �  �  �  �     �  �               �t�bhhK ��h��R�(KK��h�C�  	     �t�bhhK ��h��R�(KK��h�C8#   !               (      
   @   �   F         �t�bhhK ��h��R�(KK��h�C8�  �        O          �     �  �         �t�bhhK ��h��R�(KK��h�C,/      )   ;         �     �        �t�bhhK ��h��R�(KK��h�CD         �  "   �      (        -   z         X        �t�bhhK ��h��R�(KK��h�Ct   r  '     �     �  �      +   e  
   �   |      �     h   �   �            .   h   %   �	        �t�bhhK ��h��R�(KK��h�C<�   �   +   x      B   
  :      �        S         �t�bhhK ��h��R�(KK��h�C*         %         �t�bhhK ��h��R�(KK��h�CH         .   �  (   {         �        =        �        �t�bhhK ��h��R�(KK��h�C)     �t�bhhK ��h��R�(KK	��h�C$         �   �              �t�bhhK ��h��R�(KK��h�C8   $   �  &           8   4      �  �        �t�bhhK ��h��R�(KK��h�C4�     /      �   '   �         �  �        �t�bhhK ��h��R�(KK��h�C      0   �        �t�bhhK ��h��R�(KK��h�C<#   !      �   �   z        ?      9   �   �         �t�bhhK ��h��R�(KK��h�C
     �t�bhhK ��h��R�(KK��h�CP      U      W       i                 m      �     �        �t�bhhK ��h��R�(KK��h�CH1   #         }     o   
   3   6   7  }     o               �t�bhhK ��h��R�(KK��h�CP�      �       �  7      U   �       �  O     �  �           �t�bhhK ��h��R�(KK��h�C      	     �t�bhhK ��h��R�(KK��h�C8=  �     J         )   �  `   �     �        �t�bhhK ��h��R�(KK��h�C<   �  �      }     �     h  �	  �     �        �t�bhhK ��h��R�(KK
��h�C(�      r     v        �        �t�bhhK ��h��R�(KK��h�C�        	         �t�bhhK ��h��R�(KK	��h�C$   �  �  .   
   c  X         �t�bhhK ��h��R�(KK��h�CD#   !         =      �  4   ?      
   3   6   �  4         �t�bhhK ��h��R�(KK��h�C@^      �        =         n   "   -     .  �        �t�bhhK ��h��R�(KK��h�C<      �      �      L   G   �                  �t�bhhK ��h��R�(KK��h�C    4  '   -   H            �t�bhhK ��h��R�(KK��h�C       #                �t�bhhK ��h��R�(KK��h�CL         �           �   >      v                  �        �t�bhhK ��h��R�(KK��h�C    	      	         �t�bhhK ��h��R�(KK��h�CD         .      :   ,     C  5               �        �t�bhhK ��h��R�(KK��h�Cp  �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C8   �  �      �        a      �             �t�bhhK ��h��R�(KK��h�C
     �t�bhhK ��h��R�(KK��h�Ci     �t�bhhK ��h��R�(KK��h�C4
   3   6   �  '   #   !      �   k  �        �t�bhhK ��h��R�(KK��h�C8#   !      �  (      
   3   6   9     	        �t�bhhK ��h��R�(KK��h�CH%   �  �  ~         �     �        n      %   �  �        �t�bhhK ��h��R�(KK��h�Cp         $   8     �     B   _  z    �      .   9               �  _            4         �t�bhhK ��h��R�(KK��h�C@D      )   0   �                          �
        �t�bhhK ��h��R�(KK ��h�C�      �  8   /      V     5   �          D         .   *      &   $  �            U                     �t�bhhK ��h��R�(KK��h�C4y   �  L  &      e       A     �        �t�bhhK ��h��R�(KK	��h�C$#   !   (      
   u  F         �t�bhhK ��h��R�(KK��h�Cx                          L   �        /   9   -  &      M   �      4     8   �                 �t�bhhK ��h��R�(KK��h�CT�  /   5      .  �  q     j            �              B            �t�bhhK ��h��R�(KK
��h�C(4  L  �                       �t�bhhK ��h��R�(KK��h�CX*      &   �  �      8  (      [      .         i        Z  "           �t�bhhK ��h��R�(KK��h�C�
        �t�bhhK ��h��R�(KK��h�CX   $   �     �  ~   �                  0   4         
   _      �        �t�bhhK ��h��R�(KK��h�C   "   E     �t�bhhK ��h��R�(KK��h�C�
  V   �   �	     �t�bhhK ��h��R�(KK��h�CD   �         �        #        i     "  �   n         �t�bhhK ��h��R�(KK��h�C     Q   
  r  C      �t�bhhK ��h��R�(KK��h�C0      �   �  ^   �     
   �   F         �t�bhhK ��h��R�(KK��h�C<      �  �            �         �     #        �t�bhhK ��h��R�(KK��h�C    !  �                 �t�bhhK ��h��R�(KK��h�C8      )   z   �   A   }      �        �         �t�bhhK ��h��R�(KK��h�C0   &   �  W      �        l  �         �t�bhhK ��h��R�(KK��h�C T         �  �  w         �t�bhhK ��h��R�(KK��h�C<'  �   �        �  ^                          �t�bhhK ��h��R�(KK+��h�C�         O         Y      Q         Q     Q      x        �      %     z           ;      �      9   $            5   7  �  �               �t�bhhK ��h��R�(KK��h�Cd      R  4            �         `   8     �     ]             �
  �   O         �t�bhhK ��h��R�(KK-��h�C�         w      O         Y      Q      �     x  �   �     4              t        Y      O      >      =      2        t        Y      O         �t�bhhK ��h��R�(KK	��h�C$%   �  �           6        �t�bhhK ��h��R�(KK��h�Cd            
         �  �  (   �  �         &      b   x   "                     �t�bhhK ��h��R�(KK��h�CD   �     e  N      �   �        +     �   �            �t�bhhK ��h��R�(KK��h�C0�   l  �      y  T   D   �  P  7         �t�bhhK ��h��R�(KK��h�Cb     p      /      �t�bhhK ��h��R�(KK��h�C     ^     �t�bhhK ��h��R�(KK��h�C      	      	         �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C}     �t�bhhK ��h��R�(KK
��h�C(   5   7  �  �        �        �t�bhhK ��h��R�(KK��h�C,H     (      �  =                 �t�bhhK ��h��R�(KK
��h�C(�                    *        �t�bhhK ��h��R�(KK��h�Ch�   �  �     �   D   '  w  9   b                 J   �  �  D      m  �  �   �        �t�bhhK ��h��R�(KK
��h�C(2           <      �   m         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C      �         �t�bhhK ��h��R�(KK��h�C4R        �  	      	      	   K   	   �      �t�bhhK ��h��R�(KK��h�C   �     N      �t�bhhK ��h��R�(KK
��h�C(   R           <     �        �t�bhhK ��h��R�(KK��h�C8
   k  (      !      �           8   �        �t�bhhK ��h��R�(KK��h�CH      (      !      .   :   q      �     �     �	           �t�bhhK ��h��R�(KK��h�CZ         z        �t�bhhK ��h��R�(KK��h�C      9  	         �t�bhhK ��h��R�(KK��h�CD           '     �   x      \      &   $  `   �         �t�bhhK ��h��R�(KK��h�CT   (   #   !         #              e  /   
   3   6      e  /         �t�bhhK ��h��R�(KK��h�C�  ;     �t�bhhK ��h��R�(KK��h�CDT      %     �  �   O  �     �  �	  �     w
          �t�bhhK ��h��R�(KK	��h�C$)   �   �  ,   O      U        �t�bhhK ��h��R�(KK��h�CP      N   �  9     q  �  0  i         �              �         �t�bhhK ��h��R�(KK��h�C8�      :  I         $     	     �           �t�bhhK ��h��R�(KK��h�C4      &   �  C   &   �  N   
  "           �t�bhhK ��h��R�(KK��h�C,8   /         a      }      X        �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C@   	     %   �  #  �  �   Q
     `   b     �        �t�bhhK ��h��R�(KK��h�C    �   c  �      m        �t�bhhK ��h��R�(KK��h�C\
   �          F   '      H     %        B  �      *         �   �         �t�bhhK ��h��R�(KK��h�C      �     �     �t�bhhK ��h��R�(KK��h�C4      A     i  
        G  v  �        �t�bhhK ��h��R�(KK��h�C,�      �      +   �      �           �t�bhhK ��h��R�(KK	��h�C$@      [          u        �t�bhhK ��h��R�(KK��h�C<   �   8   .  @
  y            a  �      �        �t�bhhK ��h��R�(KK	��h�C$      -   b   �      �        �t�bhhK ��h��R�(KK��h�CD�   �      ;     l              �   f     �           �t�bhhK ��h��R�(KK��h�C�      u      �t�bhhK ��h��R�(KK��h�CX
   3   6   �     �      �  '   !      �   2      0   <      m      �        �t�bhhK ��h��R�(KK��h�C0      �   L   "   I   +  
   �   �        �t�bhhK ��h��R�(KK��h�CD   �  �   �           �      �         G              �t�bhhK ��h��R�(KK��h�Cw  �     �t�bhhK ��h��R�(KK��h�CF     �     �t�bhhK ��h��R�(KK��h�C�  	      	         �t�bhhK ��h��R�(KK��h�C<0       K         �     �  )      A   }         �t�bhhK ��h��R�(KK��h�C0H	  �   )   �   y  !      R      o        �t�bhhK ��h��R�(KK��h�C      =         �     �t�bhhK ��h��R�(KK��h�C0!         	      	      	   �   	   /     �t�bhhK ��h��R�(KK��h�C0�  ]   5         �                   �t�bhhK ��h��R�(KK��h�C8W   �   c   m  
   �   |  -      Y     �        �t�bhhK ��h��R�(KK��h�C       -      �            �t�bhhK ��h��R�(KK��h�C	     %   {
  �         �t�bhhK ��h��R�(KK
��h�C(4       P     "   �  �        �t�bhhK ��h��R�(KK��h�CP   '   �     R
     /     �   �         .     Q      �   [        �t�bhhK ��h��R�(KK��h�C\\   �        v    
   $   |     �   &      a     ]  �   �     �  7         �t�bhhK ��h��R�(KK��h�CD6  �     	  �           �  F     G     C  /         �t�bhhK ��h��R�(KK��h�C0v  R         .   	     b     �         �t�bhhK ��h��R�(KK��h�C4   8   �   �     �      �	     8   �         �t�bhhK ��h��R�(KK��h�Cp  L  
   t         �t�bhhK ��h��R�(KK��h�C@   �  C      �	  C      S  �     �   -               �t�bhhK ��h��R�(KK��h�Cx            �           *  X     -      �   �  B   R            .     K     �      -  	        �t�bhhK ��h��R�(KK��h�Cd      �  R  �     4   
   _            
   �   �   _   (   �      �   H              �t�bhhK ��h��R�(KK��h�CL   �  �   �  �   8  �   �  R     4      o     4      �	        �t�bhhK ��h��R�(KK��h�CHT            �            &      F  +           <        �t�bhhK ��h��R�(KK��h�Ch"   m   G   /      -  (   2   <   G                                                   �t�bhhK ��h��R�(KK
��h�C(�  �   -   h            Q	        �t�bhhK ��h��R�(KK ��h�C�      J   �     �        -           �        �                x      .   "   \           1        �t�bhhK ��h��R�(KK��h�C,   <        o      �     \
        �t�bhhK ��h��R�(KK��h�C�	     �t�bhhK ��h��R�(KK��h�CL         J   �  !     �  �  �     �     �     �  u        �t�bhhK ��h��R�(KK0��h�C�  ^     �   �      ,   "     ^        X  h   �                       �      ^  u           -      z   ,   h   �      :          �     "     ^           �t�bhhK ��h��R�(KK��h�C   �  �          �t�bhhK ��h��R�(KK��h�C1   #       �         �t�bhhK ��h��R�(KK��h�C	         �t�bhhK ��h��R�(KK��h�CLD     �     v   �  *      $        �      �  
               �t�bhhK ��h��R�(KK��h�C0�      �                             �t�bhhK ��h��R�(KK	��h�C$         L	                 �t�bhhK ��h��R�(KK��h�C<a  '      @   
   �     9                      �t�bhhK ��h��R�(KK��h�C1     +         �t�bhhK ��h��R�(KK
��h�C(�         (   w   �  �   d        �t�bhhK ��h��R�(KK��h�C@U   �  �         "     r          Z     %        �t�bhhK ��h��R�(KK��h�C\            2      �     �       A   |        (           
  L         �t�bhhK ��h��R�(KK��h�C<      5   <   �  &      I        *      j        �t�bhhK ��h��R�(KK��h�C4                 �  �     �  �        �t�bhhK ��h��R�(KK��h�CZ   c     �t�bhhK ��h��R�(KK��h�C8#   !      ]   '   
   3   6      �               �t�bhhK ��h��R�(KK��h�CT               �  G      o  �     (   �  q       �   :   P        �t�bhhK ��h��R�(KK��h�CT            ;      �   %   �              P   +         �   �        �t�bhhK ��h��R�(KK
��h�C(#   !   ?      
   X   �   F         �t�bhhK ��h��R�(KK��h�C   }     �t�bhhK ��h��R�(KK��h�C      1  	         �t�bhhK ��h��R�(KK��h�C8�   "     �   �   *                  �          �t�bhhK ��h��R�(KK��h�CDV                    �  �         �   f     �        �t�bhhK ��h��R�(KK��h�CH        �         �
     6  C         �  i      A         �t�bhhK ��h��R�(KK��h�C[      �     �t�bhhK ��h��R�(KK��h�C b      `  "   $            �t�bhhK ��h��R�(KK	��h�C$      �   "   T     :        �t�bhhK ��h��R�(KK��h�C0      N      .   �                    �t�bhhK ��h��R�(KK��h�CD      5   \  �       M   �      @                   �t�bhhK ��h��R�(KK��h�C�
  =  �  �     �t�bhhK ��h��R�(KK��h�CX     �t�bhhK ��h��R�(KK��h�C<7     �     �   �     
   �           �         �t�bhhK ��h��R�(KK��h�C\@   �   �   �      	  "   �     �     '  	     /         	  i   s   7         �t�bhhK ��h��R�(KK��h�CD      ,     R      $   �   x           k               �t�bhhK ��h��R�(KK��h�C4h  ?      
   3   6         b      x         �t�bhhK ��h��R�(KK��h�C    �      Q  :   W         �t�bhhK ��h��R�(KK��h�C          	      	         �t�bhhK ��h��R�(KK��h�Cp      -   �   L   G      �	     �   B  *      �  �     �        �      �     �     8        �t�bhhK ��h��R�(KK��h�C4!      1     �  ?      
   3   6   	        �t�bhhK ��h��R�(KK	��h�C$   "     �  	      	         �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6            �t�bhhK ��h��R�(KK	��h�C$�  �       	      	         �t�bhhK ��h��R�(KK��h�CDK     �     :   �          m  �      �     9        �t�bhhK ��h��R�(KK��h�C�   �     �t�bhhK ��h��R�(KK��h�CX   �   n  "   �     �   d  �      "   %   	     �           �           �t�bhhK ��h��R�(KK��h�C$   k      X      �t�bhhK ��h��R�(KK��h�Cx!      Y        	      	      	   �   	   �   	   I  	   /  	   s  	   )  	   �  	   �  	   �  	   �     �t�bhhK ��h��R�(KK��h�C�   "   |     �t�bhhK ��h��R�(KK��h�CL            �
        .         �        w                  �t�bhhK ��h��R�(KK��h�C             I  �        �t�bhhK ��h��R�(KK	��h�C$      '   #  `             �t�bhhK ��h��R�(KK��h�C �   �     N      .          �t�bhhK ��h��R�(KK��h�C8      "  c   �      �   �   9   A  s   7         �t�bhhK ��h��R�(KK
��h�C(
      �  '                     �t�bhhK ��h��R�(KK��h�C8�            .  %   M           A   ?        �t�bhhK ��h��R�(KK��h�C8     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�
  	         �t�bhhK ��h��R�(KK��h�C<      �   j  j      )               �	           �t�bhhK ��h��R�(KK��h�CLg     �        �        
  Q      Y      Q   5      {	        �t�bhhK ��h��R�(KK��h�CP             $   n      �     �           |  c      L         �t�bhhK ��h��R�(KK��h�C0h   5    )   �      ,      A   }         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C5     A      	         �t�bhhK ��h��R�(KK	��h�C$�  �  �      �              �t�bhhK ��h��R�(KK��h�C@W   	        B         �     �      ~               �t�bhhK ��h��R�(KK	��h�C$   �    
   �      D
        �t�bhhK ��h��R�(KK��h�Cx3         �             2                     4
        �     3          	  �
              �t�bhhK ��h��R�(KK��h�C b   #   "   $   �   �        �t�bhhK ��h��R�(KK��h�CI      ;               �t�bhhK ��h��R�(KK��h�CD      �            8   �     4         >   �   u        �t�bhhK ��h��R�(KK��h�Cp     �        �t�bhhK ��h��R�(KK��h�C<      )   J     �                 v            �t�bhhK ��h��R�(KK	��h�C$�        ;      o           �t�bhhK ��h��R�(KK��h�C1   #       `     �t�bhhK ��h��R�(KK��h�C8�  �   -   !      V
       Q        �         �t�bhhK ��h��R�(KK
��h�C(      0        	     
        �t�bhhK ��h��R�(KK��h�C8�     �
  �     ;     #          �        �t�bhhK ��h��R�(KK��h�CT      0   �  !      B           �  p     B   3     2              �t�bhhK ��h��R�(KK��h�CT         f       g   {      &      )  +      �  G   |      �         �t�bhhK ��h��R�(KK��h�C0>        '   9      �  
               �t�bhhK ��h��R�(KK��h�CTS     �        j      �            a   ;      �  �  �              �t�bhhK ��h��R�(KK��h�CP�   '      5           #           �   5     �   �     �         �t�bhhK ��h��R�(KK��h�Cw     x        �t�bhhK ��h��R�(KK��h�Cw  l     E        �t�bhhK ��h��R�(KK
��h�C(   @   '            �   �
        �t�bhhK ��h��R�(KK��h�C[         w  �     �t�bhhK ��h��R�(KK��h�C`"   t         0      �   ~                 �	     ]                 4         �t�bhhK ��h��R�(KK��h�C,      J     �   �     �  G        �t�bhhK ��h��R�(KK��h�C,#   !      P  '   
   �  �  F         �t�bhhK ��h��R�(KK��h�Cl   �         �            I     *      $  @     �        �           z              �t�bhhK ��h��R�(KK��h�C4      .                  �
             �t�bhhK ��h��R�(KK��h�C@�     �    �  8   /      
  y   �   W              �t�bhhK ��h��R�(KK��h�C4�   J  �   /      w  �      �     {        �t�bhhK ��h��R�(KK��h�CP      �       G  S     D   5                        >        �t�bhhK ��h��R�(KK��h�C4�         �         
   z        �        �t�bhhK ��h��R�(KK
��h�C(   �     �      �     |        �t�bhhK ��h��R�(KK��h�C   L  
   7        �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C\�  "   Q  �       a  �      O                   �      �             �t�bhhK ��h��R�(KK��h�CD   e   '      {     �
     V   ^     �         �        �t�bhhK ��h��R�(KK��h�CD%     8              :                     T        �t�bhhK ��h��R�(KK��h�C g              �        �t�bhhK ��h��R�(KK��h�C<   0   �	  �           �      a	           	     �t�bhhK ��h��R�(KK��h�C0�  0     �  �     %   H  �     �      �t�bhhK ��h��R�(KK��h�C      �        �t�bhhK ��h��R�(KK��h�C    �  �  :        �     �t�bhhK ��h��R�(KK��h�C   �         �t�bhhK ��h��R�(KK��h�C4s
           �     @      �     M        �t�bhhK ��h��R�(KK��h�ChO         Y      Q      #     $           x     )  C      �  ^   |      <  �        �t�bhhK ��h��R�(KK��h�C0   �  �        $  H      �   =        �t�bhhK ��h��R�(KK��h�C@   �   '                  �      x                  �t�bhhK ��h��R�(KK��h�C�	  �  �  "   t         �t�bhhK ��h��R�(KK%��h�C�               Y      Q         Q     Q      x        m                 &   $   �   �  &     �   
     +   "   �        �t�bhhK ��h��R�(KK��h�C       M  	      	         �t�bhhK ��h��R�(KK��h�C�  �        �t�bhhK ��h��R�(KK��h�CP      =      	              �           $        	          �t�bhhK ��h��R�(KK��h�C0   �  �   +   :   8   �   j      �       �t�bhhK ��h��R�(KK	��h�C$�                           �t�bhhK ��h��R�(KK��h�CX         �              �         a   ;      �   %   �                 �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�C�     _     �t�bhhK ��h��R�(KK��h�C8         k               ,  %   �           �t�bhhK ��h��R�(KK
��h�C(   ?   �        
      F         �t�bhhK ��h��R�(KK��h�C !      8     �           �t�bhhK ��h��R�(KK��h�CE      p      �t�bhhK ��h��R�(KK��h�C      0   o  �      �t�bhhK ��h��R�(KK��h�C    �
  �  �     �        �t�bhhK ��h��R�(KK
��h�C(#   !   ?      "   �      (        �t�bhhK ��h��R�(KK��h�Ch      �   :   �   S   Q               z   5         =  Z  y         0   4               �t�bhhK ��h��R�(KK��h�C=     	      	         �t�bhhK ��h��R�(KK��h�C01     �   Z  ?         .   
   &        �t�bhhK ��h��R�(KK ��h�C�      �   :      Y      Q         Q     Q      x              z         ;      y  ^        N  �        �t�bhhK ��h��R�(KK
��h�C(�      (  �	     )     N   >     �t�bhhK ��h��R�(KK��h�C<U        8   �  �  *      �        �  /         �t�bhhK ��h��R�(KK��h�ClN  �     �     K     �           ,   	      	   K   	   �   	     	   �   	   �  	   �     �t�bhhK ��h��R�(KK$��h�C�   0  J         U              �	        >   �   �     �  g  �  �  7   g      x     �     0  
   P     �  8        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C1   #          �t�bhhK ��h��R�(KK��h�CH]           %     3  �           -   �     8   �        �t�bhhK ��h��R�(KK��h�C R      r  	      	         �t�bhhK ��h��R�(KK&��h�C�   
      	      	      	   K   	   �   	   �   	   I  	   �  	   U  	   �  	   �   	   /  	     	   s  	   )  	   �  	   �  	   �     �t�bhhK ��h��R�(KK��h�CDV        >      �        �     [  �  Y               �t�bhhK ��h��R�(KK��h�C8      �           F     �  i      �        �t�bhhK ��h��R�(KK��h�Ct      ~  @   �     �t�bhhK ��h��R�(KK��h�Cx         .   c       "        .     �  �     �      R  9      >	        =  �     �  4         �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C@     1     \      �   ~        \      J  +         �t�bhhK ��h��R�(KK��h�C]   L        �t�bhhK ��h��R�(KK��h�C<�	                    �   [      !   �            �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C0      �  k            A  �   7         �t�bhhK ��h��R�(KK��h�C,-   @  �
  �   T  "   m      @        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�CD�  >      =      4      n     Y      �  �     D         �t�bhhK ��h��R�(KK��h�C<W      �  �  $                       �         �t�bhhK ��h��R�(KK��h�C8%      �  �  \   �   <      &   �     �        �t�bhhK ��h��R�(KK��h�CH   8   S              �   '  )                 �         �t�bhhK ��h��R�(KK��h�C\      )   )  +      �  �      }                   (   :   $   �   �        �t�bhhK ��h��R�(KK��h�C4  :         �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK��h�C@     �         �t�bhhK ��h��R�(KK��h�Cd      +                  ;     �  +      %   �  �                   �         �t�bhhK ��h��R�(KK	��h�C$l  E      �     �  	         �t�bhhK ��h��R�(KK��h�CP      =      �     �               O        p      �  O        �t�bhhK ��h��R�(KK��h�CH�  :   O        �
  �     ,            X        A   }      �t�bhhK ��h��R�(KK��h�C          	      	         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C �  �  ~  
   �   }          �t�bhhK ��h��R�(KK��h�C8`     ;     I   p        �     W  7         �t�bhhK ��h��R�(KK��h�C,T         �                        �t�bhhK ��h��R�(KK��h�C      '               �t�bhhK ��h��R�(KK	��h�C$  1  ?      
      F         �t�bhhK ��h��R�(KK��h�C      �     �     �t�bhhK ��h��R�(KK��h�CHw  �  (   #   !      ]   �   s     
   �  F         e        �t�bhhK ��h��R�(KK��h�C4   @   �                    �
  
         �t�bhhK ��h��R�(KK��h�C1   #       p     �     �t�bhhK ��h��R�(KK��h�CLT      `   U     $        8   X     8   �        �           �t�bhhK ��h��R�(KK��h�CT#   !      �  �  %   B   u  �     %  (      
   u          F         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK	��h�C$      )   R  �  
            �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C8�      (     |      s	     �        R        �t�bhhK ��h��R�(KK
��h�C(1   #      T  
   3   6            �t�bhhK ��h��R�(KK��h�C4      w   �        �  n      +   w         �t�bhhK ��h��R�(KK	��h�C$I  �     2        	         �t�bhhK ��h��R�(KK��h�C@     e  
   �     -      �  �   ^   �      �
        �t�bhhK ��h��R�(KK��h�CP     �   �  $   �      U     4  8   h  	              �         �t�bhhK ��h��R�(KK��h�CP                       P        �	        J   6     �	        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C4   r  '  L  "   �      (     "   <        �t�bhhK ��h��R�(KK��h�C�	  �           �t�bhhK ��h��R�(KK��h�CPW      v   
                 f  �            G        <        �t�bhhK ��h��R�(KK��h�C8      �  �  �      ,      A   �      n        �t�bhhK ��h��R�(KK��h�C\            P        �   r                    �   S  �       V        �t�bhhK ��h��R�(KK��h�Ch#   !      4      �            Z     v        0   4   (      
   �     �     F         �t�bhhK ��h��R�(KK��h�C V         "   >  �        �t�bhhK ��h��R�(KK��h�C   �  �      J  #     �t�bhhK ��h��R�(KK��h�C0E      4      �     �	     s   q         �t�bhhK ��h��R�(KK��h�C,         l  �     �     b        �t�bhhK ��h��R�(KK��h�CH      9   �   %  +      B   3     d  
   #     J   z         �t�bhhK ��h��R�(KK��h�C8�        �  �   �  �     =                  �t�bhhK ��h��R�(KK
��h�C(
   ,   Z     �     �           �t�bhhK ��h��R�(KK��h�C@*  I
     d   �     2     .            �   �         �t�bhhK ��h��R�(KK	��h�C$h         n  s         R     �t�bhhK ��h��R�(KK��h�C@   I   �        "     �  -   �   n     9            �t�bhhK ��h��R�(KK��h�C�  �      �t�bhhK ��h��R�(KK	��h�C$   �          �          �t�bhhK ��h��R�(KK��h�C1   #               �t�bhhK ��h��R�(KK��h�C0g  
   +           E  
   ,            �t�bhhK ��h��R�(KK	��h�C$2      4  �   ,   �      2      �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK��h�C      �    7   �     �t�bhhK ��h��R�(KK��h�C@      M  	      	      	   K   	     	   �   	   �     �t�bhhK ��h��R�(KK��h�C@         �           8            Z  �   s   7      �t�bhhK ��h��R�(KK��h�CT*      J   �   L          &      �   X                 $   k         �t�bhhK ��h��R�(KK��h�C�  �  �     �t�bhhK ��h��R�(KK��h�C4      P         �  
   }                 �t�bhhK ��h��R�(KK��h�CL           �  �        �      �     �           �         �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6   j        �t�bhhK ��h��R�(KK	��h�C$         2      �           �t�bhhK ��h��R�(KK��h�Ch        �      �      +   w            =               }	  /            l           �t�bhhK ��h��R�(KK��h�C             �t�bhhK ��h��R�(KK��h�C0  :   �  �	  �        :   �           �t�bhhK ��h��R�(KK	��h�C$     9   �       A        �t�bhhK ��h��R�(KK��h�C5                 �t�bhhK ��h��R�(KK��h�C �  &     T   E   ;        �t�bhhK ��h��R�(KK��h�CH      -   0   ;         �   �         �      �               �t�bhhK ��h��R�(KK��h�C -            1	  F
        �t�bhhK ��h��R�(KK��h�C8b   #      �         "   $   �   �              �t�bhhK ��h��R�(KK��h�Cl      �   :         Q      &   �      9   �   �      >      =            G      �   �        �t�bhhK ��h��R�(KK��h�C8�     �   �                                �t�bhhK ��h��R�(KK��h�CH         k         &      �   U   $   �   N     i           �t�bhhK ��h��R�(KK��h�C)                  �t�bhhK ��h��R�(KK��h�CG     |        �t�bhhK ��h��R�(KK��h�CH         E  �        =                 3  "           �t�bhhK ��h��R�(KK��h�C4�  $   �      $   �  s   �   y      l        �t�bhhK ��h��R�(KK��h�C,1   #   
   3   6   �
        &  r      �t�bhhK ��h��R�(KK��h�C89        i  �        �      i   
   )        �t�bhhK ��h��R�(KK
��h�C(     {         	      	         �t�bhhK ��h��R�(KK��h�C8"   �  v  �    �     p   �       u         �t�bhhK ��h��R�(KK
��h�C(              ^     �	        �t�bhhK ��h��R�(KK��h�C�     Q     �   p      �t�bhhK ��h��R�(KK��h�CT     N      .                                   4     A         �t�bhhK ��h��R�(KK��h�C   �         �t�bhhK ��h��R�(KK��h�CD   �   R      u      ~      �      A   �     �   p        �t�bhhK ��h��R�(KK��h�C<�
     
     �        �     ,   	      	         �t�bhhK ��h��R�(KK��h�C4
   1     �     �  :   A   ?              �t�bhhK ��h��R�(KK��h�C4b      >     ,   
   $   �   �              �t�bhhK ��h��R�(KK��h�C   v  	      	         �t�bhhK ��h��R�(KK��h�C               �t�bhhK ��h��R�(KK��h�CL�   L     r  �     L     u            F  C      f  �        �t�bhhK ��h��R�(KK��h�C@            �     �      V     v         �        �t�bhhK ��h��R�(KK��h�C<   >   �   a      L           5   L              �t�bhhK ��h��R�(KK��h�Cz   g   �   �         �t�bhhK ��h��R�(KK$��h�C��  `    �     C      \        �              A  �  �  
   _           �   %   H         h  %   
        �        �t�bhhK ��h��R�(KK��h�C0`      (      �       .   
   m        �t�bhhK ��h��R�(KK��h�CL   Y  
  �  �  :     
              �  y      �  f        �t�bhhK ��h��R�(KK��h�CD   ]   �   &      U   t           1     \   D   T        �t�bhhK ��h��R�(KK��h�C/     �t�bhhK ��h��R�(KK��h�C,*              U   �  
            �t�bhhK ��h��R�(KK
��h�C(b   #   "   $   �   �              �t�bhhK ��h��R�(KK��h�CT        H              ;      �     �      -  '     $           �t�bhhK ��h��R�(KK��h�C'            �t�bhhK ��h��R�(KK��h�C,�     �     z   "                �t�bhhK ��h��R�(KK��h�C8l         �   k      e      ;      �   R         �t�bhhK ��h��R�(KK��h�C8�  -  :   .        �  T      �  �   A        �t�bhhK ��h��R�(KK��h�C@1   #   
   3   �  7  �        L     �     r        �t�bhhK ��h��R�(KK��h�CT�         "     =                  !  �   �     G      �   	        �t�bhhK ��h��R�(KK	��h�C$]          �  �           �t�bhhK ��h��R�(KK
��h�C(*      L           0   j        �t�bhhK ��h��R�(KK��h�C<      N         �     �
  &      �   �   �        �t�bhhK ��h��R�(KK��h�C1   #          e  /      �t�bhhK ��h��R�(KK��h�CL               J  #           )   0   <   "   s
              �t�bhhK ��h��R�(KK��h�CT�      �        �  ]   
   �   �      �  o     Q        �           �t�bhhK ��h��R�(KK��h�C�     	      	         �t�bhhK ��h��R�(KK��h�C,T            P         d
          �t�bhhK ��h��R�(KK��h�C      k     �t�bhhK ��h��R�(KK��h�C\]     �   �  m     &   �         �  0      �   ~  j      �  $     t         �t�bhhK ��h��R�(KK��h�CL�  �  (     )        S   �  �        ;            �         �t�bhhK ��h��R�(KK��h�Cd   f   w     B  �   �        �     �  0              .              �        �t�bhhK ��h��R�(KK��h�CX      0   
                �   �         �  +  �      {   �   �
        �t�bhhK ��h��R�(KK��h�CT*              W  �     B     �
              .                  �t�bhhK ��h��R�(KK��h�CD   �  �  P     2      �	     �  T   �   ]              �t�bhhK ��h��R�(KK��h�Cp�        �   X  q
     �   
   �   B   }         .   9      �
           �   
   �  B   }         �t�bhhK ��h��R�(KK	��h�C$�      ,         �      M     �t�bhhK ��h��R�(KK��h�C4            �  b     (                  �t�bhhK ��h��R�(KK��h�C8   (   #   !   
   3   6   �
        &  r         �t�bhhK ��h��R�(KK	��h�C$�   �  >   �  Y  �  �        �t�bhhK ��h��R�(KK��h�C`      J   0      �     �     &      ;  +      G     *  <                    �t�bhhK ��h��R�(KK��h�C�           �         �t�bhhK ��h��R�(KK��h�CT         �  ^  �      �   +      B   �   9   �  T   H  <
  $   E         �t�be(hhK ��h��R�(KK��h�C8      }     E   
   &     #        W         �t�bhhK ��h��R�(KK��h�C !      �  	      	         �t�bhhK ��h��R�(KK��h�CL      5   #   !      t
     �     U   t      �     8   E        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C82   &   �      P     t   *   2                  �t�bhhK ��h��R�(KK��h�C   	  �      �        �t�bhhK ��h��R�(KK��h�Cl
   3   6   �     �      �     (      !      �         0   x   "   m      �        @        �t�bhhK ��h��R�(KK��h�C �   
      	      	         �t�bhhK ��h��R�(KK	��h�C$�     n   O        �        �t�bhhK ��h��R�(KK	��h�C$�        E     �           �t�bhhK ��h��R�(KK��h�CL         E  �                          �  �   �         �t�bhhK ��h��R�(KK��h�C �     r  	      	         �t�bhhK ��h��R�(KK��h�C,�         (   w   �  �   �   d        �t�bhhK ��h��R�(KK��h�C@2   �  �  �   �   �  D   �            �   �  '        �t�bhhK ��h��R�(KK��h�C8�     "   >  �  �          
      �        �t�bhhK ��h��R�(KK	��h�C$!         
   A   �  
   &     �t�bhhK ��h��R�(KK	��h�C$�        �  i   h          �t�bhhK ��h��R�(KK��h�C0              �
  �   �
  )            �t�bhhK ��h��R�(KK��h�C0   	      	      	   K   	   �   	   U     �t�bhhK ��h��R�(KK��h�C0   0      �  
          �           �t�bhhK ��h��R�(KK
��h�C("   �  (      !      B   J        �t�bhhK ��h��R�(KK	��h�C$�        +   -   
            �t�bhhK ��h��R�(KK��h�C,|           &   0     �	           �t�bhhK ��h��R�(KK��h�C*     �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C0   �     �      (  �  -      B        �t�bhhK ��h��R�(KK��h�C0%      �  �              A            �t�bhhK ��h��R�(KK��h�C!         	         �t�bhhK ��h��R�(KK��h�C<�     �   �  
   �                 �   �        �t�bhhK ��h��R�(KK��h�C�      u      �t�bhhK ��h��R�(KK��h�C4           �t�bhhK ��h��R�(KK��h�C      �  �        �t�bhhK ��h��R�(KK��h�CT      ,  �     �       �  |      �            0      �          �t�bhhK ��h��R�(KK��h�CD           0  %   h  �        (                    �t�bhhK ��h��R�(KK	��h�C$6  �  �  8     H  @         �t�bhhK ��h��R�(KK��h�CD         9     7            b   x         
   O        �t�bhhK ��h��R�(KK��h�C8   X   '   �  �	       %   f     g  �	        �t�bhhK ��h��R�(KK��h�C,   �                 R           �t�bhhK ��h��R�(KK��h�C8_  +   ,      <      �	  	      	   �  	   �      �t�bhhK ��h��R�(KK��h�C<q   �                 %  �                   �t�bhhK ��h��R�(KK
��h�C(!            �  	      	         �t�bhhK ��h��R�(KK��h�C,3  �     �  +         �  {        �t�bhhK ��h��R�(KK��h�CP�   �   �   I        %   �     �   �      /   9   �   7      V        �t�bhhK ��h��R�(KK��h�Cd.     N      .               R      Q        a
        B   
           �        �t�bhhK ��h��R�(KK��h�CD            �     �    (   �     �  +   
            �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6            �t�bhhK ��h��R�(KK��h�C,f  =           b	          �
     �t�bhhK ��h��R�(KK��h�CT      �      �  :   �        �     `           V  �             �t�bhhK ��h��R�(KK��h�CH�        .   �      �  �
     �     n      �      �        �t�bhhK ��h��R�(KK��h�C<   >        �      |      �   y      �  �         �t�bhhK ��h��R�(KK��h�C 1   #       {     �        �t�bhhK ��h��R�(KK��h�C4   .   :     0     �	    )      M        �t�bhhK ��h��R�(KK��h�C4�  �   {     �  7      W  
      �         �t�bhhK ��h��R�(KK��h�Cd"   e        �  #	        2      .   �  �     |     F	  �     }     B
  q        �t�bhhK ��h��R�(KK��h�CX2      w        <   G   v     �            �         �        �        �t�bhhK ��h��R�(KK��h�CH   	      	      	   K   	   �   	     	   �  	   �   	   �     �t�bhhK ��h��R�(KK��h�CX�     	                �   B        �         g     
               �t�bhhK ��h��R�(KK��h�C<I  �                 �  
     �      �        �t�bhhK ��h��R�(KK��h�C	     �      �         �t�bhhK ��h��R�(KK	��h�C$H   ?        �              �t�bhhK ��h��R�(KK
��h�C(!           �  	      	         �t�bhhK ��h��R�(KK��h�C`           �      �      W   &      �   �   $   E      �      W   y   t  l        �t�bhhK ��h��R�(KK��h�C@                                �   
   c        �t�bhhK ��h��R�(KK��h�CD%   >  �        �     @     I        J   �  �
        �t�bhhK ��h��R�(KK��h�C<   �      �        d   �      (   D   �  �         �t�bhhK ��h��R�(KK��h�C0         -  c     $   |     A         �t�bhhK ��h��R�(KK��h�C     
   �     �t�bhhK ��h��R�(KK��h�Cp�  a  C   �           $  �     �     Y	        �  %   �      �      -     �     �         �t�bhhK ��h��R�(KK��h�C 6        3      ]         �t�bhhK ��h��R�(KK��h�C<:     )   N   �     C	     �   "        �        �t�bhhK ��h��R�(KK��h�CH  N        �     �t�bhhK ��h��R�(KK��h�CX*      �   #
     8   �            �      z     �   �         �   �        �t�bhhK ��h��R�(KK��h�C b      >  �   "   �        �t�bhhK ��h��R�(KK
��h�C(*   �  {  �	           �         �t�bhhK ��h��R�(KK
��h�C(-   `   3  �      �
              �t�bhhK ��h��R�(KK��h�C`@     �     �  �  �     �   �  �           $     5   <           �        �t�bh�      hK ��h��R�(KK��h�C0i  �   "   >  �      +      `   /         �t�bhhK ��h��R�(KK��h�C@      )   �   �   e     �   T   >      w     �        �t�bhhK ��h��R�(KK��h�C1   #       �        �t�bhhK ��h��R�(KK��h�CD   �   R      u      ~      �      A   �     �   p        �t�bhhK ��h��R�(KK��h�CX�   �	     E         �  +  �   �         
     n   �        a  L         �t�bhhK ��h��R�(KK��h�CP      �     �      p	  S  %   A   T     d  
                     �t�bhhK ��h��R�(KK��h�C8     m  
   _      C                      �t�bhhK ��h��R�(KK��h�C<   "   �     �  -      *     �  c      �         �t�bhhK ��h��R�(KK��h�C       �         �	        �t�bhhK ��h��R�(KK��h�C             �            �t�bhhK ��h��R�(KK��h�CPp        C      �   �      �      �           �     U           �t�bhhK ��h��R�(KK��h�C\   
  -  C   
        �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6   N	        �t�bhhK ��h��R�(KK
��h�C(      �     7   v     �        �t�bhhK ��h��R�(KK��h�CQ          M        �t�bhhK ��h��R�(KK��h�C8�        J        v   �     %     �        �t�bhhK ��h��R�(KK��h�C1   #       �     �t�bhhK ��h��R�(KK��h�CP*      �      4   >      a      +      �        D  �  $   0        �t�bhhK ��h��R�(KK��h�CP�       0  `     �                 J    
   _              �t�bhhK ��h��R�(KK��h�C         h     �   �     �t�bhhK ��h��R�(KK��h�Cj        	         �t�bhhK ��h��R�(KK��h�C3   F               �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C�   E  	         �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   �  �             �t�bhhK ��h��R�(KK
��h�C(%  +            �  �           �t�bhhK ��h��R�(KK��h�C=         �t�bhhK ��h��R�(KK	��h�C$Z         �  )   
            �t�bhhK ��h��R�(KK��h�C,      �   z   ,      �   Y  �        �t�bhhK ��h��R�(KK��h�C1   #       j     �t�bhhK ��h��R�(KK	��h�C$     �   
                 �t�bhhK ��h��R�(KK��h�CT   X   �     "      g  �  �           �         -  T     X         �t�bhhK ��h��R�(KK��h�C0V         )         �   �      a        �t�bhhK ��h��R�(KK��h�C,               �     �  p        �t�bhhK ��h��R�(KK��h�CD         �               �     >      v      �        �t�bhhK ��h��R�(KK��h�C8*      (      �  (      �     �   �  �        �t�bhhK ��h��R�(KK#��h�C�      5   �  �         .         �  c         ]           ;      �  0   �   
   �  "      W          W  �        �t�bhhK ��h��R�(KK��h�Cp     �     �t�bhhK ��h��R�(KK��h�C0�  �      �  �  {  �   y      l        �t�bhhK ��h��R�(KK��h�C�     v  �     �     �t�bhhK ��h��R�(KK��h�C41   #         
   3   6   �  g  �   �        �t�bhhK ��h��R�(KK��h�C8      �     .   �     q     �     �        �t�bhhK ��h��R�(KK��h�C@�      �  !            V  �      O     9           �t�bhhK ��h��R�(KK��h�Cp                     �   ]  �      �      7   &      -   F  +           t      �           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C      �      �t�bhhK ��h��R�(KK��h�C89      �     �     �  �      �  h   �        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C@�      &	     �     �   S  )   �         �           �t�bhhK ��h��R�(KK��h�C               �t�bhhK ��h��R�(KK��h�C0B           �   �        c  p         �t�bhhK ��h��R�(KK��h�C,   ?   !      �   
   3   6   �	        �t�bhhK ��h��R�(KK��h�C_     �         �t�bhhK ��h��R�(KK��h�C<�   o  7        �         9     7      /         �t�bhhK ��h��R�(KK��h�C    �  �  m              �t�bhhK ��h��R�(KK��h�C`            �                 �         �   �         �   �  $   2  Y        �t�bhhK ��h��R�(KK��h�C   =  �  9     �t�bhhK ��h��R�(KK$��h�C�                                    �      �          7      O  �     �      �     y           7   �           �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�C\      	  8   /   '        2       �   �         V         A  A   �        �t�bhhK ��h��R�(KK��h�C\      P         C  E   )         �            �     �        J  E         �t�bhhK ��h��R�(KK��h�CH�  d  �                    >                 �         �t�bhhK ��h��R�(KK��h�C<      )  +   e  ^   �     �  
   |      �         �t�bhhK ��h��R�(KK��h�CT      ;      �      �     o      z            �  |     ,   O         �t�bhhK ��h��R�(KK��h�CP      �      �   �     �     �     �                        �t�bhhK ��h��R�(KK��h�CD   @	  �
     .      u  �  
               <        �t�bhhK ��h��R�(KK	��h�C$      �     "     ?	        �t�bhhK ��h��R�(KK��h�C^  |      �     �t�bhhK ��h��R�(KK��h�C0%   �  �          A      �  �         �t�bhhK ��h��R�(KK��h�C         	      	         �t�bhhK ��h��R�(KK��h�Ck  7   R        �t�bhhK ��h��R�(KK��h�C0  g     1     B      	      	         �t�bhhK ��h��R�(KK��h�C0  (   �  �           2     �         �t�bhhK ��h��R�(KK��h�C 9  �     �   S   X        �t�bhhK ��h��R�(KK��h�C   >   a   Q           �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C1   #       m      �     �t�bhhK ��h��R�(KK��h�C1   -   3   6          �t�bhhK ��h��R�(KK��h�CX'     �              %   h    z     N  �     %                     �t�bhhK ��h��R�(KK��h�C<�     R         .   �             y           �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C �        %               �t�bhhK ��h��R�(KK��h�C[           �      �t�bhhK ��h��R�(KK��h�C0   2            2   0   �  �   �        �t�bhhK ��h��R�(KK
��h�C(!      x         	      	         �t�bhhK ��h��R�(KK��h�CT%   �   �     �   E     �  :   �  d  2   %   E     �  ~              �t�bhhK ��h��R�(KK��h�C\      �         �     5                  �         "   e      @   �         �t�bhhK ��h��R�(KK
��h�C(v   �                t        �t�bhhK ��h��R�(KK��h�CL      �        5   !      G     S        U   $   �   N        �t�bhhK ��h��R�(KK��h�C0           D        �               �t�bhhK ��h��R�(KK	��h�C$   �	     -   N   !  �        �t�bhhK ��h��R�(KK��h�C4�          .                           �t�bhhK ��h��R�(KK��h�C4�   �   w       �   +   !      �   R         �t�bhhK ��h��R�(KK��h�C<      �  �     �     x	     P     %   w	        �t�bhhK ��h��R�(KK��h�CL      �  
   X   �         X   �        �     
   �  �        �t�bhhK ��h��R�(KK��h�C   D     l  �      �t�bhhK ��h��R�(KK��h�C0      C     �  "     '  O  7         �t�bhhK ��h��R�(KK��h�C<k     �  �   �      �  
   �     ^   F  F         �t�bhhK ��h��R�(KK��h�C@      J   �  L         Z  &      M   �               �t�bhhK ��h��R�(KK��h�Cm      �      �t�bhhK ��h��R�(KK��h�C�  :   M     �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C   :   n     �t�bhhK ��h��R�(KK��h�C!         I  	         �t�bhhK ��h��R�(KK��h�Ct   5   �   �      ;     \              
           �               �  !  +      8            �t�bhhK ��h��R�(KK��h�C%   �  O     �t�bhhK ��h��R�(KK��h�C             �t�bhhK ��h��R�(KK��h�C      �  	         �t�bhhK ��h��R�(KK
��h�C(�         ;      2              �t�bhhK ��h��R�(KK��h�C �
              �         �t�bhhK ��h��R�(KK��h�C`M      +   �     %   5     v     E   *      �  �   $   E   "         �  �        �t�bhhK ��h��R�(KK	��h�C$               J  +         �t�bhhK ��h��R�(KK��h�C d        �              �t�bhhK ��h��R�(KK��h�C<-      %   A         @   �         /      �         �t�bhhK ��h��R�(KK��h�CH      5   �  �   
   `
           U   T   �     �           �t�bhhK ��h��R�(KK��h�C   (             �t�bhhK ��h��R�(KK��h�CD
   3   6   �     X   ?      !      �     /      X         �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CT         $   �  �   �     �              =      �   �   q   7        �t�bhhK ��h��R�(KK��h�Cd
         2               S         �  �   �     �     
     �                  �t�bhhK ��h��R�(KK��h�CT   �   �  b     ,        -   U   �     �        p
                 �t�bhhK ��h��R�(KK��h�C8�   �        �      
  X  �	  	      	         �t�bhhK ��h��R�(KK��h�CL  ^  -  �        �      X                                �t�bhhK ��h��R�(KK��h�C*                  �t�bhhK ��h��R�(KK��h�C8/               w               
   �
        �t�bhhK ��h��R�(KK��h�C8   H   ?  �  �   �  �            �   \        �t�bhhK ��h��R�(KK��h�C b   #   G   $   �   �        �t�bhhK ��h��R�(KK��h�C0#   !   ?      
   3   6   �             �t�bhhK ��h��R�(KK��h�C`�     -   l                 �   f  a   ;      �  :   W      b   #   G   W         �t�bhhK ��h��R�(KK��h�CT                  �  �     (   �           =      @  G   W         �t�bhhK ��h��R�(KK��h�C    e   '   -   �   �        �t�bhhK ��h��R�(KK��h�C       5  	      	         �t�bhhK ��h��R�(KK��h�CD`   �     0      n   �     8   5
     `   6
     b        �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C0B  �                  
  ;           �t�bhhK ��h��R�(KK
��h�C(      I  ,                     �t�bhhK ��h��R�(KK��h�C4�              ,     �        �        �t�bhhK ��h��R�(KK��h�C08  4
     8   o   S  y      |  �        �t�bhhK ��h��R�(KK��h�C<         ;      Q        =      Q  G   W         �t�bhhK ��h��R�(KK��h�Cl         �	     �         .           `   �        ]   �	     �        0   o  �         �t�bhhK ��h��R�(KK��h�Cp�  �   )   �      �   B   }         S   ,                  /     �      K      I     �        �t�bhhK ��h��R�(KK��h�C:          �t�bhhK ��h��R�(KK��h�C8[  �  5     �  �   !      D         K        �t�bhhK ��h��R�(KK��h�C4   �  �   �     �      P        �         �t�bhhK ��h��R�(KK��h�C    	      	      	   K      �t�bhhK ��h��R�(KK��h�C{  b     �t�bhhK ��h��R�(KK��h�C           �t�bhhK ��h��R�(KK��h�CP      �   �         9      /            0   �        :           �t�bhhK ��h��R�(KK��h�CL      �  �  
        W  �     �  B  8   �        t        �t�bhhK ��h��R�(KK	��h�C$%   �     )      �  �         �t�bhhK ��h��R�(KK��h�C8   i  #     /   9     7         �     s     �t�bhhK ��h��R�(KK��h�C,�   h  �  �  �  �      A   !        �t�bhhK ��h��R�(KK��h�C4
     (      1        �  F     �        �t�bhhK ��h��R�(KK��h�C,l   9     7   &   a   �      �        �t�bhhK ��h��R�(KK��h�Cl*      �  �      �  [        .   "   �      (     ~  �  �              �   6	  �         �t�bhhK ��h��R�(KK��h�C0'  �  
   ,            K               �t�bhhK ��h��R�(KK ��h�C�            �                     f   w  �  a   ;      w  {          �   �         �     ,  ]        �t�bhhK ��h��R�(KK��h�C8f   �  �  �  '  G   %   /           �        �t�bhhK ��h��R�(KK
��h�C(�        :   �  	      	         �t�bhhK ��h��R�(KK��h�CH      �
        �           S                 �
        �t�bhhK ��h��R�(KK��h�C �     �        �         �t�bhhK ��h��R�(KK
��h�C(I      *     �  "      ]        �t�bhhK ��h��R�(KK��h�C         �     �t�bhhK ��h��R�(KK��h�C8     '   �     5     �   5     �   �        �t�bhhK ��h��R�(KK ��h�C�   $   �  �   �  �   8  �   �     �  H     �     �  �      M    
     �         �   �  W              �t�bhhK ��h��R�(KK��h�C0�        "   >  U   �                 �t�bhhK ��h��R�(KK��h�C0�     �     �  �   *      �  �        �t�bhhK ��h��R�(KK��h�CP   &      �         �  E     V   �     �             �        �t�bhhK ��h��R�(KK��h�CD�   �  �  �
  w     |                             �t�bhhK ��h��R�(KK	��h�C$            �      �        �t�bhhK ��h��R�(KK��h�CD   X   '   �   �     �   9     �  �     /      �         �t�bhhK ��h��R�(KK��h�C "   �        �   p        �t�bhhK ��h��R�(KK��h�C�     �     I         �t�bhhK ��h��R�(KK��h�C8�  J  �            /   9     7               �t�bhhK ��h��R�(KK��h�CD      �                    �  &                    �t�bhhK ��h��R�(KK��h�CD@   �   �      u      @      �     �  I   u      T        �t�bhhK ��h��R�(KK��h�C4/         �      
  X  �	  	      	         �t�bhhK ��h��R�(KK��h�CX      J   6     �	     e         P        �	          �     :        �t�bhhK ��h��R�(KK��h�C0K  �   �     �  c           C         �t�bhhK ��h��R�(KK��h�Ch*      t  5      <      	     �  �     %     '      �     0   [           <        �t�bhhK ��h��R�(KK��h�CL      P         c  c        J   �      �   "   T     �         �t�bhhK ��h��R�(KK��h�CT      J   =      �     @      e      X      &      �   �     U
        �t�bhhK ��h��R�(KK��h�CT      '   )   H   �     �   �         �     �           I           �t�bhhK ��h��R�(KK��h�C`%   �     �   �     v           ;      �               8   �   �               �t�bhhK ��h��R�(KK��h�C8      H  %           `        B            �t�bhhK ��h��R�(KK��h�C8^            �  �      s     ?     4        �t�bhhK ��h��R�(KK��h�C4o  (      �  c   �   D      �  s   7         �t�bhhK ��h��R�(KK��h�C    �   
        �        �t�bhhK ��h��R�(KK��h�CH      5   <      �      -     �             U            �t�bhhK ��h��R�(KK��h�C4B  �  "         V      J      �  �         �t�bhhK ��h��R�(KK��h�CX�   �          �      �          �  �    �	  �
     &              �t�bhhK ��h��R�(KK��h�Cd�        }        	      	      	   K   	   �   	   �   	     	   �  	   U  	   �      �t�bhhK ��h��R�(KK��h�CL            �  �  �  :   �   �   �          $   �           �t�bhhK ��h��R�(KK��h�C�      �	  	         �t�bhhK ��h��R�(KK��h�C�
     !      �t�bhhK ��h��R�(KK
��h�C(
   �  F   '   �   !      4         �t�bhhK ��h��R�(KK��h�C,   e   �   �           e           �t�bhhK ��h��R�(KK��h�C     M     �      �t�bhhK ��h��R�(KK��h�C      �     �t�bhhK ��h��R�(KK
��h�C(c     |  �      q             �t�bhhK ��h��R�(KK��h�CX      l  �  *        �                 .                           �t�bhhK ��h��R�(KK��h�C      �     7   v     �t�bhhK ��h��R�(KK��h�C\
   T  '   !      %   w  T      �  a   ;         �   �     |  C   
   �         �t�bhhK ��h��R�(KK��h�CXS   3  V   8   �   �              O         Y      Q         
  Q         �t�bhhK ��h��R�(KK��h�C   V           �t�bhhK ��h��R�(KK��h�C[   9        �t�bhhK ��h��R�(KK��h�C<   �        �  
   �     U   �     8           �t�bhhK ��h��R�(KK��h�C0�      M  	      	   K   	     	   �      �t�bhhK ��h��R�(KK��h�CT
      F         P   �
  �   �   
         ,      *    �     �        �t�bhhK ��h��R�(KK��h�C<!      �      -     	      	      	   K   	   �      �t�bhhK ��h��R�(KK��h�C46  �   
   T        %  +      l	  F         �t�bhhK ��h��R�(KK��h�C 1     �  	      	         �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK
��h�C(         p        �           �t�bhhK ��h��R�(KK��h�CH      4      -   �     %   �  
     B  o     
  $        �t�bhhK ��h��R�(KK��h�C0   �  �            �  �     $   �     �t�bhhK ��h��R�(KK��h�CT     �  1     x         �   �                 �      $          �t�bhhK ��h��R�(KK��h�C -         �     k        �t�bhhK ��h��R�(KK��h�C`                #          &      U      "      y                       �t�bhhK ��h��R�(KK��h�C1   #       �          �t�bhhK ��h��R�(KK��h�C   �    �          �t�bhhK ��h��R�(KK��h�C8   e   '   H   B   j        .         �        �t�bhhK ��h��R�(KK��h�C�  �  �         �t�bhhK ��h��R�(KK��h�C8"   m      $  /      -  �      .   /  i        �t�bhhK ��h��R�(KK��h�CP�      �         .      v   c      �    i   #     �     �        �t�bhhK ��h��R�(KK��h�CH�      &  J  �   �   u         �      �        �   �         �t�bhhK ��h��R�(KK��h�C�  (      "   2        �t�bhhK ��h��R�(KK��h�C   �  �                �t�bhhK ��h��R�(KK��h�C,         {         	      	         �t�bhhK ��h��R�(KK��h�C                   �t�bhhK ��h��R�(KK��h�C@g  
   g           E  
   ,                  B     �t�bhhK ��h��R�(KK��h�C@�         ]  �     �      �	     �   4	     �        �t�bhhK ��h��R�(KK��h�CH]      �            A   �           �        (   Q        �t�bhhK ��h��R�(KK��h�C 1     |         	         �t�bhhK ��h��R�(KK��h�C    =      �    	         �t�bhhK ��h��R�(KK��h�Ci  n      �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�CD~        �	     �              
   A     e           �t�bhhK ��h��R�(KK��h�C �     .   
   8   �        �t�bhhK ��h��R�(KK��h�C�     [     �t�bhhK ��h��R�(KK��h�C               �t�bhhK ��h��R�(KK#��h�C�2      0   �  �   g         �  �                       J   �  g            �     �     �   �  �  9      7         �t�bhhK ��h��R�(KK��h�C|      <  R      �t�bhhK ��h��R�(KK
��h�C(               �              �t�bhhK ��h��R�(KK��h�CP
   f   �     2   i  F        2      �   
         �
     �        �t�bhhK ��h��R�(KK��h�C    
      	      	         �t�bhhK ��h��R�(KK	��h�C$�  ;                       �t�bhhK ��h��R�(KK��h�C�  E      �   �        �t�bhhK ��h��R�(KK
��h�C(        @            4        �t�bhhK ��h��R�(KK��h�C<   �      �  "      �        V         �        �t�bhhK ��h��R�(KK	��h�C$
     L   *         P         �t�bhhK ��h��R�(KK��h�C<;      �           �     �           S   Q      �t�bhhK ��h��R�(KK��h�C�  �      S        �t�bhhK ��h��R�(KK��h�C         .            �t�bhhK ��h��R�(KK)��h�C��              t  b     �         u  �                    �         m   9   �        �         �  �     "   >        �  �         �t�bhhK ��h��R�(KK��h�C8�   '         �     p     	        �         �t�bhhK ��h��R�(KK��h�C,   y	  L  �   >   )   y	  N            �t�bhhK ��h��R�(KK��h�C@�       �     �  �  �     ?          �        �t�bhhK ��h��R�(KK��h�CL   S  5         �  u  V   8   �   �     �           Z        �t�bhhK ��h��R�(KK��h�C
     '   H            �t�bhhK ��h��R�(KK
��h�C(      �              �        �t�bhhK ��h��R�(KK��h�C�     �   '   "         �t�bhhK ��h��R�(KK��h�CH      )   =         ~        "   t      2  
   $   �        �t�bhhK ��h��R�(KK��h�C`�     *     @            .      X      e                 �  i      @         �t�bhhK ��h��R�(KK��h�C      *
  r      �t�bhhK ��h��R�(KK��h�C,      )   0              �
        �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C�  
   ,             �t�bhhK ��h��R�(KK��h�C0�      �  /     =         "   W         �t�bhhK ��h��R�(KK��h�C!      �
  �  	   K      �t�bhhK ��h��R�(KK��h�C8�  +            t       �   7  
            �t�bhhK ��h��R�(KK��h�C t      ~     �     @      �t�bhhK ��h��R�(KK��h�C   �   �  �          �t�bhhK ��h��R�(KK��h�C,�   �   >   2   �  K  A     �        �t�bhhK ��h��R�(KK��h�C`9   �  (   2   �      �   9   %   s   �           "        9   s   �  g   �        �t�bhhK ��h��R�(KK��h�Cd�  �  �      .                                    %   R            �        �t�bhhK ��h��R�(KK��h�C<�	        m      �      0   <   ^   �   �  P        �t�bhhK ��h��R�(KK��h�C,                 �     F
        �t�bhhK ��h��R�(KK��h�C�  �     �  �     �t�bhhK ��h��R�(KK��h�C      �     �t�bhhK ��h��R�(KK
��h�C(�   �           �   �            �t�bhhK ��h��R�(KK��h�Cx�                 4      �  
        �     �                  �     .   �      �  8   4         �t�bhhK ��h��R�(KK��h�CT      $        �      T   $   �                 J   b      x         �t�bhhK ��h��R�(KK
��h�C(D  �   �      �         &        �t�bhhK ��h��R�(KK��h�C`%        	      	      	   �   	   �   	   I  	   �  	   /  	   s  	   )  	   �     �t�bhhK ��h��R�(KK��h�C\Y  3        �                       �   %         $  
   3  >            �t�bhhK ��h��R�(KK��h�CX�     �  	      	      	   K   	   �   	   �   	     	   I  	   U  	   �      �t�bhhK ��h��R�(KK��h�C8  >   A  )        �  �   �  h   �   �         �t�bhhK ��h��R�(KK��h�C    �  R  \   �  -        �t�bhhK ��h��R�(KK��h�C<      !  �     �t�bhhK ��h��R�(KK��h�C0_  #      �  R   
   3   6      �         �t�bhhK ��h��R�(KK��h�C0�   :   &
     =               r
        �t�bhhK ��h��R�(KK��h�C�  B  �  �         �t�bhhK ��h��R�(KK��h�CP      }     E   
   &     �        W   �   s     \  �   c	        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C �
        	      	         �t�bhhK ��h��R�(KK��h�C@      '   �        .                 &   a         �t�bhhK ��h��R�(KK
��h�C(   �  )         H   l  �         �t�bhhK ��h��R�(KK��h�C0M   �      �              $   k         �t�bhhK ��h��R�(KK��h�C4   5     �             ;   j          �t�bhhK ��h��R�(KK��h�Cd   f   �   �   W      .   [     �     f   ?  )   T            u     �      7         �t�bhhK ��h��R�(KK
��h�C(1   #      �  
   3   6   �        �t�bhhK ��h��R�(KK	��h�C$1   #   
   3   6   	  �         �t�bhhK ��h��R�(KK��h�Cl                     �   (      �   ;      �   �  9   $   2     )   *   $   2     X
        �t�bhhK ��h��R�(KK��h�C         	         �t�bhhK ��h��R�(KK��h�Cj  g       �t�bhhK ��h��R�(KK��h�C4  8         t   *      �  +              �t�bhhK ��h��R�(KK��h�CL�   n     7  �
        �        7  �	     �                  �t�bhhK ��h��R�(KK��h�C      /      a     �t�bhhK ��h��R�(KK��h�C�  F      �t�bhhK ��h��R�(KK��h�C<   <                  .   +
  H      
   y        �t�bhhK ��h��R�(KK
��h�C(      a  m  �      �            �t�bhhK ��h��R�(KK��h�C   "     n      �t�bhhK ��h��R�(KK��h�C4         m      -  �
        U            �t�bhhK ��h��R�(KK��h�Cd      b   x   
   �   )   
   y  �      }                (      �   �     s        �t�bhhK ��h��R�(KK��h�C�  �      �t�bhhK ��h��R�(KK��h�C,�  �   +   <      [         w        �t�bhhK ��h��R�(KK��h�C<�  �  (  G   t      �        �     �           �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C4"   �     T   D   �           C           �t�bhhK ��h��R�(KK��h�C�     	      	         �t�bhhK ��h��R�(KK��h�C4      )  8   /                          �t�bhhK ��h��R�(KK
��h�C(  �      S   H  �              �t�bhhK ��h��R�(KK��h�C@                    )   U   @     �     e         �t�bhhK ��h��R�(KK��h�CL   �   J   a        �   &   �   �  �      P     G     t         �t�bhhK ��h��R�(KK��h�C\   ?   �      �  r      �t�bhhK ��h��R�(KK��h�C1   #       ,        �t�bhhK ��h��R�(KK��h�C 1   #     �   �            �t�bhhK ��h��R�(KK��h�C8T   ,     �  _     (   
   �    �          �t�bhhK ��h��R�(KK��h�C8      �  �   *   2      V  �                �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�CD-      @   '           `  V   2      z   h   H   �        �t�bhhK ��h��R�(KK��h�CT   �              �           %         v     �  �     ,         �t�bhhK ��h��R�(KK��h�C0                           �         �t�bhhK ��h��R�(KK��h�Cl      \  |      �               )  +      �  
   y              O      �   S   Q         �t�bhhK ��h��R�(KK%��h�C�         O      �   Q           Y                  �      5      e     4      �         4      m        4      �        �t�bhhK ��h��R�(KK��h�C        �      r      �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK
��h�C(>     �        �      I         �t�bhhK ��h��R�(KK��h�C    >   w   �  K  �        �t�bhhK ��h��R�(KK
��h�C(�   �  >      K  A     �        �t�bhhK ��h��R�(KK	��h�C$
       d   �      
        �t�bhhK ��h��R�(KK��h�C<�  (      L            N        �     N        �t�bhhK ��h��R�(KK��h�C8      )  +      �	  �   �   �      ^           �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C{     �t�bhhK ��h��R�(KK��h�Cf     g  /     �t�bhhK ��h��R�(KK��h�C     �        �     �t�bhhK ��h��R�(KK��h�CM     �t�bhhK ��h��R�(KK��h�CXP        L     �   P     L     %     �       �                    �t�bhhK ��h��R�(KK��h�C07     �     �        @              �t�bhhK ��h��R�(KK��h�CX
  $   |  �      �      \   �         v      "              0            �t�bhhK ��h��R�(KK
��h�C(   �     �  +      �  n         �t�bhhK ��h��R�(KK��h�C,1   #       [      �      /      V     �t�bhhK ��h��R�(KK��h�C #   !   '   
      F         �t�bhhK ��h��R�(KK��h�C8   �        �  -   �      P   H              �t�bhhK ��h��R�(KK
��h�C(]     
   %  x     ~            �t�bhhK ��h��R�(KK��h�C<                 �   �  7      �     �         �t�bhhK ��h��R�(KK��h�C`      �   �  A     �  �         �      �  �  �     �  g            �        �t�bhhK ��h��R�(KK��h�CX"   m      @     �   (   2   )   <      C  "   X   (     g                 �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C0:        �   �  
      �     �        �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�CT�  �   �	  �              /   9     7      )      %      ~   �         �t�bhhK ��h��R�(KK��h�Cd"   t      �     
   $   �            M     
            ;         k               �t�bhhK ��h��R�(KK��h�C1   #               �t�bhhK ��h��R�(KK��h�C4!      1     n   ?      
   3   6           �t�bhhK ��h��R�(KK��h�C       �     �   �        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK
��h�C(      A    �                  �t�bhhK ��h��R�(KK��h�C<   	     �t�bhhK ��h��R�(KK'��h�C�      =      |
                �   �                             S   �     Q     Q      x           _  �      "           �t�bhhK ��h��R�(KK��h�C@   I   o      l      �   <      �  �      .           �t�bhhK ��h��R�(KK��h�Cn      ]     �t�bhhK ��h��R�(KK	��h�C$   �     �      .            �t�bhhK ��h��R�(KK��h�CT
   3   6   �     /   �        '   #   !      8  O  /   �              �t�bhhK ��h��R�(KK��h�C81   #               
   3   6                  �t�bhhK ��h��R�(KK��h�Cd   �  	      	         �t�bhhK ��h��R�(KK��h�CT
     ?         *      �  "  n  o  "     u  �         p           �t�bhhK ��h��R�(KK��h�C  �   �      �t�bhhK ��h��R�(KK��h�C0      @                    :
        �t�bhhK ��h��R�(KK
��h�C(      �   L   
     �   �         �t�bhhK ��h��R�(KK��h�CT   (   �   j        �  �  V   �     �      �     
        �        �t�bhhK ��h��R�(KK��h�C<3   6     �           �  !                     �t�bhhK ��h��R�(KK��h�C         q            �t�bhhK ��h��R�(KK��h�C4   �   �  �  I      �   ~      �   n         �t�bhhK ��h��R�(KK��h�C4%   N
  �  [            %   c     �        �t�bhhK ��h��R�(KK
��h�C(`     �	  �            �
        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C\   '   )        �        �           [      9         |                 �t�bhhK ��h��R�(KK��h�CL      a                 3
     �
     %      a  j   �        �t�bhhK ��h��R�(KK��h�C9     �t�bhhK ��h��R�(KK��h�CO  7      �t�bhhK ��h��R�(KK��h�Cn     %        �t�bhhK ��h��R�(KK
��h�C(      1	  2	                  �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C,   &   �  �   �   $   E      e         �t�bhhK ��h��R�(KK��h�C�  N        ?     �t�bhhK ��h��R�(KK��h�C �     E      �   *        �t�bhhK ��h��R�(KK��h�C[      �  	         �t�bhhK ��h��R�(KK	��h�C$�   !      9  	      	         �t�bhhK ��h��R�(KK��h�CX   $   k                  �      )   h   %   �  .        .   
           �t�bhhK ��h��R�(KK��h�C 3   F   h     @   �         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CR      m     �      �t�bhhK ��h��R�(KK��h�C�            �t�bhhK ��h��R�(KK��h�C<   �        
   ]        �  �        U	        �t�bhhK ��h��R�(KK��h�C,      '   H   �                   �t�bhhK ��h��R�(KK��h�CH      \  �  j   �     �      O           �      L         �t�bhhK ��h��R�(KK��h�CT   �      A      ,     C   w      �  �     C   w      %   �   $        �t�bhhK ��h��R�(KK��h�C,              \
        0
        �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C0
      ]  T  '   !      .     �         �t�bhhK ��h��R�(KK��h�C�   
          �	     �t�bhhK ��h��R�(KK��h�C<   X   �   �     .   "   X   E	     g             �t�bhhK ��h��R�(KK��h�CH      �  �  j      R           &      +   :   $   \        �t�bhhK ��h��R�(KK��h�C<   (      
   �   �     A      ~         �         �t�bhhK ��h��R�(KK��h�C   �      c       �t�bhhK ��h��R�(KK��h�C!         l      �t�bhhK ��h��R�(KK��h�C,�      ,         I  	      	   K      �t�bhhK ��h��R�(KK��h�C�        �        �t�bhhK ��h��R�(KK��h�CD         �       �        z  N   �
  T   Q  �        �t�bhhK ��h��R�(KK��h�C\"   �  �  �   �        �  �      u   
   ,            K      �      �         �t�bhhK ��h��R�(KK��h�CP      &   z         
  i   �  _  5         4   
   _      �         �t�bhhK ��h��R�(KK��h�CT�          �  /      p  �   C  �     0   <   G   �                 �t�bhhK ��h��R�(KK��h�C�   �  �  7        �t�bhhK ��h��R�(KK��h�Ch         �        �     5   [                 0   �        j  ^   |      �         �t�bhhK ��h��R�(KK
��h�C(      )   �   *  *      �        �t�bhhK ��h��R�(KK
��h�C(      �      �  �     s        �t�bhhK ��h��R�(KK��h�CD
   3   6   �        ?      !      A   �  �              �t�bhhK ��h��R�(KK��h�CP            "     .   
   _      d           �  �      �        �t�bhhK ��h��R�(KK��h�Cl      �               �         �   >      �     8   {      $   �     +      �  o        �t�bhhK ��h��R�(KK��h�C@!                 �              	      	   K      �t�bhhK ��h��R�(KK	��h�C$�      y     |      �        �t�bhhK ��h��R�(KK��h�CLI   k  �     �                    j                       �t�bhhK ��h��R�(KK��h�C<m  �  �     k     #     9  �     A   X        �t�bhhK ��h��R�(KK��h�C@
   C  _        )     �     w  
   ,               �t�bhhK ��h��R�(KK��h�Ca
     	      	         �t�bhhK ��h��R�(KK��h�C@"         2     ,  N   A           L   x  �        �t�bhhK ��h��R�(KK��h�C@d  �   +   )   �  !      �       0  `     �        �t�bhhK ��h��R�(KK	��h�C$   >   =   �     �  ;         �t�bhhK ��h��R�(KK
��h�C(.  "   �  "     |     8        �t�bhhK ��h��R�(KK��h�C0               �t�bhhK ��h��R�(KK��h�CE      2     �t�bhhK ��h��R�(KK��h�C\   H     �
           f   �   =         G   >  H                          �t�bhhK ��h��R�(KK��h�Ch      H        �  :
  �	           �	                       "            �         �t�bhhK ��h��R�(KK��h�C      L  !           �t�bhhK ��h��R�(KK��h�CL   e          �   �
     �       +     )   �     �        �t�bhhK ��h��R�(KK��h�C!  �     �t�bhhK ��h��R�(KK��h�C,         /         �               �t�bhhK ��h��R�(KK��h�Cd                       �        �   L   G   �  e  
        
      �   D        �t�bhhK ��h��R�(KK��h�C\   Q   h   6  �     Y            Q   h      6          Q        x        �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�CD      �  I  �   s     �      �     t      8   �        �t�bhhK ��h��R�(KK��h�C`
   �   �  '   -   A   �                 �        �     s     %   e           �t�bhhK ��h��R�(KK��h�C8�      u   	     ^   �        	      	         �t�bhhK ��h��R�(KK��h�C4�  �  �        '              �         �t�bhhK ��h��R�(KK��h�CH
   �  (   2      $  �   �   �     j   ]   >   �  �  g	        �t�bhhK ��h��R�(KK��h�C,C  �  /   9     7      C  8        �t�bhhK ��h��R�(KK��h�CD      5   &        
          &        "            �t�bhhK ��h��R�(KK��h�C       '   �  R  e        �t�bhhK ��h��R�(KK��h�CD�      N      .   
     �     �       U     �        �t�bhhK ��h��R�(KK��h�C01   #   
   3   6   �     /               �t�bhhK ��h��R�(KK��h�C<�   &   *               0       
   �        �t�bhhK ��h��R�(KK��h�CD     �  8   4               �  4   
   _      �        �t�bhhK ��h��R�(KK��h�C   �   B     �t�bhhK ��h��R�(KK��h�Ch      P         d
             E  �        �   �         �     �     �   �         �t�bhhK ��h��R�(KK��h�C      �     �t�bhhK ��h��R�(KK��h�CD!      �     �  m   '   -   
   3   6   �     �  m         �t�bhhK ��h��R�(KK��h�CH�   *  o  �   G   +     �      �   �         
     �        �t�bhhK ��h��R�(KK��h�C        	         �t�bhhK ��h��R�(KK	��h�C$z  �               W         �t�bhhK ��h��R�(KK��h�Cm
     6  �            �t�bhhK ��h��R�(KK��h�CL
   Z        R  �     �          �     	     �   S         �t�bhhK ��h��R�(KK��h�C8              �   �  7      �     �         �t�bhhK ��h��R�(KK��h�CH   z  �	  �            �t�bhhK ��h��R�(KK��h�CH         .         L   �  �     �   
   �     �   �        �t�bhhK ��h��R�(KK	��h�C$   R  �         �  �        �t�bhhK ��h��R�(KK��h�C       B    "   >        �t�bhhK ��h��R�(KK��h�C09   �  L   (      �  m                 �t�bhhK ��h��R�(KK��h�C4�        �      
  X  �	  	      	         �t�bhhK ��h��R�(KK��h�Cm         �       �t�bhhK ��h��R�(KK��h�C84  �   R      �      �      %      �   B        �t�bhhK ��h��R�(KK��h�C          �      	         �t�bhhK ��h��R�(KK��h�C'  �  /         �t�bhhK ��h��R�(KK��h�C               �t�bhhK ��h��R�(KK��h�Cl      -      A   ?     G              .      �                   �   �               �t�bhhK ��h��R�(KK��h�C4   �     %      �          
   3        �t�bhhK ��h��R�(KK��h�C<      D  z         *	  &      a   E  0  p        �t�bhhK ��h��R�(KK��h�C,            �  �     �           �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C8�  ]   '      H   �        �                 �t�bhhK ��h��R�(KK��h�C@   |     �     '      M       �   �  O  "   �      �t�bhhK ��h��R�(KK	��h�C$�     N   e                �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�Ch�  ;     -   {  �     %  2   
                 =      ;  &   2   a         �        �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C�          �t�bhhK ��h��R�(KK��h�C   {     �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK
��h�C(<      �        	      	         �t�bhhK ��h��R�(KK��h�C@                  
  (      �      k               �t�bhhK ��h��R�(KK��h�C<      �          �t�bhhK ��h��R�(KK��h�CH�  �   ~     �     	  l      5   [      <      �   �         �t�bhhK ��h��R�(KK��h�C,   f                  �  7         �t�bhhK ��h��R�(KK��h�C�      (     �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C      	      	         �t�bhhK ��h��R�(KK��h�C\)      �  �   �     �        0   4         �      �           �  �        �t�bhhK ��h��R�(KK��h�C@N        �      �        �
     ,   	      	   K      �t�bhhK ��h��R�(KK��h�Cp      0   y  �               o   
   ,                  K      �      �      /     �        �t�bhhK ��h��R�(KK
��h�C(/         �    	      	         �t�bhhK ��h��R�(KK��h�C@      �   �   "   �   �
  �     (                    �t�bhhK ��h��R�(KK��h�CD      5   !        V           U      O	     �        �t�bhhK ��h��R�(KK��h�C8I         �                �  �   7        �t�bhhK ��h��R�(KK��h�CP            ;      %   �              P   <   
      �   D        �t�bhhK ��h��R�(KK��h�CH         �
     v   �     $   n   &      M   �      �        �t�bhhK ��h��R�(KK��h�C8   s      �     e   '      �                 �t�bhhK ��h��R�(KK
��h�C(     B        �     p        �t�bhhK ��h��R�(KK��h�C8   `   b     �        =      �              �t�bhhK ��h��R�(KK
��h�C(
        �   H   B   �           �t�bhhK ��h��R�(KK��h�C5     �t�bhhK ��h��R�(KK��h�C   �           �t�bhhK ��h��R�(KK��h�Cz  {  |     �	     �t�bhhK ��h��R�(KK��h�Cl
   T  �     /   �        '   �  !      %   �  �         >   M   �      *   D      �        �t�bhhK ��h��R�(KK��h�CP�  �  u      �               �      �      �  +     �  �        �t�bhhK ��h��R�(KK��h�C      r     �t�bhhK ��h��R�(KK��h�C@   c     �  B  
   m                    7         �t�bhhK ��h��R�(KK��h�C�     ?	     �t�bhhK ��h��R�(KK
��h�C(T   r  �  K     �  
   �        �t�bhhK ��h��R�(KK��h�C8         �              Y  H   �  K        �t�bhhK ��h��R�(KK��h�CtN  �  	      	      	   �   	   �   	   I  	   /  	   s  	   )  	   �  	   �	  	   �  	   �  	   �     �t�bhhK ��h��R�(KK��h�CH   �      (   ^     �  V        >   �     �              �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK
��h�C(      w  (     �     {        �t�bhhK ��h��R�(KK��h�C�     �      �        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C1   #       j     �t�bhhK ��h��R�(KK��h�CH1  5     v           �  W  
        Q        L        �t�bhhK ��h��R�(KK��h�C4p  :   e      -   P      �     A           �t�bhhK ��h��R�(KK��h�CL�
     U  "      �    S     +   �   s  z     �  �   n        �t�bhhK ��h��R�(KK
��h�C(      �   >      h   #  �         �t�bhhK ��h��R�(KK��h�C<�  �  d            D      �   !      ;   g        �t�bhhK ��h��R�(KK��h�C<         �      �      )      l   9   �  7         �t�bhhK ��h��R�(KK��h�C0      5         �           <        �t�bhhK ��h��R�(KK��h�C)     u      �t�bhhK ��h��R�(KK
��h�C(%      "   >  +   �     ~
        �t�bhhK ��h��R�(KK	��h�C$H   �   �  )                  �t�bhhK ��h��R�(KK��h�CD
   3   6   )  ?   �   �   r   ?      !      ?              �t�bhhK ��h��R�(KK��h�CP
   =  �	        �
  `   ,
  :   O        (            �  �         �t�bhhK ��h��R�(KK��h�C0$   0        :      �	                 �t�bhhK ��h��R�(KK��h�C4+           �   +            c         �t�bhhK ��h��R�(KK��h�C �  Z       �     @      �t�bhhK ��h��R�(KK��h�CD�   (      v              �  i   #          �        �t�bhhK ��h��R�(KK��h�C �  �                    �t�bhhK ��h��R�(KK��h�CT   G     3            �       �  �        '         �   }         �t�bhhK ��h��R�(KK��h�CD      =      �        �  5  ^   &           �        �t�bhhK ��h��R�(KK��h�CD      =      �   �  )      $   �     �     J   �        �t�bhhK ��h��R�(KK��h�C�     �  	         �t�bhhK ��h��R�(KK��h�CW      �t�bhhK ��h��R�(KK��h�CZ   t        �t�bhhK ��h��R�(KK
��h�C(      )   �      c  
            �t�bhhK ��h��R�(KK��h�C,�	        0   �        S             �t�bhhK ��h��R�(KK��h�CD         C   
     �     �                   �
     �t�bhhK ��h��R�(KK��h�C1   #       m  �      �t�bhhK ��h��R�(KK��h�C@
   3   6      (      !      \         �     +        �t�bhhK ��h��R�(KK��h�C�      �     �t�bhhK ��h��R�(KK��h�C�     4      �      �t�bhhK ��h��R�(KK+��h�C�   �  ?      �  !   
   8   �   }                 �     �      �      ,         �      p      �  �     �     R      �     G  w     x        �t�bhhK ��h��R�(KK��h�C�  "      �t�bhhK ��h��R�(KK	��h�C$      �      6  �  �        �t�bhhK ��h��R�(KK��h�C<)   �      �   L   G   �     0      �     �        �t�bhhK ��h��R�(KK��h�C�  O	         �t�bhhK ��h��R�(KK��h�CL�        "   @               m	  0              @           �t�bhhK ��h��R�(KK��h�C      �   �  �        �t�bhhK ��h��R�(KK��h�C<         �  �     �t�bhhK ��h��R�(KK��h�CP   �  G     Y   U     �         %     z        �     J
        �t�bhhK ��h��R�(KK��h�C,H   3  �     E     X      @         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�
  O  �     �t�bhhK ��h��R�(KK��h�C*         c      �t�bhhK ��h��R�(KK��h�C@
   3   6            ?      #   !      4      m        �t�bhhK ��h��R�(KK��h�C   0         �t�bhhK ��h��R�(KK��h�C4   p     �  �	        �                 �t�bhhK ��h��R�(KK��h�CH         f     �     :      .   �     �            �      �t�bhhK ��h��R�(KK��h�C1   #   
      F         �t�bhhK ��h��R�(KK��h�C�  �  �     $   �     �t�bhhK ��h��R�(KK��h�C<   Y  
  R     �        <  V         G        �t�bhhK ��h��R�(KK��h�C8      P                  >  ^   �   n        �t�bhhK ��h��R�(KK��h�C   v   �     L         �t�bhhK ��h��R�(KK��h�C�   	
  2   (           �t�bhhK ��h��R�(KK	��h�C$   x           �  	         �t�bhhK ��h��R�(KK��h�CH�  &         �  9       �  g   �     �        W         �t�bhhK ��h��R�(KK��h�C4      J   z         5         D  ,         �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK	��h�C$          	      	         �t�bhhK ��h��R�(KK��h�C �      2   
     &  r      �t�bhhK ��h��R�(KK��h�C4V      )   C
           �     )  �        �t�bhhK ��h��R�(KK��h�C4%   (   -   [      `  Z	  "   �  
   �        �t�bhhK ��h��R�(KK��h�CT   ?   �  !      \         P         c  c  
   3   6         p         �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C,         I   �     0   R  [
        �t�bhhK ��h��R�(KK��h�CP         4      k               ;      �   %   R      <  h        �t�bhhK ��h��R�(KK��h�C 1        	      	         �t�bhhK ��h��R�(KK��h�C@      J   �                    �  B      �        �t�bhhK ��h��R�(KK��h�C4�      ;
                              �t�bhhK ��h��R�(KK��h�C45        |     �      -  D      �         �t�bhhK ��h��R�(KK��h�C�  E      �t�bhhK ��h��R�(KK
��h�C('     T   �         �     V     �t�bhhK ��h��R�(KK��h�C�   R      �     �t�bhhK ��h��R�(KK��h�C     q     �t�bhhK ��h��R�(KK��h�C8b      $   k        �   �   
         <        �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C,�     /   �           �  �  r      �t�bhhK ��h��R�(KK��h�CH      N   �  
      �      �      �     �     �  �        �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C   �    
          �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CD   /              �     q          �     �        �t�bhhK ��h��R�(KK��h�CLM   �            C  8   >     [           R   �  $   |        �t�bhhK ��h��R�(KK��h�C0�	  P     �  �  �     �   �   S        �t�bhhK ��h��R�(KK��h�C<1   #         N   �   
   3   6           �        �t�bhhK ��h��R�(KK��h�CP!      A   �     z   ,         ?         3   �  �        �         �t�bhhK ��h��R�(KK��h�C1   #       x        �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6   c        �t�bhhK ��h��R�(KK��h�CB       	         �t�bhhK ��h��R�(KK��h�C   �          {     �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK$��h�C�   $   �        Y  #   i   �   �   j   �  &      =      n     �     Y      O      �   �        
   �     �     �        �t�bhhK ��h��R�(KK��h�C    �   �   �      �        �t�bhhK ��h��R�(KK��h�C@)   �
  �        �     �  +        c   8   �        �t�bhhK ��h��R�(KK	��h�C$9   �     �     K           �t�bhhK ��h��R�(KK��h�C0   �              i      P           �t�bhhK ��h��R�(KK��h�C\      �   
   _      �   �     �   \  )   d    R      	        �  "        �t�bhhK ��h��R�(KK��h�C4�
  
      �  �     m        A     �     �t�bhhK ��h��R�(KK��h�C8T   ,     �  _     (   
   �    �          �t�bhhK ��h��R�(KK��h�CP_        �  �     ]          �     �   �      �     u         �t�bhhK ��h��R�(KK��h�C<�           �   ;     l            C           �t�bhhK ��h��R�(KK
��h�C(%   �   .     �  i   %   �         �t�bhhK ��h��R�(KK��h�CD         t        �   O      5   $   �     N   �        �t�bhhK ��h��R�(KK��h�Cp`  '      A   �        X         .   	     �           H           �                    �t�bhhK ��h��R�(KK��h�C`           m      �     C      +      �   �   v   �     �  A         `        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C4�   �      r     �  �  �     �   �         �t�bhhK ��h��R�(KK��h�C@�  �	     $   E      4      �        �     H        �t�bhhK ��h��R�(KK��h�C          	   �   	   �     �t�bhhK ��h��R�(KK��h�C09  �   .     d   :     �    �        �t�bhhK ��h��R�(KK��h�C �   '   
   ,               �t�bhhK ��h��R�(KK��h�C4         P   H        
      ,   �        �t�bhhK ��h��R�(KK��h�Cd
                   �   �               ;      �   �        ~   �               �t�bhhK ��h��R�(KK��h�C8#   !      W        E   ?      
     F         �t�bhhK ��h��R�(KK��h�CT      �      �  C         �   +     "  g            �              �t�bhhK ��h��R�(KK��h�C8            �     $   �   �  �  $   �        �t�bhhK ��h��R�(KK��h�CH      �  �   �   �  
         X      e           @         �t�bhhK ��h��R�(KK��h�CD      (         �   
   $   �                H        �t�bhhK ��h��R�(KK��h�Ct$     �     �	        �  n        �         �  O         l           0      4               �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C4)      �  �   �     �        0   4         �t�bhhK ��h��R�(KK��h�CP      5   x      �   �  �  Q              �      L   G   C        �t�bhhK ��h��R�(KK
��h�C(   #     I	  �     8   S        �t�bhhK ��h��R�(KK
��h�C(   @   '   �   �
     �           �t�bhhK ��h��R�(KK��h�CD�  0  D      �  >   T	     .         �     �  <        �t�bhhK ��h��R�(KK��h�C8#   !   (      
   3   6   �     �      �        �t�bhhK ��h��R�(KK��h�C8�     T  �   �  �   y   D   &   �     5        �t�bhhK ��h��R�(KK��h�C,   S   �   >      v                  �t�bhhK ��h��R�(KK��h�Ct
     �     �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C0              {     U   �  �         �t�bhhK ��h��R�(KK��h�CP      �   �  
                      (      t      
            �t�bhhK ��h��R�(KK��h�C1   #       �     �t�bhhK ��h��R�(KK��h�C@$   K     �              W     $   8     �   �     �t�bhhK ��h��R�(KK��h�C,�  �  �     ?        �   o         �t�bhhK ��h��R�(KK	��h�C$#   !   ?      
   w
  F         �t�bhhK ��h��R�(KK	��h�C$h  �                      �t�bhhK ��h��R�(KK
��h�C(      ;      0      r  �        �t�bhhK ��h��R�(KK��h�Cl            ;      
     �  �     �           �   �                  =      -
        �t�bhhK ��h��R�(KK
��h�C(#   !   (      :   8   A
  �        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C<<      V     �     �        �
     ,   	         �t�bhhK ��h��R�(KK��h�C`      �         �     �   E      p
                 %     )   �      T        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CQ  -     �        �t�bhhK ��h��R�(KK��h�C4:   �  �  (      -   <         �           �t�bhhK ��h��R�(KK��h�CH                  ;      �         j   4   :   �  F         �t�bhhK ��h��R�(KK��h�C@                              0   R      o        �t�bhhK ��h��R�(KK��h�Cu     !     �t�bhhK ��h��R�(KK��h�Ct   h	       p      u      2   z      ,   �         ,   f           �  C   �        �   �        �t�bhhK ��h��R�(KK��h�C9  	         �t�bhhK ��h��R�(KK��h�C0�      +      �   �           J   �      �t�bhhK ��h��R�(KK��h�C          	      	         �t�bhhK ��h��R�(KK��h�CH      g  �            �   "      �        �              �t�bhhK ��h��R�(KK��h�C    �  �   �	  G   t         �t�bhhK ��h��R�(KK��h�C\      J         )           �  
              N   
        
   �        �t�bhhK ��h��R�(KK��h�C8F     �      8   E           �  +            �t�bhhK ��h��R�(KK
��h�C(H  �   x      �      -  �          �t�bhhK ��h��R�(KK��h�Cd      �           %   h                 �  �     �   S   &     e              �t�bhhK ��h��R�(KK ��h�C��         �  "   �      (     |      �      a        r  �        L     �           �  +      �        �t�bhhK ��h��R�(KK��h�CT	  l      a   �     �        �  �  
   _      �   �     �   \        �t�bhhK ��h��R�(KK
��h�C(@   �   I  �   +   !               �t�bhhK ��h��R�(KK��h�C !        	      	         �t�bhhK ��h��R�(KK��h�C8!      R      /      p     �  	      	         �t�bhhK ��h��R�(KK��h�C0      =      �   =     �   �           �t�bhhK ��h��R�(KK��h�C,�  $   �     �  %        E         �t�bhhK ��h��R�(KK��h�CP]   P     �   �  �     �   �  �   C      �  �   �  �      �         �t�bhhK ��h��R�(KK��h�C N     �                  �t�bhhK ��h��R�(KK��h�CH   �  E  :   H   ?        �       �     :      f        �t�bhhK ��h��R�(KK��h�CP                        8   S  &      �            ^   �         �t�bhhK ��h��R�(KK��h�C0      �      E      �  
   �   I        �t�bhhK ��h��R�(KK
��h�C(   W        @      X   �        �t�bhhK ��h��R�(KK��h�C\         �         �   �         U            6  �                       �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C,   >        w   v   �     	        �t�bhhK ��h��R�(KK��h�CG     �     �t�bhhK ��h��R�(KK��h�C41   #   
   3   6   (  O      Y      O         �t�bhhK ��h��R�(KK��h�C       �           �      �t�bhhK ��h��R�(KK
��h�C(      �  U
     �   B   ?        �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�CxW        �     �     {  �     ,   	      	      	   K   	   �   	     	   �  	   �   	   �  	   �     �t�bhhK ��h��R�(KK��h�C@      /   9   9  7   '      ~     
   d     @         �t�bhhK ��h��R�(KK��h�C<)      9	     [     i  N   �                    �t�bhhK ��h��R�(KK��h�C<            �     �  9     �  �  �   �
        �t�bhhK ��h��R�(KK��h�CD�      �  �    9      _     '  :   ]      �   w         �t�bhhK ��h��R�(KK��h�C4�     �  \          �  
   A   }         �t�bhhK ��h��R�(KK��h�C@   D   ;         �   �        
   �      6            �t�bhhK ��h��R�(KK��h�C,%         �      :         �        �t�bhhK ��h��R�(KK��h�C   �   '      u        �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C !         �   �      c     �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C<     �t�bhhK ��h��R�(KK��h�C   R      �t�bhhK ��h��R�(KK��h�C      �     �t�bhhK ��h��R�(KK	��h�C$#   !   ?      
   �  F         �t�bhhK ��h��R�(KK��h�C<      �  F  +   
   �   `	           j            �t�bhhK ��h��R�(KK��h�C         �        �t�bhhK ��h��R�(KK��h�C@�   �          +      [           a     �  �     �t�bhhK ��h��R�(KK��h�CD      �      %  H  �   5      �                        �t�bhhK ��h��R�(KK��h�C   +     �t�bhhK ��h��R�(KK��h�C0      �   �  �     ,         �         �t�bhhK ��h��R�(KK��h�CD,   O      f        �     !  �           .           �t�bhhK ��h��R�(KK��h�C,      0   �   �                    �t�bhhK ��h��R�(KK��h�C<�     {     
   _         �           �        �t�bhhK ��h��R�(KK��h�C42   �
  -   �  2      �        �   �        �t�bhhK ��h��R�(KK��h�C4      M     
      
   c  
      F         �t�bhhK ��h��R�(KK��h�C4�     �  $          4  '  O  7         �t�bhhK ��h��R�(KK��h�CD      �        �  ]   �      �        +      �        �t�bhhK ��h��R�(KK��h�CX2   �        �     �   
   J  �     I   �  D  "      2   �             �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C0.  M        �     
   ,               �t�bhhK ��h��R�(KK��h�C<   �   �   	        �   D   '     (      �	        �t�bhhK ��h��R�(KK��h�C<   ]   �            $   Z       �   �           �t�bhhK ��h��R�(KK��h�C1   #       �        �t�bhhK ��h��R�(KK��h�C0
   ]   1  8   �   �      {               �t�bhhK ��h��R�(KK
��h�C(T  :         �                 �t�bhhK ��h��R�(KK��h�C4n     )   c         *     %   �  c         �t�bhhK ��h��R�(KK��h�CP      )   6     X   �     g  	        6  �        	           �t�bhhK ��h��R�(KK��h�CH   x  )      �     =              �           k        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK	��h�C$�       �      N     �     �t�bhhK ��h��R�(KK	��h�C$      U  &   ]  �  A        �t�bhhK ��h��R�(KK��h�C@      )   =      �  4   
   �   _   i         3  B     �t�bhhK ��h��R�(KK��h�ClU  &   N   �      ;     �        7  �	  '            �      �  �   �     7   �           �t�bhhK ��h��R�(KK��h�CT      �  �  =     $   E      �   ]      �  ^   8   �        t        �t�bhhK ��h��R�(KK
��h�C(!   
   B   }      m  �   
         �t�bhhK ��h��R�(KK
��h�C(h   v     d   b     >           �t�bhhK ��h��R�(KK��h�C
     �t�bhhK ��h��R�(KK��h�CT              �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C      �   O      �t�bhhK ��h��R�(KK��h�CD      �
  �                  )      
   _               �t�bhhK ��h��R�(KK��h�C`   �         �     C                �  d   �     �
  �     I   d   �        �t�bhhK ��h��R�(KK��h�C,   *        )   `      �  �        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C@   (      �  8   �        �  �        S           �t�bhhK ��h��R�(KK��h�Cl*   �      �  �        �   3  5   �      �   �  u                P     �  �   �         �t�bhhK ��h��R�(KK��h�C<�  �   '      �   �                    e         �t�bhhK ��h��R�(KK��h�Cg  �   �     �t�bhhK ��h��R�(KK��h�CTW   �   c   :     �   /      ~                    �   �               �t�bhhK ��h��R�(KK��h�C<�  
        �   
      b
  l      ~      �         �t�bhhK ��h��R�(KK��h�C8      0   o  �   �   u	                       �t�bhhK ��h��R�(KK
��h�C(1   #          J  C      !        �t�bhhK ��h��R�(KK��h�C         �  �        �t�bhhK ��h��R�(KK
��h�C(x         	      	      	   I     �t�bhhK ��h��R�(KK��h�CH   $   k      X            0      n   ^      �              �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   �                 �t�bhhK ��h��R�(KK��h�C[      E     �t�bhhK ��h��R�(KK��h�C0"   m      $  /   9   -     U   T        �t�bhhK ��h��R�(KK��h�C`D      )   �  �   �   X     2      �  �   S   }   i   ,            X     D         �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�Cl   �   (   %   �   <                     �                                            �t�bhhK ��h��R�(KK��h�C,     "   �  �   -   J     �         �t�bhhK ��h��R�(KK��h�C[
     �t�bhhK ��h��R�(KK��h�CL      ~   
   "        C     &      �   v                     �t�bhhK ��h��R�(KK��h�CT   b  �      �     �         �    7      (   w   5     �   d        �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C<"   e         �           /      �   z   �        �t�bhhK ��h��R�(KK��h�CH
   u  F   ?         �  �   �  �     %   [       �         �t�bhhK ��h��R�(KK��h�C   �     �
     �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�CH�  '   �      Q     y        �    -            �         �t�bhhK ��h��R�(KK��h�C8         .      �  �              �         �t�bhhK ��h��R�(KK��h�C,"        2   z      H   B   ^	        �t�bhhK ��h��R�(KK��h�CT     �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK
��h�C(�    �   
   �  *      �        �t�bhhK ��h��R�(KK��h�C`   �  �
        �t�bhhK ��h��R�(KK
��h�C(   �                           �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK
��h�C(l  �         C     �           �t�bhhK ��h��R�(KK��h�C@   f               :   �        �  ^              �t�bhhK ��h��R�(KK��h�C0:  
   �     N   �     �     Y        �t�bhhK ��h��R�(KK��h�C�  �         �t�bhhK ��h��R�(KK��h�C8         A  $                    �        �t�bhhK ��h��R�(KK��h�C4)   /      �     0   R      l      �        �t�bhhK ��h��R�(KK��h�CD   (   )        \      	  �      �      4      m        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C    X   '   �  �  `        �t�bhhK ��h��R�(KK��h�Cm      @     �t�bhhK ��h��R�(KK��h�C      �
  �   O         �t�b��      hhK ��h��R�(KK��h�CHd  -            �  �           8  \      &   �  ;        �t�bhhK ��h��R�(KK��h�C�             �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CP      J             �   �     �           �  �     �         �t�bhhK ��h��R�(KK��h�C �
    
   m              �t�bhhK ��h��R�(KK��h�CT      _  C   D   I  ,      �        �     V      D   A  A   /         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C �      M  	      	   K      �t�bhhK ��h��R�(KK��h�CT      |  z   ,   "   $   �   �     '      �      ,   "   H   A   �        �t�bhhK ��h��R�(KK��h�C�  �     4        �t�bhhK ��h��R�(KK��h�C<`       ^                 �         R         �t�bhhK ��h��R�(KK
��h�C(�  a  �     �  9   �  �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CE            �t�bhhK ��h��R�(KK��h�C          	      	         �t�bhhK ��h��R�(KK��h�C4      '   )   H      �        F  =        �t�bhhK ��h��R�(KK��h�C\   �  ^          Y  �  �  y      �  f     
     �     
  9            �t�bhhK ��h��R�(KK��h�CD�  j           �        �        .                 �t�bhhK ��h��R�(KK��h�C,   (      �   
         j            �t�bhhK ��h��R�(KK��h�C<      :  "      .  (      -                     �t�bhhK ��h��R�(KK��h�CP         4   
   _      �           ;      �      z               �t�bhhK ��h��R�(KK��h�CL      P         c  c  -            E     +        p        �t�bhhK ��h��R�(KK��h�C�      �     �t�bhhK ��h��R�(KK��h�C`"   e        �  #	           z      .   }      	     �     2     �  q        �t�bhhK ��h��R�(KK��h�C4�       Y  �           2              �t�bhhK ��h��R�(KK��h�C|            �   E   
           D  \   2   a           -   �   �            5  "   q   �  x  +         �t�bhhK ��h��R�(KK��h�C@^   �   �  ?           !         5                 �t�bhhK ��h��R�(KK��h�C8!         	      	   K   	     	   �   	   �     �t�bhhK ��h��R�(KK��h�CD"      �     2   �   p     �	           @     	        �t�bhhK ��h��R�(KK��h�C      l               �t�bhhK ��h��R�(KK	��h�C$�        �  
  i            �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�C   �      	         �t�bhhK ��h��R�(KK��h�C<u                     &  �        '  (        �t�bhhK ��h��R�(KK��h�CT�      ;     �      J   z   
   �     �   O  �        �     �        �t�bhhK ��h��R�(KK��h�C    �
  c         Z        �t�bhhK ��h��R�(KK��h�CD�  &   N            t   &   D  �  �   `   3             �t�bhhK ��h��R�(KK��h�C    �  ]      $   �        �t�bhhK ��h��R�(KK��h�C`      J   �               &      U      .            R  `	  "   $   �   �        �t�bhhK ��h��R�(KK��h�C4           i            p     �        �t�bhhK ��h��R�(KK
��h�C(d   A   K     N      
   �        �t�bhhK ��h��R�(KK��h�C 2         i     �        �t�bhhK ��h��R�(KK��h�C4�  3     �  '   
   3   6   3              �t�bhhK ��h��R�(KK��h�C�  p      �     �t�bhhK ��h��R�(KK��h�CD�     �     <  �  )   A   R   �     	     V           �t�bhhK ��h��R�(KK��h�C,�  �            
   ,               �t�bhhK ��h��R�(KK��h�Cd   f   �         �      $   ;         �   �         )         G  �   �      7         �t�bhhK ��h��R�(KK��h�C,   �      ,  ~  l         �  �      �t�bhhK ��h��R�(KK��h�CH/      �      2     �   �           �     �     �
        �t�bhhK ��h��R�(KK��h�CT         ;      0     m     A   U     &      =      �   "   W         �t�bhhK ��h��R�(KK��h�C@      (      4         T     �        ,           �t�bhhK ��h��R�(KK��h�CH1   #               +        .         
   3   6            �t�bhhK ��h��R�(KK��h�C      d   �     �t�bhhK ��h��R�(KK��h�CH-   !       l            o  �         }     "	          �t�bhhK ��h��R�(KK��h�CZ  	      	         �t�bhhK ��h��R�(KK	��h�C$   e   '   �                  �t�bhhK ��h��R�(KK��h�CT3    >      F  C      �     j   %      )      j      a   �  C         �t�bhhK ��h��R�(KK��h�C �        ;      �        �t�bhhK ��h��R�(KK��h�C8   e   '   �  6        �	  9     �	           �t�bhhK ��h��R�(KK��h�C      �   |      �     �t�bhhK ��h��R�(KK��h�C`G      �            6       0      n      �   �     N   �  i      �   =        �t�bhhK ��h��R�(KK��h�C n     �  	      	         �t�bhhK ��h��R�(KK!��h�C��
     b     �      �        �     ,   	      	      	   K   	   �   	   �   	   I  	   U  	   �  	   �   	   s     �t�bhhK ��h��R�(KK��h�CTp     �      �              ,   	      	   K   	     	   �   	   �     �t�bhhK ��h��R�(KK��h�CL�     4      �     $  q   �     �  �        �  $   0        �t�bhhK ��h��R�(KK��h�C@   �     �  g   O        .        �             �t�bhhK ��h��R�(KK��h�CH�   �                   h   Y      �        �            �t�bhhK ��h��R�(KK��h�C<   �     �          Q     �  0  B   ?        �t�bhhK ��h��R�(KK��h�C    ;  �                �t�bhhK ��h��R�(KK	��h�C$|      �   a     r  '        �t�bhhK ��h��R�(KK��h�CT         ;           8   E           )   0      �                 �t�bhhK ��h��R�(KK��h�C�   �     �t�bhhK ��h��R�(KK	��h�C$[      �      	      	         �t�bhhK ��h��R�(KK��h�CD               P   <         0   [         �          �t�bhhK ��h��R�(KK��h�C0      N               M               �t�bhhK ��h��R�(KK��h�CL   �   {     0  �   f     �      �   =      �  e  :   �        �t�bhhK ��h��R�(KK��h�CT@      z             �     k     ,      �  �           X        �t�bhhK ��h��R�(KK	��h�C$   >   =      �     w        �t�bhhK ��h��R�(KK��h�CH         �   �        P                 �   �  �         �t�bhhK ��h��R�(KK��h�C4         0      0  �   
        �         �t�bhhK ��h��R�(KK��h�CD   X   '   )         �     V   2      �   O  
            �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C8!        	      	      	   K   	   �   	   �      �t�bhhK ��h��R�(KK��h�CX         Y      O         =      +  �  *                 �  7         �t�bhhK ��h��R�(KK��h�C �            j   v        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�Ce   �   �           �t�bhhK ��h��R�(KK��h�Ch     �t�bhhK ��h��R�(KK��h�C R     ;     �  �        �t�bhhK ��h��R�(KK
��h�C(   ^  �        �     T
        �t�bhhK ��h��R�(KK��h�C<   `   �         �  A  �   �   5      7  4         �t�bhhK ��h��R�(KK��h�C0*        A  &      U   �  "            �t�bhhK ��h��R�(KK��h�C    �   	  �     ~        �t�bhhK ��h��R�(KK��h�CTi        �        K        ~      D   �         2     d            �t�bhhK ��h��R�(KK��h�CL         O         Y      Q      (            H              �t�bhhK ��h��R�(KK��h�C8I   (   �  �  �   �     J  C   -              �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C          �t�be.