Grundläggande information
Historia
Trafik
Religion
Beslutsfattande och påverkan
Grundläggande information
Karleby finns i Mellersta Österbotten invid Bottniska viken.
Karleby stad är grundad 1620 och hette då Gamlakarleby.
Senare blev Kokkola stadens finska namn.
Vid Karleby centrum finns en av landets mest omfattande historiska trästadshelheter.
Stadsplanen är från 1650-talet.
Den omfattar 12 kvarter med hundratals trähus och gårdsbyggnader.
De äldsta av dessa är från 1600-talet.
Karleby är en kulturstad med mycket att se och uppleva.
Karleby hamn ligger i stadsdelen Yxpila och är en av Finlands mest trafikerade godshamnar.
Grunden för näringslivet i Karleby är den internationella storindustrin.
I Karleby är den kemiska industrin och industri i anslutning till denna särskilt viktig.
Karleby är även en betydande handelsstad.
Information om Karlebyfinska _ svenska _ engelska
Historia
Redan under medeltiden fanns det hamn, båtbygge och handelsplats i Karleby.
Landhöjningen har varit en central faktor i Karlebys historia.
Den har format omgivningen i hög grad och bland annat påverkat utvecklingen av hamnverksamheten och handeln.
Handel bedrevs längs med Bottniska vikens kust och jordbruk, jakt, fiske och sälfångst var även viktiga näringar.
Exporten av tjära, som blev mycket viktig för Karlebys historia, inleddes redan på 1500-talet.
Den sjunde september 1620 undertecknade Sveriges kung Gustav II Adolf en handling som gav den lilla jordbruks- och fiskebyn vid Ristrand status som stad.
Dagens stadssund var då en smal havsvik som sträckte sig ända till Kyrkbacken.
Sakta men säkert blev Karleby en viktig stad för sjöfart och skeppsbygge.
Skeppsvarv fanns bland annat i Kaustarviken, Svartskär och Soldatskär.
Inledningsvis seglade man endast till Åbo och Stockholm, eftersom Karleby som s.k. uppstad inte fick bedriva utrikeshandel.
År 1765 erhöll staden stapelrättigheter, dvs. rätt till fri utrikeshandel, främst tack vare den aktiva kyrkoherden och lantdagsmannen Anders Chydenius.
Karleby blev snabbt en förmögen stad i början av 1800-talet tack vare just handeln med tjära och rederiverksamheten.
Stadens borgare köpte tjära av bönder och exporterade den, ofta till hamnar vid Medelhavet och i England.
Karleby handelsflotta var under perioder Finlands största.
Den snabba ekonomiska utvecklingen avtog i mitten av 1800-talet, men tog ny fart i slutet av århundradet tack vare industrialiseringen.
Karleby blev en viktig industristad främst tack vare läder- och metallindustrin.
Karlebys historiafinska _ svenska _ engelska
Trafik
Karleby har goda trafikförbindelser.
Via Karleby löper riksväg 8 och 13.
Järnvägsstationen finns i stadens centrum.
Restiden med tåg till Helsingfors är cirka fyra timmar.
Flygplatsen finns i Kronoby på endast 22 kilometers avstånd från Karleby centrum.
Stadsborna erbjuds även ett tryggt, omfattande, fungerande och trivsamt nätverk för den lätta trafiken.
Karleby har satsat på att förbättra förhållandena för cyklister.
Lokalbussarna trafikerar de olika delarna av staden på vardagar.
Läs mer: Trafik.
Gator och trafikfinska _ svenska
Kollektivtrafikfinska _ svenska
linkkiVR:
Tågtidtabellerfinska _ svenska _ engelska _ ryska
Busstidtabellerfinska _ svenska _ engelska
Flyg från Karleby-Jakobstad flygplatsfinska _ svenska _ engelska
Religion
I Karleby finns flera olika religiösa samfund.
I tjänsten Uskonnot Suomessa (Religioner i Finland) finns information om religiösa samfund enligt ort.
Den evangelisk-lutherska kyrkan har fyra finskspråkiga församlingar och en svenskspråkig församling i Karleby.
Läs mer på Karleby kyrkliga samfällighets webbplats.
I Karleby finns en ortodox kyrka.
Mer information om den ortodoxa församlingens verksamhet i Karleby finns på Vasa ortodoxa församlings webbplats.
Läs mer: Kulturer och religioner i Finland.
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiVasa ortodoxa församling:
Vasa ortodoxa församlingfinska _ engelska _ ryska
Beslutsfattande och påverkan
Den högsta beslutsfattande makten i Karleby stad innehas av stadsfullmäktige.
Fullmäktigeledamöterna och deras suppleanter väljs vid kommunalval vart fjärde år.
På stadens webbplats finns information om stadsfullmäktige och dess beslut.
Invånarna kan påverka stadens beslutsfattande redan då beslut bereds.
Information om olika sätt att delta och påverka finns på stadens webbplats.
Kommunens invånare har enligt kommunallagen rätt att lämna in motioner till kommunen i ärenden som gäller dess verksamhet.
I Karleby finns ungdomsfullmäktige, äldre- och handikappråd samt ett råd för kulturell mångfald.
Läs mer: Finlands förvaltning, Val och röstning i Finland
Beslutsfattandefinska _ svenska _ engelska
Grundläggande information
Historia
Trafik
Religion
Beslutsfattande och påverkan
Grundläggande information
Karleby finns i Mellersta Österbotten invid Bottniska viken.
Karleby stad är grundad 1620 och hette då Gamlakarleby.
Senare blev Kokkola stadens finska namn.
Vid Karleby centrum finns en av landets mest omfattande historiska trästadshelheter.
Stadsplanen är från 1650-talet.
Den omfattar 12 kvarter med hundratals trähus och gårdsbyggnader.
De äldsta av dessa är från 1600-talet.
Karleby är en kulturstad med mycket att se och uppleva.
Karleby hamn ligger i stadsdelen Yxpila och är en av Finlands mest trafikerade godshamnar.
Grunden för näringslivet i Karleby är den internationella storindustrin.
I Karleby är den kemiska industrin och industri i anslutning till denna särskilt viktig.
Karleby är även en betydande handelsstad.
Information om Karlebyfinska _ svenska _ engelska
Historia
Redan under medeltiden fanns det hamn, båtbygge och handelsplats i Karleby.
Landhöjningen har varit en central faktor i Karlebys historia.
Den har format omgivningen i hög grad och bland annat påverkat utvecklingen av hamnverksamheten och handeln.
Handel bedrevs längs med Bottniska vikens kust och jordbruk, jakt, fiske och sälfångst var även viktiga näringar.
Exporten av tjära, som blev mycket viktig för Karlebys historia, inleddes redan på 1500-talet.
Den sjunde september 1620 undertecknade Sveriges kung Gustav II Adolf en handling som gav den lilla jordbruks- och fiskebyn vid Ristrand status som stad.
Dagens stadssund var då en smal havsvik som sträckte sig ända till Kyrkbacken.
Sakta men säkert blev Karleby en viktig stad för sjöfart och skeppsbygge.
Skeppsvarv fanns bland annat i Kaustarviken, Svartskär och Soldatskär.
Inledningsvis seglade man endast till Åbo och Stockholm, eftersom Karleby som s.k. uppstad inte fick bedriva utrikeshandel.
År 1765 erhöll staden stapelrättigheter, dvs. rätt till fri utrikeshandel, främst tack vare den aktiva kyrkoherden och lantdagsmannen Anders Chydenius.
Karleby blev snabbt en förmögen stad i början av 1800-talet tack vare just handeln med tjära och rederiverksamheten.
Stadens borgare köpte tjära av bönder och exporterade den, ofta till hamnar vid Medelhavet och i England.
Karleby handelsflotta var under perioder Finlands största.
Den snabba ekonomiska utvecklingen avtog i mitten av 1800-talet, men tog ny fart i slutet av århundradet tack vare industrialiseringen.
Karleby blev en viktig industristad främst tack vare läder- och metallindustrin.
Karlebys historiafinska _ svenska _ engelska
Trafik
Karleby har goda trafikförbindelser.
Via Karleby löper riksväg 8 och 13.
Järnvägsstationen finns i stadens centrum.
Restiden med tåg till Helsingfors är cirka fyra timmar.
Flygplatsen finns i Kronoby på endast 22 kilometers avstånd från Karleby centrum.
Stadsborna erbjuds även ett tryggt, omfattande, fungerande och trivsamt nätverk för den lätta trafiken.
Karleby har satsat på att förbättra förhållandena för cyklister.
Lokalbussarna trafikerar de olika delarna av staden på vardagar.
Läs mer: Trafik.
Gator och trafikfinska _ svenska
Kollektivtrafikfinska _ svenska
linkkiVR:
Tågtidtabellerfinska _ svenska _ engelska _ ryska
Busstidtabellerfinska _ svenska _ engelska
Flyg från Karleby-Jakobstad flygplatsfinska _ svenska _ engelska
Religion
I Karleby finns flera olika religiösa samfund.
I tjänsten Uskonnot Suomessa (Religioner i Finland) finns information om religiösa samfund enligt ort.
Den evangelisk-lutherska kyrkan har fyra finskspråkiga församlingar och en svenskspråkig församling i Karleby.
Läs mer på Karleby kyrkliga samfällighets webbplats.
I Karleby finns en ortodox kyrka.
Mer information om den ortodoxa församlingens verksamhet i Karleby finns på Vasa ortodoxa församlings webbplats.
Läs mer: Kulturer och religioner i Finland.
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiVasa ortodoxa församling:
Vasa ortodoxa församlingfinska _ engelska _ ryska
Beslutsfattande och påverkan
Den högsta beslutsfattande makten i Karleby stad innehas av stadsfullmäktige.
Fullmäktigeledamöterna och deras suppleanter väljs vid kommunalval vart fjärde år.
På stadens webbplats finns information om stadsfullmäktige och dess beslut.
Invånarna kan påverka stadens beslutsfattande redan då beslut bereds.
Information om olika sätt att delta och påverka finns på stadens webbplats.
Kommunens invånare har enligt kommunallagen rätt att lämna in motioner till kommunen i ärenden som gäller dess verksamhet.
I Karleby finns ungdomsfullmäktige, äldre- och handikappråd samt ett råd för kulturell mångfald.
Läs mer: Finlands förvaltning, Val och röstning i Finland
Beslutsfattandefinska _ svenska _ engelska
Grundläggande information
Historia
Trafik
Religion
Beslutsfattande och påverkan
Grundläggande information
Karleby finns i Mellersta Österbotten invid Bottniska viken.
Karleby stad är grundad 1620 och hette då Gamlakarleby.
Senare blev Kokkola stadens finska namn.
Vid Karleby centrum finns en av landets mest omfattande historiska trästadshelheter.
Stadsplanen är från 1650-talet.
Den omfattar 12 kvarter med hundratals trähus och gårdsbyggnader.
De äldsta av dessa är från 1600-talet.
Karleby är en kulturstad med mycket att se och uppleva.
Karleby hamn ligger i stadsdelen Yxpila och är en av Finlands mest trafikerade godshamnar.
Grunden för näringslivet i Karleby är den internationella storindustrin.
I Karleby är den kemiska industrin och industri i anslutning till denna särskilt viktig.
Karleby är även en betydande handelsstad.
Information om Karlebyfinska _ svenska _ engelska
Historia
Redan under medeltiden fanns det hamn, båtbygge och handelsplats i Karleby.
Landhöjningen har varit en central faktor i Karlebys historia.
Den har format omgivningen i hög grad och bland annat påverkat utvecklingen av hamnverksamheten och handeln.
Handel bedrevs längs med Bottniska vikens kust och jordbruk, jakt, fiske och sälfångst var även viktiga näringar.
Exporten av tjära, som blev mycket viktig för Karlebys historia, inleddes redan på 1500-talet.
Den sjunde september 1620 undertecknade Sveriges kung Gustav II Adolf en handling som gav den lilla jordbruks- och fiskebyn vid Ristrand status som stad.
Dagens stadssund var då en smal havsvik som sträckte sig ända till Kyrkbacken.
Sakta men säkert blev Karleby en viktig stad för sjöfart och skeppsbygge.
Skeppsvarv fanns bland annat i Kaustarviken, Svartskär och Soldatskär.
Inledningsvis seglade man endast till Åbo och Stockholm, eftersom Karleby som s.k. uppstad inte fick bedriva utrikeshandel.
År 1765 erhöll staden stapelrättigheter, dvs. rätt till fri utrikeshandel, främst tack vare den aktiva kyrkoherden och lantdagsmannen Anders Chydenius.
Karleby blev snabbt en förmögen stad i början av 1800-talet tack vare just handeln med tjära och rederiverksamheten.
Stadens borgare köpte tjära av bönder och exporterade den, ofta till hamnar vid Medelhavet och i England.
Karleby handelsflotta var under perioder Finlands största.
Den snabba ekonomiska utvecklingen avtog i mitten av 1800-talet, men tog ny fart i slutet av århundradet tack vare industrialiseringen.
Karleby blev en viktig industristad främst tack vare läder- och metallindustrin.
Karlebys historiafinska _ svenska _ engelska
Trafik
Karleby har goda trafikförbindelser.
Via Karleby löper riksväg 8 och 13.
Järnvägsstationen finns i stadens centrum.
Restiden med tåg till Helsingfors är cirka fyra timmar.
Flygplatsen finns i Kronoby på endast 22 kilometers avstånd från Karleby centrum.
Stadsborna erbjuds även ett tryggt, omfattande, fungerande och trivsamt nätverk för den lätta trafiken.
Karleby har satsat på att förbättra förhållandena för cyklister.
Lokalbussarna trafikerar de olika delarna av staden på vardagar.
Läs mer: Trafik.
Gator och trafikfinska _ svenska
Kollektivtrafikfinska _ svenska
linkkiVR:
Tågtidtabellerfinska _ svenska _ engelska _ ryska
Busstidtabellerfinska _ svenska _ engelska
Flyg från Karleby-Jakobstad flygplatsfinska _ svenska _ engelska
Religion
I Karleby finns flera olika religiösa samfund.
I tjänsten Uskonnot Suomessa (Religioner i Finland) finns information om religiösa samfund enligt ort.
Den evangelisk-lutherska kyrkan har fyra finskspråkiga församlingar och en svenskspråkig församling i Karleby.
Läs mer på Karleby kyrkliga samfällighets webbplats.
I Karleby finns en ortodox kyrka.
Mer information om den ortodoxa församlingens verksamhet i Karleby finns på Vasa ortodoxa församlings webbplats.
Läs mer: Kulturer och religioner i Finland.
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiVasa ortodoxa församling:
Vasa ortodoxa församlingfinska _ engelska _ ryska
Beslutsfattande och påverkan
Den högsta beslutsfattande makten i Karleby stad innehas av stadsfullmäktige.
Fullmäktigeledamöterna och deras suppleanter väljs vid kommunalval vart fjärde år.
På stadens webbplats finns information om stadsfullmäktige och dess beslut.
Invånarna kan påverka stadens beslutsfattande redan då beslut bereds.
Information om olika sätt att delta och påverka finns på stadens webbplats.
Kommunens invånare har enligt kommunallagen rätt att lämna in motioner till kommunen i ärenden som gäller dess verksamhet.
I Karleby finns ungdomsfullmäktige, äldre- och handikappråd samt ett råd för kulturell mångfald.
Läs mer: Finlands förvaltning, Val och röstning i Finland
Beslutsfattandefinska _ svenska _ engelska
Detta innehåll finns inte på det språk som du har valt.
Välj något annat språk.
Finska
Detta innehåll finns inte på det språk som du har valt.
Välj något annat språk.
Finska
Detta innehåll finns inte på det språk som du har valt.
Välj något annat språk.
Finska
Bibliotek
Motion
Att röra sig i naturen
Teater och film
Museer
Hobbyer för barn och unga
Föreningar
Karleby är en gammal sjöstad som erbjuder mångsidiga möjligheter för utfärder och friluftsliv.
Personer ntresserad av friluftsliv bör läsa mer om allemansrätten under rubriken ”Att röra sig i naturen” i denna tjänst.
Flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet.
Föreningar och organisationer samt hobbygrupper och kommunala institut erbjuder kurser i idrott och kultur samt bl.a. språk och hantverk.
I Snellman-salen och i stadens övriga kulturlokaler erbjuds kulturevenemang av varierande slag.
Årliga evenemang i Karleby är bland annat Veneziansk afton i slutet av sommaren, Kokkola Cup för fotbollsjuniorer, Stadsfestivalen Karleby sommarveckor, Lochteå kyrkomusikfest samt Vinterdans i Karleby och festivalen Karleby Vinterharmonika.
Mer information om fritidstjänsterna i Karleby finns på Karleby stads webbplats.
På stadens webbplats finns även en länk till Evenemangskalendern med daglig information om stadens kultur- och motionsevenemang.
Läs mer: Fritid.
Evenemangskalenderfinska
Kulturtjänsterfinska _ svenska _ engelska
Idrottstjänsterfinska _ svenska _ engelska
Bibliotek
Karleby stadsbibliotek finns i stadens centrum.
Närbiblioteken finns i Björkhagen, Kelviå, Lochteå samt Ullava kyrkby och Rahkonen.
Information om bibliotekets öppettider och tjänster finns på dess webbplats.
Biblioteket finns även på nätet.
Där kan kunderna bläddra i bibliotekets samlingar, reservera material, förnya sina lån, beställa fjärrlån och låna e-böcker under alla tider på dygnet.
Tack vare det effektiva biblioteksnätverket i Finland är nästan alla finländska biblioteks samlingar tillgängliga för bibliotekskunderna i Karleby.
Karleby stadsbibliotek/huvudbiblioteket
Storgatan 3, 67100 Karleby
Telefon: 040 806 5124, 040 806 5133
Läs mer: Bibliotek.
Bibliotekstjänsterfinska _ svenska _ engelska
Motion
I Karleby finns mångsidiga motionsmöjligheter året runt.
Staden anordnar ledda aktiviteter i Simcentret VesiVeijari och motionshallarna.
Dessutom finns det gym av flera olika slag.
Gym anpassade för äldre finns i Furuåsens aktivitetscenter och Kuusikumpu servicehus.
Staden underhåller cykelvägar, motionsrutter, joggingbanor, skidspår, badstränder, bollplaner och skridskobanor samt platser för närmotion.
I Karlebynejdens instituts nättjänst finns information om institutets mångsidiga motionsutbud.
I Karleby finns nära på hundra idrottsföreningar för olika grenar samt föreningar som arrangerar övrig motion.
Mer information om motionsmöjligheter i Karleby finns på Karleby stads webbplats.
Läs mer:
Motion.
Idrottstjänsterfinska _ svenska _ engelska
Motionsplatserfinska _ svenska
Gym för äldrefinska
Karlebynejdens institutfinska _ svenska
Att röra sig i naturen
Att röra sig i naturen är en traditionell och populär form av avkoppling för finländarna under alla årstider.
I Finland kan man med stöd av allemansrätten plocka bär och svamp i skogen och röra sig till fots, med cykel eller skidor vintertid.
Det är inte tillåtet att beträda folks gårdar utan lov.
För fiske krävs fiskelov, med undantag för mete och pilkning.
Även jakt fordrar jakttillstånd.
Allemansrätten ger inte rätt att skräpa ner i naturen, skada träd eller växter, störa eller skada fågelbon eller fågelungar, köra motorfordon utan markägarens tillstånd eller bygga ens tillfälliga byggen.
Mer information om motionsrutterna, rastplatser, möjligheter till fiske och båtliv samt exempelvis fågeltorn i Karleby finns på stadens webbplats.
Rutterna för camping, paddling, vandring, cykling och övriga rutter i Karleby finns i karttjänsten på nätet.
I karttjänsten visas även var största delen av motionsplatserna finns.
Du kan köpa friluftskartor över Karleby hos Karleby Turism: Salutorget 5, 67100 Karleby.
Läs mer: Att röra sig i naturen.
linkkiMiljöförvaltningen:
Allemansrättenfinska _ svenska _ engelska _ ryska
Motionskarta över Karlebyfinska _ svenska
Motionsrutter i Karlebyfinska _ svenska
Teater och film
Karleby är en teaterstad med långa anor, som erbjuder scenkonst på hög nivå framförd av både proffs och amatörer.
Karleby stadsteater finns i det stämningsfulla Vartiolinna (Torggatan 48).
Du kan läsa mer om amatörteatrarnas verksamhet på deras webbplats och i evenemangskalendern.
I Karleby finns biografen Bio Rex, vars två salar använder digital- och 3D-teknik.
Bio Rex program finns under länken här intill.
Läs mer: Teater och film.
Stadsteaternfinska
Biograffinska
Teater och danskonst i Karlebyfinska _ svenska _ engelska
Evenemangskalenderfinska
Museer
I hjärtat av staden, i det anrika Rooska gården, finns K.H.Renlunds museum.
Karleby stad grundade museet 1909 utgående från en testamentsgåva av affärsmannen Karl Herman Renlund (1850–1908) .
På museet finns Renlunds samling av finländsk konst från guldåldern och tillfälliga utställningar i en kulturhistorisk miljö.
Även i museikvarterens övriga byggnader finns utställningar om stadens kulturhistoria och utställningar med ITE-konst.
På K.H.Renlunds museums webbplats finns mer information om museets tjänster, utställningar samt aktuell verksamhet.
Utöver K.H.Renlunds museum lönar det sig att besöka det naturhistoriska museet Kieppi (Kieppi är stängt tills vidare på grund av brand) samt de många hembygdsmuseerna och övriga de historiska resmålen i regionen.
Exempelvis i Konst-Vionoja-centret presenteras konstnären Veikko Vionojas verk.
I Kelviå, ca 10 km norrut från Karleby, finns Toivonen djurpark och drängmuseum.
Mer information om dessa museer finns under länkarna här intill.
Läs mer: Museer.
Museer och traditionsarbetefinska _ svenska _ engelska
K.H. Renlunds museum - Mellersta Österbottens landskapsmuseumfinska _ svenska _ engelska
Kieppi, Karleby naturvetenskapliga museumfinska _ svenska _ engelska
linkkiToivonens djurpark och drängmuseum :
Toivonens djurpark och drängmuseum finska _ svenska _ engelska
Konst Vionojafinska
Hobbyer för barn och unga
Flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet.
Flera olika föreningar samt kommunala institut ger unga möjlighet att studera idrott och kultur samt bl.a. språk och hantverk.
Barn och unga kan delta i grundläggande undervisning i musik, dans, bildkonst och hantverk.
Dessutom erbjuder stadens ungdomstjänster en rockskola.
Stadens ungdomstjänster driver sju ungdomsgårdar runt om i Karleby.
De rusmedels- och rökfria ungdomslokalerna erbjuder handledd verksamhet för barn i årskurserna 3–6 och unga i åldern 13–17 år i olika delar av Karleby.
Information om hobbyverksamheter för barn och unga finns på stadens webbplats.
Rådgivningen vid Ungdomsgården Vinge ger aktuell information om bl.a. internationalisering, studier, arbetsliv, hälsa, hobbyverksamhet och boende.
Karlebynejdens institut erbjuder barn och unga olika former av hobbyverksamhet, exempelvis i konstämnen och musik.
Kontrollera vilka kurser som är aktuella i institutets webbtjänst.
Karleby evangelisk-lutherska församlingar erbjuder även hobbyverksamhet för barn och unga, såsom lekparksträffar, klubbar, musikverksamhet och läger.
Mer information om verksamheten finns på Karleby församlingssammanslutnings webbplats.
Ungdomsgården Vinge
67100 Karleby
Läs mer: Hobbyer för barn och unga.
Övrig undervisning i Karlebyfinska _ svenska
Ungdomstjänsterfinska _ svenska _ engelska
Karlebynejdens institutfinska _ svenska
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
Föreningar
Karleby har ett aktivt och mångsidigt föreningsliv för invånare i alla åldrar.
Läs mer: Föreningar.
Bibliotek
Motion
Att röra sig i naturen
Teater och film
Museer
Hobbyer för barn och unga
Föreningar
Karleby är en gammal sjöstad som erbjuder mångsidiga möjligheter för utfärder och friluftsliv.
Personer ntresserad av friluftsliv bör läsa mer om allemansrätten under rubriken ”Att röra sig i naturen” i denna tjänst.
Flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet.
Föreningar och organisationer samt hobbygrupper och kommunala institut erbjuder kurser i idrott och kultur samt bl.a. språk och hantverk.
I Snellman-salen och i stadens övriga kulturlokaler erbjuds kulturevenemang av varierande slag.
Årliga evenemang i Karleby är bland annat Veneziansk afton i slutet av sommaren, Kokkola Cup för fotbollsjuniorer, Stadsfestivalen Karleby sommarveckor, Lochteå kyrkomusikfest samt Vinterdans i Karleby och festivalen Karleby Vinterharmonika.
Mer information om fritidstjänsterna i Karleby finns på Karleby stads webbplats.
På stadens webbplats finns även en länk till Evenemangskalendern med daglig information om stadens kultur- och motionsevenemang.
Läs mer: Fritid.
Evenemangskalenderfinska
Kulturtjänsterfinska _ svenska _ engelska
Idrottstjänsterfinska _ svenska _ engelska
Bibliotek
Karleby stadsbibliotek finns i stadens centrum.
Närbiblioteken finns i Björkhagen, Kelviå, Lochteå samt Ullava kyrkby och Rahkonen.
Information om bibliotekets öppettider och tjänster finns på dess webbplats.
Biblioteket finns även på nätet.
Där kan kunderna bläddra i bibliotekets samlingar, reservera material, förnya sina lån, beställa fjärrlån och låna e-böcker under alla tider på dygnet.
Tack vare det effektiva biblioteksnätverket i Finland är nästan alla finländska biblioteks samlingar tillgängliga för bibliotekskunderna i Karleby.
Karleby stadsbibliotek/huvudbiblioteket
Storgatan 3, 67100 Karleby
Telefon: 040 806 5124, 040 806 5133
Läs mer: Bibliotek.
Bibliotekstjänsterfinska _ svenska _ engelska
Motion
I Karleby finns mångsidiga motionsmöjligheter året runt.
Staden anordnar ledda aktiviteter i Simcentret VesiVeijari och motionshallarna.
Dessutom finns det gym av flera olika slag.
Gym anpassade för äldre finns i Furuåsens aktivitetscenter och Kuusikumpu servicehus.
Staden underhåller cykelvägar, motionsrutter, joggingbanor, skidspår, badstränder, bollplaner och skridskobanor samt platser för närmotion.
I Karlebynejdens instituts nättjänst finns information om institutets mångsidiga motionsutbud.
I Karleby finns nära på hundra idrottsföreningar för olika grenar samt föreningar som arrangerar övrig motion.
Mer information om motionsmöjligheter i Karleby finns på Karleby stads webbplats.
Läs mer:
Motion.
Idrottstjänsterfinska _ svenska _ engelska
Motionsplatserfinska _ svenska
Gym för äldrefinska
Karlebynejdens institutfinska _ svenska
Att röra sig i naturen
Att röra sig i naturen är en traditionell och populär form av avkoppling för finländarna under alla årstider.
I Finland kan man med stöd av allemansrätten plocka bär och svamp i skogen och röra sig till fots, med cykel eller skidor vintertid.
Det är inte tillåtet att beträda folks gårdar utan lov.
För fiske krävs fiskelov, med undantag för mete och pilkning.
Även jakt fordrar jakttillstånd.
Allemansrätten ger inte rätt att skräpa ner i naturen, skada träd eller växter, störa eller skada fågelbon eller fågelungar, köra motorfordon utan markägarens tillstånd eller bygga ens tillfälliga byggen.
Mer information om motionsrutterna, rastplatser, möjligheter till fiske och båtliv samt exempelvis fågeltorn i Karleby finns på stadens webbplats.
Rutterna för camping, paddling, vandring, cykling och övriga rutter i Karleby finns i karttjänsten på nätet.
I karttjänsten visas även var största delen av motionsplatserna finns.
Du kan köpa friluftskartor över Karleby hos Karleby Turism: Salutorget 5, 67100 Karleby.
Läs mer: Att röra sig i naturen.
linkkiMiljöförvaltningen:
Allemansrättenfinska _ svenska _ engelska _ ryska
Motionskarta över Karlebyfinska _ svenska
Motionsrutter i Karlebyfinska _ svenska
Teater och film
Karleby är en teaterstad med långa anor, som erbjuder scenkonst på hög nivå framförd av både proffs och amatörer.
Karleby stadsteater finns i det stämningsfulla Vartiolinna (Torggatan 48).
Du kan läsa mer om amatörteatrarnas verksamhet på deras webbplats och i evenemangskalendern.
I Karleby finns biografen Bio Rex, vars två salar använder digital- och 3D-teknik.
Bio Rex program finns under länken här intill.
Läs mer: Teater och film.
Stadsteaternfinska
Biograffinska
Teater och danskonst i Karlebyfinska _ svenska _ engelska
Evenemangskalenderfinska
Museer
I hjärtat av staden, i det anrika Rooska gården, finns K.H.Renlunds museum.
Karleby stad grundade museet 1909 utgående från en testamentsgåva av affärsmannen Karl Herman Renlund (1850–1908) .
På museet finns Renlunds samling av finländsk konst från guldåldern och tillfälliga utställningar i en kulturhistorisk miljö.
Även i museikvarterens övriga byggnader finns utställningar om stadens kulturhistoria och utställningar med ITE-konst.
På K.H.Renlunds museums webbplats finns mer information om museets tjänster, utställningar samt aktuell verksamhet.
Utöver K.H.Renlunds museum lönar det sig att besöka det naturhistoriska museet Kieppi (Kieppi är stängt tills vidare på grund av brand) samt de många hembygdsmuseerna och övriga de historiska resmålen i regionen.
Exempelvis i Konst-Vionoja-centret presenteras konstnären Veikko Vionojas verk.
I Kelviå, ca 10 km norrut från Karleby, finns Toivonen djurpark och drängmuseum.
Mer information om dessa museer finns under länkarna här intill.
Läs mer: Museer.
Museer och traditionsarbetefinska _ svenska _ engelska
K.H. Renlunds museum - Mellersta Österbottens landskapsmuseumfinska _ svenska _ engelska
Kieppi, Karleby naturvetenskapliga museumfinska _ svenska _ engelska
linkkiToivonens djurpark och drängmuseum :
Toivonens djurpark och drängmuseum finska _ svenska _ engelska
Konst Vionojafinska
Hobbyer för barn och unga
Flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet.
Flera olika föreningar samt kommunala institut ger unga möjlighet att studera idrott och kultur samt bl.a. språk och hantverk.
Barn och unga kan delta i grundläggande undervisning i musik, dans, bildkonst och hantverk.
Dessutom erbjuder stadens ungdomstjänster en rockskola.
Stadens ungdomstjänster driver sju ungdomsgårdar runt om i Karleby.
De rusmedels- och rökfria ungdomslokalerna erbjuder handledd verksamhet för barn i årskurserna 3–6 och unga i åldern 13–17 år i olika delar av Karleby.
Information om hobbyverksamheter för barn och unga finns på stadens webbplats.
Rådgivningen vid Ungdomsgården Vinge ger aktuell information om bl.a. internationalisering, studier, arbetsliv, hälsa, hobbyverksamhet och boende.
Karlebynejdens institut erbjuder barn och unga olika former av hobbyverksamhet, exempelvis i konstämnen och musik.
Kontrollera vilka kurser som är aktuella i institutets webbtjänst.
Karleby evangelisk-lutherska församlingar erbjuder även hobbyverksamhet för barn och unga, såsom lekparksträffar, klubbar, musikverksamhet och läger.
Mer information om verksamheten finns på Karleby församlingssammanslutnings webbplats.
Ungdomsgården Vinge
67100 Karleby
Läs mer: Hobbyer för barn och unga.
Övrig undervisning i Karlebyfinska _ svenska
Ungdomstjänsterfinska _ svenska _ engelska
Karlebynejdens institutfinska _ svenska
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
Föreningar
Karleby har ett aktivt och mångsidigt föreningsliv för invånare i alla åldrar.
Läs mer: Föreningar.
Bibliotek
Motion
Att röra sig i naturen
Teater och film
Museer
Hobbyer för barn och unga
Föreningar
Karleby är en gammal sjöstad som erbjuder mångsidiga möjligheter för utfärder och friluftsliv.
Personer ntresserad av friluftsliv bör läsa mer om allemansrätten under rubriken ”Att röra sig i naturen” i denna tjänst.
Flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet.
Föreningar och organisationer samt hobbygrupper och kommunala institut erbjuder kurser i idrott och kultur samt bl.a. språk och hantverk.
I Snellman-salen och i stadens övriga kulturlokaler erbjuds kulturevenemang av varierande slag.
Årliga evenemang i Karleby är bland annat Veneziansk afton i slutet av sommaren, Kokkola Cup för fotbollsjuniorer, Stadsfestivalen Karleby sommarveckor, Lochteå kyrkomusikfest samt Vinterdans i Karleby och festivalen Karleby Vinterharmonika.
Mer information om fritidstjänsterna i Karleby finns på Karleby stads webbplats.
På stadens webbplats finns även en länk till Evenemangskalendern med daglig information om stadens kultur- och motionsevenemang.
Läs mer: Fritid.
Evenemangskalenderfinska
Kulturtjänsterfinska _ svenska _ engelska
Idrottstjänsterfinska _ svenska _ engelska
Bibliotek
Karleby stadsbibliotek finns i stadens centrum.
Närbiblioteken finns i Björkhagen, Kelviå, Lochteå samt Ullava kyrkby och Rahkonen.
Information om bibliotekets öppettider och tjänster finns på dess webbplats.
Biblioteket finns även på nätet.
Där kan kunderna bläddra i bibliotekets samlingar, reservera material, förnya sina lån, beställa fjärrlån och låna e-böcker under alla tider på dygnet.
Tack vare det effektiva biblioteksnätverket i Finland är nästan alla finländska biblioteks samlingar tillgängliga för bibliotekskunderna i Karleby.
Karleby stadsbibliotek/huvudbiblioteket
Storgatan 3, 67100 Karleby
Telefon: 040 806 5124, 040 806 5133
Läs mer: Bibliotek.
Bibliotekstjänsterfinska _ svenska _ engelska
Motion
I Karleby finns mångsidiga motionsmöjligheter året runt.
Staden anordnar ledda aktiviteter i Simcentret VesiVeijari och motionshallarna.
Dessutom finns det gym av flera olika slag.
Gym anpassade för äldre finns i Furuåsens aktivitetscenter och Kuusikumpu servicehus.
Staden underhåller cykelvägar, motionsrutter, joggingbanor, skidspår, badstränder, bollplaner och skridskobanor samt platser för närmotion.
I Karlebynejdens instituts nättjänst finns information om institutets mångsidiga motionsutbud.
I Karleby finns nära på hundra idrottsföreningar för olika grenar samt föreningar som arrangerar övrig motion.
Mer information om motionsmöjligheter i Karleby finns på Karleby stads webbplats.
Läs mer:
Motion.
Idrottstjänsterfinska _ svenska _ engelska
Motionsplatserfinska _ svenska
Gym för äldrefinska
Karlebynejdens institutfinska _ svenska
Att röra sig i naturen
Att röra sig i naturen är en traditionell och populär form av avkoppling för finländarna under alla årstider.
I Finland kan man med stöd av allemansrätten plocka bär och svamp i skogen och röra sig till fots, med cykel eller skidor vintertid.
Det är inte tillåtet att beträda folks gårdar utan lov.
För fiske krävs fiskelov, med undantag för mete och pilkning.
Även jakt fordrar jakttillstånd.
Allemansrätten ger inte rätt att skräpa ner i naturen, skada träd eller växter, störa eller skada fågelbon eller fågelungar, köra motorfordon utan markägarens tillstånd eller bygga ens tillfälliga byggen.
Mer information om motionsrutterna, rastplatser, möjligheter till fiske och båtliv samt exempelvis fågeltorn i Karleby finns på stadens webbplats.
Rutterna för camping, paddling, vandring, cykling och övriga rutter i Karleby finns i karttjänsten på nätet.
I karttjänsten visas även var största delen av motionsplatserna finns.
Du kan köpa friluftskartor över Karleby hos Karleby Turism: Salutorget 5, 67100 Karleby.
Läs mer: Att röra sig i naturen.
linkkiMiljöförvaltningen:
Allemansrättenfinska _ svenska _ engelska _ ryska
Motionskarta över Karlebyfinska _ svenska
Motionsrutter i Karlebyfinska _ svenska
Teater och film
Karleby är en teaterstad med långa anor, som erbjuder scenkonst på hög nivå framförd av både proffs och amatörer.
Karleby stadsteater finns i det stämningsfulla Vartiolinna (Torggatan 48).
Du kan läsa mer om amatörteatrarnas verksamhet på deras webbplats och i evenemangskalendern.
I Karleby finns biografen Bio Rex, vars två salar använder digital- och 3D-teknik.
Bio Rex program finns under länken här intill.
Läs mer: Teater och film.
Stadsteaternfinska
Biograffinska
Teater och danskonst i Karlebyfinska _ svenska _ engelska
Evenemangskalenderfinska
Museer
I hjärtat av staden, i det anrika Rooska gården, finns K.H.Renlunds museum.
Karleby stad grundade museet 1909 utgående från en testamentsgåva av affärsmannen Karl Herman Renlund (1850–1908) .
På museet finns Renlunds samling av finländsk konst från guldåldern och tillfälliga utställningar i en kulturhistorisk miljö.
Även i museikvarterens övriga byggnader finns utställningar om stadens kulturhistoria och utställningar med ITE-konst.
På K.H.Renlunds museums webbplats finns mer information om museets tjänster, utställningar samt aktuell verksamhet.
Utöver K.H.Renlunds museum lönar det sig att besöka det naturhistoriska museet Kieppi (Kieppi är stängt tills vidare på grund av brand) samt de många hembygdsmuseerna och övriga de historiska resmålen i regionen.
Exempelvis i Konst-Vionoja-centret presenteras konstnären Veikko Vionojas verk.
I Kelviå, ca 10 km norrut från Karleby, finns Toivonen djurpark och drängmuseum.
Mer information om dessa museer finns under länkarna här intill.
Läs mer: Museer.
Museer och traditionsarbetefinska _ svenska _ engelska
K.H. Renlunds museum - Mellersta Österbottens landskapsmuseumfinska _ svenska _ engelska
Kieppi, Karleby naturvetenskapliga museumfinska _ svenska _ engelska
linkkiToivonens djurpark och drängmuseum :
Toivonens djurpark och drängmuseum finska _ svenska _ engelska
Konst Vionojafinska
Hobbyer för barn och unga
Flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet.
Flera olika föreningar samt kommunala institut ger unga möjlighet att studera idrott och kultur samt bl.a. språk och hantverk.
Barn och unga kan delta i grundläggande undervisning i musik, dans, bildkonst och hantverk.
Dessutom erbjuder stadens ungdomstjänster en rockskola.
Stadens ungdomstjänster driver sju ungdomsgårdar runt om i Karleby.
De rusmedels- och rökfria ungdomslokalerna erbjuder handledd verksamhet för barn i årskurserna 3–6 och unga i åldern 13–17 år i olika delar av Karleby.
Information om hobbyverksamheter för barn och unga finns på stadens webbplats.
Rådgivningen vid Ungdomsgården Vinge ger aktuell information om bl.a. internationalisering, studier, arbetsliv, hälsa, hobbyverksamhet och boende.
Karlebynejdens institut erbjuder barn och unga olika former av hobbyverksamhet, exempelvis i konstämnen och musik.
Kontrollera vilka kurser som är aktuella i institutets webbtjänst.
Karleby evangelisk-lutherska församlingar erbjuder även hobbyverksamhet för barn och unga, såsom lekparksträffar, klubbar, musikverksamhet och läger.
Mer information om verksamheten finns på Karleby församlingssammanslutnings webbplats.
Ungdomsgården Vinge
67100 Karleby
Läs mer: Hobbyer för barn och unga.
Övrig undervisning i Karlebyfinska _ svenska
Ungdomstjänsterfinska _ svenska _ engelska
Karlebynejdens institutfinska _ svenska
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
Föreningar
Karleby har ett aktivt och mångsidigt föreningsliv för invånare i alla åldrar.
Läs mer: Föreningar.
Problem med uppehållstillstånd
Brott
Våld
Diskriminering och rasism
Behöver du en jurist?
Död
Problem i äktenskap eller parförhållande
Skilsmässa
Problem med den mentala hälsan
Missbruksproblem
I en krissituation kan du ringa nödcentralen på numret 112.
De slussar vid behov dig vidare till socialjouren.
Du ska endast ringa nödcentralen i brådskande nödsituationer, där liv, egendom eller miljön är i fara.
Problem med uppehållstillstånd
Om du har problem eller oklarheter med ditt uppehållstillstånd kan du kontakta Migrationsverket.
Migrationsverket
Korsholmsesplanaden 45
Vasa
Läs mer: Problem med uppehållstillstånd.
Brott
Om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112.
Ring inte nödnumret om det inte är fråga om en nödsituation.
Du kan göra en polisanmälan på nätet.
Mer information finns på Polisens webbplats.
Du kan även skriva ut anmälningsblanketten på nätet och lämna in den till polisstationen.
Karleby polisstation
Karlebygatan 74
67100 Karleby
Läs mer: Brott.
Tidsbokningfinska _ svenska _ engelska
Polisamälanfinska _ svenska _ engelska
Våld
Om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112.
Läs mer: Våld.
Diskriminering och rasism
Om du misstänker att du blivit utsatt för diskriminering då du sökt arbete eller på arbetsplatsen ska du först ta upp detta på din arbetsplats.
Om saken inte kan lösas på arbetsplatsen ska du kontakta arbetarskyddet vid Regionförvaltningsverket i Västra och Inre Finland.
Besöksadress:
Regionförvaltningsverket i Västra och Inre Finland
Wollfskavägen 35
65101 Vasa
Telefon: 0295 018 450
Om du utsätts för diskriminering kan du be om hjälp av Diskrimineringsombudsmannen.
Om du fallit offer för ett rasistiskt motiverat brott kan du göra en polisanmälan på nätet eller polisstationen.
Läs mer: Diskriminering och rasism.
linkkiRegionförvaltningsverket i Västra och Inre Finland:
Regionförvaltningsverket i Västra och Inre Finlandfinska _ svenska _ engelska
Hjälp och information för personer som drabbats av etnisk diskrimineringfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Behöver du en jurist?
Juridiska tjänster är avgiftsbelagda men om du har små eller medelstora inkomster, kan du få helt eller delvis avgiftsfri rättshjälp från statens rättshjälpsbyrå.
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
Besöksadress: Ämbetshuset, Torggatan 40, 67100 Karleby
Telefon: 029 566 1270
Information om enskilda jurister finns bland annat på Finlands Advokatförbunds webbplats.
Läs mer:
Behöver du en jurist?
linkkiFinlands advokatförbund:
Finlands advokatförbundfinska _ svenska _ engelska
Död
Den evangelisk-lutherska kyrkans församlingars begravningsplatser fungerar som allmänna begravningsplatser.
Där kan även avlidna som inte är medlemmar i kyrkan begravas.
De är alltså avsedda för alla invånare i staden.
Mer information finns på Karleby kyrkliga samfällighets webbplats.
Om en närstående plötsligt dör kan du söka krishjälp vid din egen hälsostation, eller utanför tjänstetid vid samjouren för Mellersta Österbottens centralsjukhus.
De evangelisk-lutherska församlingarna i Karlebynejden erbjuder även sorggrupper.
Även församlingarnas diakonimottagningar erbjuder samtalshjälp för sorgearbetet.
Läs mer: Död.
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Problem i äktenskap eller parförhållande
Vid problem i äktenskap eller parförhållande får du hjälp av Mellersta Österbottens familjerådgivningscentral som underhålls av Karleby kyrkliga samfällighets och Mellersta Österbottens social- och hälsovårdssamkommun Soites familjerådgivning.
Familjerågivningscentralen
Telefon: 050 3147 464.
Karleby familjerådgivning
67100 Karleby
tel. 044 730 7640
Läs mer: Problem i äktenskap eller parförhållande.
linkkiMellersta Österbottens Familjerådgivningscentral:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
Skilsmässa
Skilsmässa kan sökas av kvinnan, av mannen eller av båda makarna tillsammans.
Man ansöker om skilsmässa i tingsrätten.
Till att börja med görs en skriftlig skilsmässoansökan.
Österbottens tingsrätt Karleby kansli
Besöksadress: Karlebygatan 27, 67100 Karleby
Telefon: 029 56 49294
Läs mer: Skilsmässa.
Hälsovårdaren på barnrådgivningsbyrån ger råd i frågor som gäller små barns hälsa, tillväxt och utveckling.
Barnrådgivningsbyrån ger information om platser som erbjuder hjälp vid behov.
Vid problem hos unga i skolåldern hjälper exempelvis skolans hälsovårdare eller skolkuratorn.
Läs mer: Barns och ungas problem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Skolhälsovårdfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barnrådgivningarfinska _ svenska
Du kan ta upp problem med hälsovårdaren på skolan eller studieplatsen eller vuxna på ungdomsgården.
Mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats.
Föräldrar eller unga själva kan kontakta familjerådgivningen.
Där kan man tala om problem och få hjälp och stöd.
Mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats.
Familjerådgivningens telefonnummer: 044 730 7640.
Läs mer: Barns och ungas problem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Studerandehälsovårdfinska _ svenska
Ungdomsgårdar och -lokaler finska _ svenska
Problem med den mentala hälsan
Om du behöver hjälp och stöd för din mentala hälsa kan du boka en läkartid vid hälsostationen.
Läkaren bedömer situationen.
Vid behov skriver läkaren en remiss till psykiatrisk specialsjukvård.
Läs mer: Mental hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Mentalvårdstjänsterfinska _ svenska
Om du har ekonomiska problem kan du be om råd hos Mellersta Österbottens social- och hälsovårdssamkommun Soites enheter för socialarbete eller utkomststöd, tfn 040 806 5095 eller tjänstestyrningen, tfn 040 806 5093.
Om du har problem med skulder, kontakta rättshjälpsbyrån.
Du kan anlita vilken som helst rättshjälpsbyrå oberoende av din hemkommun.
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
Telefon: 029 566 1270
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Servicehandledningfinska _ svenska
Missbruksproblem
Om du har problem med alkohol, droger, läkemedel eller hasardspel kan du få vård och rehabilitering vid Porten, Mellersta Österbottens social- och hälsovårdssamkommun Soites center för missbruksproblem.
Du kan ta upp problemet med proffs inom hälsovården eller företagshälsovården, som kan slussa dig vidare i vårdsystemet, eller direkt kontakta Soites missbrukstjänster, tfn 040 8068 101.
För tillnyktrings- och avgiftningsvård debiteras en patientavgift liksom även för korttidsrehabilitering, öppen rehabilitering är gratis.
Även Karleby evangelisk-lutherska församlingssammanslutnings specialdiakoner erbjuder samtalshjälp vid missbruksproblem.
Kontaktuppgifter
Hälsovägen 4
67200 Karleby
Telefon: 040 806 8101
Läs mer: Missbruksproblem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Service för missbrukarefinska _ svenska
linkkiKarleby evangelisk-lutherska församlingssammansutning:
Karleby evangelisk-lutherska församlings arbete bland missbrukarefinska _ svenska
Problem med uppehållstillstånd
Brott
Våld
Diskriminering och rasism
Behöver du en jurist?
Död
Problem i äktenskap eller parförhållande
Skilsmässa
Problem med den mentala hälsan
Missbruksproblem
I en krissituation kan du ringa nödcentralen på numret 112.
De slussar vid behov dig vidare till socialjouren.
Du ska endast ringa nödcentralen i brådskande nödsituationer, där liv, egendom eller miljön är i fara.
Problem med uppehållstillstånd
Om du har problem eller oklarheter med ditt uppehållstillstånd kan du kontakta Migrationsverket.
Migrationsverket
Korsholmsesplanaden 45
Vasa
Läs mer: Problem med uppehållstillstånd.
Brott
Om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112.
Ring inte nödnumret om det inte är fråga om en nödsituation.
Du kan göra en polisanmälan på nätet.
Mer information finns på Polisens webbplats.
Du kan även skriva ut anmälningsblanketten på nätet och lämna in den till polisstationen.
Karleby polisstation
Karlebygatan 74
67100 Karleby
Läs mer: Brott.
Tidsbokningfinska _ svenska _ engelska
Polisamälanfinska _ svenska _ engelska
Våld
Om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112.
Läs mer: Våld.
Diskriminering och rasism
Om du misstänker att du blivit utsatt för diskriminering då du sökt arbete eller på arbetsplatsen ska du först ta upp detta på din arbetsplats.
Om saken inte kan lösas på arbetsplatsen ska du kontakta arbetarskyddet vid Regionförvaltningsverket i Västra och Inre Finland.
Besöksadress:
Regionförvaltningsverket i Västra och Inre Finland
Wollfskavägen 35
65101 Vasa
Telefon: 0295 018 450
Om du utsätts för diskriminering kan du be om hjälp av Diskrimineringsombudsmannen.
Om du fallit offer för ett rasistiskt motiverat brott kan du göra en polisanmälan på nätet eller polisstationen.
Läs mer: Diskriminering och rasism.
linkkiRegionförvaltningsverket i Västra och Inre Finland:
Regionförvaltningsverket i Västra och Inre Finlandfinska _ svenska _ engelska
Hjälp och information för personer som drabbats av etnisk diskrimineringfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Behöver du en jurist?
Juridiska tjänster är avgiftsbelagda men om du har små eller medelstora inkomster, kan du få helt eller delvis avgiftsfri rättshjälp från statens rättshjälpsbyrå.
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
Besöksadress: Ämbetshuset, Torggatan 40, 67100 Karleby
Telefon: 029 566 1270
Information om enskilda jurister finns bland annat på Finlands Advokatförbunds webbplats.
Läs mer:
Behöver du en jurist?
linkkiFinlands advokatförbund:
Finlands advokatförbundfinska _ svenska _ engelska
Död
Den evangelisk-lutherska kyrkans församlingars begravningsplatser fungerar som allmänna begravningsplatser.
Där kan även avlidna som inte är medlemmar i kyrkan begravas.
De är alltså avsedda för alla invånare i staden.
Mer information finns på Karleby kyrkliga samfällighets webbplats.
Om en närstående plötsligt dör kan du söka krishjälp vid din egen hälsostation, eller utanför tjänstetid vid samjouren för Mellersta Österbottens centralsjukhus.
De evangelisk-lutherska församlingarna i Karlebynejden erbjuder även sorggrupper.
Även församlingarnas diakonimottagningar erbjuder samtalshjälp för sorgearbetet.
Läs mer: Död.
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Problem i äktenskap eller parförhållande
Vid problem i äktenskap eller parförhållande får du hjälp av Mellersta Österbottens familjerådgivningscentral som underhålls av Karleby kyrkliga samfällighets och Mellersta Österbottens social- och hälsovårdssamkommun Soites familjerådgivning.
Familjerågivningscentralen
Telefon: 050 3147 464.
Karleby familjerådgivning
67100 Karleby
tel. 044 730 7640
Läs mer: Problem i äktenskap eller parförhållande.
linkkiMellersta Österbottens Familjerådgivningscentral:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
Skilsmässa
Skilsmässa kan sökas av kvinnan, av mannen eller av båda makarna tillsammans.
Man ansöker om skilsmässa i tingsrätten.
Till att börja med görs en skriftlig skilsmässoansökan.
Österbottens tingsrätt Karleby kansli
Besöksadress: Karlebygatan 27, 67100 Karleby
Telefon: 029 56 49294
Läs mer: Skilsmässa.
Hälsovårdaren på barnrådgivningsbyrån ger råd i frågor som gäller små barns hälsa, tillväxt och utveckling.
Barnrådgivningsbyrån ger information om platser som erbjuder hjälp vid behov.
Vid problem hos unga i skolåldern hjälper exempelvis skolans hälsovårdare eller skolkuratorn.
Läs mer: Barns och ungas problem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Skolhälsovårdfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barnrådgivningarfinska _ svenska
Du kan ta upp problem med hälsovårdaren på skolan eller studieplatsen eller vuxna på ungdomsgården.
Mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats.
Föräldrar eller unga själva kan kontakta familjerådgivningen.
Där kan man tala om problem och få hjälp och stöd.
Mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats.
Familjerådgivningens telefonnummer: 044 730 7640.
Läs mer: Barns och ungas problem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Studerandehälsovårdfinska _ svenska
Ungdomsgårdar och -lokaler finska _ svenska
Problem med den mentala hälsan
Om du behöver hjälp och stöd för din mentala hälsa kan du boka en läkartid vid hälsostationen.
Läkaren bedömer situationen.
Vid behov skriver läkaren en remiss till psykiatrisk specialsjukvård.
Läs mer: Mental hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Mentalvårdstjänsterfinska _ svenska
Om du har ekonomiska problem kan du be om råd hos Mellersta Österbottens social- och hälsovårdssamkommun Soites enheter för socialarbete eller utkomststöd, tfn 040 806 5095 eller tjänstestyrningen, tfn 040 806 5093.
Om du har problem med skulder, kontakta rättshjälpsbyrån.
Du kan anlita vilken som helst rättshjälpsbyrå oberoende av din hemkommun.
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
Telefon: 029 566 1270
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Servicehandledningfinska _ svenska
Missbruksproblem
Om du har problem med alkohol, droger, läkemedel eller hasardspel kan du få vård och rehabilitering vid Porten, Mellersta Österbottens social- och hälsovårdssamkommun Soites center för missbruksproblem.
Du kan ta upp problemet med proffs inom hälsovården eller företagshälsovården, som kan slussa dig vidare i vårdsystemet, eller direkt kontakta Soites missbrukstjänster, tfn 040 8068 101.
För tillnyktrings- och avgiftningsvård debiteras en patientavgift liksom även för korttidsrehabilitering, öppen rehabilitering är gratis.
Även Karleby evangelisk-lutherska församlingssammanslutnings specialdiakoner erbjuder samtalshjälp vid missbruksproblem.
Kontaktuppgifter
Hälsovägen 4
67200 Karleby
Telefon: 040 806 8101
Läs mer: Missbruksproblem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Service för missbrukarefinska _ svenska
linkkiKarleby evangelisk-lutherska församlingssammansutning:
Karleby evangelisk-lutherska församlings arbete bland missbrukarefinska _ svenska
Problem med uppehållstillstånd
Brott
Våld
Diskriminering och rasism
Behöver du en jurist?
Död
Problem i äktenskap eller parförhållande
Skilsmässa
Problem med den mentala hälsan
Missbruksproblem
I en krissituation kan du ringa nödcentralen på numret 112.
De slussar vid behov dig vidare till socialjouren.
Du ska endast ringa nödcentralen i brådskande nödsituationer, där liv, egendom eller miljön är i fara.
Problem med uppehållstillstånd
Om du har problem eller oklarheter med ditt uppehållstillstånd kan du kontakta Migrationsverket.
Migrationsverket
Korsholmsesplanaden 45
Vasa
Läs mer: Problem med uppehållstillstånd.
Brott
Om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112.
Ring inte nödnumret om det inte är fråga om en nödsituation.
Du kan göra en polisanmälan på nätet.
Mer information finns på Polisens webbplats.
Du kan även skriva ut anmälningsblanketten på nätet och lämna in den till polisstationen.
Karleby polisstation
Karlebygatan 74
67100 Karleby
Läs mer: Brott.
Tidsbokningfinska _ svenska _ engelska
Polisamälanfinska _ svenska _ engelska
Våld
Om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112.
Läs mer: Våld.
Diskriminering och rasism
Om du misstänker att du blivit utsatt för diskriminering då du sökt arbete eller på arbetsplatsen ska du först ta upp detta på din arbetsplats.
Om saken inte kan lösas på arbetsplatsen ska du kontakta arbetarskyddet vid Regionförvaltningsverket i Västra och Inre Finland.
Besöksadress:
Regionförvaltningsverket i Västra och Inre Finland
Wollfskavägen 35
65101 Vasa
Telefon: 0295 018 450
Om du utsätts för diskriminering kan du be om hjälp av Diskrimineringsombudsmannen.
Om du fallit offer för ett rasistiskt motiverat brott kan du göra en polisanmälan på nätet eller polisstationen.
Läs mer: Diskriminering och rasism.
linkkiRegionförvaltningsverket i Västra och Inre Finland:
Regionförvaltningsverket i Västra och Inre Finlandfinska _ svenska _ engelska
Hjälp och information för personer som drabbats av etnisk diskrimineringfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Behöver du en jurist?
Juridiska tjänster är avgiftsbelagda men om du har små eller medelstora inkomster, kan du få helt eller delvis avgiftsfri rättshjälp från statens rättshjälpsbyrå.
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
Besöksadress: Ämbetshuset, Torggatan 40, 67100 Karleby
Telefon: 029 566 1270
Information om enskilda jurister finns bland annat på Finlands Advokatförbunds webbplats.
Läs mer:
Behöver du en jurist?
linkkiFinlands advokatförbund:
Finlands advokatförbundfinska _ svenska _ engelska
Död
Den evangelisk-lutherska kyrkans församlingars begravningsplatser fungerar som allmänna begravningsplatser.
Där kan även avlidna som inte är medlemmar i kyrkan begravas.
De är alltså avsedda för alla invånare i staden.
Mer information finns på Karleby kyrkliga samfällighets webbplats.
Om en närstående plötsligt dör kan du söka krishjälp vid din egen hälsostation, eller utanför tjänstetid vid samjouren för Mellersta Österbottens centralsjukhus.
De evangelisk-lutherska församlingarna i Karlebynejden erbjuder även sorggrupper.
Även församlingarnas diakonimottagningar erbjuder samtalshjälp för sorgearbetet.
Läs mer: Död.
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Problem i äktenskap eller parförhållande
Vid problem i äktenskap eller parförhållande får du hjälp av Mellersta Österbottens familjerådgivningscentral som underhålls av Karleby kyrkliga samfällighets och Mellersta Österbottens social- och hälsovårdssamkommun Soites familjerådgivning.
Familjerågivningscentralen
Telefon: 050 3147 464.
Karleby familjerådgivning
67100 Karleby
tel. 044 730 7640
Läs mer: Problem i äktenskap eller parförhållande.
linkkiMellersta Österbottens Familjerådgivningscentral:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
Skilsmässa
Skilsmässa kan sökas av kvinnan, av mannen eller av båda makarna tillsammans.
Man ansöker om skilsmässa i tingsrätten.
Till att börja med görs en skriftlig skilsmässoansökan.
Österbottens tingsrätt Karleby kansli
Besöksadress: Karlebygatan 27, 67100 Karleby
Telefon: 029 56 49294
Läs mer: Skilsmässa.
Hälsovårdaren på barnrådgivningsbyrån ger råd i frågor som gäller små barns hälsa, tillväxt och utveckling.
Barnrådgivningsbyrån ger information om platser som erbjuder hjälp vid behov.
Vid problem hos unga i skolåldern hjälper exempelvis skolans hälsovårdare eller skolkuratorn.
Läs mer: Barns och ungas problem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Skolhälsovårdfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barnrådgivningarfinska _ svenska
Du kan ta upp problem med hälsovårdaren på skolan eller studieplatsen eller vuxna på ungdomsgården.
Mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats.
Föräldrar eller unga själva kan kontakta familjerådgivningen.
Där kan man tala om problem och få hjälp och stöd.
Mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats.
Familjerådgivningens telefonnummer: 044 730 7640.
Läs mer: Barns och ungas problem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Studerandehälsovårdfinska _ svenska
Ungdomsgårdar och -lokaler finska _ svenska
Problem med den mentala hälsan
Om du behöver hjälp och stöd för din mentala hälsa kan du boka en läkartid vid hälsostationen.
Läkaren bedömer situationen.
Vid behov skriver läkaren en remiss till psykiatrisk specialsjukvård.
Läs mer: Mental hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Mentalvårdstjänsterfinska _ svenska
Om du har ekonomiska problem kan du be om råd hos Mellersta Österbottens social- och hälsovårdssamkommun Soites enheter för socialarbete eller utkomststöd, tfn 040 806 5095 eller tjänstestyrningen, tfn 040 806 5093.
Om du har problem med skulder, kontakta rättshjälpsbyrån.
Du kan anlita vilken som helst rättshjälpsbyrå oberoende av din hemkommun.
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
Telefon: 029 566 1270
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Servicehandledningfinska _ svenska
Missbruksproblem
Om du har problem med alkohol, droger, läkemedel eller hasardspel kan du få vård och rehabilitering vid Porten, Mellersta Österbottens social- och hälsovårdssamkommun Soites center för missbruksproblem.
Du kan ta upp problemet med proffs inom hälsovården eller företagshälsovården, som kan slussa dig vidare i vårdsystemet, eller direkt kontakta Soites missbrukstjänster, tfn 040 8068 101.
För tillnyktrings- och avgiftningsvård debiteras en patientavgift liksom även för korttidsrehabilitering, öppen rehabilitering är gratis.
Även Karleby evangelisk-lutherska församlingssammanslutnings specialdiakoner erbjuder samtalshjälp vid missbruksproblem.
Kontaktuppgifter
Hälsovägen 4
67200 Karleby
Telefon: 040 806 8101
Läs mer: Missbruksproblem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Service för missbrukarefinska _ svenska
linkkiKarleby evangelisk-lutherska församlingssammansutning:
Karleby evangelisk-lutherska församlings arbete bland missbrukarefinska _ svenska
Äktenskap
Skilsmässa
Barn vid skilsmässa
När du väntar barn
Vård av barnet
Vård av barnet i hemmet
Äktenskap
Innan äktenskapet ingås ska du skriftligen be om prövning av äktenskapshinder.
Prövningen görs vid magistraten. Du kan lämna in ansökan om prövning vid vilken magistrat som helst.
Civilvigsel äger rum vid magistraten.
Magistraten i Västra Finland
Karleby enhet
Karlebygatan 27, PB 581
67701 Karleby
Telefon: 029 553 9451
Läs mer:
Äktenskap.
Skilsmässa
Skilsmässa kan sökas av kvinnan, av mannen eller av båda makarna tillsammans.
Man ansöker om skilsmässa i tingsrätten.
Till att börja med görs en skriftlig skilsmässoansökan.
Österbottens tingsrätt Karleby kansli
Besöksadress: Karlebygatan 27, 67100 Karleby
Telefon: 029 56 49294
Läs mer: Skilsmässa.
Barn vid skilsmässa
Om du har barn och går igenom en skilsmässa ska du ta kontakt med barnatillsyningsmannen.
Barnatillsyningsmannen bekräftar överenskommelsen om var barnen ska bo, vården av barnen, umgängesrätt och underhållsbidrag.
Barnatillsyningsmannen
67100 Karleby
Telefontid och tidsbokning
tel. 06 826 4111
Läs mer: Barn vid skilsmässa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barnatillsyningsmannenfinska _ svenska
När du väntar barn
Ta kontakt med rådgivningen då du märker att du är gravid.
På rådgivningen följer man med moderns, barnets och hela familjens välmående under graviditeten.
Du kan be om råd per telefon (06) 826 4477.
Läs mer:
När du väntar barn.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Mödrarådgivningfinska _ svenska
Vård av barnet
I Karleby finns stadens daghem, gruppfamiljedaghem, familjedagvårdare samt barnklubbar.
Dessutom finns det daghem som köptjänst (svenskspråkiga), ett privat daghem och privata familjedagvårdare i Karleby.
Du kan ansöka om plats inom småbarnspedagogiken för ditt barn elektroniskt via tjänsten suomi.fi eller med en blankett på stadens webbplats (ansökan om småbarnspedagogik).
Ansökan ska lämnas in fyra månader innan du behöver plats inom småbarnspedagogiken.
Det är möjligt att få en plats snabbare om den behövs för att du exempelvis erhållit arbete eller studieplats.
Ansökan kan returneras till platsen för småbarnspedagogik, kontorstjänster för småbarnspedagogik eller lämnas i brevlådan i den nedre aulan i Bildningscentralen.
Du kan ansöka om en plats i stadens barnklubbar med blanketten som finns på stadens webbplats.
Ansökan kan även skickas per post till följande adress:
Bildningscentralen
Tjänster för småbarnspedagogik
Strandgatan16
67100 Karleby
Läs mer:
Daghem och andra dagvårdsplatserfinska _ svenska
Gruppfamiljedaghemfinska _ svenska
Dagvårdsblanketterfinska _ svenska
Att ansöka om kommunal dagvårdfinska _ svenska
Vård av barnet i hemmet
Om familjens yngsta barn är yngre än tre år kan föräldern få hemvårdsstöd för vård av barnet i hemmet.
Om du har rätt till stödet kan du ansöka om stödet hos FPA.
Du kan fylla i ansökan på nätet eller skicka den per post till FPA.
Du kan även besöka FPA:s kontor.
Karleby stad betalar extra Karlebystöd för de familjer som tar hand om barn under tre år i hemmet.
Du kan ansöka om Karlebystödet om den ena av föräldrarna vårdar samtliga av familjens barn under skolåldern i hemmet.
Om din familj fyller villkoren, beviljas Karlebystödet i samband med beviljandet av vårdnadsbidraget.
Läs mer:
Stöd för vård av barn i hemmet.
Karlebystödfinska _ svenska
Information om FPA:s hemvårdsstödfinska _ svenska _ engelska
FPA kontaktuppgifterfinska _ svenska _ engelska
Äktenskap
Skilsmässa
Barn vid skilsmässa
När du väntar barn
Vård av barnet
Vård av barnet i hemmet
Äktenskap
Innan äktenskapet ingås ska du skriftligen be om prövning av äktenskapshinder.
Prövningen görs vid magistraten. Du kan lämna in ansökan om prövning vid vilken magistrat som helst.
Civilvigsel äger rum vid magistraten.
Magistraten i Västra Finland
Karleby enhet
Karlebygatan 27, PB 581
67701 Karleby
Telefon: 029 553 9451
Läs mer:
Äktenskap.
Skilsmässa
Skilsmässa kan sökas av kvinnan, av mannen eller av båda makarna tillsammans.
Man ansöker om skilsmässa i tingsrätten.
Till att börja med görs en skriftlig skilsmässoansökan.
Österbottens tingsrätt Karleby kansli
Besöksadress: Karlebygatan 27, 67100 Karleby
Telefon: 029 56 49294
Läs mer: Skilsmässa.
Barn vid skilsmässa
Om du har barn och går igenom en skilsmässa ska du ta kontakt med barnatillsyningsmannen.
Barnatillsyningsmannen bekräftar överenskommelsen om var barnen ska bo, vården av barnen, umgängesrätt och underhållsbidrag.
Barnatillsyningsmannen
67100 Karleby
Telefontid och tidsbokning
tel. 06 826 4111
Läs mer: Barn vid skilsmässa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barnatillsyningsmannenfinska _ svenska
När du väntar barn
Ta kontakt med rådgivningen då du märker att du är gravid.
På rådgivningen följer man med moderns, barnets och hela familjens välmående under graviditeten.
Du kan be om råd per telefon (06) 826 4477.
Läs mer:
När du väntar barn.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Mödrarådgivningfinska _ svenska
Vård av barnet
I Karleby finns stadens daghem, gruppfamiljedaghem, familjedagvårdare samt barnklubbar.
Dessutom finns det daghem som köptjänst (svenskspråkiga), ett privat daghem och privata familjedagvårdare i Karleby.
Du kan ansöka om plats inom småbarnspedagogiken för ditt barn elektroniskt via tjänsten suomi.fi eller med en blankett på stadens webbplats (ansökan om småbarnspedagogik).
Ansökan ska lämnas in fyra månader innan du behöver plats inom småbarnspedagogiken.
Det är möjligt att få en plats snabbare om den behövs för att du exempelvis erhållit arbete eller studieplats.
Ansökan kan returneras till platsen för småbarnspedagogik, kontorstjänster för småbarnspedagogik eller lämnas i brevlådan i den nedre aulan i Bildningscentralen.
Du kan ansöka om en plats i stadens barnklubbar med blanketten som finns på stadens webbplats.
Ansökan kan även skickas per post till följande adress:
Bildningscentralen
Tjänster för småbarnspedagogik
Strandgatan16
67100 Karleby
Läs mer:
Daghem och andra dagvårdsplatserfinska _ svenska
Gruppfamiljedaghemfinska _ svenska
Dagvårdsblanketterfinska _ svenska
Att ansöka om kommunal dagvårdfinska _ svenska
Vård av barnet i hemmet
Om familjens yngsta barn är yngre än tre år kan föräldern få hemvårdsstöd för vård av barnet i hemmet.
Om du har rätt till stödet kan du ansöka om stödet hos FPA.
Du kan fylla i ansökan på nätet eller skicka den per post till FPA.
Du kan även besöka FPA:s kontor.
Karleby stad betalar extra Karlebystöd för de familjer som tar hand om barn under tre år i hemmet.
Du kan ansöka om Karlebystödet om den ena av föräldrarna vårdar samtliga av familjens barn under skolåldern i hemmet.
Om din familj fyller villkoren, beviljas Karlebystödet i samband med beviljandet av vårdnadsbidraget.
Läs mer:
Stöd för vård av barn i hemmet.
Karlebystödfinska _ svenska
Information om FPA:s hemvårdsstödfinska _ svenska _ engelska
FPA kontaktuppgifterfinska _ svenska _ engelska
Äktenskap
Skilsmässa
Barn vid skilsmässa
När du väntar barn
Vård av barnet
Vård av barnet i hemmet
Äktenskap
Innan äktenskapet ingås ska du skriftligen be om prövning av äktenskapshinder.
Prövningen görs vid magistraten. Du kan lämna in ansökan om prövning vid vilken magistrat som helst.
Civilvigsel äger rum vid magistraten.
Magistraten i Västra Finland
Karleby enhet
Karlebygatan 27, PB 581
67701 Karleby
Telefon: 029 553 9451
Läs mer:
Äktenskap.
Skilsmässa
Skilsmässa kan sökas av kvinnan, av mannen eller av båda makarna tillsammans.
Man ansöker om skilsmässa i tingsrätten.
Till att börja med görs en skriftlig skilsmässoansökan.
Österbottens tingsrätt Karleby kansli
Besöksadress: Karlebygatan 27, 67100 Karleby
Telefon: 029 56 49294
Läs mer: Skilsmässa.
Barn vid skilsmässa
Om du har barn och går igenom en skilsmässa ska du ta kontakt med barnatillsyningsmannen.
Barnatillsyningsmannen bekräftar överenskommelsen om var barnen ska bo, vården av barnen, umgängesrätt och underhållsbidrag.
Barnatillsyningsmannen
67100 Karleby
Telefontid och tidsbokning
tel. 06 826 4111
Läs mer: Barn vid skilsmässa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barnatillsyningsmannenfinska _ svenska
När du väntar barn
Ta kontakt med rådgivningen då du märker att du är gravid.
På rådgivningen följer man med moderns, barnets och hela familjens välmående under graviditeten.
Du kan be om råd per telefon (06) 826 4477.
Läs mer: Graviditet och förlossning.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Mödrarådgivningfinska _ svenska
Vård av barnet
I Karleby finns stadens daghem, gruppfamiljedaghem, familjedagvårdare samt barnklubbar.
Dessutom finns det daghem som köptjänst (svenskspråkiga), ett privat daghem och privata familjedagvårdare i Karleby.
Du kan ansöka om plats inom småbarnspedagogiken för ditt barn elektroniskt via tjänsten suomi.fi eller med en blankett på stadens webbplats (ansökan om småbarnspedagogik).
Ansökan ska lämnas in fyra månader innan du behöver plats inom småbarnspedagogiken.
Det är möjligt att få en plats snabbare om den behövs för att du exempelvis erhållit arbete eller studieplats.
Ansökan kan returneras till platsen för småbarnspedagogik, kontorstjänster för småbarnspedagogik eller lämnas i brevlådan i den nedre aulan i Bildningscentralen.
Du kan ansöka om en plats i stadens barnklubbar med blanketten som finns på stadens webbplats.
Ansökan kan även skickas per post till följande adress:
Bildningscentralen
Tjänster för småbarnspedagogik
Strandgatan16
67100 Karleby
Läs mer:
Vård av barnet.
Daghem och andra dagvårdsplatserfinska _ svenska
Gruppfamiljedaghemfinska _ svenska
Dagvårdsblanketterfinska _ svenska
Att ansöka om kommunal dagvårdfinska _ svenska
Vård av barnet i hemmet
Om familjens yngsta barn är yngre än tre år kan föräldern få hemvårdsstöd för vård av barnet i hemmet.
Om du har rätt till stödet kan du ansöka om stödet hos FPA.
Du kan fylla i ansökan på nätet eller skicka den per post till FPA.
Du kan även besöka FPA:s kontor.
Karleby stad betalar extra Karlebystöd för de familjer som tar hand om barn under tre år i hemmet.
Du kan ansöka om Karlebystödet om den ena av föräldrarna vårdar samtliga av familjens barn under skolåldern i hemmet.
Om din familj fyller villkoren, beviljas Karlebystödet i samband med beviljandet av vårdnadsbidraget.
Läs mer:
Stöd för vård av barn i hemmet.
Karlebystödfinska _ svenska
Information om FPA:s hemvårdsstödfinska _ svenska _ engelska
FPA kontaktuppgifterfinska _ svenska _ engelska
Hälsovårdstjänster i Karleby
Äldre människors hälsa
Tandvård
Mental hälsa
Sexuell hälsa
När du väntar barn
Förlossning
Läkemedel
Handikappade personer
Ett handikappat barn
Hälsovårdstjänster i Karleby
I Karleby finns hälsostationer i olika delar av staden.
Varje hälsostation har ett eget telefonnummer för tidsbokning, som man kan ringa för att boka tid till sjukskötare eller läkare.
Kontaktuppgifter:
Karleby huvudhälsostation
Mariegatan 28
67200 Karleby
Telefon: (06) 8287 580
På Karleby huvudhälsostationen styrs patienterna till mottagningen på basis av hur akuta deras symptom är.
Klienten får en tid till akutvården, mottagningen eller Min Soite-mottagningen.
Samtal till huvudhälsostationen styrs till ett och samma telefonnummer, (06) 8287 310.
67800 Karleby
Telefon: (06) 8287 580
Mottagning /Kelviå
Ellfolkgatan 5
68300 Kelviå
Telefon: (06) 8287 701
Mottagning /Lochteå
Telefon: (06) 8287 750
Mottagning /Ullava
Ullavavägen 701
68370 Ullava
Telefon: (06) 8287 639
Om du kommer som flykting till Finland ska du komma överens om en hälsokontroll med Utlänningsbyrån.
Läs mer: Hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
Under kvällar och helger är hälsostationerna stängda.
Då hanteras plötsliga sjukdomar och olyckor vid jouren.
Jouren är avsedd för patienter vars sjukdom kräver brådskande bedömning och vård.
I livshotande situationer ska du ringa nödnumret 112.
Om du besöker jouren kvällstid eller under helger ska du först ringa jourens telefonrådgivning (06) 826 4500.
Samjourens adress:
Mellersta Österbottens centralsjukhus
Mariegatan 16–20 (l-flygeln, ingång B1)
67200 Karleby
Läs mer: Hälsovårdstjänster i Finland
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barns hälsa
Om ditt barn insjuknar ska du kontakta hälsostationen vid behov.
ådgivningarna erbjuder tjänster för gravida och barn under skolåldern.
Vid rådgivningarna utförs vaccinationer av barn och vuxna.
Du kan kontakta rådgivningen via den centraliserade telefontjänsten (06) 826 4477.
Genom regelbundna besök på barnrådgivningsbyrån följs barnets hälsa, tillväxt och utveckling upp.
På rådgivningen vårdas inte barn som insjuknar plötsligt, men du kan be om råd via den centraliserade telefontjänsten (06) 826 4477.
Skolhälsovårdaren har hand om skolelevers hälsa.
Mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats.
Läs mer: Barns hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barnrådgivningarfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Rådgivningarfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Skolhälsovårdfinska _ svenska
Äldre människors hälsa
Vid hälsopunkten Daalia ges vägledning och rådgivning för personer över 65 år om diet, motion och livsstil.
Vaccinering av personer över 65 år utförs vid seniorrådgivning.
Läs mer:
Äldre människors hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Seniorernas hälsopunkterfinska _ svenska
Tandvård
Om du behöver icke-brådskande tandvård ska du ringa munhälsans centraliserade tidsbokningen.
Centraliserad tidsbokning per telefon: (06) 8287 400
Huvudhälsostationens tandklinik
Mariegatan 28, 67200 Karleby
Björkhagens tandklinik
Storkisbackens tandklinik
Korpvägen 11, 67100 Karleby
Kelviå tandklinik
Ellfolkgatan 5, 68300, Kelviå
Lochteå tandklinik
Ullava tandklinik
Ullavavägen 701, 68370 Ullava
Vardagar kan tider till smärtjouren bokas enligt överenskommelse vid samtliga tandkliniker.
Brådskande tandvård/första hjälpen (kvälls-, vardags-, helg- och nattjour):
Vid smärtjouren får du första hjälpen vid plötslig tandvärk och tandolyckor.
Tandläkarjouren (kvälls-, vardags- och helgjour) ordnas vid polikliniken för tand- och munsjukdomar vid Mellersta Österbottens social- och hälsovårdssamkommun Soite, Mariegatan 16–20, 67200 Karleby (vån 1, del D), vardagkvällar kl. 16.00–21.00 samt veckoslut och helgdagar kl. 8.00–21.00.
Du kan i regel komma till jourmottagningen genom att först kontakta jouren via telefon.
För frågor gällande jouren ring tel. (06) 828 7450.
När du kommer till jourmottagningen ska du ta en kölapp, såvida du inte har en bokad tid.
Brådskande tandvård/första hjälpen (nattjour):
Allvarliga fall i samjour Uleåborgs universitetssjukhus (Oulun yliopistollinen sairaala OYS) kl. 21.00−8.00, tel. (08) 315 2655
Läs mer: Tandvård.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Munhälsovårdenfinska _ svenska
Mental hälsa
Vid problem med din mentala hälsa ska du i första hand kontakta din egen hälsostation eller företagshälsovårdens mottagning.
Vid brådskande problem, kontakta hälsovårdcentralens jour.
Läs mer: Mental hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
Sexuell hälsa
Om du känner att du behöver information om familjeplanering och prevention kan du kontakta din egen hälsostation.
Boka tid till hälsostationen om du behöver preventivmedel, överväger att göra en abort eller misstänker att du lider av en könssjukdom.
Du kan även boka en tid hos en allmänläkare för en gynekologisk eller urologisk undersökning.
I preventionsfrågor kan du kontakta den centraliserade telefontjänsten (06) 826 4477.
Läs mer:
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Preventivrådgivningfinska _ svenska
När du väntar barn
Ta kontakt med rådgivningen då du märker att du är gravid.
På rådgivningen följer man med moderns, barnets och hela familjens välmående under graviditeten.
Läs mer:
När du väntar barn.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Mödrarådgivningfinska _ svenska
Förlossning
Förlossningsavdelningen är öppen dygnet runt.
Om du önskar kan du ringa förlossningsavdelning då din förlossning satt igång eller om du vill fråga om råd.
Då du kommer till sjukhuset ska du använda centralsjukhusets huvudingång kl. 7–20 och övriga tider bör du använda den gemensamma jourens/poliklinikens dörr.
Kontaktuppgifter för förlossningsavdelningen:
Mariegatan 16–20,
67200 Karleby
Telefon: (06) 8264355.
Läs mer: Förlossning.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Förlossningarfinska _ svenska
Läkemedel
Du kan köpa läkemedel på apoteket.
Du kan besöka vilket apotek som helst.
Du kan även besöka apotek som inte finns i din egen kommun.
Läs mer: Läkemedel.
Handikappade personer
En handikappad person bosatt i Karleby har rätt att erhålla de tjänster han eller hon behöver på samma grunder som de övriga invånarna i kommunen.
Personen kan dock på grund av sitt handikapp eller sin sjukdom även behöva särskilda tjänster för handikappade för att klara vardagen.
För tjänsterna för handikappade i Karleby svarar Mellersta Österbottens social- och hälsovårdssamkommun Soite, där man kan ansöka om tjänster och stödfunktioner.
Tjänster av flera olika slag erbjuds även för personer med gravt handikapp.
Dessa tjänster inkluderar bland annat:
transporttjänster
ombyggnad och nödvändig utrustning för hemmet
maskiner och utrustning
personlig hjälp och dagverksamhet
stödboende
stöd för närståendevård av personer under 65 och arbetsverksamhet.
Dessutom är det möjligt att ansöka om specialboende, korttidsvård eller tillfällig vård samt handledning hos den öppna vården.
Mer information om tjänster för handikappade får du från Mellersta Österbottens social- och hälsovårdssamkommun Soites handikapptjänster per telefon: 040 804 2122.
Läs mer: Handikappade personer.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Tjänster för handikappadefinska _ svenska
Specialpedagogik i förskolanfinska _ svenska
Kontaktuppgifter för den grundläggande utbildningenfinska
Ett handikappat barn
Särskilt stöd erbjuds barn med handikapp inom småbarnspedagogiken och skolan.
Kontakta Karleby stads förskoleundervisning för information om specialsmåbarnspedagogiken.
Du kan be undervisningsväsendet om mer information om tjänster som skolan erbjuder.
Bildningscentralen
Strandgatan 16 (våning 5 och 6)
67100 Karleby
Telefon: 040 8065 149
Läs mer: Ett handikappat barn.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Tjänster för handikappadefinska _ svenska
Specialpedagogik i förskolanfinska _ svenska
Kontaktuppgifter för den grundläggande utbildningenfinska
Hälsovårdstjänster i Karleby
Äldre människors hälsa
Tandvård
Mental hälsa
Sexuell hälsa
När du väntar barn
Förlossning
Läkemedel
Handikappade personer
Ett handikappat barn
Hälsovårdstjänster i Karleby
I Karleby finns hälsostationer i olika delar av staden.
Varje hälsostation har ett eget telefonnummer för tidsbokning, som man kan ringa för att boka tid till sjukskötare eller läkare.
Kontaktuppgifter:
Karleby huvudhälsostation
Mariegatan 28
67200 Karleby
Telefon: (06) 8287 580
På Karleby huvudhälsostationen styrs patienterna till mottagningen på basis av hur akuta deras symptom är.
Klienten får en tid till akutvården, mottagningen eller Min Soite-mottagningen.
Samtal till huvudhälsostationen styrs till ett och samma telefonnummer, (06) 8287 310.
67800 Karleby
Telefon: (06) 8287 580
Mottagning /Kelviå
Ellfolkgatan 5
68300 Kelviå
Telefon: (06) 8287 701
Mottagning /Lochteå
Telefon: (06) 8287 750
Mottagning /Ullava
Ullavavägen 701
68370 Ullava
Telefon: (06) 8287 639
Om du kommer som flykting till Finland ska du komma överens om en hälsokontroll med Utlänningsbyrån.
Läs mer: Hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
Under kvällar och helger är hälsostationerna stängda.
Då hanteras plötsliga sjukdomar och olyckor vid jouren.
Jouren är avsedd för patienter vars sjukdom kräver brådskande bedömning och vård.
I livshotande situationer ska du ringa nödnumret 112.
Om du besöker jouren kvällstid eller under helger ska du först ringa jourens telefonrådgivning (06) 826 4500.
Samjourens adress:
Mellersta Österbottens centralsjukhus
Mariegatan 16–20 (l-flygeln, ingång B1)
67200 Karleby
Läs mer: Hälsovårdstjänster i Finland
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barns hälsa
Om ditt barn insjuknar ska du kontakta hälsostationen vid behov.
ådgivningarna erbjuder tjänster för gravida och barn under skolåldern.
Vid rådgivningarna utförs vaccinationer av barn och vuxna.
Du kan kontakta rådgivningen via den centraliserade telefontjänsten (06) 826 4477.
Genom regelbundna besök på barnrådgivningsbyrån följs barnets hälsa, tillväxt och utveckling upp.
På rådgivningen vårdas inte barn som insjuknar plötsligt, men du kan be om råd via den centraliserade telefontjänsten (06) 826 4477.
Skolhälsovårdaren har hand om skolelevers hälsa.
Mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats.
Läs mer: Barns hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barnrådgivningarfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Rådgivningarfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Skolhälsovårdfinska _ svenska
Äldre människors hälsa
Vid hälsopunkten Daalia ges vägledning och rådgivning för personer över 65 år om diet, motion och livsstil.
Vaccinering av personer över 65 år utförs vid seniorrådgivning.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Seniorernas hälsopunkterfinska _ svenska
Tandvård
Om du behöver icke-brådskande tandvård ska du ringa munhälsans centraliserade tidsbokningen.
Centraliserad tidsbokning per telefon: (06) 8287 400
Huvudhälsostationens tandklinik
Mariegatan 28, 67200 Karleby
Björkhagens tandklinik
Storkisbackens tandklinik
Korpvägen 11, 67100 Karleby
Kelviå tandklinik
Ellfolkgatan 5, 68300, Kelviå
Lochteå tandklinik
Ullava tandklinik
Ullavavägen 701, 68370 Ullava
Vardagar kan tider till smärtjouren bokas enligt överenskommelse vid samtliga tandkliniker.
Brådskande tandvård/första hjälpen (kvälls-, vardags-, helg- och nattjour):
Vid smärtjouren får du första hjälpen vid plötslig tandvärk och tandolyckor.
Tandläkarjouren (kvälls-, vardags- och helgjour) ordnas vid polikliniken för tand- och munsjukdomar vid Mellersta Österbottens social- och hälsovårdssamkommun Soite, Mariegatan 16–20, 67200 Karleby (vån 1, del D), vardagkvällar kl. 16.00–21.00 samt veckoslut och helgdagar kl. 8.00–21.00.
Du kan i regel komma till jourmottagningen genom att först kontakta jouren via telefon.
För frågor gällande jouren ring tel. (06) 828 7450.
När du kommer till jourmottagningen ska du ta en kölapp, såvida du inte har en bokad tid.
Brådskande tandvård/första hjälpen (nattjour):
Allvarliga fall i samjour Uleåborgs universitetssjukhus (Oulun yliopistollinen sairaala OYS) kl. 21.00−8.00, tel. (08) 315 2655
Läs mer: Tandvård.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Munhälsovårdenfinska _ svenska
Mental hälsa
Vid problem med din mentala hälsa ska du i första hand kontakta din egen hälsostation eller företagshälsovårdens mottagning.
Vid brådskande problem, kontakta hälsovårdcentralens jour.
Läs mer: Mental hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
Sexuell hälsa
Om du känner att du behöver information om familjeplanering och prevention kan du kontakta din egen hälsostation.
Boka tid till hälsostationen om du behöver preventivmedel, överväger att göra en abort eller misstänker att du lider av en könssjukdom.
Du kan även boka en tid hos en allmänläkare för en gynekologisk eller urologisk undersökning.
I preventionsfrågor kan du kontakta den centraliserade telefontjänsten (06) 826 4477.
Läs mer:
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Preventivrådgivningfinska _ svenska
När du väntar barn
Ta kontakt med rådgivningen då du märker att du är gravid.
På rådgivningen följer man med moderns, barnets och hela familjens välmående under graviditeten.
Läs mer:
När du väntar barn.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Mödrarådgivningfinska _ svenska
Förlossning
Förlossningsavdelningen är öppen dygnet runt.
Om du önskar kan du ringa förlossningsavdelning då din förlossning satt igång eller om du vill fråga om råd.
Då du kommer till sjukhuset ska du använda centralsjukhusets huvudingång kl. 7–20 och övriga tider bör du använda den gemensamma jourens/poliklinikens dörr.
Kontaktuppgifter för förlossningsavdelningen:
Mariegatan 16–20,
67200 Karleby
Telefon: (06) 8264355.
Läs mer: Förlossning.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Förlossningarfinska _ svenska
Läkemedel
Du kan köpa läkemedel på apoteket.
Du kan besöka vilket apotek som helst.
Du kan även besöka apotek som inte finns i din egen kommun.
Läs mer: Läkemedel.
Handikappade personer
En handikappad person bosatt i Karleby har rätt att erhålla de tjänster han eller hon behöver på samma grunder som de övriga invånarna i kommunen.
Personen kan dock på grund av sitt handikapp eller sin sjukdom även behöva särskilda tjänster för handikappade för att klara vardagen.
För tjänsterna för handikappade i Karleby svarar Mellersta Österbottens social- och hälsovårdssamkommun Soite, där man kan ansöka om tjänster och stödfunktioner.
Tjänster av flera olika slag erbjuds även för personer med gravt handikapp.
Dessa tjänster inkluderar bland annat:
transporttjänster
ombyggnad och nödvändig utrustning för hemmet
maskiner och utrustning
personlig hjälp och dagverksamhet
stödboende
stöd för närståendevård av personer under 65 och arbetsverksamhet.
Dessutom är det möjligt att ansöka om specialboende, korttidsvård eller tillfällig vård samt handledning hos den öppna vården.
Mer information om tjänster för handikappade får du från Mellersta Österbottens social- och hälsovårdssamkommun Soites handikapptjänster per telefon: 040 804 2122.
Läs mer: Handikappade personer.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Tjänster för handikappadefinska _ svenska
Specialpedagogik i förskolanfinska _ svenska
Kontaktuppgifter för den grundläggande utbildningenfinska
Ett handikappat barn
Särskilt stöd erbjuds barn med handikapp inom småbarnspedagogiken och skolan.
Kontakta Karleby stads förskoleundervisning för information om specialsmåbarnspedagogiken.
Du kan be undervisningsväsendet om mer information om tjänster som skolan erbjuder.
Bildningscentralen
Strandgatan 16 (våning 5 och 6)
67100 Karleby
Telefon: 040 8065 149
Läs mer: Ett handikappat barn.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Tjänster för handikappadefinska _ svenska
Specialpedagogik i förskolanfinska _ svenska
Kontaktuppgifter för den grundläggande utbildningenfinska
Hälsovårdstjänster i Karleby
Äldre människors hälsa
Tandvård
Mental hälsa
Sexuell hälsa
När du väntar barn
Förlossning
Läkemedel
Handikappade personer
Ett handikappat barn
Hälsovårdstjänster i Karleby
I Karleby finns hälsostationer i olika delar av staden.
Varje hälsostation har ett eget telefonnummer för tidsbokning, som man kan ringa för att boka tid till sjukskötare eller läkare.
Kontaktuppgifter:
Karleby huvudhälsostation
Mariegatan 28
67200 Karleby
Telefon: (06) 8287 580
På Karleby huvudhälsostationen styrs patienterna till mottagningen på basis av hur akuta deras symptom är.
Klienten får en tid till akutvården, mottagningen eller Min Soite-mottagningen.
Samtal till huvudhälsostationen styrs till ett och samma telefonnummer, (06) 8287 310.
67800 Karleby
Telefon: (06) 8287 580
Mottagning /Kelviå
Ellfolkgatan 5
68300 Kelviå
Telefon: (06) 8287 701
Mottagning /Lochteå
Telefon: (06) 8287 750
Mottagning /Ullava
Ullavavägen 701
68370 Ullava
Telefon: (06) 8287 639
Om du kommer som flykting till Finland ska du komma överens om en hälsokontroll med Utlänningsbyrån.
Läs mer: Hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
Under kvällar och helger är hälsostationerna stängda.
Då hanteras plötsliga sjukdomar och olyckor vid jouren.
Jouren är avsedd för patienter vars sjukdom kräver brådskande bedömning och vård.
I livshotande situationer ska du ringa nödnumret 112.
Om du besöker jouren kvällstid eller under helger ska du först ringa jourens telefonrådgivning (06) 826 4500.
Samjourens adress:
Mellersta Österbottens centralsjukhus
Mariegatan 16–20 (l-flygeln, ingång B1)
67200 Karleby
Läs mer: Hälsovårdstjänster i Finland
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barns hälsa
Om ditt barn insjuknar ska du kontakta hälsostationen vid behov.
ådgivningarna erbjuder tjänster för gravida och barn under skolåldern.
Vid rådgivningarna utförs vaccinationer av barn och vuxna.
Du kan kontakta rådgivningen via den centraliserade telefontjänsten (06) 826 4477.
Genom regelbundna besök på barnrådgivningsbyrån följs barnets hälsa, tillväxt och utveckling upp.
På rådgivningen vårdas inte barn som insjuknar plötsligt, men du kan be om råd via den centraliserade telefontjänsten (06) 826 4477.
Skolhälsovårdaren har hand om skolelevers hälsa.
Mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats.
Läs mer: Barns hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barnrådgivningarfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Rådgivningarfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Skolhälsovårdfinska _ svenska
Äldre människors hälsa
Vid hälsopunkten Daalia ges vägledning och rådgivning för personer över 65 år om diet, motion och livsstil.
Vaccinering av personer över 65 år utförs vid seniorrådgivning.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Seniorernas hälsopunkterfinska _ svenska
Tandvård
Om du behöver icke-brådskande tandvård ska du ringa munhälsans centraliserade tidsbokningen.
Centraliserad tidsbokning per telefon: (06) 8287 400
Huvudhälsostationens tandklinik
Mariegatan 28, 67200 Karleby
Björkhagens tandklinik
Storkisbackens tandklinik
Korpvägen 11, 67100 Karleby
Kelviå tandklinik
Ellfolkgatan 5, 68300, Kelviå
Lochteå tandklinik
Ullava tandklinik
Ullavavägen 701, 68370 Ullava
Vardagar kan tider till smärtjouren bokas enligt överenskommelse vid samtliga tandkliniker.
Brådskande tandvård/första hjälpen (kvälls-, vardags-, helg- och nattjour):
Vid smärtjouren får du första hjälpen vid plötslig tandvärk och tandolyckor.
Tandläkarjouren (kvälls-, vardags- och helgjour) ordnas vid polikliniken för tand- och munsjukdomar vid Mellersta Österbottens social- och hälsovårdssamkommun Soite, Mariegatan 16–20, 67200 Karleby (vån 1, del D), vardagkvällar kl. 16.00–21.00 samt veckoslut och helgdagar kl. 8.00–21.00.
Du kan i regel komma till jourmottagningen genom att först kontakta jouren via telefon.
För frågor gällande jouren ring tel. (06) 828 7450.
När du kommer till jourmottagningen ska du ta en kölapp, såvida du inte har en bokad tid.
Brådskande tandvård/första hjälpen (nattjour):
Allvarliga fall i samjour Uleåborgs universitetssjukhus (Oulun yliopistollinen sairaala OYS) kl. 21.00−8.00, tel. (08) 315 2655
Läs mer: Tandvård.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Munhälsovårdenfinska _ svenska
Mental hälsa
Vid problem med din mentala hälsa ska du i första hand kontakta din egen hälsostation eller företagshälsovårdens mottagning.
Vid brådskande problem, kontakta hälsovårdcentralens jour.
Läs mer: Mental hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
Sexuell hälsa
Om du känner att du behöver information om familjeplanering och prevention kan du kontakta din egen hälsostation.
Boka tid till hälsostationen om du behöver preventivmedel, överväger att göra en abort eller misstänker att du lider av en könssjukdom.
Du kan även boka en tid hos en allmänläkare för en gynekologisk eller urologisk undersökning.
I preventionsfrågor kan du kontakta den centraliserade telefontjänsten (06) 826 4477.
Läs mer:
Sexuell hälsa och prevention.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Preventivrådgivningfinska _ svenska
När du väntar barn
Ta kontakt med rådgivningen då du märker att du är gravid.
På rådgivningen följer man med moderns, barnets och hela familjens välmående under graviditeten.
Läs mer: Graviditet och förlossning.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Mödrarådgivningfinska _ svenska
Förlossning
Förlossningsavdelningen är öppen dygnet runt.
Om du önskar kan du ringa förlossningsavdelning då din förlossning satt igång eller om du vill fråga om råd.
Då du kommer till sjukhuset ska du använda centralsjukhusets huvudingång kl. 7–20 och övriga tider bör du använda den gemensamma jourens/poliklinikens dörr.
Kontaktuppgifter för förlossningsavdelningen:
Mariegatan 16–20,
67200 Karleby
Telefon: (06) 8264355.
Läs mer: Graviditet och förlossning.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Förlossningarfinska _ svenska
Läkemedel
Du kan köpa läkemedel på apoteket.
Du kan besöka vilket apotek som helst.
Du kan även besöka apotek som inte finns i din egen kommun.
Läs mer: Läkemedel.
Handikappade personer
En handikappad person bosatt i Karleby har rätt att erhålla de tjänster han eller hon behöver på samma grunder som de övriga invånarna i kommunen.
Personen kan dock på grund av sitt handikapp eller sin sjukdom även behöva särskilda tjänster för handikappade för att klara vardagen.
För tjänsterna för handikappade i Karleby svarar Mellersta Österbottens social- och hälsovårdssamkommun Soite, där man kan ansöka om tjänster och stödfunktioner.
Tjänster av flera olika slag erbjuds även för personer med gravt handikapp.
Dessa tjänster inkluderar bland annat:
transporttjänster
ombyggnad och nödvändig utrustning för hemmet
maskiner och utrustning
personlig hjälp och dagverksamhet
stödboende
stöd för närståendevård av personer under 65 och arbetsverksamhet.
Dessutom är det möjligt att ansöka om specialboende, korttidsvård eller tillfällig vård samt handledning hos den öppna vården.
Mer information om tjänster för handikappade får du från Mellersta Österbottens social- och hälsovårdssamkommun Soites handikapptjänster per telefon: 040 804 2122.
Läs mer: Handikappade personer.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Tjänster för handikappadefinska _ svenska
Specialpedagogik i förskolanfinska _ svenska
Kontaktuppgifter för den grundläggande utbildningenfinska
Ett handikappat barn
Särskilt stöd erbjuds barn med handikapp inom småbarnspedagogiken och skolan.
Kontakta Karleby stads förskoleundervisning för information om specialsmåbarnspedagogiken.
Du kan be undervisningsväsendet om mer information om tjänster som skolan erbjuder.
Bildningscentralen
Strandgatan 16 (våning 5 och 6)
67100 Karleby
Telefon: 040 8065 149
Läs mer: Ett handikappat barn.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Tjänster för handikappadefinska _ svenska
Specialpedagogik i förskolanfinska _ svenska
Kontaktuppgifter för den grundläggande utbildningenfinska
Småbarnspedagogik
Förskoleundervisning
Grundläggande utbildning
Undervisning i det egna modersmålet för invandrare
Yrkesutbildning
Gymnasium
Unga utan studieplats
Högskoleutbildning
Andra studiemöjligheter
Småbarnspedagogik
I Karleby finns stadens egna daghem, gruppfamiljedaghem, familjedagvårdare samt barnklubbar.
Dessutom finns det daghem som köptjänst (svenskspråkiga), ett privat daghem och privata familjedagvårdare i Karleby.
Du kan ansöka om plats inom småbarnspedagogiken för ditt barn elektroniskt via tjänsten Suomi.fi eller med en blankett på stadens webbplats (ansökan till småbarnspedagogiken).
Ansökan ska lämnas in fyra månader innan du behöver plats inom småbarnspedagogiken.
Det är möjligt att få en plats snabbare om den behövs för att du exempelvis erhållit arbete eller studieplats.
Ansökan kan returneras till platsen för småbarnspedagogik, kontorstjänster för småbarnspedagogik eller lämnas i brevlådan i den nedre aulan i Bildningscentralen.
Du kan ansöka om en plats i stadens barnklubbar med blanketten som finns på stadens webbplats.
Ansökan kan även skickas per post till följande adress:
Bildningscentralen
Tjänster för småbarnspedagogik
Strandgatan16
67100 Karleby
Läs mer:
Daghem och andra dagvårdsplatserfinska _ svenska
Gruppfamiljedaghemfinska _ svenska
Dagvårdsblanketterfinska _ svenska
Att ansöka om kommunal dagvårdfinska _ svenska
Förskoleundervisning
Karleby stad erbjuder gratis förskoleundervisning för alla 6 år fyllda barn.
Förskoleundervisningen ges av lärare med utbildning i pedagogik i minst 700 timmar om året, dvs. cirka fyra timmar om dagen, enligt skolans arbetstider.
Förskoleundervisningen är gratis.
Om barnet dessutom behöver avgiftsbelagd småbarnspedagogisk verksamhet arrangeras denna på samma ställe som förskoleundervisningen, dock med undantag för skiftesvård.
Anmälningar till förskoleundervisningen sker i januari–februari.
Detta meddelas i lokaltidningarna och på stadens webbplats.
Om du inte fått ett brev om förskoleplats eller ansöker om förskoleplats under annan tid på året, ta kontakt med kontorstjänster för småbarnspedagogik per telefon på numret 040 806 5089.
Läs mer: Förskoleundervisning.
Förskoleundervisningfinska _ svenska
Grundläggande utbildning
I Finland har alla barn som fyllt 7 år läroplikt, vilket innebär att de måste delta i den grundläggande utbildningen.
Läroplikten upphör i slutet av det läsår då barnet fyller 17.
Det är föräldrarna som har ansvaret för att barnet går i skolan.
Anmälan till grundskolan sker i början av året.
På stadens webbplats finns skolornas kontaktuppgifter och mer information om anmälan.
Om du har frågor om den grundläggande utbildningen kan du även kontakta stadens undervisningstjänster.
Varje barn och ung person har rätt att gå i skola.
Om barnet flyttar till Karleby under läsåret kan han eller hon genast börja i skolan.
Om barnet saknar tillräckliga färdigheter i finska eller svenska för att delta i undervisningen i klassen inleder han eller hon studierna i förberedande undervisning i en egen grupp eller i klassen enligt det egna studieprogrammet.
I Karleby finns grupper för den förberedande utbildningen i lågstadiet i Hollihaan koulu och Koivuhaan koulu och i högstadiet i Stenängens skola.
Övergången till den vanliga undervisningen sker steg för steg enligt elevens förutsättningar.
Undervisning i enlighet med lärokursen finska som andra språk och litteratur stödjer en helhetsmässig utveckling av språket.
Stöd för lärande arrangeras i mån av möjlighet på elevens eget modersmål i skolan.
Mer information om den förberedande undervisningen för invandrare får du av stadens undervisningstjänster.
Läs mer: Grundläggande utbildning.
Kontaktuppgifter för den grundläggande utbildningenfinska
Undervisning i det egna modersmålet för invandrare
Undervisning i elevens eget modersmål arrangeras i Karleby på flera olika språk, till exempel under läsåret 2017–2018 arrangerades undervisning på nio olika språk.
Undervisningsgruppen ska ha minst fyra elever.
Undervisningen sker vanligtvis i de skolor där det finns flest elever som talar språket i fråga.
Som elevens egen religion undervisas bland annat islam, buddhism och ortodox religion, beroende på antalet elever.
Information om undervisning i elevens eget modersmål och religion får du av koordinatoren för undervisningen för olika språk- och kulturgrupper:
Tfn 040 489 2129
Utbildning för invandrarefinska
Yrkesutbildning
Mellersta Österbottens yrkesinstitut erbjuder yrkesutbildning i Karleby, Kelviå, Kannus, Kaustby, Perho och Jakobstad.
Yrkesinstitutet anordnar även handledande utbildning för grundläggande yrkesutbildning, dvs. VALMA-utbildning samt förberedande utbildningar för vuxna invandrare vid Mellersta Österbottens folkhögskola i Kelviå.
Läs mer: Yrkesutbildning.
linkkiMellersta Österbottens utbildningskoncern:
Mellersta Österbottens utbildningskoncernfinska _ engelska
linkkiMellersta Österbottens utbildningskoncern:
Utbildning för invandrarefinska _ engelska
linkkiMellersta Österbottens folkhögskola:
Folkhögskolans invandrarlinjefinska
Gymnasium
I Karleby ges gymnasieutbildning för ungdomar vid Karleby finska gymnasium och Karleby svenska gymnasium, samt för vuxna vid Karleby vuxengymnasium.
Till gymnasieutbildning för ungdomar ansöker man under våren via gemensam ansökning för gymnasierna och man kan bli antagen om man i slutbetyget från grundskolan har tillräckligt högt snittbetyg i läsämnena.
Du kan ansöka till vuxenutbildningen direkt hos vuxengymnasiet året runt.
Karleby finska gymnasium erbjuder förberedande undervisning för gymnasiet även för invandrare.
Den förberedande undervisningen för gymnasiet är ett läsår och målet med den är att förbättra möjligheterna för elever med ett annat modersmål att klara av gymnasiestudierna.
Varje år fattas ett skilt beslut om undervisningens start.
För varje studerande utarbetas ett eget studieprogram.
Man ansöker till förberedande undervisning för gymnasiet under sommaren på webbsidan Opintopolku.fi.
Undervisningsspråket i vid Karleby finska gymnasium och Karleby vuxengymnasium är finska och svenska vid Karleby svenska gymnasium.
Vid Karleby finska gymnasium anordnas undervisning i finska som andraspråk för invandrare invandrare.
Målet är att invandrarna ska klara av gymnasiestudierna och efter gymnasiet kunna söka sig till fortsatta studier.
Mer information om gymnasieskolorna och den förberedande undervisningen för gymnasiet fås av stadens undervisningstjänster.
Kontaktuppgifterna för gymnasierna finns på stadens undervisningstjänsters webbplats.
Bildningscentralen
Strandgatan 16 (våning 5 och 6)
67100 Karleby
Telefon: 044 756 7673
Läs mer:
Gymnasium.
Gymnasie- och yrkesutbildningfinska _ svenska
Unga utan studieplats
Unga som saknar studieplats eller arbete kan få hjälp av det uppsökande ungdomsarbetet.
Det uppsökande ungdomsarbetet hjälper unga i åldern 15–28 år hitta rätt tjänster till stöd för utbildning, arbete och utkomst.
De anställda inom uppsökande ungdomsarbete hjälper med att klara upp den ungas livssituation, hantera praktiska ärenden, såsom besök hos olika myndigheter, och ger personlig handledning enligt den ungas önskemål.
Uppsökande ungdomsarbetefinska _ svenska
Högskoleutbildning
Vid Centria yrkeshögskola kan man avlägga högskoleexamen i teknik, företagsekonomi, social- och hälsovård.
Man kan även avlägga en examen inom musikpedagogik och samhällspedagogik.
Det är dessutom möjligt att studera vid den öppna yrkeshögskolan.
Vid Karleby universitetscenter Chydenius kan man avlägga såväl högre högskoleexamen som doktorsexamen.
Vid Chydenius anordnas även vuxenutbildning och vetenskaplig forskning bedrivs.
Läs mer: Högskoleutbildning.
Högskole- och universitetsutbildningfinska
linkkiCentria yrkeshögskola:
Centria yrkeshögskolafinska _ svenska _ engelska
Universitetscentret Chydeniusfinska _ svenska _ engelska
Andra studiemöjligheter
Karlebynejdens institut, som ägs och drivs av Karleby stad, är ett tvåspråkigt (finska och svenska) medborgarinstitut.
Institutet erbjuder undervisning i datateknik, musik, idrott och dans, konstämnen, hantverk, matlagning och första hjälpen.
Institutet erbjuder även undervisning i flera olika språk, bland annat finska, svenska, engelska, tyska, franska, ryska, spanska och italienska.
Undervisningsutbudet varierar från år till år, så det lönar sig att kontrollera aktuella kurser på institutets webbplats.
Invandrare ges rabatt på vissa kurser.
I kursuppgifterna anges om det är möjligt att få rabatt på kursen.
Kontrollera på institutets webbplats vilka kurser som är aktuella.
Vasavägen 7
67100 Karleby
Telefon: 040 8065 169, 040 8065 168
Vid Mellersta Österbottens sommaruniversitet kan du läsa kurser på universitetsnivå vid det öppna universitetet, delta i kompletterande yrkesutbildning samt läsa språk- och kulturkurser.
Under sommaren är det möjligt att repetera gymnasiestudier vid sommaruniversitetet.
Dessutom är det även möjligt att läsa normala gymnasiekurser vid sommaruniversitetets sommargymnasium.
Sommaruniversitets kurser är avgiftsbelagda för deltagarna.
Läs mer:
Studier som hobby, Arbetskraftsutbildning
Karlebynejdens institutfinska _ svenska
linkkiArbets- och näringsbyråns tjänster:
Offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiMellersta Österbottens sommaruniversitet:
Mellersta Österbottens sommaruniversitetfinska
Övrig undervisning i Karlebyfinska _ svenska
Småbarnspedagogik
Förskoleundervisning
Grundläggande utbildning
Undervisning i det egna modersmålet för invandrare
Yrkesutbildning
Gymnasium
Unga utan studieplats
Högskoleutbildning
Andra studiemöjligheter
Småbarnspedagogik
I Karleby finns stadens egna daghem, gruppfamiljedaghem, familjedagvårdare samt barnklubbar.
Dessutom finns det daghem som köptjänst (svenskspråkiga), ett privat daghem och privata familjedagvårdare i Karleby.
Du kan ansöka om plats inom småbarnspedagogiken för ditt barn elektroniskt via tjänsten Suomi.fi eller med en blankett på stadens webbplats (ansökan till småbarnspedagogiken).
Ansökan ska lämnas in fyra månader innan du behöver plats inom småbarnspedagogiken.
Det är möjligt att få en plats snabbare om den behövs för att du exempelvis erhållit arbete eller studieplats.
Ansökan kan returneras till platsen för småbarnspedagogik, kontorstjänster för småbarnspedagogik eller lämnas i brevlådan i den nedre aulan i Bildningscentralen.
Du kan ansöka om en plats i stadens barnklubbar med blanketten som finns på stadens webbplats.
Ansökan kan även skickas per post till följande adress:
Bildningscentralen
Tjänster för småbarnspedagogik
Strandgatan16
67100 Karleby
Läs mer:
Daghem och andra dagvårdsplatserfinska _ svenska
Gruppfamiljedaghemfinska _ svenska
Dagvårdsblanketterfinska _ svenska
Att ansöka om kommunal dagvårdfinska _ svenska
Förskoleundervisning
Karleby stad erbjuder gratis förskoleundervisning för alla 6 år fyllda barn.
Förskoleundervisningen ges av lärare med utbildning i pedagogik i minst 700 timmar om året, dvs. cirka fyra timmar om dagen, enligt skolans arbetstider.
Förskoleundervisningen är gratis.
Om barnet dessutom behöver avgiftsbelagd småbarnspedagogisk verksamhet arrangeras denna på samma ställe som förskoleundervisningen, dock med undantag för skiftesvård.
Anmälningar till förskoleundervisningen sker i januari–februari.
Detta meddelas i lokaltidningarna och på stadens webbplats.
Om du inte fått ett brev om förskoleplats eller ansöker om förskoleplats under annan tid på året, ta kontakt med kontorstjänster för småbarnspedagogik per telefon på numret 040 806 5089.
Läs mer: Förskoleundervisning.
Förskoleundervisningfinska _ svenska
Grundläggande utbildning
I Finland har alla barn som fyllt 7 år läroplikt, vilket innebär att de måste delta i den grundläggande utbildningen.
Läroplikten upphör i slutet av det läsår då barnet fyller 17.
Det är föräldrarna som har ansvaret för att barnet går i skolan.
Anmälan till grundskolan sker i början av året.
På stadens webbplats finns skolornas kontaktuppgifter och mer information om anmälan.
Om du har frågor om den grundläggande utbildningen kan du även kontakta stadens undervisningstjänster.
Varje barn och ung person har rätt att gå i skola.
Om barnet flyttar till Karleby under läsåret kan han eller hon genast börja i skolan.
Om barnet saknar tillräckliga färdigheter i finska eller svenska för att delta i undervisningen i klassen inleder han eller hon studierna i förberedande undervisning i en egen grupp eller i klassen enligt det egna studieprogrammet.
I Karleby finns grupper för den förberedande utbildningen i lågstadiet i Hollihaan koulu och Koivuhaan koulu och i högstadiet i Stenängens skola.
Övergången till den vanliga undervisningen sker steg för steg enligt elevens förutsättningar.
Undervisning i enlighet med lärokursen finska som andra språk och litteratur stödjer en helhetsmässig utveckling av språket.
Stöd för lärande arrangeras i mån av möjlighet på elevens eget modersmål i skolan.
Mer information om den förberedande undervisningen för invandrare får du av stadens undervisningstjänster.
Läs mer: Grundläggande utbildning.
Kontaktuppgifter för den grundläggande utbildningenfinska
Undervisning i det egna modersmålet för invandrare
Undervisning i elevens eget modersmål arrangeras i Karleby på flera olika språk, till exempel under läsåret 2017–2018 arrangerades undervisning på nio olika språk.
Undervisningsgruppen ska ha minst fyra elever.
Undervisningen sker vanligtvis i de skolor där det finns flest elever som talar språket i fråga.
Som elevens egen religion undervisas bland annat islam, buddhism och ortodox religion, beroende på antalet elever.
Information om undervisning i elevens eget modersmål och religion får du av koordinatoren för undervisningen för olika språk- och kulturgrupper:
Tfn 040 489 2129
Utbildning för invandrarefinska
Yrkesutbildning
Mellersta Österbottens yrkesinstitut erbjuder yrkesutbildning i Karleby, Kelviå, Kannus, Kaustby, Perho och Jakobstad.
Yrkesinstitutet anordnar även handledande utbildning för grundläggande yrkesutbildning, dvs. VALMA-utbildning samt förberedande utbildningar för vuxna invandrare vid Mellersta Österbottens folkhögskola i Kelviå.
Läs mer: Yrkesutbildning.
linkkiMellersta Österbottens utbildningskoncern:
Mellersta Österbottens utbildningskoncernfinska _ engelska
linkkiMellersta Österbottens utbildningskoncern:
Utbildning för invandrarefinska _ engelska
linkkiMellersta Österbottens folkhögskola:
Folkhögskolans invandrarlinjefinska
Gymnasium
I Karleby ges gymnasieutbildning för ungdomar vid Karleby finska gymnasium och Karleby svenska gymnasium, samt för vuxna vid Karleby vuxengymnasium.
Till gymnasieutbildning för ungdomar ansöker man under våren via gemensam ansökning för gymnasierna och man kan bli antagen om man i slutbetyget från grundskolan har tillräckligt högt snittbetyg i läsämnena.
Du kan ansöka till vuxenutbildningen direkt hos vuxengymnasiet året runt.
Karleby finska gymnasium erbjuder förberedande undervisning för gymnasiet även för invandrare.
Den förberedande undervisningen för gymnasiet är ett läsår och målet med den är att förbättra möjligheterna för elever med ett annat modersmål att klara av gymnasiestudierna.
Varje år fattas ett skilt beslut om undervisningens start.
För varje studerande utarbetas ett eget studieprogram.
Man ansöker till förberedande undervisning för gymnasiet under sommaren på webbsidan Opintopolku.fi.
Undervisningsspråket i vid Karleby finska gymnasium och Karleby vuxengymnasium är finska och svenska vid Karleby svenska gymnasium.
Vid Karleby finska gymnasium anordnas undervisning i finska som andraspråk för invandrare invandrare.
Målet är att invandrarna ska klara av gymnasiestudierna och efter gymnasiet kunna söka sig till fortsatta studier.
Mer information om gymnasieskolorna och den förberedande undervisningen för gymnasiet fås av stadens undervisningstjänster.
Kontaktuppgifterna för gymnasierna finns på stadens undervisningstjänsters webbplats.
Bildningscentralen
Strandgatan 16 (våning 5 och 6)
67100 Karleby
Telefon: 044 756 7673
Läs mer:
Gymnasium.
Gymnasie- och yrkesutbildningfinska _ svenska
Unga utan studieplats
Unga som saknar studieplats eller arbete kan få hjälp av det uppsökande ungdomsarbetet.
Det uppsökande ungdomsarbetet hjälper unga i åldern 15–28 år hitta rätt tjänster till stöd för utbildning, arbete och utkomst.
De anställda inom uppsökande ungdomsarbete hjälper med att klara upp den ungas livssituation, hantera praktiska ärenden, såsom besök hos olika myndigheter, och ger personlig handledning enligt den ungas önskemål.
Uppsökande ungdomsarbetefinska _ svenska
Högskoleutbildning
Vid Centria yrkeshögskola kan man avlägga högskoleexamen i teknik, företagsekonomi, social- och hälsovård.
Man kan även avlägga en examen inom musikpedagogik och samhällspedagogik.
Det är dessutom möjligt att studera vid den öppna yrkeshögskolan.
Vid Karleby universitetscenter Chydenius kan man avlägga såväl högre högskoleexamen som doktorsexamen.
Vid Chydenius anordnas även vuxenutbildning och vetenskaplig forskning bedrivs.
Läs mer: Högskoleutbildning.
Högskole- och universitetsutbildningfinska
linkkiCentria yrkeshögskola:
Centria yrkeshögskolafinska _ svenska _ engelska
Universitetscentret Chydeniusfinska _ svenska _ engelska
Andra studiemöjligheter
Karlebynejdens institut, som ägs och drivs av Karleby stad, är ett tvåspråkigt (finska och svenska) medborgarinstitut.
Institutet erbjuder undervisning i datateknik, musik, idrott och dans, konstämnen, hantverk, matlagning och första hjälpen.
Institutet erbjuder även undervisning i flera olika språk, bland annat finska, svenska, engelska, tyska, franska, ryska, spanska och italienska.
Undervisningsutbudet varierar från år till år, så det lönar sig att kontrollera aktuella kurser på institutets webbplats.
Invandrare ges rabatt på vissa kurser.
I kursuppgifterna anges om det är möjligt att få rabatt på kursen.
Kontrollera på institutets webbplats vilka kurser som är aktuella.
Vasavägen 7
67100 Karleby
Telefon: 040 8065 169, 040 8065 168
Vid Mellersta Österbottens sommaruniversitet kan du läsa kurser på universitetsnivå vid det öppna universitetet, delta i kompletterande yrkesutbildning samt läsa språk- och kulturkurser.
Under sommaren är det möjligt att repetera gymnasiestudier vid sommaruniversitetet.
Dessutom är det även möjligt att läsa normala gymnasiekurser vid sommaruniversitetets sommargymnasium.
Sommaruniversitets kurser är avgiftsbelagda för deltagarna.
Läs mer:
Studier som hobby, Arbetskraftsutbildning
Karlebynejdens institutfinska _ svenska
linkkiArbets- och näringsbyråns tjänster:
Offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiMellersta Österbottens sommaruniversitet:
Mellersta Österbottens sommaruniversitetfinska
Övrig undervisning i Karlebyfinska _ svenska
Småbarnspedagogik
Förskoleundervisning
Grundläggande utbildning
Undervisning i det egna modersmålet för invandrare
Yrkesutbildning
Gymnasium
Unga utan studieplats
Högskoleutbildning
Andra studiemöjligheter
Småbarnspedagogik
I Karleby finns stadens egna daghem, gruppfamiljedaghem, familjedagvårdare samt barnklubbar.
Dessutom finns det daghem som köptjänst (svenskspråkiga), ett privat daghem och privata familjedagvårdare i Karleby.
Du kan ansöka om plats inom småbarnspedagogiken för ditt barn elektroniskt via tjänsten Suomi.fi eller med en blankett på stadens webbplats (ansökan till småbarnspedagogiken).
Ansökan ska lämnas in fyra månader innan du behöver plats inom småbarnspedagogiken.
Det är möjligt att få en plats snabbare om den behövs för att du exempelvis erhållit arbete eller studieplats.
Ansökan kan returneras till platsen för småbarnspedagogik, kontorstjänster för småbarnspedagogik eller lämnas i brevlådan i den nedre aulan i Bildningscentralen.
Du kan ansöka om en plats i stadens barnklubbar med blanketten som finns på stadens webbplats.
Ansökan kan även skickas per post till följande adress:
Bildningscentralen
Tjänster för småbarnspedagogik
Strandgatan16
67100 Karleby
Läs mer:
Småbarnspedagogik.
Daghem och andra dagvårdsplatserfinska _ svenska
Gruppfamiljedaghemfinska _ svenska
Dagvårdsblanketterfinska _ svenska
Att ansöka om kommunal dagvårdfinska _ svenska
Förskoleundervisning
Karleby stad erbjuder gratis förskoleundervisning för alla 6 år fyllda barn.
Förskoleundervisningen ges av lärare med utbildning i pedagogik i minst 700 timmar om året, dvs. cirka fyra timmar om dagen, enligt skolans arbetstider.
Förskoleundervisningen är gratis.
Om barnet dessutom behöver avgiftsbelagd småbarnspedagogisk verksamhet arrangeras denna på samma ställe som förskoleundervisningen, dock med undantag för skiftesvård.
Anmälningar till förskoleundervisningen sker i januari–februari.
Detta meddelas i lokaltidningarna och på stadens webbplats.
Om du inte fått ett brev om förskoleplats eller ansöker om förskoleplats under annan tid på året, ta kontakt med kontorstjänster för småbarnspedagogik per telefon på numret 040 806 5089.
Läs mer: Förskoleundervisning.
Förskoleundervisningfinska _ svenska
Grundläggande utbildning
I Finland har alla barn som fyllt 7 år läroplikt, vilket innebär att de måste delta i den grundläggande utbildningen.
Läroplikten upphör i slutet av det läsår då barnet fyller 17.
Det är föräldrarna som har ansvaret för att barnet går i skolan.
Anmälan till grundskolan sker i början av året.
På stadens webbplats finns skolornas kontaktuppgifter och mer information om anmälan.
Om du har frågor om den grundläggande utbildningen kan du även kontakta stadens undervisningstjänster.
Varje barn och ung person har rätt att gå i skola.
Om barnet flyttar till Karleby under läsåret kan han eller hon genast börja i skolan.
Om barnet saknar tillräckliga färdigheter i finska eller svenska för att delta i undervisningen i klassen inleder han eller hon studierna i förberedande undervisning i en egen grupp eller i klassen enligt det egna studieprogrammet.
I Karleby finns grupper för den förberedande utbildningen i lågstadiet i Hollihaan koulu och Koivuhaan koulu och i högstadiet i Stenängens skola.
Övergången till den vanliga undervisningen sker steg för steg enligt elevens förutsättningar.
Undervisning i enlighet med lärokursen finska som andra språk och litteratur stödjer en helhetsmässig utveckling av språket.
Stöd för lärande arrangeras i mån av möjlighet på elevens eget modersmål i skolan.
Mer information om den förberedande undervisningen för invandrare får du av stadens undervisningstjänster.
Läs mer: Grundläggande utbildning.
Kontaktuppgifter för den grundläggande utbildningenfinska
Undervisning i det egna modersmålet för invandrare
Undervisning i elevens eget modersmål arrangeras i Karleby på flera olika språk, till exempel under läsåret 2017–2018 arrangerades undervisning på nio olika språk.
Undervisningsgruppen ska ha minst fyra elever.
Undervisningen sker vanligtvis i de skolor där det finns flest elever som talar språket i fråga.
Som elevens egen religion undervisas bland annat islam, buddhism och ortodox religion, beroende på antalet elever.
Information om undervisning i elevens eget modersmål och religion får du av koordinatoren för undervisningen för olika språk- och kulturgrupper:
Tfn 040 489 2129
Utbildning för invandrarefinska
Yrkesutbildning
Mellersta Österbottens yrkesinstitut erbjuder yrkesutbildning i Karleby, Kelviå, Kannus, Kaustby, Perho och Jakobstad.
Yrkesinstitutet anordnar även handledande utbildning för grundläggande yrkesutbildning, dvs. VALMA-utbildning samt förberedande utbildningar för vuxna invandrare vid Mellersta Österbottens folkhögskola i Kelviå.
Läs mer: Yrkesutbildning.
linkkiMellersta Österbottens utbildningskoncern:
Mellersta Österbottens utbildningskoncernfinska _ engelska
linkkiMellersta Österbottens utbildningskoncern:
Utbildning för invandrarefinska _ engelska
linkkiMellersta Österbottens folkhögskola:
Folkhögskolans invandrarlinjefinska
Gymnasium
I Karleby ges gymnasieutbildning för ungdomar vid Karleby finska gymnasium och Karleby svenska gymnasium, samt för vuxna vid Karleby vuxengymnasium.
Till gymnasieutbildning för ungdomar ansöker man under våren via gemensam ansökning för gymnasierna och man kan bli antagen om man i slutbetyget från grundskolan har tillräckligt högt snittbetyg i läsämnena.
Du kan ansöka till vuxenutbildningen direkt hos vuxengymnasiet året runt.
Karleby finska gymnasium erbjuder förberedande undervisning för gymnasiet även för invandrare.
Den förberedande undervisningen för gymnasiet är ett läsår och målet med den är att förbättra möjligheterna för elever med ett annat modersmål att klara av gymnasiestudierna.
Varje år fattas ett skilt beslut om undervisningens start.
För varje studerande utarbetas ett eget studieprogram.
Man ansöker till förberedande undervisning för gymnasiet under sommaren på webbsidan Opintopolku.fi.
Undervisningsspråket i vid Karleby finska gymnasium och Karleby vuxengymnasium är finska och svenska vid Karleby svenska gymnasium.
Vid Karleby finska gymnasium anordnas undervisning i finska som andraspråk för invandrare invandrare.
Målet är att invandrarna ska klara av gymnasiestudierna och efter gymnasiet kunna söka sig till fortsatta studier.
Mer information om gymnasieskolorna och den förberedande undervisningen för gymnasiet fås av stadens undervisningstjänster.
Kontaktuppgifterna för gymnasierna finns på stadens undervisningstjänsters webbplats.
Bildningscentralen
Strandgatan 16 (våning 5 och 6)
67100 Karleby
Telefon: 044 756 7673
Läs mer:
Gymnasium.
Gymnasie- och yrkesutbildningfinska _ svenska
Unga utan studieplats
Unga som saknar studieplats eller arbete kan få hjälp av det uppsökande ungdomsarbetet.
Det uppsökande ungdomsarbetet hjälper unga i åldern 15–28 år hitta rätt tjänster till stöd för utbildning, arbete och utkomst.
De anställda inom uppsökande ungdomsarbete hjälper med att klara upp den ungas livssituation, hantera praktiska ärenden, såsom besök hos olika myndigheter, och ger personlig handledning enligt den ungas önskemål.
Uppsökande ungdomsarbetefinska _ svenska
Högskoleutbildning
Vid Centria yrkeshögskola kan man avlägga högskoleexamen i teknik, företagsekonomi, social- och hälsovård.
Man kan även avlägga en examen inom musikpedagogik och samhällspedagogik.
Det är dessutom möjligt att studera vid den öppna yrkeshögskolan.
Vid Karleby universitetscenter Chydenius kan man avlägga såväl högre högskoleexamen som doktorsexamen.
Vid Chydenius anordnas även vuxenutbildning och vetenskaplig forskning bedrivs.
Läs mer:
Yrkeshögskolor, Universitet.
Högskole- och universitetsutbildningfinska
linkkiCentria yrkeshögskola:
Centria yrkeshögskolafinska _ svenska _ engelska
Universitetscentret Chydeniusfinska _ svenska _ engelska
Andra studiemöjligheter
Karlebynejdens institut, som ägs och drivs av Karleby stad, är ett tvåspråkigt (finska och svenska) medborgarinstitut.
Institutet erbjuder undervisning i datateknik, musik, idrott och dans, konstämnen, hantverk, matlagning och första hjälpen.
Institutet erbjuder även undervisning i flera olika språk, bland annat finska, svenska, engelska, tyska, franska, ryska, spanska och italienska.
Undervisningsutbudet varierar från år till år, så det lönar sig att kontrollera aktuella kurser på institutets webbplats.
Invandrare ges rabatt på vissa kurser.
I kursuppgifterna anges om det är möjligt att få rabatt på kursen.
Kontrollera på institutets webbplats vilka kurser som är aktuella.
Vasavägen 7
67100 Karleby
Telefon: 040 8065 169, 040 8065 168
Vid Mellersta Österbottens sommaruniversitet kan du läsa kurser på universitetsnivå vid det öppna universitetet, delta i kompletterande yrkesutbildning samt läsa språk- och kulturkurser.
Under sommaren är det möjligt att repetera gymnasiestudier vid sommaruniversitetet.
Dessutom är det även möjligt att läsa normala gymnasiekurser vid sommaruniversitetets sommargymnasium.
Sommaruniversitets kurser är avgiftsbelagda för deltagarna.
Läs mer:
Studier som hobby, Arbetskraftsutbildning
Karlebynejdens institutfinska _ svenska
linkkiArbets- och näringsbyråns tjänster:
Offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiMellersta Österbottens sommaruniversitet:
Mellersta Österbottens sommaruniversitetfinska
Övrig undervisning i Karlebyfinska _ svenska
Hyresbostad
Ägarbostad
Tillfälligt boende
Stöd- och serviceboende
Bostadslöshet
Avfallshantering för bostaden
Hyresbostad
Karleby stads blankett för ansökan om hyresbostad kan fyllas i och skickas in på nätet.
Bilagor till ansökningen ska tillhandahållas då bostad erbjuds, men kan även lämnas in tidigare.
Man kan även lämna in bostadsansökan på papper.
Ansökningsblanketterna kan hämtas från och lämnas in till Kokkolan Vuokra Asunnot Oy:s verksamhetsställen.
67800 Karleby
Telefon: 040 1817 400
Studiebostäder hyrs ut av Kiinteistöyhtiö Tankkari, som erbjuder möblerade kollektivbostäder samt familjebostäder i olika storlek.
En familjebostad är en omöblerad lägenhet som endast hyrs ut till personer i samma hushåll.
Såväl individer som sambor/gifta par kan ansöka om en hyresetta.
Bondegatan 2
67100 Karleby
Telefon: 040 193 6468
Läs mer:
Hyresbostad.
Hyresbostäderfinska _ svenska
Ansökan om Karleby stads hyresbostadfinska _ svenska _ engelska
Hyresbostäder enligt stadsdelfinska _ svenska
Studiebostäderfinska _ engelska
Privata hyresbostäderfinska _ svenska
Ägarbostad
De flesta finländarna bor i en ägarbostad, alltså i en bostad som de själva äger.
På lång sikt är det ofta förmånligare att köpa sin egen bostad än att hyra.
Bland annat hos bostadsförmedlingen, på internet och i lokala tidningar finns annonser om bostäder som är till salu.
Läs mer:
Ägarbostad.
Tillfälligt boende
I Karlebynejden erbjuds olika inkvarteringsalternativ.
Kontaktuppgifterna finns under länkarna nedan.
Läs mer:
Tillfälligt boende.
Övernattningsalternativ i Karlebyfinska _ svenska _ engelska
Om du saknar boende på grund av kris eller olycka ska du kontakta Kokkolan Vuokra Asunnot Oy eller bostadsbyrån.
Om din bostad har skadats, till exempel till följd av brand eller vattenskada, kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
Kontakta ditt försäkringsbolag direkt när skadan har inträffat.
Om en familjemedlem är våldsam eller hotar med våld, ta kontakt med Karleby mödra- och skyddshem.
Du kan ringa skyddshemmet under alla tider på dygnet.
Du behöver inte uppge ditt namn då du ringer.
Karleby mödra- och skyddshem
Telefon: 044 336 0056
Hyresbostäderfinska _ svenska
Karleby mödra- och skyddshemfinska
Stöd- och serviceboende
Äldre människor erbjuds boendeservice anordnad av Mellersta Österbottens social- och hälsovårdssamkommun Soite samt privata servicebostäder.
Serviceboende för äldre är avsett för personer över 65 år som behöver vård och omsorg dygnet runt.
Serviceboende är lämpat för personer som inte längre klarar sig på egen hand med tjänster som tillhandahålls i hemmet.
Mer information om boendeservice anordnad av Mellersta Österbottens social- och hälsovårdssamkommun Soite får du av bland annat samkommunens servicestyrcentral, tfn 040 806 5093.
För handikappade och personer som återhämtar sig från mentala problem erbjuds bostäder som beaktar invånarnas särskilda behov.
Hemvårdens stödtjänster erbjuds personer som har svårigheter med att klara vardagen utan hjälp, såsom äldre och handikappade personer.
Tjänster av detta slag är bland annat måltidstjänst och transporttjänst.
Målet med hemvården är att erbjuda trygg vård och omsorg samt främja invånarnas ork, handlingskraft och företagsamhet.
Läs mer:
Stöd- och serviceboende.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Servicehandledningscentretfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Seniorernas tjänster, hemvårdfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Seniorernas tjänster, serviceboendet och anstaltsvårdenfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Boendetjänster för utvecklingsstörda och handikappadefinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Socialrådgivningfinska _ svenska
Bostadslöshet
Om du blir bostadslös bör du kontakta Kokkolan Vuokra Asunnot Oy eller bostadsbyrån.
Hyresbostäderfinska _ svenska
Avfallshantering för bostaden
Med bioavfall avses bl.a.:
matrester
skämda och torra livsmedel
skal från frukt och grönsaker
Separat insamlat bioavfall packas i en papperspåse, en påse vikt av en dagstidning eller en plastkasse. Kassen eller påsen får vara högst 30l stor.
En full sopsäck ska tillslutas noggrant.
Med energiavfall avses bl.a.:
bakplåtspapper, hushållspapper och våtservetter
kläder (inte skor, regnställ eller läderplagg)
små plastleksaker och bruksföremål i plast såsom disk- och tandborstar.
Separat insamlat energiavfall ska packas i plastkasse eller papperspåsar.
Kassen eller påsen får vara högst 30 l stor.
Påsen tillsluts noga.
Avfall som inte får läggas i det egna husets sopbehållare kan föras till återvinningsstationer.
Kontrollera på förhand vilken typ av avfall stationen tar emot.
Mer information om avfallshanteringen i Karlebynejden finns på Karleby stads och på Ab Ekorosk Oy:s (kommunalt avfallshanteringsbolag) webbplats.
Läs mer: Avfallshantering och återvinning.
Avfallshantering för bostaden finska _ svenska
Ett kommunalt avfallshanteringsbolagfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ vietnamesiska _ polska _ kroatiska
Hyresbostad
Köpa bostad
Tillfälligt boende
Stöd- och serviceboende
Bostadslöshet
Avfallshantering för bostaden
Hyresbostad
Karleby stads blankett för ansökan om hyresbostad kan fyllas i och skickas in på nätet.
Bilagor till ansökningen ska tillhandahållas då bostad erbjuds, men kan även lämnas in tidigare.
Man kan även lämna in bostadsansökan på papper.
Ansökningsblanketterna kan hämtas från och lämnas in till Kokkolan Vuokra Asunnot Oy:s verksamhetsställen.
67800 Karleby
Telefon: 040 1817 400
Studiebostäder hyrs ut av Kiinteistöyhtiö Tankkari, som erbjuder möblerade kollektivbostäder samt familjebostäder i olika storlek.
En familjebostad är en omöblerad lägenhet som endast hyrs ut till personer i samma hushåll.
Såväl individer som sambor/gifta par kan ansöka om en hyresetta.
Bondegatan 2
67100 Karleby
Telefon: 040 193 6468
Läs mer: Hyresbostad.
Hyresbostäderfinska _ svenska
Ansökan om Karleby stads hyresbostadfinska _ svenska _ engelska
Hyresbostäder enligt stadsdelfinska _ svenska
Studiebostäderfinska _ engelska
Privata hyresbostäderfinska _ svenska
Köpa bostad
De flesta finländarna bor i en ägarbostad, alltså i en bostad som de själva äger.
På lång sikt är det ofta förmånligare att köpa sin egen bostad än att hyra.
Bland annat hos bostadsförmedlingen, på internet och i lokala tidningar finns annonser om bostäder som är till salu.
Läs mer: Köpa bostad.
Tillfälligt boende
I Karlebynejden erbjuds olika inkvarteringsalternativ.
Kontaktuppgifterna finns under länkarna nedan.
Läs mer:
Tillfälligt boende.
Övernattningsalternativ i Karlebyfinska _ svenska _ engelska
Om du saknar boende på grund av kris eller olycka ska du kontakta Kokkolan Vuokra Asunnot Oy eller bostadsbyrån.
Om din bostad har skadats, till exempel till följd av brand eller vattenskada, kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
Kontakta ditt försäkringsbolag direkt när skadan har inträffat.
Om en familjemedlem är våldsam eller hotar med våld, ta kontakt med Karleby mödra- och skyddshem.
Du kan ringa skyddshemmet under alla tider på dygnet.
Du behöver inte uppge ditt namn då du ringer.
Karleby mödra- och skyddshem
Telefon: 044 336 0056
Läs mer: Boende.
Hyresbostäderfinska _ svenska
Karleby mödra- och skyddshemfinska
Stöd- och serviceboende
Äldre människor erbjuds boendeservice anordnad av Mellersta Österbottens social- och hälsovårdssamkommun Soite samt privata servicebostäder.
Serviceboende för äldre är avsett för personer över 65 år som behöver vård och omsorg dygnet runt.
Serviceboende är lämpat för personer som inte längre klarar sig på egen hand med tjänster som tillhandahålls i hemmet.
Mer information om boendeservice anordnad av Mellersta Österbottens social- och hälsovårdssamkommun Soite får du av bland annat samkommunens servicestyrcentral, tfn 040 806 5093.
För handikappade och personer som återhämtar sig från mentala problem erbjuds bostäder som beaktar invånarnas särskilda behov.
Hemvårdens stödtjänster erbjuds personer som har svårigheter med att klara vardagen utan hjälp, såsom äldre och handikappade personer.
Tjänster av detta slag är bland annat måltidstjänst och transporttjänst.
Målet med hemvården är att erbjuda trygg vård och omsorg samt främja invånarnas ork, handlingskraft och företagsamhet.
Läs mer:
Stöd- och serviceboende.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Servicehandledningscentretfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Seniorernas tjänster, hemvårdfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Seniorernas tjänster, serviceboendet och anstaltsvårdenfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Boendetjänster för utvecklingsstörda och handikappadefinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Socialrådgivningfinska _ svenska
Bostadslöshet
Om du blir bostadslös bör du kontakta Kokkolan Vuokra Asunnot Oy eller bostadsbyrån.
Läs mer: Bostadslöshet.
Hyresbostäderfinska _ svenska
Avfallshantering för bostaden
Med bioavfall avses bl.a.:
matrester
skämda och torra livsmedel
skal från frukt och grönsaker
Separat insamlat bioavfall packas i en papperspåse, en påse vikt av en dagstidning eller en plastkasse. Kassen eller påsen får vara högst 30l stor.
En full sopsäck ska tillslutas noggrant.
Med energiavfall avses bl.a.:
bakplåtspapper, hushållspapper och våtservetter
kläder (inte skor, regnställ eller läderplagg)
små plastleksaker och bruksföremål i plast såsom disk- och tandborstar.
Separat insamlat energiavfall ska packas i plastkasse eller papperspåsar.
Kassen eller påsen får vara högst 30 l stor.
Påsen tillsluts noga.
Avfall som inte får läggas i det egna husets sopbehållare kan föras till återvinningsstationer.
Kontrollera på förhand vilken typ av avfall stationen tar emot.
Mer information om avfallshanteringen i Karlebynejden finns på Karleby stads och på Ab Ekorosk Oy:s (kommunalt avfallshanteringsbolag) webbplats.
Läs mer: Avfallshantering och återvinning.
Avfallshantering för bostaden finska _ svenska
Ett kommunalt avfallshanteringsbolagfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ vietnamesiska _ polska _ kroatiska
Hyresbostad
Köpa bostad
Tillfälligt boende
Stöd- och serviceboende
Bostadslöshet
Avfallshantering för bostaden
Hyresbostad
Karleby stads blankett för ansökan om hyresbostad kan fyllas i och skickas in på nätet.
Bilagor till ansökningen ska tillhandahållas då bostad erbjuds, men kan även lämnas in tidigare.
Man kan även lämna in bostadsansökan på papper.
Ansökningsblanketterna kan hämtas från och lämnas in till Kokkolan Vuokra Asunnot Oy:s verksamhetsställen.
67800 Karleby
Telefon: 040 1817 400
Studiebostäder hyrs ut av Kiinteistöyhtiö Tankkari, som erbjuder möblerade kollektivbostäder samt familjebostäder i olika storlek.
En familjebostad är en omöblerad lägenhet som endast hyrs ut till personer i samma hushåll.
Såväl individer som sambor/gifta par kan ansöka om en hyresetta.
Bondegatan 2
67100 Karleby
Telefon: 040 193 6468
Läs mer: Hyresbostad.
Hyresbostäderfinska _ svenska
Ansökan om Karleby stads hyresbostadfinska _ svenska _ engelska
Hyresbostäder enligt stadsdelfinska _ svenska
Studiebostäderfinska _ engelska
Privata hyresbostäderfinska _ svenska
Köpa bostad
De flesta finländarna bor i en ägarbostad, alltså i en bostad som de själva äger.
På lång sikt är det ofta förmånligare att köpa sin egen bostad än att hyra.
Bland annat hos bostadsförmedlingen, på internet och i lokala tidningar finns annonser om bostäder som är till salu.
Läs mer: Köpa bostad.
Tillfälligt boende
I Karlebynejden erbjuds olika inkvarteringsalternativ.
Kontaktuppgifterna finns under länkarna nedan.
Läs mer:
Tillfälligt boende.
Övernattningsalternativ i Karlebyfinska _ svenska _ engelska
Om du saknar boende på grund av kris eller olycka ska du kontakta Kokkolan Vuokra Asunnot Oy eller bostadsbyrån.
Om din bostad har skadats, till exempel till följd av brand eller vattenskada, kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
Kontakta ditt försäkringsbolag direkt när skadan har inträffat.
Om en familjemedlem är våldsam eller hotar med våld, ta kontakt med Karleby mödra- och skyddshem.
Du kan ringa skyddshemmet under alla tider på dygnet.
Du behöver inte uppge ditt namn då du ringer.
Karleby mödra- och skyddshem
Telefon: 044 336 0056
Läs mer: Boende.
Hyresbostäderfinska _ svenska
Karleby mödra- och skyddshemfinska
Stöd- och serviceboende
Äldre människor erbjuds boendeservice anordnad av Mellersta Österbottens social- och hälsovårdssamkommun Soite samt privata servicebostäder.
Serviceboende för äldre är avsett för personer över 65 år som behöver vård och omsorg dygnet runt.
Serviceboende är lämpat för personer som inte längre klarar sig på egen hand med tjänster som tillhandahålls i hemmet.
Mer information om boendeservice anordnad av Mellersta Österbottens social- och hälsovårdssamkommun Soite får du av bland annat samkommunens servicestyrcentral, tfn 040 806 5093.
För handikappade och personer som återhämtar sig från mentala problem erbjuds bostäder som beaktar invånarnas särskilda behov.
Hemvårdens stödtjänster erbjuds personer som har svårigheter med att klara vardagen utan hjälp, såsom äldre och handikappade personer.
Tjänster av detta slag är bland annat måltidstjänst och transporttjänst.
Målet med hemvården är att erbjuda trygg vård och omsorg samt främja invånarnas ork, handlingskraft och företagsamhet.
Läs mer:
Stöd- och serviceboende.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Servicehandledningscentretfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Seniorernas tjänster, hemvårdfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Seniorernas tjänster, serviceboendet och anstaltsvårdenfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Boendetjänster för utvecklingsstörda och handikappadefinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Socialrådgivningfinska _ svenska
Bostadslöshet
Om du blir bostadslös bör du kontakta Kokkolan Vuokra Asunnot Oy eller bostadsbyrån.
Läs mer: Bostadslöshet.
Hyresbostäderfinska _ svenska
Avfallshantering för bostaden
Med bioavfall avses bl.a.:
matrester
skämda och torra livsmedel
skal från frukt och grönsaker
Separat insamlat bioavfall packas i en papperspåse, en påse vikt av en dagstidning eller en plastkasse. Kassen eller påsen får vara högst 30l stor.
En full sopsäck ska tillslutas noggrant.
Med energiavfall avses bl.a.:
bakplåtspapper, hushållspapper och våtservetter
kläder (inte skor, regnställ eller läderplagg)
små plastleksaker och bruksföremål i plast såsom disk- och tandborstar.
Separat insamlat energiavfall ska packas i plastkasse eller papperspåsar.
Kassen eller påsen får vara högst 30 l stor.
Påsen tillsluts noga.
Avfall som inte får läggas i det egna husets sopbehållare kan föras till återvinningsstationer.
Kontrollera på förhand vilken typ av avfall stationen tar emot.
Mer information om avfallshanteringen i Karlebynejden finns på Karleby stads och på Ab Ekorosk Oy:s (kommunalt avfallshanteringsbolag) webbplats.
Läs mer: Avfallshantering och återvinning.
Avfallshantering för bostaden finska _ svenska
Ett kommunalt avfallshanteringsbolagfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ vietnamesiska _ polska _ kroatiska
Möjligheter att studera finska eller svenska
Karlebynejdens institut erbjuder undervisning i finska och svenska från grundnivå.
Mellersta Österbottens utbildningskoncern erbjuder kurser i finska vid Mellersta Österbottens folkhögskola i Kelviå inom utbildningen i läs- och skrivfärdigheter och den förberedande utbildningen för vuxna invandrare. Det går också att studera finska inom utbildningen som handleder för yrkesutbildning (VALMA) vid Mellersta Österbottens Vuxeninstitut.
Vuxenutbildningen anordnar även förberedande utbildning för vuxna invandrare vid Mellersta Österbottens folkhögskola i Kelviå.
Vid Kronoby folkhögskola kan du studera finska och svenska på grund- och påbyggnadsnivå.
Om du är berättigad till integrationsstöd ska du kontakta TE-byrån innan du ansöker.
Du kan be om information om undervisning i finska och svenska för invandrare hos utlänningsbyrån.
Läs mer: Finska och svenska språket
Karlebynejdens institutfinska _ svenska
linkkiMellersta Österbottens utbildningskoncern:
Utbildning för invandrarefinska _ engelska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Utlänningsbyrånfinska _ svenska
linkkiKronoby folkhögskola:
Kronoby folkhögskolafinska _ svenska _ engelska
Möjligheter att studera finska eller svenska
Karlebynejdens institut erbjuder undervisning i finska och svenska från grundnivå.
Mellersta Österbottens utbildningskoncern erbjuder kurser i finska vid Mellersta Österbottens folkhögskola i Kelviå inom utbildningen i läs- och skrivfärdigheter och den förberedande utbildningen för vuxna invandrare. Det går också att studera finska inom utbildningen som handleder för yrkesutbildning (VALMA) vid Mellersta Österbottens Vuxeninstitut.
Vuxenutbildningen anordnar även förberedande utbildning för vuxna invandrare vid Mellersta Österbottens folkhögskola i Kelviå.
Vid Kronoby folkhögskola kan du studera finska och svenska på grund- och påbyggnadsnivå.
Om du är berättigad till integrationsstöd ska du kontakta TE-byrån innan du ansöker.
Du kan be om information om undervisning i finska och svenska för invandrare hos utlänningsbyrån.
Läs mer: Finska och svenska språket
Karlebynejdens institutfinska _ svenska
linkkiMellersta Österbottens utbildningskoncern:
Utbildning för invandrarefinska _ engelska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Utlänningsbyrånfinska _ svenska
linkkiKronoby folkhögskola:
Kronoby folkhögskolafinska _ svenska _ engelska
Möjligheter att studera finska eller svenska
Karlebynejdens institut erbjuder undervisning i finska och svenska från grundnivå.
Mellersta Österbottens utbildningskoncern erbjuder kurser i finska vid Mellersta Österbottens folkhögskola i Kelviå inom utbildningen i läs- och skrivfärdigheter och den förberedande utbildningen för vuxna invandrare. Det går också att studera finska inom utbildningen som handleder för yrkesutbildning (VALMA) vid Mellersta Österbottens Vuxeninstitut.
Vuxenutbildningen anordnar även förberedande utbildning för vuxna invandrare vid Mellersta Österbottens folkhögskola i Kelviå.
Vid Kronoby folkhögskola kan du studera finska och svenska på grund- och påbyggnadsnivå.
Om du är berättigad till integrationsstöd ska du kontakta TE-byrån innan du ansöker.
Du kan be om information om undervisning i finska och svenska för invandrare hos utlänningsbyrån.
Läs mer: Finska och svenska språket
Karlebynejdens institutfinska _ svenska
linkkiMellersta Österbottens utbildningskoncern:
Utbildning för invandrarefinska _ engelska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Utlänningsbyrånfinska _ svenska
linkkiKronoby folkhögskola:
Kronoby folkhögskolafinska _ svenska _ engelska
Var hittar jag jobb?
Att grunda ett företag
Beskattning
Om du blir arbetslös
Var hittar jag jobb?
Du kan söka arbetsplatser på internet och i tidningar.
På internet hittar du jobbsajter när du skriver ”avoimet työpaikat” (lediga jobb) i sökmotorns textfält.
På många jobbsajter kan du spara din jobbansökan och meritförteckning (CV) så att arbetsgivaren kan läsa dem.
Vid Österbottens TE-byrå (arbets- och näringsbyrå) får du hjälp med att hitta en arbetsplats.
Du behöver inte alltid boka tid för att besöka TE-byrån.
I Mina e-tjänster på nätet kan du bl.a. ändra dina uppgifter som arbetssökande och kontrollera giltighetstiden för jobbsökningen och utlåtandet om arbetslöshetsförsäkring.
Om du behöver boka en tid till TE-byrån ska du kontakta TE-byrån direkt per telefon eller boka en tid på plats.
Var även direkt i kontakt med TE-byrån om du önskar ändra en tidsbokning.
Du kan ringa TE-telefonservice då du behöver information om TE-byråns tjänster eller vägledning i tjänsterna på nätet.
Telefonnumret till TE-telefonservice är 0295 025 500 på finska, 0295 025 510 på svenska, 0295 020 713 på engelska och 0295 020 715 på ryska.
TE-byrån i Österbotten betjänar i Karleby, Kaustby, Jakobstad, Närpes, Kristinestad och Vasa.
Du kan fritt välja vilken TE-byrå du besöker.
Adressen för TE-byrån i Karleby är
67100 Karleby.
På TE-byråns jobbsajt finns tusentals arbetsplatser runt om i Finland.
Du hittar lediga arbetsplatser i din kommun genom att skriva kommunens namn i sökfältet ”Region”.
Läs mer:
Var hittar jag jobb?
linkkiArbets- och näringsbyråns tjänster:
Offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiArbets- och näringsbyråns tjänster:
Österbottens TE-byråfinska _ svenska
linkkiArbets- och näringsbyråns tjänster:
TE-telefonservicefinska _ svenska _ engelska _ ryska
linkkiArbets- och näringsbyråns tjänster:
Arbets- och näringsbyråns arbetsplatssajtfinska _ svenska
Att grunda ett företag
KOSEK (Karlebynejdens Utveckling Ab) erbjuder tjänster som nyttar företaget under hela dess livscykel, från och med att starta företagsverksamhet.
KOSEKs experter hjälper bland annat med att utarbeta en affärsverksamhetsplan och att ansöka startpeng.
Tjänsterna är avgiftsfria.
Verksamheten av Mellersta Österbottens Nyföretagarcentral FIRMAXI fortsätter som en del av KOSEKs tjänster.
Du kan besöka Karlebynejdens Utveckling Ab om du behöver information om att grunda ett företag.
Detta kan exempelvis inkludera
företagsfinansiering
rekrytering av anställda
samarbetsnätverk
verksamhetslokaler
Läs mer:
Att grunda ett företag.
linkkiNyföretagarcentralen Firmaxi:
Nyföretagarcentralen Firmaxifinska
Karlebynejdens Utveckling Abfinska _ svenska _ engelska
Beskattning
Om du behöver ett skattekort eller skattenummer kan du besöka Västra Finlands skattebyrå.
Skattebyråns kontaktuppgifter:
PB 1002, 67101 Karleby
Besöksadress: Karlebygatan 27, Karleby
Skatteförvaltningens riksomfattande telefontjänst: 029 497 050
Läs mer: Beskattning.
Om du blir arbetslös
Medborgare i EU- och EES-länderna kan anmäla sig som arbetslösa på nätet i TE-byråns ”Mina e-tjänster”.
Du kan besöka TE-byrån om du inte kan anmäla dig som arbetssökande på nätet eller om du är medborgare i något annat land.
Du kan ringa till riksomfattande servicenummer om du behöver hjälp med att använda e-tjänsterna eller mer information om TE-byråns tjänster.
Det riksomfattande servicenumret är 0295 025 500 på finska, 0295 025 510 på svenska, 0295 020 713 på engelska och 0295 020 715 på ryska.
TE-byrån i Österbotten betjänar i Karleby, Kaustby, Jakobstad, Närpes, Kristinestad och Vasa.
Du kan fritt välja vilken TE-byrå du besöker.
TE-byråns adress i Karleby
Läs mer: Arbetslöshetsförsäkring.
linkkiArbets- och näringsbyråns tjänster:
Offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiArbets- och näringsbyråns tjänster:
Österbottens TE-byråfinska _ svenska
linkkiArbets- och näringsbyråns tjänster:
TE-telefonservicefinska _ svenska _ engelska _ ryska
Fennovoima bygger kärnkraftverksenheten Hanhikivi 1 i Pyhäjoki.
Kärnkraftverket levereras av RAOS Project Oy, ett bolag som ingår i den ryska Rosatom-koncernen.
Enligt den överenskomna tidtabellen kommer kärnkraftverket att producera el år 2024.
Planeringen och konstruktionen av kärnkraftverket är ett omfattande projekt som tar cirka 10 år att slutföra.
Under tiden kärnkraftverket uppförs kommer som mest upp till 3 000–4 000 personer att arbeta på området.
Arbetsgivaren arrangerar logi för merparten av arbetstagarna, och man strävar efter att ordna inkvartering så nära bygget som möjligt.
I kärnkraftverkets omedelbara närhet byggs ett inkvarteringsområde för 1 000 personer.
I Pyhäjoki och det omgivande området har man förberett sig på kärnkraftverksprojektet redan i flera års tid.
Information om området har sammanställts bl.a. i Hanhikivi-guiden som publicerats på finska, engelska, svenska och ryska.
Elektroniska versioner av guiden finns på storprojektets webbplats.
Den tryckta guiden finns i företagsservicecentralerna i kommunerna på området.
Som en del av förberedelserna för kärnkraftverksprojektet finns information samlad om tjänsterna på området på dessa lokala InfoFinland-sidor.
Mer information om Fennovoimas kärnkraftverksprojekt i Pyhäjoki:
Fennovoima Oyfinska _ engelska
linkkiBrahestadsregionens företagstjänster:
Information om storprojekt som förverkligas i regionen och förberedelserna för dessafinska _ engelska _ ryska
Karlebynejdens Utveckling Abfinska _ svenska _ engelska
linkkiPyhäjoki kommun:
Pyhäjoki kommunfinska _ svenska _ engelska
Information om verksamhetsmiljön för kärnkraftverksprojektetfinska _ svenska _ engelska _ ryska
Var hittar jag jobb?
Att grunda ett företag
Beskattning
Om du blir arbetslös
Var hittar jag jobb?
Du kan söka arbetsplatser på internet och i tidningar.
På internet hittar du jobbsajter när du skriver ”avoimet työpaikat” (lediga jobb) i sökmotorns textfält.
På många jobbsajter kan du spara din jobbansökan och meritförteckning (CV) så att arbetsgivaren kan läsa dem.
Vid Österbottens TE-byrå (arbets- och näringsbyrå) får du hjälp med att hitta en arbetsplats.
Du behöver inte alltid boka tid för att besöka TE-byrån.
I Mina e-tjänster på nätet kan du bl.a. ändra dina uppgifter som arbetssökande och kontrollera giltighetstiden för jobbsökningen och utlåtandet om arbetslöshetsförsäkring.
Om du behöver boka en tid till TE-byrån ska du kontakta TE-byrån direkt per telefon eller boka en tid på plats.
Var även direkt i kontakt med TE-byrån om du önskar ändra en tidsbokning.
Du kan ringa TE-telefonservice då du behöver information om TE-byråns tjänster eller vägledning i tjänsterna på nätet.
Telefonnumret till TE-telefonservice är 0295 025 500 på finska, 0295 025 510 på svenska, 0295 020 713 på engelska och 0295 020 715 på ryska.
TE-byrån i Österbotten betjänar i Karleby, Kaustby, Jakobstad, Närpes, Kristinestad och Vasa.
Du kan fritt välja vilken TE-byrå du besöker.
Adressen för TE-byrån i Karleby är
67100 Karleby.
På TE-byråns jobbsajt finns tusentals arbetsplatser runt om i Finland.
Du hittar lediga arbetsplatser i din kommun genom att skriva kommunens namn i sökfältet ”Region”.
Läs mer:
Var hittar jag jobb?
linkkiArbets- och näringsbyråns tjänster:
Offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiArbets- och näringsbyråns tjänster:
Österbottens TE-byråfinska _ svenska
linkkiArbets- och näringsbyråns tjänster:
TE-telefonservicefinska _ svenska _ engelska _ ryska
linkkiArbets- och näringsbyråns tjänster:
Arbets- och näringsbyråns arbetsplatssajtfinska _ svenska
Att grunda ett företag
KOSEK (Karlebynejdens Utveckling Ab) erbjuder tjänster som nyttar företaget under hela dess livscykel, från och med att starta företagsverksamhet.
KOSEKs experter hjälper bland annat med att utarbeta en affärsverksamhetsplan och att ansöka startpeng.
Tjänsterna är avgiftsfria.
Verksamheten av Mellersta Österbottens Nyföretagarcentral FIRMAXI fortsätter som en del av KOSEKs tjänster.
Du kan besöka Karlebynejdens Utveckling Ab om du behöver information om att grunda ett företag.
Detta kan exempelvis inkludera
företagsfinansiering
rekrytering av anställda
samarbetsnätverk
verksamhetslokaler
Läs mer:
Att grunda ett företag.
linkkiNyföretagarcentralen Firmaxi:
Nyföretagarcentralen Firmaxifinska
Karlebynejdens Utveckling Abfinska _ svenska _ engelska
Beskattning
Om du behöver ett skattekort eller skattenummer kan du besöka Västra Finlands skattebyrå.
Skattebyråns kontaktuppgifter:
PB 1002, 67101 Karleby
Besöksadress: Karlebygatan 27, Karleby
Skatteförvaltningens riksomfattande telefontjänst: 029 497 050
Läs mer: Beskattning.
Om du blir arbetslös
Medborgare i EU- och EES-länderna kan anmäla sig som arbetslösa på nätet i TE-byråns ”Mina e-tjänster”.
Du kan besöka TE-byrån om du inte kan anmäla dig som arbetssökande på nätet eller om du är medborgare i något annat land.
Du kan ringa till riksomfattande servicenummer om du behöver hjälp med att använda e-tjänsterna eller mer information om TE-byråns tjänster.
Det riksomfattande servicenumret är 0295 025 500 på finska, 0295 025 510 på svenska, 0295 020 713 på engelska och 0295 020 715 på ryska.
TE-byrån i Österbotten betjänar i Karleby, Kaustby, Jakobstad, Närpes, Kristinestad och Vasa.
Du kan fritt välja vilken TE-byrå du besöker.
TE-byråns adress i Karleby
Läs mer: Arbetslöshetsförsäkring.
linkkiArbets- och näringsbyråns tjänster:
Offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiArbets- och näringsbyråns tjänster:
Österbottens TE-byråfinska _ svenska
linkkiArbets- och näringsbyråns tjänster:
TE-telefonservicefinska _ svenska _ engelska _ ryska
Fennovoima bygger kärnkraftverksenheten Hanhikivi 1 i Pyhäjoki.
Kärnkraftverket levereras av RAOS Project Oy, ett bolag som ingår i den ryska Rosatom-koncernen.
Enligt den överenskomna tidtabellen kommer kärnkraftverket att producera el år 2024.
Planeringen och konstruktionen av kärnkraftverket är ett omfattande projekt som tar cirka 10 år att slutföra.
Under tiden kärnkraftverket uppförs kommer som mest upp till 3 000–4 000 personer att arbeta på området.
Arbetsgivaren arrangerar logi för merparten av arbetstagarna, och man strävar efter att ordna inkvartering så nära bygget som möjligt.
I kärnkraftverkets omedelbara närhet byggs ett inkvarteringsområde för 1 000 personer.
I Pyhäjoki och det omgivande området har man förberett sig på kärnkraftverksprojektet redan i flera års tid.
Information om området har sammanställts bl.a. i Hanhikivi-guiden som publicerats på finska, engelska, svenska och ryska.
Elektroniska versioner av guiden finns på storprojektets webbplats.
Den tryckta guiden finns i företagsservicecentralerna i kommunerna på området.
Som en del av förberedelserna för kärnkraftverksprojektet finns information samlad om tjänsterna på området på dessa lokala InfoFinland-sidor.
Mer information om Fennovoimas kärnkraftverksprojekt i Pyhäjoki:
Fennovoima Oyfinska _ engelska
linkkiBrahestadsregionens företagstjänster:
Information om storprojekt som förverkligas i regionen och förberedelserna för dessafinska _ engelska _ ryska
Karlebynejdens Utveckling Abfinska _ svenska _ engelska
linkkiPyhäjoki kommun:
Pyhäjoki kommunfinska _ svenska _ engelska
Information om verksamhetsmiljön för kärnkraftverksprojektetfinska _ svenska _ engelska _ ryska
Var hittar jag jobb?
Att grunda ett företag
Beskattning
Om du blir arbetslös
Var hittar jag jobb?
Du kan söka arbetsplatser på internet och i tidningar.
På internet hittar du jobbsajter när du skriver ”avoimet työpaikat” (lediga jobb) i sökmotorns textfält.
På många jobbsajter kan du spara din jobbansökan och meritförteckning (CV) så att arbetsgivaren kan läsa dem.
Vid Österbottens TE-byrå (arbets- och näringsbyrå) får du hjälp med att hitta en arbetsplats.
Du behöver inte alltid boka tid för att besöka TE-byrån.
I Mina e-tjänster på nätet kan du bl.a. ändra dina uppgifter som arbetssökande och kontrollera giltighetstiden för jobbsökningen och utlåtandet om arbetslöshetsförsäkring.
Om du behöver boka en tid till TE-byrån ska du kontakta TE-byrån direkt per telefon eller boka en tid på plats.
Var även direkt i kontakt med TE-byrån om du önskar ändra en tidsbokning.
Du kan ringa TE-telefonservice då du behöver information om TE-byråns tjänster eller vägledning i tjänsterna på nätet.
Telefonnumret till TE-telefonservice är 0295 025 500 på finska, 0295 025 510 på svenska, 0295 020 713 på engelska och 0295 020 715 på ryska.
TE-byrån i Österbotten betjänar i Karleby, Kaustby, Jakobstad, Närpes, Kristinestad och Vasa.
Du kan fritt välja vilken TE-byrå du besöker.
Adressen för TE-byrån i Karleby är
67100 Karleby.
På TE-byråns jobbsajt finns tusentals arbetsplatser runt om i Finland.
Du hittar lediga arbetsplatser i din kommun genom att skriva kommunens namn i sökfältet ”Region”.
Läs mer:
Var hittar jag jobb?
linkkiArbets- och näringsbyråns tjänster:
Offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiArbets- och näringsbyråns tjänster:
Österbottens TE-byråfinska _ svenska
linkkiArbets- och näringsbyråns tjänster:
TE-telefonservicefinska _ svenska _ engelska _ ryska
linkkiArbets- och näringsbyråns tjänster:
Arbets- och näringsbyråns arbetsplatssajtfinska _ svenska
Att grunda ett företag
KOSEK (Karlebynejdens Utveckling Ab) erbjuder tjänster som nyttar företaget under hela dess livscykel, från och med att starta företagsverksamhet.
KOSEKs experter hjälper bland annat med att utarbeta en affärsverksamhetsplan och att ansöka startpeng.
Tjänsterna är avgiftsfria.
Verksamheten av Mellersta Österbottens Nyföretagarcentral FIRMAXI fortsätter som en del av KOSEKs tjänster.
Du kan besöka Karlebynejdens Utveckling Ab om du behöver information om att grunda ett företag.
Detta kan exempelvis inkludera
företagsfinansiering
rekrytering av anställda
samarbetsnätverk
verksamhetslokaler
Läs mer:
Att grunda ett företag.
linkkiNyföretagarcentralen Firmaxi:
Nyföretagarcentralen Firmaxifinska
Karlebynejdens Utveckling Abfinska _ svenska _ engelska
Beskattning
Om du behöver ett skattekort eller skattenummer kan du besöka Västra Finlands skattebyrå.
Skattebyråns kontaktuppgifter:
PB 1002, 67101 Karleby
Besöksadress: Karlebygatan 27, Karleby
Skatteförvaltningens riksomfattande telefontjänst: 029 497 050
Läs mer: Beskattning.
Om du blir arbetslös
Medborgare i EU- och EES-länderna kan anmäla sig som arbetslösa på nätet i TE-byråns ”Mina e-tjänster”.
Du kan besöka TE-byrån om du inte kan anmäla dig som arbetssökande på nätet eller om du är medborgare i något annat land.
Du kan ringa till riksomfattande servicenummer om du behöver hjälp med att använda e-tjänsterna eller mer information om TE-byråns tjänster.
Det riksomfattande servicenumret är 0295 025 500 på finska, 0295 025 510 på svenska, 0295 020 713 på engelska och 0295 020 715 på ryska.
TE-byrån i Österbotten betjänar i Karleby, Kaustby, Jakobstad, Närpes, Kristinestad och Vasa.
Du kan fritt välja vilken TE-byrå du besöker.
TE-byråns adress i Karleby
Läs mer: Arbetslöshetsförsäkring.
linkkiArbets- och näringsbyråns tjänster:
Offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
linkkiArbets- och näringsbyråns tjänster:
Österbottens TE-byråfinska _ svenska
linkkiArbets- och näringsbyråns tjänster:
TE-telefonservicefinska _ svenska _ engelska _ ryska
Fennovoima bygger kärnkraftverksenheten Hanhikivi 1 i Pyhäjoki.
Kärnkraftverket levereras av RAOS Project Oy, ett bolag som ingår i den ryska Rosatom-koncernen.
Enligt den överenskomna tidtabellen kommer kärnkraftverket att producera el år 2024.
Planeringen och konstruktionen av kärnkraftverket är ett omfattande projekt som tar cirka 10 år att slutföra.
Under tiden kärnkraftverket uppförs kommer som mest upp till 3 000–4 000 personer att arbeta på området.
Arbetsgivaren arrangerar logi för merparten av arbetstagarna, och man strävar efter att ordna inkvartering så nära bygget som möjligt.
I kärnkraftverkets omedelbara närhet byggs ett inkvarteringsområde för 1 000 personer.
I Pyhäjoki och det omgivande området har man förberett sig på kärnkraftverksprojektet redan i flera års tid.
Information om området har sammanställts bl.a. i Hanhikivi-guiden som publicerats på finska, engelska, svenska och ryska.
Elektroniska versioner av guiden finns på storprojektets webbplats.
Den tryckta guiden finns i företagsservicecentralerna i kommunerna på området.
Som en del av förberedelserna för kärnkraftverksprojektet finns information samlad om tjänsterna på området på dessa lokala InfoFinland-sidor.
Mer information om Fennovoimas kärnkraftverksprojekt i Pyhäjoki:
Fennovoima Oyfinska _ engelska
linkkiBrahestadsregionens företagstjänster:
Information om storprojekt som förverkligas i regionen och förberedelserna för dessafinska _ engelska _ ryska
Karlebynejdens Utveckling Abfinska _ svenska _ engelska
linkkiPyhäjoki kommun:
Pyhäjoki kommunfinska _ svenska _ engelska
Information om verksamhetsmiljön för kärnkraftverksprojektetfinska _ svenska _ engelska _ ryska
Rådgivning och integration för invandrare
Inledande kartläggning och integrationsplan
Behöver du en tolk?
Rådgivning och integration för invandrare
Då du flyttar till Finland kan du använda dig av TE-byråns (arbets- och näringsbyrån) tjänster som hjälper dig att göra dig hemmastadd i Finland och hitta en arbetsplats.
Tjänster särskilt avsedda för invandrare är:
handledning och rådgivning för invandrare
inledande kartläggning
integrationsutbildning
Österbottens TE-byrå
67100 Karleby
Telefonväxel: 0295 025 500
Karleby evangelisk-lutherska församlingssammanslutnings invandrararbete stöder invandrares integrering i det finländska samhället.
linkkiArbets- och näringsbyråns tjänster:
Offentliga arbets- och näringstjänsterfinska _ svenska
linkkiArbets- och näringsministeriet:
Guiden Välkommen till Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
linkkiKarleby evangelisk-lutherska församlingssammansutning:
Karleby evangelisk-lutherska församlings invandrararbetefinska _ svenska _ engelska _ ryska
Inledande kartläggning och integrationsplan
En inledande kartläggning och integrationsplan utarbetas för dig i arbets- och näringsbyrån. Om du kommit till
Finland som flykting utarbetas en inledande kartläggning och integrationsplan för dig vid utlänningsbyrån.
Du kan fråga mer om kartläggningen och integrationsplanen vid utlänningsbyrån eller TE-byrån.
Utlänningsbyrån
Vasavägen 6 C
67100 Karleby
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Utlänningsbyrånfinska _ svenska
Behöver du en tolk?
Om du måste sköta ärenden med finländska myndigheter, men inte kan finska eller svenska och det inte heller finns något annat språk som både du och myndigheten talar, kan du i vissa fall ha rätt till tolkning.
Myndigheten beställer tolken om du på förhand uppgett att du behöver en tolk.
I detta fall är det gratis för dig att använda dig av tolk.
Du kan använda tolken när du själv önskar om du betalar kostnaderna och beställer tolken själv.
Läs mer:
Behöver du en tolk?
Rådgivning och integration för invandrare
Inledande kartläggning och integrationsplan
Behöver du en tolk?
Rådgivning och integration för invandrare
Då du flyttar till Finland kan du använda dig av TE-byråns (arbets- och näringsbyrån) tjänster som hjälper dig att göra dig hemmastadd i Finland och hitta en arbetsplats.
Tjänster särskilt avsedda för invandrare är:
handledning och rådgivning för invandrare
inledande kartläggning
integrationsutbildning
Österbottens TE-byrå
67100 Karleby
Telefonväxel: 0295 025 500
Karleby evangelisk-lutherska församlingssammanslutnings invandrararbete stöder invandrares integrering i det finländska samhället.
linkkiArbets- och näringsbyråns tjänster:
Offentliga arbets- och näringstjänsterfinska _ svenska
linkkiArbets- och näringsministeriet:
Guiden Välkommen till Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
linkkiKarleby evangelisk-lutherska församlingssammansutning:
Karleby evangelisk-lutherska församlings invandrararbetefinska _ svenska _ engelska _ ryska
Inledande kartläggning och integrationsplan
En inledande kartläggning och integrationsplan utarbetas för dig i arbets- och näringsbyrån. Om du kommit till
Finland som flykting utarbetas en inledande kartläggning och integrationsplan för dig vid utlänningsbyrån.
Du kan fråga mer om kartläggningen och integrationsplanen vid utlänningsbyrån eller TE-byrån.
Utlänningsbyrån
Vasavägen 6 C
67100 Karleby
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Utlänningsbyrånfinska _ svenska
Behöver du en tolk?
Om du måste sköta ärenden med finländska myndigheter, men inte kan finska eller svenska och det inte heller finns något annat språk som både du och myndigheten talar, kan du i vissa fall ha rätt till tolkning.
Myndigheten beställer tolken om du på förhand uppgett att du behöver en tolk.
I detta fall är det gratis för dig att använda dig av tolk.
Du kan använda tolken när du själv önskar om du betalar kostnaderna och beställer tolken själv.
Läs mer:
Behöver du en tolk?
Rådgivning och integration för invandrare
Inledande kartläggning och integrationsplan
Behöver du en tolk?
Rådgivning och integration för invandrare
Då du flyttar till Finland kan du använda dig av TE-byråns (arbets- och näringsbyrån) tjänster som hjälper dig att göra dig hemmastadd i Finland och hitta en arbetsplats.
Tjänster särskilt avsedda för invandrare är:
handledning och rådgivning för invandrare
inledande kartläggning
integrationsutbildning
Österbottens TE-byrå
67100 Karleby
Telefonväxel: 0295 025 500
Karleby evangelisk-lutherska församlingssammanslutnings invandrararbete stöder invandrares integrering i det finländska samhället.
linkkiArbets- och näringsbyråns tjänster:
Offentliga arbets- och näringstjänsterfinska _ svenska
linkkiArbets- och näringsministeriet:
Guiden Välkommen till Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
linkkiKarleby evangelisk-lutherska församlingssammansutning:
Karleby evangelisk-lutherska församlings invandrararbetefinska _ svenska _ engelska _ ryska
Inledande kartläggning och integrationsplan
En inledande kartläggning och integrationsplan utarbetas för dig i arbets- och näringsbyrån. Om du kommit till
Finland som flykting utarbetas en inledande kartläggning och integrationsplan för dig vid utlänningsbyrån.
Du kan fråga mer om kartläggningen och integrationsplanen vid utlänningsbyrån eller TE-byrån.
Utlänningsbyrån
Vasavägen 6 C
67100 Karleby
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Utlänningsbyrånfinska _ svenska
Behöver du en tolk?
Om du måste sköta ärenden med finländska myndigheter, men inte kan finska eller svenska och det inte heller finns något annat språk som både du och myndigheten talar, kan du i vissa fall ha rätt till tolkning.
Myndigheten beställer tolken om du på förhand uppgett att du behöver en tolk.
I detta fall är det gratis för dig att använda dig av tolk.
Du kan använda tolken när du själv önskar om du betalar kostnaderna och beställer tolken själv.
Läs mer:
Behöver du en tolk?
Registrering som invånare
Om du vill flytta till Finland behöver du vanligtvis ett uppehållstillstånd.
Uppehållstillståndsärenden hanteras av Finlands beskickningar i utlandet och Migrationsverket.
Läs mer: Flytta till Finland.
Då du flyttar till Karleby (Kokkola) ska du registrera dig som invånare i kommunen.
Du kan personligen registrera dig på Karleby enheten för Magistraten i Västra Finland:
Magistraten i Västra Finland
Karleby enhet
Karlebygatan 27
67701 Karleby
Telefon: 029 553 9451
När du går till magistraten ska du ta med dig
uppehållstillstånd och uppehållskort (om du behöver ett uppehållstillstånd i Finland)
registreringsintyget över uppehållsrätt för EU-medborgare (om du är EU-medborgare)
äktenskapsbevis
födelseattester för dina barn
Observera att officiella handlingar som tagits med från utlandet ska vara legaliserade och i original samt översatta till finska, svenska eller engelska.
Mer information om legalisering av handlingar får du hos magistraten eller hos ditt lands beskickning i Finland.
Läs mer:
Registrering som invånare.
Magistratens kontaktuppgifterfinska _ svenska _ engelska
Fortsatt uppehållstillstånd
Du ska ansöka om fortsatt uppehållstillstånd innan ditt tidigare uppehållstillstånd går ut.
Du ansöker om tillståndet vid Migrationsverkets servicesställen.
Du kan endast ansöka om fortsatt uppehållstillstånd i Finland.
Migrationsverket
Korsholmsesplanaden 45
Vasa
Läs mer: Fortsatt uppehållstillstånd.
Registrering som invånare
Om du vill flytta till Finland behöver du vanligtvis ett uppehållstillstånd.
Uppehållstillståndsärenden hanteras av Finlands beskickningar i utlandet och Migrationsverket.
Läs mer: Flytta till Finland.
Då du flyttar till Karleby (Kokkola) ska du registrera dig som invånare i kommunen.
Du kan personligen registrera dig på Karleby enheten för Magistraten i Västra Finland:
Magistraten i Västra Finland
Karleby enhet
Karlebygatan 27
67701 Karleby
Telefon: 029 553 9451
När du går till magistraten ska du ta med dig
uppehållstillstånd och uppehållskort (om du behöver ett uppehållstillstånd i Finland)
registreringsintyget över uppehållsrätt för EU-medborgare (om du är EU-medborgare)
äktenskapsbevis
födelseattester för dina barn
Observera att officiella handlingar som tagits med från utlandet ska vara legaliserade och i original samt översatta till finska, svenska eller engelska.
Mer information om legalisering av handlingar får du hos magistraten eller hos ditt lands beskickning i Finland.
Läs mer:
Registrering som invånare.
Magistratens kontaktuppgifterfinska _ svenska _ engelska
Fortsatt uppehållstillstånd
Du ska ansöka om fortsatt uppehållstillstånd innan ditt tidigare uppehållstillstånd går ut.
Du ansöker om tillståndet vid Migrationsverkets servicesställen.
Du kan endast ansöka om fortsatt uppehållstillstånd i Finland.
Migrationsverket
Korsholmsesplanaden 45
Vasa
Läs mer: Fortsatt uppehållstillstånd.
Registrering som invånare
Om du vill flytta till Finland behöver du vanligtvis ett uppehållstillstånd.
Uppehållstillståndsärenden hanteras av Finlands beskickningar i utlandet och Migrationsverket.
Läs mer: Flytta till Finland.
Då du flyttar till Karleby (Kokkola) ska du registrera dig som invånare i kommunen.
Du kan personligen registrera dig på Karleby enheten för Magistraten i Västra Finland:
Magistraten i Västra Finland
Karleby enhet
Karlebygatan 27
67701 Karleby
Telefon: 029 553 9451
När du går till magistraten ska du ta med dig
uppehållstillstånd och uppehållskort (om du behöver ett uppehållstillstånd i Finland)
registreringsintyget över uppehållsrätt för EU-medborgare (om du är EU-medborgare)
äktenskapsbevis
födelseattester för dina barn
Observera att officiella handlingar som tagits med från utlandet ska vara legaliserade och i original samt översatta till finska, svenska eller engelska.
Mer information om legalisering av handlingar får du hos magistraten eller hos ditt lands beskickning i Finland.
Läs mer:
Registrering som invånare.
Magistratens kontaktuppgifterfinska _ svenska _ engelska
Fortsatt uppehållstillstånd
Du ska ansöka om fortsatt uppehållstillstånd innan ditt tidigare uppehållstillstånd går ut.
Du ansöker om tillståndet vid Migrationsverkets servicesställen.
Du kan endast ansöka om fortsatt uppehållstillstånd i Finland.
Migrationsverket
Korsholmsesplanaden 45
Vasa
Läs mer: Fortsatt uppehållstillstånd.
InfoFinland finansieras av Samarbetskommunerna och staten.
Åren 2017–2020 var statens finansiärer arbets- och näringsministeriet, undervisnings- och kulturministeriet, miljöministeriet, FPA och Skatteförvaltningen.
InfoFinland utvecklas i samarbete med finansiärerna.
Den som planerar att flytta till Finland med hjälp av Infobanken hittar lätt information om att leva, bo, arbeta och studera i Finland på många olika språk.
Staten
Arbets- och näringsministeriet
Arbets- och näringsministeriet svarar för beredningen av ärenden i anslutning till integrationen av invandrare i Finland.
Kompetenscentret för integration av invandrare stöder arbete som främjar integrationen av invandrare lokalt, regionalt och riksomfattande.
linkkiArbets- och näringsministeriet :
Integration av invandrarefinska _ svenska _ engelska
Undervisnings- och kulturministeriet
Undervisnings- och kulturministeriet svarar för utvecklingen av och det internationella samarbetet inom utbildnings-, vetenskaps-, kultur-, motions- och ungdomspolitiken.
linkkiUndervisnings- och kulturministeriet:
Webbsidorfinska _ svenska _ engelska
Miljöministeriet
linkkiMiljöministeriet:
Webbsidorfinska _ svenska _ engelska
FPA
FPA sköter grundtryggheten i olika skeden av livet för dem som bor i Finland.
FPA:s kunder är alla personer som bor i Finland och utomlands och som omfattas av socialskyddet i Finland.
FPA och Skatteförvaltningen erbjuder information till utländska anställda på servicestället In To Finland i Helsingfors.
Flyttning till eller från Finlandfinska _ svenska _ engelska
Skatteförvaltningen
linkkiSkatteförvaltningen:
Webbsidorfinska _ svenska _ engelska
Kommunerna
Helsingfors stad
Publicerar och administrerar InfoFinland.
Kommuner som är med i samarbetsavtalet
InfoFinlands samarbetsavtal
InfoFinlands finansiärer har ingått ett samarbetsavtal med vilket man överenskommit om principerna för genomförandet och finansieringen av nättjänsten InfoFinland (tidigare Infobanken) för åren 2017–2020.
Samarbetet möjliggör riksomfattande webbinformation för invandrare och personer som planerar att flytta till Finland och för myndigheter inom invandrarsektorn på ett sätt som också stöder behovet av information i kommunerna.
Det är lätt att på ett pålitligt sätt hitta väsentlig information om integration av invandrare och om att bo i Finland på ett ställe, www.infofinland.fi.
Avtalsparterna driver och utvecklar tjänsten tillsammans.
De vill dessutom stärka InfoFinlands riksomfattande ställning, så att det är möjligt för nya kommuner och andra organisationer att ansluta sig till tjänsten också i fortsättningen.
Kommunernas finansieringsandelar fastställs utgående från antalet invånare.
Genomförandet av avtalet följs upp av en styrgrupp.
Nya aktörer är välkomna att utveckla den flerspråkiga informationen till invandrare och ansluta sig till InfoFinlands samarbetsavtal.
Närmare information om hur man ansluter sig till avtalet ger InfoFinlands chefredaktör Eija Kyllönen-Saarnio, eija.kyllonen-saarnio(snabel-a)hel.fi, tfn 050 363 3285.
InfoFinland finansieras av Samarbetskommunerna och staten.
Åren 2017–2020 var statens finansiärer arbets- och näringsministeriet, undervisnings- och kulturministeriet, miljöministeriet, FPA och Skatteförvaltningen.
InfoFinland utvecklas i samarbete med finansiärerna.
Den som planerar att flytta till Finland med hjälp av Infobanken hittar lätt information om att leva, bo, arbeta och studera i Finland på många olika språk.
Staten
Arbets- och näringsministeriet
Arbets- och näringsministeriet svarar för beredningen av ärenden i anslutning till integrationen av invandrare i Finland.
Kompetenscentret för integration av invandrare stöder arbete som främjar integrationen av invandrare lokalt, regionalt och riksomfattande.
linkkiArbets- och näringsministeriet :
Integration av invandrarefinska _ svenska _ engelska
Undervisnings- och kulturministeriet
Undervisnings- och kulturministeriet svarar för utvecklingen av och det internationella samarbetet inom utbildnings-, vetenskaps-, kultur-, motions- och ungdomspolitiken.
linkkiUndervisnings- och kulturministeriet:
Webbsidorfinska _ svenska _ engelska
Miljöministeriet
linkkiMiljöministeriet:
Webbsidorfinska _ svenska _ engelska
FPA
FPA sköter grundtryggheten i olika skeden av livet för dem som bor i Finland.
FPA:s kunder är alla personer som bor i Finland och utomlands och som omfattas av socialskyddet i Finland.
FPA och Skatteförvaltningen erbjuder information till utländska anställda på servicestället In To Finland i Helsingfors.
Flyttning till eller från Finlandfinska _ svenska _ engelska
Skatteförvaltningen
linkkiSkatteförvaltningen:
Webbsidorfinska _ svenska _ engelska
Kommunerna
Helsingfors stad
Publicerar och administrerar InfoFinland.
Kommuner som är med i samarbetsavtalet
InfoFinlands samarbetsavtal
InfoFinlands finansiärer har ingått ett samarbetsavtal med vilket man överenskommit om principerna för genomförandet och finansieringen av nättjänsten InfoFinland (tidigare Infobanken) för åren 2017–2020.
Samarbetet möjliggör riksomfattande webbinformation för invandrare och personer som planerar att flytta till Finland och för myndigheter inom invandrarsektorn på ett sätt som också stöder behovet av information i kommunerna.
Det är lätt att på ett pålitligt sätt hitta väsentlig information om integration av invandrare och om att bo i Finland på ett ställe, www.infofinland.fi.
Avtalsparterna driver och utvecklar tjänsten tillsammans.
De vill dessutom stärka InfoFinlands riksomfattande ställning, så att det är möjligt för nya kommuner och andra organisationer att ansluta sig till tjänsten också i fortsättningen.
Kommunernas finansieringsandelar fastställs utgående från antalet invånare.
Genomförandet av avtalet följs upp av en styrgrupp.
Nya aktörer är välkomna att utveckla den flerspråkiga informationen till invandrare och ansluta sig till InfoFinlands samarbetsavtal.
Närmare information om hur man ansluter sig till avtalet ger InfoFinlands chefredaktör Eija Kyllönen-Saarnio, eija.kyllonen-saarnio(snabel-a)hel.fi, tfn 050 363 3285.
InfoFinland finansieras av Samarbetskommunerna och staten.
Åren 2017–2020 var statens finansiärer arbets- och näringsministeriet, undervisnings- och kulturministeriet, miljöministeriet, FPA och Skatteförvaltningen.
InfoFinland utvecklas i samarbete med finansiärerna.
Den som planerar att flytta till Finland med hjälp av Infobanken hittar lätt information om att leva, bo, arbeta och studera i Finland på många olika språk.
Staten
Arbets- och näringsministeriet
Arbets- och näringsministeriet svarar för beredningen av ärenden i anslutning till integrationen av invandrare i Finland.
Kompetenscentret för integration av invandrare stöder arbete som främjar integrationen av invandrare lokalt, regionalt och riksomfattande.
linkkiArbets- och näringsministeriet :
Integration av invandrarefinska _ svenska _ engelska
Undervisnings- och kulturministeriet
Undervisnings- och kulturministeriet svarar för utvecklingen av och det internationella samarbetet inom utbildnings-, vetenskaps-, kultur-, motions- och ungdomspolitiken.
linkkiUndervisnings- och kulturministeriet:
Webbsidorfinska _ svenska _ engelska
Miljöministeriet
linkkiMiljöministeriet:
Webbsidorfinska _ svenska _ engelska
FPA
FPA sköter grundtryggheten i olika skeden av livet för dem som bor i Finland.
FPA:s kunder är alla personer som bor i Finland och utomlands och som omfattas av socialskyddet i Finland.
FPA och Skatteförvaltningen erbjuder information till utländska anställda på servicestället In To Finland i Helsingfors.
Flyttning till eller från Finlandfinska _ svenska _ engelska
Skatteförvaltningen
linkkiSkatteförvaltningen:
Webbsidorfinska _ svenska _ engelska
Kommunerna
Helsingfors stad
Publicerar och administrerar InfoFinland.
Kommuner som är med i samarbetsavtalet
InfoFinlands samarbetsavtal
InfoFinlands finansiärer har ingått ett samarbetsavtal med vilket man överenskommit om principerna för genomförandet och finansieringen av nättjänsten InfoFinland (tidigare Infobanken) för åren 2017–2020.
Samarbetet möjliggör riksomfattande webbinformation för invandrare och personer som planerar att flytta till Finland och för myndigheter inom invandrarsektorn på ett sätt som också stöder behovet av information i kommunerna.
Det är lätt att på ett pålitligt sätt hitta väsentlig information om integration av invandrare och om att bo i Finland på ett ställe, www.infofinland.fi.
Avtalsparterna driver och utvecklar tjänsten tillsammans.
De vill dessutom stärka InfoFinlands riksomfattande ställning, så att det är möjligt för nya kommuner och andra organisationer att ansluta sig till tjänsten också i fortsättningen.
Kommunernas finansieringsandelar fastställs utgående från antalet invånare.
Genomförandet av avtalet följs upp av en styrgrupp.
Nya aktörer är välkomna att utveckla den flerspråkiga informationen till invandrare och ansluta sig till InfoFinlands samarbetsavtal.
Närmare information om hur man ansluter sig till avtalet ger InfoFinlands chefredaktör Eija Kyllönen-Saarnio, eija.kyllonen-saarnio(snabel-a)hel.fi, tfn 050 363 3285.
Alla texter som publicerats på InfoFinlands webbplats på alla språk är fritt tillgängliga i enlighet med licensen Creative Commons Erkännande 4.0.
Du har tillstånd att:
Dela – kopiera och vidaredistribuera materialet oavsett medium eller format
Bearbeta – remixa, transformera, och bygga vidare på materialet för alla ändamål, även kommersiellt.
På följande villkor:
Erkännande (BY) – Du måste nämna källan InfoFinland.fi.
Ange en länk till webbplatsen InfoFinland.fi och nämn licensen CC BY 4.0.
Ange om bearbetningar är gjorda.
Du behöver göra så i enlighet med god sed, och inte på ett sätt som ger en bild av att InfoFinland stödjer dig eller ditt användande.
Inga ytterligare begränsningar – Du får inte tillämpa lagliga begränsningar eller teknologiska metoder som juridiskt begränsar andra från att gör något som licensen tillåter.
Erkännande 4.0 Internationellfinska _ svenska _ engelska _ ryska _ franska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ japanska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ grekiska
_ tjeckiska
Öppet programmeringsgränssnitt (API)
Vi erbjuder allt textinnehåll i InfoFinland via ett öppet programmeringsgränssnitt (API).
Med hjälp av gränssnittet kan du visa InfoFinlands innehåll på andra webbplatser eller skapa olika applikationer.
Information om gränssnittetfinska _ engelska
Öppet programmeringsgränssnittfinska
Alla texter som publicerats på InfoFinlands webbplats på alla språk är fritt tillgängliga i enlighet med licensen Creative Commons Erkännande 4.0.
Du har tillstånd att:
Dela – kopiera och vidaredistribuera materialet oavsett medium eller format
Bearbeta – remixa, transformera, och bygga vidare på materialet för alla ändamål, även kommersiellt.
På följande villkor:
Erkännande (BY) – Du måste nämna källan InfoFinland.fi.
Ange en länk till webbplatsen InfoFinland.fi och nämn licensen CC BY 4.0.
Ange om bearbetningar är gjorda.
Du behöver göra så i enlighet med god sed, och inte på ett sätt som ger en bild av att InfoFinland stödjer dig eller ditt användande.
Inga ytterligare begränsningar – Du får inte tillämpa lagliga begränsningar eller teknologiska metoder som juridiskt begränsar andra från att gör något som licensen tillåter.
Erkännande 4.0 Internationellfinska _ svenska _ engelska _ ryska _ franska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ japanska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ grekiska
_ tjeckiska
Öppet programmeringsgränssnitt (API)
Vi erbjuder allt textinnehåll i InfoFinland via ett öppet programmeringsgränssnitt (API).
Med hjälp av gränssnittet kan du visa InfoFinlands innehåll på andra webbplatser eller skapa olika applikationer.
Information om gränssnittetfinska _ engelska
Öppet programmeringsgränssnittfinska
Användning av InfoFinland-texterna på andra ställen
Texterna ur webbtjänsten InfoFinland.fi används i följande tjänster:
linkkiArbets- och näringsministeriet:
Guiden Välkommen till Finland(pdf, 3,40 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
Alla texter som publicerats på InfoFinlands webbplats på alla språk är fritt tillgängliga i enlighet med licensen Creative Commons Erkännande 4.0.
Du har tillstånd att:
Dela – kopiera och vidaredistribuera materialet oavsett medium eller format
Bearbeta – remixa, transformera, och bygga vidare på materialet för alla ändamål, även kommersiellt.
På följande villkor:
Erkännande (BY) – Du måste nämna källan InfoFinland.fi.
Ange en länk till webbplatsen InfoFinland.fi och nämn licensen CC BY 4.0.
Ange om bearbetningar är gjorda.
Du behöver göra så i enlighet med god sed, och inte på ett sätt som ger en bild av att InfoFinland stödjer dig eller ditt användande.
Inga ytterligare begränsningar – Du får inte tillämpa lagliga begränsningar eller teknologiska metoder som juridiskt begränsar andra från att gör något som licensen tillåter.
Erkännande 4.0 Internationellfinska _ svenska _ engelska _ ryska _ franska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ tyska _ portugisiska _ polska _ norska
_ holländska _ kroatiska _ rumänska _ ungerska _ japanska _ italienska
_ lettiska
_ litauiska
_ danska
_ isländska
_ grekiska
_ tjeckiska
Öppet programmeringsgränssnitt (API)
Vi erbjuder allt textinnehåll i InfoFinland via ett öppet programmeringsgränssnitt (API).
Med hjälp av gränssnittet kan du visa InfoFinlands innehåll på andra webbplatser eller skapa olika applikationer.
Information om gränssnittetfinska _ engelska
Öppet programmeringsgränssnittfinska
Användning av InfoFinland-texterna på andra ställen
Texterna ur webbtjänsten InfoFinland.fi används i följande tjänster:
linkkiArbets- och näringsministeriet:
Guiden Välkommen till Finland(pdf, 3,40 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
Medlemskommunerna har själv hand om översättningen av de övriga kommunsidorna.
Översättningsanvisning:
Översättningsanvisningen är på finska.
Översättningsanvisning:
Översättningsanvisningen är på finska.
Översättningsanvisning:
Översättningsanvisningen är på finska.
Trafik
Beslutsfattande och påverkan
Religion
Grundläggande information
Historia
Trafik
Huvudstadsregionen har goda kollektivtrafikförbindelser.
I Grankulla finns en järnvägsstation och i staden finns många busslinjer.
Du kan söka information om rutterna i tjänsten Reseplaneraren.
Tjänsten ger dig förslag på olika kollektivtrafikförbindelser från ett ställe till ett annat.
Reseplanerarefinska _ svenska _ engelska _ ryska
Inom kollektivtrafiken kan du betala med kontanter eller resekort.
I närtågen måste du köpa biljetten i förväg.
Du kan köpa resekortet på Grankulla stadshus.
Du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat.
Stadshuset
Grankullavägen 10
Mån–fre kl. 8.00–15.00; tis, ons, tors även kl. 17.00–19.30
Den närmaste flygstationen är Helsingfors–Vanda flygplats.
Flygplatsenfinska _ svenska _ engelska _ ryska _ kinesiska
Läs mer:
Trafiken i Finland.
Beslutsfattande och påverkan
I Grankulla beslutas ärenden av stadsfullmäktige.
I stadsfullmäktige sitter 35 ledamöter som representerar olika politiska grupper.
Fullmäktige väljs var fjärde år genom kommunalval.
På Grankulla stads webbplats kan du skicka respons till förvaltningen.
Du kan också lämna initiativ och ställa frågor samt kommentera ärenden på finska och på svenska.
Även engelskspråkiga frågor besvaras.
Delta och påverkafinska _ svenska
Religion
Många religiösa samfund är verksamma i Esbo och Helsingfors.
I tjänsten Uskonnot Suomessa kan du söka information enligt det religiösa samfundet och orten.
Religiösa samfundfinska _ engelska
linkkiHelsingfors ortodoxa församling:
Ortodoxa församlingenfinska _ ryska
I Grankulla finns en evangelisk-luthersk kyrka med två församlingar, en finskspråkig och en svenskspråkig.
Församlingarfinska _ svenska
Läs mer: Kulturer och religioner i Finland.
Grundläggande information
Grankulla är en av de fyra kommunerna i huvudstadsregionen.
Den ligger mitt i Esbo, 15 kilometer västerut från Helsingfors.
Grankulla har cirka 9 600 invånare, varav 60 procent har finska, 36 procent svenska och 4 procent ett annat språk som modersmål.
Grankullas areal är 6,0 km2.
Information om stadenfinska _ svenska _ engelska
Historia
År 1906 grundades ett aktiebolag i Grankulla som sålde villatomter till invånarna i huvudstadsregionen.
Området hade en direkt förbindelse till Helsingfors.
År 1920 blev villasamhället en köping.
Till en början var största delen av invånarna svenskspråkiga.
År 1972 fick köpingen stadsrättigheter.
Nätmuseetfinska _ svenska
Trafik
Beslutsfattande och påverkan
Religion
Grundläggande information
Historia
Trafik
Huvudstadsregionen har goda kollektivtrafikförbindelser.
I Grankulla finns en järnvägsstation och i staden finns många busslinjer.
Du kan söka information om rutterna i tjänsten Reseplaneraren.
Tjänsten ger dig förslag på olika kollektivtrafikförbindelser från ett ställe till ett annat.
Reseplanerarefinska _ svenska _ engelska _ ryska
Inom kollektivtrafiken kan du betala med kontanter eller resekort.
I närtågen måste du köpa biljetten i förväg.
Du kan köpa resekortet på Grankulla stadshus.
Du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat.
Stadshuset
Grankullavägen 10
Mån–fre kl. 8.00–15.00; tis, ons, tors även kl. 17.00–19.30
Den närmaste flygstationen är Helsingfors–Vanda flygplats.
Flygplatsenfinska _ svenska _ engelska _ ryska _ kinesiska
Läs mer:
Trafiken i Finland.
Beslutsfattande och påverkan
I Grankulla beslutas ärenden av stadsfullmäktige.
I stadsfullmäktige sitter 35 ledamöter som representerar olika politiska grupper.
Fullmäktige väljs var fjärde år genom kommunalval.
På Grankulla stads webbplats kan du skicka respons till förvaltningen.
Du kan också lämna initiativ och ställa frågor samt kommentera ärenden på finska och på svenska.
Även engelskspråkiga frågor besvaras.
Delta och påverkafinska _ svenska
Religion
Många religiösa samfund är verksamma i Esbo och Helsingfors.
I tjänsten Uskonnot Suomessa kan du söka information enligt det religiösa samfundet och orten.
Religiösa samfundfinska _ engelska
linkkiHelsingfors ortodoxa församling:
Ortodoxa församlingenfinska _ ryska
I Grankulla finns en evangelisk-luthersk kyrka med två församlingar, en finskspråkig och en svenskspråkig.
Församlingarfinska _ svenska
Läs mer: Kulturer och religioner i Finland.
Grundläggande information
Grankulla är en av de fyra kommunerna i huvudstadsregionen.
Den ligger mitt i Esbo, 15 kilometer västerut från Helsingfors.
Grankulla har cirka 9 600 invånare, varav 60 procent har finska, 36 procent svenska och 4 procent ett annat språk som modersmål.
Grankullas areal är 6,0 km2.
Information om stadenfinska _ svenska _ engelska
Historia
År 1906 grundades ett aktiebolag i Grankulla som sålde villatomter till invånarna i huvudstadsregionen.
Området hade en direkt förbindelse till Helsingfors.
År 1920 blev villasamhället en köping.
Till en början var största delen av invånarna svenskspråkiga.
År 1972 fick köpingen stadsrättigheter.
Nätmuseetfinska _ svenska
Trafik
Beslutsfattande och påverkan
Religion
Grundläggande information
Historia
Trafik
Huvudstadsregionen har goda kollektivtrafikförbindelser.
I Grankulla finns en järnvägsstation och i staden finns många busslinjer.
Du kan söka information om rutterna i tjänsten Reseplaneraren.
Tjänsten ger dig förslag på olika kollektivtrafikförbindelser från ett ställe till ett annat.
Reseplanerarefinska _ svenska _ engelska
Inom kollektivtrafiken kan du betala med kontanter eller resekort.
I närtågen måste du köpa biljetten i förväg.
Du kan köpa resekortet på Grankulla stadshus.
Du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat.
Stadshuset
Grankullavägen 10
Mån–fre kl. 8.00–15.00; tis, ons, tors även kl. 17.00–19.30
Den närmaste flygstationen är Helsingfors–Vanda flygplats.
Flygplatsenfinska _ svenska _ engelska _ ryska _ kinesiska
Läs mer:
Trafiken i Finland.
Beslutsfattande och påverkan
I Grankulla beslutas ärenden av stadsfullmäktige.
I stadsfullmäktige sitter 35 ledamöter som representerar olika politiska grupper.
Fullmäktige väljs var fjärde år genom kommunalval.
På Grankulla stads webbplats kan du skicka respons till förvaltningen.
Du kan också lämna initiativ och ställa frågor samt kommentera ärenden på finska och på svenska.
Även engelskspråkiga frågor besvaras.
Delta och påverkafinska _ svenska
Religion
Många religiösa samfund är verksamma i Esbo och Helsingfors.
I tjänsten Uskonnot Suomessa kan du söka information enligt det religiösa samfundet och orten.
Religiösa samfundfinska _ engelska
linkkiHelsingfors ortodoxa församling:
Ortodoxa församlingenfinska _ ryska
I Grankulla finns en evangelisk-luthersk kyrka med två församlingar, en finskspråkig och en svenskspråkig.
Församlingarfinska _ svenska
Läs mer: Kulturer och religioner i Finland.
Grundläggande information
Grankulla är en av de fyra kommunerna i huvudstadsregionen.
Den ligger mitt i Esbo, 15 kilometer västerut från Helsingfors.
Grankulla har cirka 9 600 invånare, varav 60 procent har finska, 36 procent svenska och 4 procent ett annat språk som modersmål.
Grankullas areal är 6,0 km2.
Information om stadenfinska _ svenska _ engelska
Historia
År 1906 grundades ett aktiebolag i Grankulla som sålde villatomter till invånarna i huvudstadsregionen.
Området hade en direkt förbindelse till Helsingfors.
År 1920 blev villasamhället en köping.
Till en början var största delen av invånarna svenskspråkiga.
År 1972 fick köpingen stadsrättigheter.
Nätmuseetfinska _ svenska
Evenemang
Bibliotek
Fritidsverksamhet för barn och unga
Föreningar
Evenemang
Evenemang i Grankullafinska _ svenska _ engelska
Vid medborgarinstitutet kan man till exempel skapa konst, göra handarbeten, laga mat, dansa eller motionera.
Man kan även studera språk.
Medborgarinstitutetfinska _ svenska _ engelska
Vid musikinstitutet kan man musicera.
Information om Musikinstitutetfinska _ svenska
Grankulla stad ordnar mångsidig kulturverksamhet.
Kulturtjänsterfinska _ svenska _ engelska
I staden finns också många idrottsmöjligheter.
Idrottstjänsterfinska _ svenska _ engelska
Det finns en biograf i Grankulla.
linkkiBio Grani:
Biograffinska
Läs mer: Fritid.
Bibliotek
På Grankulla stadsbibliotek kan du låna böcker, tidningar, musik, filmer, spel och mycket annat.
I biblioteket kan du också använda dator.
Stadsbiblioteketfinska _ svenska _ engelska
Huvudstadsregionens gemensamma bibliotekstjänstfinska _ svenska _ engelska _ somaliska _ persiska _ arabiska
Läs mer: Bibliotek
Flerspråkiga biblioteket
Flerspråkiga biblioteket ligger i Böle i Helsingfors
Här finns böcker, musik, tidningar och tidskrifter samt ljudböcker på flera olika språk.
Du kan åka till Böle eller beställa material till ditt eget närbibliotek.
linkkiHelsingfors stadsbibliotek:
Flerspråkiga biblioteketfinska _ svenska _ engelska
Hobbyer för barn och unga
Barn och ungdomar kan studera musik vid Grankulla musikinstitut och bildkonst vid Grankulla konstskola.
I Grankulla kan man också motionera på många olika sätt.
På Grankulla ungdomsgård ordnas många olika slags verksamheter.
Ungdomsgårdenfinska _ svenska _ engelska
Läs mer: Hobbyer för barn och unga
Föreningar
I Grankulla finns många olika föreningar, till exempel kulturföreningar och idrottsklubbar.
Föreningarfinska _ svenska
Läs mer: Föreningar.
Läs mer: Fritid i Esbo
Evenemang
Bibliotek
Fritidsverksamhet för barn och unga
Föreningar
Evenemang
Evenemang i Grankullafinska _ svenska _ engelska
Vid medborgarinstitutet kan man till exempel skapa konst, göra handarbeten, laga mat, dansa eller motionera.
Man kan även studera språk.
Medborgarinstitutetfinska _ svenska _ engelska
Vid musikinstitutet kan man musicera.
Information om Musikinstitutetfinska _ svenska
Grankulla stad ordnar mångsidig kulturverksamhet.
Kulturtjänsterfinska _ svenska _ engelska
I staden finns också många idrottsmöjligheter.
Idrottstjänsterfinska _ svenska _ engelska
Det finns en biograf i Grankulla.
linkkiBio Grani:
Biograffinska
Läs mer: Fritid.
Bibliotek
På Grankulla stadsbibliotek kan du låna böcker, tidningar, musik, filmer, spel och mycket annat.
I biblioteket kan du också använda dator.
Stadsbiblioteketfinska _ svenska _ engelska
Huvudstadsregionens gemensamma bibliotekstjänstfinska _ svenska _ engelska _ somaliska _ persiska _ arabiska
Läs mer: Bibliotek
Flerspråkiga biblioteket
Flerspråkiga biblioteket ligger i Böle i Helsingfors
Här finns böcker, musik, tidningar och tidskrifter samt ljudböcker på flera olika språk.
Du kan åka till Böle eller beställa material till ditt eget närbibliotek.
linkkiHelsingfors stadsbibliotek:
Flerspråkiga biblioteketfinska _ svenska _ engelska
Hobbyer för barn och unga
Barn och ungdomar kan studera musik vid Grankulla musikinstitut och bildkonst vid Grankulla konstskola.
I Grankulla kan man också motionera på många olika sätt.
På Grankulla ungdomsgård ordnas många olika slags verksamheter.
Ungdomsgårdenfinska _ svenska _ engelska
Läs mer: Hobbyer för barn och unga
Föreningar
I Grankulla finns många olika föreningar, till exempel kulturföreningar och idrottsklubbar.
Föreningarfinska _ svenska
Läs mer: Föreningar.
Läs mer: Fritid i Esbo
Evenemang
Bibliotek
Fritidsverksamhet för barn och unga
Föreningar
Evenemang
Evenemang i Grankullafinska _ svenska _ engelska
Vid medborgarinstitutet kan man till exempel skapa konst, göra handarbeten, laga mat, dansa eller motionera.
Man kan även studera språk.
Medborgarinstitutetfinska _ svenska _ engelska
Vid musikinstitutet kan man musicera.
Information om Musikinstitutetfinska _ svenska
Grankulla stad ordnar mångsidig kulturverksamhet.
Kulturtjänsterfinska _ svenska _ engelska
I staden finns också många idrottsmöjligheter.
Idrottstjänsterfinska _ svenska _ engelska
Det finns en biograf i Grankulla.
linkkiBio Grani:
Biograffinska
Läs mer: Fritid.
Bibliotek
På Grankulla stadsbibliotek kan du låna böcker, tidningar, musik, filmer, spel och mycket annat.
I biblioteket kan du också använda dator.
Stadsbiblioteketfinska _ svenska _ engelska
Huvudstadsregionens gemensamma bibliotekstjänstfinska _ svenska _ engelska _ somaliska _ persiska _ arabiska
Läs mer: Bibliotek
Flerspråkiga biblioteket
Flerspråkiga biblioteket ligger i Böle i Helsingfors
Här finns böcker, musik, tidningar och tidskrifter samt ljudböcker på flera olika språk.
Du kan åka till Böle eller beställa material till ditt eget närbibliotek.
linkkiHelsingfors stadsbibliotek:
Flerspråkiga biblioteketfinska _ svenska _ engelska
Hobbyer för barn och unga
Barn och ungdomar kan studera musik vid Grankulla musikinstitut och bildkonst vid Grankulla konstskola.
I Grankulla kan man också motionera på många olika sätt.
På Grankulla ungdomsgård ordnas många olika slags verksamheter.
Ungdomsgårdenfinska _ svenska _ engelska
Läs mer: Hobbyer för barn och unga
Föreningar
I Grankulla finns många olika föreningar, till exempel kulturföreningar och idrottsklubbar.
Föreningarfinska _ svenska
Läs mer: Föreningar.
Läs mer: Fritid i Esbo
Social- och krisjouren
Problem med uppehållstillstånd
Brott
Våld
Problem i äktenskap och parförhållande
Behöver du juristhjälp? Barns och ungas problem
Död
Ring nödnumret 112 om det är fråga om en nödsituation.
Via nödnumret kan du tillkalla polis, ambulans eller brandkår.
Ring inte nödnumret om det inte är en nödsituation.
Social- och krisjouren
Social- och krisjouren vid Jorv sjukhus i Esbo hjälper dygnet runt om du eller din familj behöver hjälp i en akut krissituation, till exempel vid våld, problem med barnen eller psykiska problem.
I krissituationer kan du ringa eller åka till jouren.
Esbo social- och krisjour
Jorv sjukhus, Åbovägen 150, Esbo
Tfn (09) 816 42439
Vardagar kl. 15–08, fre–sön och helgdagar dygnet runt
linkkiEsbo stad:
Social- och krisjourenfinska _ svenska _ engelska
linkkiFöreningen för mental hälsa i Finland:
Krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Problem med uppehållstillstånd
Om du har problem med eller det råder oklarheter kring uppehållstillståndet kan du ta kontakt med Migrationsverket, Flyktingrådgivningen eller Helsingfors stads Helsinki-info.
Läs mer: Problem med uppehållstillstånd
Information om uppehållstillståndfinska _ svenska _ engelska
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Helsingfors-infofinska _ svenska _ engelska
Brott
Om du blir utsatt för ett brott, gör en brottsanmälan hos polisen.
Du kan göra brottsanmälan på internet.
Du kan även fylla i en blankett och lämna den till Esbo huvudpolisstation.
Esbo huvudpolisstation
Knektbrovägen 4
Läs mer: Brott
Kontaktuppgifterfinska _ svenska _ engelska
Elektronisk polisanmälanfinska _ svenska _ engelska
Behöver du en jurist?
Västra Nylands rättshjälpsbyrå betjänar invånarna i Grankulla.
Västra Nylands rättshjälpsbyrå
Östanvindsvägen 1 A
Tfn 029 56 61820.
linkkiVästra Nylands rättshjälpsbyrå:
Läs mer:
Behöver du en jurist?
Våld
Om du behöver brådskande hjälp av polisen i nödsituationer, ring nödnumret 112.
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kontakta ett skyddshem.
Tfn (09) 4777 180 (24h)
Hjälp till offer för familjevåldfinska
Föreningen Monika-Naiset Liitto har en jourtelefon för invandrarkvinnor som blivit utsatta för våld.
Tfn 0800 05058
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Invandrarmän som har problem med våld kan få hjälp via tjänsten Miehen linja.
Tfn (09) 276 62899
Hjälp för invandrarmänfinska _ engelska
Läs mer: Våld
Problem i äktenskap och parförhållande
Vid problem i äktenskap och parförhållande kan du få hjälp vid familjerådgivningen.
Familjerådgivningen betjänar invånarna i Grankulla.
Familjerådgivningen
Tfn (09) 5056 297
Familjerådgivningfinska _ svenska
Problem i äktenskap och parförhållande
Barns och ungas problem
Vid problem som gäller barn under skolåldern, kontakta barnrådgivningen.
Barnrådgivningen
Tfn (09) 5056 357 eller (09) 5056 358
Rådgivningsbyråerfinska _ svenska _ engelska
Vid problem som gäller barn i skolåldern hjälper till exempel skolans hälsovårdare.
Skolhälsovårdenfinska _ svenska
Om du behöver råd i frågor kring barns psykiska tillväxt och utveckling, kan du boka en tid hos familjerådgivningen.
Familjerådgivningfinska _ svenska
Du kan prata om dina problem med skolans eller läroanstaltens hälsovårdare eller de vuxna vid ungdomsgården.
Den unga själv eller föräldrarna kan också kontakta familjerådgivningen.
En ung som inte är trygg i sitt eget hem kan kontakta Finlands Röda Kors De ungas skyddshus.
Skyddshuset finns i Stensvik.
De ungas skyddshus
Tfn (09) 8195 5360
linkkiFinlands Röda Kors:
De ungas skyddshusfinska
Läs mer: Barns och ungas problem
Död
Om en nära anhörig till dig avlider oväntat, kan du få stöd av Grankullas grupp för krisbearbetning, tfn 050 344 6652.
Grankulla stad har en egen begravningsplats i Kasabergsområdet.
Den är avsedd för stadens invånare.
Läs mer: Död
Social- och krisjouren
Problem med uppehållstillstånd
Brott
Våld
Problem i äktenskap och parförhållande
Behöver du juristhjälp? Barns och ungas problem
Död
Ring nödnumret 112 om det är fråga om en nödsituation.
Via nödnumret kan du tillkalla polis, ambulans eller brandkår.
Ring inte nödnumret om det inte är en nödsituation.
Social- och krisjouren
Social- och krisjouren vid Jorv sjukhus i Esbo hjälper dygnet runt om du eller din familj behöver hjälp i en akut krissituation, till exempel vid våld, problem med barnen eller psykiska problem.
I krissituationer kan du ringa eller åka till jouren.
Esbo social- och krisjour
Jorv sjukhus, Åbovägen 150, Esbo
Tfn (09) 816 42439
Vardagar kl. 15–08, fre–sön och helgdagar dygnet runt
linkkiEsbo stad:
Social- och krisjourenfinska _ svenska _ engelska
linkkiFöreningen för mental hälsa i Finland:
Krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Problem med uppehållstillstånd
Om du har problem med eller det råder oklarheter kring uppehållstillståndet kan du ta kontakt med Migrationsverket, Flyktingrådgivningen eller Helsingfors stads Helsinki-info.
Läs mer: Problem med uppehållstillstånd
Information om uppehållstillståndfinska _ svenska _ engelska
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Helsingfors-infofinska _ svenska _ engelska
Brott
Om du blir utsatt för ett brott, gör en brottsanmälan hos polisen.
Du kan göra brottsanmälan på internet.
Du kan även fylla i en blankett och lämna den till Esbo huvudpolisstation.
Esbo huvudpolisstation
Knektbrovägen 4
Läs mer: Brott
Kontaktuppgifterfinska _ svenska _ engelska
Elektronisk polisanmälanfinska _ svenska _ engelska
Behöver du en jurist?
Västra Nylands rättshjälpsbyrå betjänar invånarna i Grankulla.
Västra Nylands rättshjälpsbyrå
Östanvindsvägen 1 A
Tfn 029 56 61820.
linkkiVästra Nylands rättshjälpsbyrå:
Läs mer:
Behöver du en jurist?
Våld
Om du behöver brådskande hjälp av polisen i nödsituationer, ring nödnumret 112.
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kontakta ett skyddshem.
Tfn (09) 4777 180 (24h)
Hjälp till offer för familjevåldfinska
Föreningen Monika-Naiset Liitto har en jourtelefon för invandrarkvinnor som blivit utsatta för våld.
Tfn 0800 05058
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Invandrarmän som har problem med våld kan få hjälp via tjänsten Miehen linja.
Tfn (09) 276 62899
Hjälp för invandrarmänfinska _ engelska
Läs mer: Våld
Problem i äktenskap och parförhållande
Vid problem i äktenskap och parförhållande kan du få hjälp vid familjerådgivningen.
Familjerådgivningen betjänar invånarna i Grankulla.
Familjerådgivningen
Tfn (09) 5056 297
Familjerådgivningfinska _ svenska
Problem i äktenskap och parförhållande
Barns och ungas problem
Vid problem som gäller barn under skolåldern, kontakta barnrådgivningen.
Barnrådgivningen
Tfn (09) 5056 357 eller (09) 5056 358
Rådgivningsbyråerfinska _ svenska _ engelska
Vid problem som gäller barn i skolåldern hjälper till exempel skolans hälsovårdare.
Skolhälsovårdenfinska _ svenska
Om du behöver råd i frågor kring barns psykiska tillväxt och utveckling, kan du boka en tid hos familjerådgivningen.
Familjerådgivningfinska _ svenska
Du kan prata om dina problem med skolans eller läroanstaltens hälsovårdare eller de vuxna vid ungdomsgården.
Den unga själv eller föräldrarna kan också kontakta familjerådgivningen.
En ung som inte är trygg i sitt eget hem kan kontakta Finlands Röda Kors De ungas skyddshus.
Skyddshuset finns i Stensvik.
De ungas skyddshus
Tfn (09) 8195 5360
linkkiFinlands Röda Kors:
De ungas skyddshusfinska
Läs mer: Barns och ungas problem
Död
Om en nära anhörig till dig avlider oväntat, kan du få stöd av Grankullas grupp för krisbearbetning, tfn 050 344 6652.
Grankulla stad har en egen begravningsplats i Kasabergsområdet.
Den är avsedd för stadens invånare.
Läs mer: Död
Social- och krisjouren
Problem med uppehållstillstånd
Brott
Våld
Problem i äktenskap och parförhållande
Behöver du juristhjälp? Barns och ungas problem
Död
Ring nödnumret 112 om det är fråga om en nödsituation.
Via nödnumret kan du tillkalla polis, ambulans eller brandkår.
Ring inte nödnumret om det inte är en nödsituation.
Social- och krisjouren
Social- och krisjouren vid Jorv sjukhus i Esbo hjälper dygnet runt om du eller din familj behöver hjälp i en akut krissituation, till exempel vid våld, problem med barnen eller psykiska problem.
I krissituationer kan du ringa eller åka till jouren.
Esbo social- och krisjour
Jorv sjukhus, Åbovägen 150, Esbo
Tfn (09) 816 42439
Vardagar kl. 15–08, fre–sön och helgdagar dygnet runt
linkkiEsbo stad:
Social- och krisjourenfinska _ svenska _ engelska
linkkiFöreningen för mental hälsa i Finland:
Krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Problem med uppehållstillstånd
Om du har problem med eller det råder oklarheter kring uppehållstillståndet kan du ta kontakt med Migrationsverket, Flyktingrådgivningen eller Helsingfors stads Helsinki-info.
Läs mer: Problem med uppehållstillstånd
Information om uppehållstillståndfinska _ svenska _ engelska
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Helsingfors-infofinska _ svenska _ engelska
Brott
Om du blir utsatt för ett brott, gör en brottsanmälan hos polisen.
Du kan göra brottsanmälan på internet.
Du kan även fylla i en blankett och lämna den till Esbo huvudpolisstation.
Esbo huvudpolisstation
Knektbrovägen 4
Läs mer: Brott
Kontaktuppgifterfinska _ svenska _ engelska
Elektronisk polisanmälanfinska _ svenska _ engelska
Behöver du en jurist?
Västra Nylands rättshjälpsbyrå betjänar invånarna i Grankulla.
Västra Nylands rättshjälpsbyrå
Östanvindsvägen 1 A
Tfn 029 56 61820.
linkkiVästra Nylands rättshjälpsbyrå:
Läs mer:
Behöver du en jurist?
Våld
Om du behöver brådskande hjälp av polisen i nödsituationer, ring nödnumret 112.
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kontakta ett skyddshem.
Tfn (09) 4777 180 (24h)
Hjälp till offer för familjevåldfinska
Föreningen Monika-Naiset Liitto har en jourtelefon för invandrarkvinnor som blivit utsatta för våld.
Tfn 0800 05058
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Invandrarmän som har problem med våld kan få hjälp via tjänsten Miehen linja.
Tfn (09) 276 62899
Hjälp för invandrarmänfinska _ engelska
Läs mer: Våld
Problem i äktenskap och parförhållande
Vid problem i äktenskap och parförhållande kan du få hjälp vid familjerådgivningen.
Familjerådgivningen betjänar invånarna i Grankulla.
Familjerådgivningen
Tfn (09) 5056 297
Familjerådgivningfinska _ svenska
Problem i äktenskap och parförhållande
Barns och ungas problem
Vid problem som gäller barn under skolåldern, kontakta barnrådgivningen.
Barnrådgivningen
Tfn (09) 5056 357 eller (09) 5056 358
Rådgivningsbyråerfinska _ svenska _ engelska
Vid problem som gäller barn i skolåldern hjälper till exempel skolans hälsovårdare.
Skolhälsovårdenfinska _ svenska
Om du behöver råd i frågor kring barns psykiska tillväxt och utveckling, kan du boka en tid hos familjerådgivningen.
Familjerådgivningfinska _ svenska
Du kan prata om dina problem med skolans eller läroanstaltens hälsovårdare eller de vuxna vid ungdomsgården.
Den unga själv eller föräldrarna kan också kontakta familjerådgivningen.
En ung som inte är trygg i sitt eget hem kan kontakta Finlands Röda Kors De ungas skyddshus.
Skyddshuset finns i Stensvik.
De ungas skyddshus
Tfn (09) 8195 5360
linkkiFinlands Röda Kors:
De ungas skyddshusfinska
Läs mer: Barns och ungas problem
Död
Om en nära anhörig till dig avlider oväntat, kan du få stöd av Grankullas grupp för krisbearbetning, tfn 050 344 6652.
Grankulla stad har en egen begravningsplats i Kasabergsområdet.
Den är avsedd för stadens invånare.
Läs mer: Död
Äktenskap
Skilsmässa
Barn vid skilsmässa
Vård av barnet
Äktenskap
Före äktenskapet ska du skriftligt begära prövning av hinder mot äktenskap.
Hindersprövningen görs i magistraten.
Läs mer: Prövning av hinder mot äktenskap, Äktenskap
Kontaktuppgifter till magistratfinska _ svenska _ engelska
Skilsmässa
Kvinnan eller mannen kan lämna in skilsmässoansökan i Västra Nylands tingsrätts kansli.
Du kan också söka skilsmässa ensam, utan din makes eller makas samtycke.
Du kan skicka in ansökan till tingsrättens kansli per post, fax eller via e-post.
Västra Nylands tingsrätt
Tfn 029 5645 000
Läs mer: Skilsmässa
linkkiVästra Nylands tingsrätt:
Kontaktuppgifterfinska _ svenska
Barn vid skilsmässa
Om du har barn och ska skilja dig, ta kontakt med barnatillsyningsmannen.
Socialväsendet bekräftar ett avtal om barnens boende, vårdnad, umgängesrätt och underhållsbidrag.
Läs mer: Barn vid skilsmässa
Vårdnad om barn och umgängesrättfinska _ svenska
Vård av barnet
På InfoFinlands sida Utbildning i Grankulla finns information om dagvård för barn.
Vård av barnet i hemmet
Om du sköter ditt barn hemma kan du delta i Grankulla stads öppna familjeverksamhet. Där kan du träffa andra barnfamiljer.
Läs mer: Stöd för vård av barn i hemmet
Öppen familjeverksamhetfinska _ svenska
Stöd för hemvård av barnfinska _ svenska
Äktenskap
Skilsmässa
Barn vid skilsmässa
Vård av barnet
Äktenskap
Före äktenskapet ska du skriftligt begära prövning av hinder mot äktenskap.
Hindersprövningen görs i magistraten.
Läs mer: Prövning av hinder mot äktenskap, Äktenskap
Kontaktuppgifter till magistratfinska _ svenska _ engelska
Skilsmässa
Kvinnan eller mannen kan lämna in skilsmässoansökan i Västra Nylands tingsrätts kansli.
Du kan också söka skilsmässa ensam, utan din makes eller makas samtycke.
Du kan skicka in ansökan till tingsrättens kansli per post, fax eller via e-post.
Västra Nylands tingsrätt
Tfn 029 5645 000
Läs mer: Skilsmässa
linkkiVästra Nylands tingsrätt:
Kontaktuppgifterfinska _ svenska
Barn vid skilsmässa
Om du har barn och ska skilja dig, ta kontakt med barnatillsyningsmannen.
Socialväsendet bekräftar ett avtal om barnens boende, vårdnad, umgängesrätt och underhållsbidrag.
Läs mer: Barn vid skilsmässa
Vårdnad om barn och umgängesrättfinska _ svenska
Vård av barnet
På InfoFinlands sida Utbildning i Grankulla finns information om dagvård för barn.
Vård av barnet i hemmet
Om du sköter ditt barn hemma kan du delta i Grankulla stads öppna familjeverksamhet. Där kan du träffa andra barnfamiljer.
Läs mer: Stöd för vård av barn i hemmet
Öppen familjeverksamhetfinska _ svenska
Stöd för hemvård av barnfinska _ svenska
Äktenskap
Skilsmässa
Barn vid skilsmässa
Vård av barnet
Äktenskap
Före äktenskapet ska du skriftligt begära prövning av hinder mot äktenskap.
Hindersprövningen görs i magistraten.
Läs mer: Prövning av hinder mot äktenskap, Äktenskap
Kontaktuppgifter till magistratfinska _ svenska _ engelska
Skilsmässa
Kvinnan eller mannen kan lämna in skilsmässoansökan i Västra Nylands tingsrätts kansli.
Du kan också söka skilsmässa ensam, utan din makes eller makas samtycke.
Du kan skicka in ansökan till tingsrättens kansli per post, fax eller via e-post.
Västra Nylands tingsrätt
Tfn 029 5645 000
Läs mer: Skilsmässa
linkkiVästra Nylands tingsrätt:
Kontaktuppgifterfinska _ svenska
Barn vid skilsmässa
Om du har barn och ska skilja dig, ta kontakt med barnatillsyningsmannen.
Socialväsendet bekräftar ett avtal om barnens boende, vårdnad, umgängesrätt och underhållsbidrag.
Läs mer: Barn vid skilsmässa
Vårdnad om barn och umgängesrättfinska _ svenska
Vård av barnet
På InfoFinlands sida Utbildning i Grankulla finns information om dagvård för barn.
Vård av barnet i hemmet
Om du sköter ditt barn hemma kan du delta i Grankulla stads öppna familjeverksamhet. Där kan du träffa andra barnfamiljer.
Läs mer: Stöd för vård av barn i hemmet
Öppen familjeverksamhetfinska _ svenska
Stöd för hemvård av barnfinska _ svenska
Hälsovårdstjänsterna i Grankulla
Barns hälsa
Äldre människors hälsa
Tandvård
Mental hälsa
Sexualhälsa
När du väntar barn
Handikappade personer
Ring nödnumret 112 om det är fråga om en brådskande nödsituation.
Ring nödnumret till exempel vid en allvarlig olycka eller när någon drabbas av en sjukdomsattack.
Ring inte nödnumret om det inte är en nödsituation.
Om du har din hemkommun i Grankulla, kan du utnyttja de offentliga hälso- och sjukvårdstjänsterna.
Offentliga hälso- och sjukvårdstjänster tillhandahålls till exempel vid hälsostationer, tandkliniker, rådgivningsbyråer och sjukhus.
Om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna, kan du söka dig till en privat läkarstation.
På en privat läkarstation måste du betala samtliga kostnader själv.
Läs mer: Hälsa
Hälsovårdstjänsterna i Grankulla
I Grankulla tillhandahålls offentliga hälso- och sjukvårdstjänster på hälsostationen.
På hälsostationen finns läkarens, sjukskötarens och hälsovårdarens mottagningar.
Hälsostationen har öppet vardagar kl. 8.00–16.00.
Om du behöver vård under samma dag ska du kontakta hälsostationen direkt på morgonen när hälsostationen öppnar.
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
Tfn (09) 8789 1300
Hälsostationenfinska _ svenska _ engelska
Privata hälsotjänster
Information om privata hälsotjänster hittar du på sidorna Hälsa i Esbo och Hälsa i Helsingfors.
Läkemedel
Du kan köpa läkemedel på apoteket.
Adressen till apoteket i Grankulla är Kyrkovägen 15, Grankulla.
Läs mer: Läkemedel.
Apotekfinska _ svenska
linkkiApotekareförbundet:
Hälsovård för papperslösa
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärvård.
Tfn 044 977 4547
Kontaktuppgifterfinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Läs mer: Hälsovårdstjänster i Finland
Kvällstid och under veckoslut har hälsostationen stängt.
Då vårdas akuta sjukdomar och olycksfall på jourmottagningen.
Den närmaste jourmottagningen finns vid Jorv sjukhus i Esbo.
Ring den kostnadsfria Jourhjälpen på tfn 116 117 innan du kommer till jourmottagningen.
Jouren vid Jorv sjukhus
Åbovägen 150
Tfn (09) 4711
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Jourfinska _ svenska _ engelska
Läs mer: Hälsovårdstjänster i Finland
Barns hälsa
I hälso- och sjukvården av barn under skolåldern får man hjälp av rådgivningens hälsovårdare och läkare.
Dem kan du fråga om råd och få stöd i föräldraskapet och fostran av barn.
På rådgivningsbyrån följs barnets hälsa och tillväxt.
Rådgivningsbyråerfinska _ svenska _ engelska
När barnet blir sjukt ska du vid behov kontakta Grankulla hälsostation.
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
Tfn (09) 8789 1300
Hälsostationenfinska _ svenska _ engelska
Skolhälsovårdaren tar hand om skolbarns hälsa.
Skolhälsovårdenfinska _ svenska
Under kvällar och veckoslut finns jourmottagningen för barn under 16 år vid Jorv sjukhus i Esbo och på Barnkliniken i Helsingfors.
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Jourmottagning för barnfinska _ svenska _ engelska
Läs mer: Barns hälsa
Äldre människors hälsa
Om du är över 65 år kan du kontakta seniorrådgivningen vid Grankulla hälsostation.
Seniorrådgivningenfinska _ svenska
Serviceguide för seniorer(pdf, 1,8 MB)finska _ svenska
Tandvård
Tidsbeställningen till tandkliniken vid Grankulla hälsostation mån–fre:
Tfn (09) 505 6379
Jourmottagningen vid Haartmanska sjukhuset har öppet vardagar kl. 14–21 och lör–sön kl. 8–21.
Tfn (09) 310 49999
Mun- och tandhälsovårdenfinska _ svenska
Privat tandvård
I Grankulla finns också privata tandläkare.
Om om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna, kan du gå till en privat tandläkare.
Privat tandvård är dyrare än offentlig tandvård.
Privat tandläkarefinska _ svenska
Läs mer: Tandvård
Mental hälsa
Om du behöver psykisk hjälp och psykiskt stöd kan du kontakta hälsostationen.
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
Tfn (09) 5056 600
Mental hälsafinska _ svenska
Esbo social- och krisjour vid Jorv sjukhus betjänar personer som bor i Grankulla.
I krissituationer kan du ringa eller åka till jouren.
Esbo social- och krisjour
Jorv sjukhus, Åbovägen 150, Esbo
Tfn (09) 816 42439
Vardagar kl. 15–08, fre–sön och helgdagar dygnet runt
Kristjänsterfinska _ svenska
Läs mer: Mental hälsa
Sexualhälsa
Vid mödra- och preventivrådgivningen får du hjälp med graviditetsprevention och familjeplanering.
Könssjukdomar behandlas på hälsostationen och på polikliniken för könssjukdomar i Helsingfors. .
Hälsostationenfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Polikliniken för könssjukdomarfinska _ svenska _ engelska
När du väntar barn
Vid mödrarådgivningen följs moderns, fostrets och hela familjens hälsotillstånd under graviditeten.
Kontakta rådgivningsbyrån när du upptäcker att du är gravid.
Tidsbokning vardagar kl. 12–13
Tfn (09) 8789 1344
Rådgivningsbyråerfinska _ svenska _ engelska
Det närmaste förlossningssjukhuset är Jorv sjukhus i Esbo.
Om du vill kan du även föda barnet på något annat sjukhus inom Helsingfors och Nylands sjukvårdsdistrikt (HNS).
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Val av förlossningssjukhusfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Läs mer: Förlossning
Handikappade personer
Grankulla stad erbjuder olika tjänster för handikappade, till exempel hjälpmedel och dagverksamhet.
Du kan fråga om tjänsterna för handikappade hos socialarbetaren för ditt område.
Tjänster inom handikappvårdenfinska _ svenska
Läs mer: Handikappade personer
Hälsovårdstjänsterna i Grankulla
Barns hälsa
Äldre människors hälsa
Tandvård
Mental hälsa
Sexualhälsa
När du väntar barn
Handikappade personer
Ring nödnumret 112 om det är fråga om en brådskande nödsituation.
Ring nödnumret till exempel vid en allvarlig olycka eller när någon drabbas av en sjukdomsattack.
Ring inte nödnumret om det inte är en nödsituation.
Om du har din hemkommun i Grankulla, kan du utnyttja de offentliga hälso- och sjukvårdstjänsterna.
Offentliga hälso- och sjukvårdstjänster tillhandahålls till exempel vid hälsostationer, tandkliniker, rådgivningsbyråer och sjukhus.
Om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna, kan du söka dig till en privat läkarstation.
På en privat läkarstation måste du betala samtliga kostnader själv.
Läs mer: Hälsa
Hälsovårdstjänsterna i Grankulla
I Grankulla tillhandahålls offentliga hälso- och sjukvårdstjänster på hälsostationen.
På hälsostationen finns läkarens, sjukskötarens och hälsovårdarens mottagningar.
Hälsostationen har öppet vardagar kl. 8.00–16.00.
Om du behöver vård under samma dag ska du kontakta hälsostationen direkt på morgonen när hälsostationen öppnar.
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
Tfn (09) 8789 1300
Hälsostationenfinska _ svenska _ engelska
Privata hälsotjänster
Information om privata hälsotjänster hittar du på sidorna Hälsa i Esbo och Hälsa i Helsingfors.
Läkemedel
Du kan köpa läkemedel på apoteket.
Adressen till apoteket i Grankulla är Kyrkovägen 15, Grankulla.
Läs mer: Läkemedel.
Apotekfinska _ svenska
linkkiApotekareförbundet:
Hälsovård för papperslösa
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärvård.
Tfn 044 977 4547
Kontaktuppgifterfinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Läs mer: Hälsovårdstjänster i Finland
Kvällstid och under veckoslut har hälsostationen stängt.
Då vårdas akuta sjukdomar och olycksfall på jourmottagningen.
Den närmaste jourmottagningen finns vid Jorv sjukhus i Esbo.
Ring den kostnadsfria Jourhjälpen på tfn 116 117 innan du kommer till jourmottagningen.
Jouren vid Jorv sjukhus
Åbovägen 150
Tfn (09) 4711
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Jourfinska _ svenska _ engelska
Läs mer: Hälsovårdstjänster i Finland
Barns hälsa
I hälso- och sjukvården av barn under skolåldern får man hjälp av rådgivningens hälsovårdare och läkare.
Dem kan du fråga om råd och få stöd i föräldraskapet och fostran av barn.
På rådgivningsbyrån följs barnets hälsa och tillväxt.
Rådgivningsbyråerfinska _ svenska _ engelska
När barnet blir sjukt ska du vid behov kontakta Grankulla hälsostation.
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
Tfn (09) 8789 1300
Hälsostationenfinska _ svenska _ engelska
Skolhälsovårdaren tar hand om skolbarns hälsa.
Skolhälsovårdenfinska _ svenska
Under kvällar och veckoslut finns jourmottagningen för barn under 16 år vid Jorv sjukhus i Esbo och på Barnkliniken i Helsingfors.
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Jourmottagning för barnfinska _ svenska _ engelska
Läs mer: Barns hälsa
Äldre människors hälsa
Om du är över 65 år kan du kontakta seniorrådgivningen vid Grankulla hälsostation.
Information om tjänster för äldrefinska _ svenska
Serviceguide för seniorer(pdf, 1,8 MB)finska _ svenska
Äldre människor
Tandvård
Tidsbeställningen till tandkliniken vid Grankulla hälsostation mån–fre:
Tfn (09) 505 6379
Jourmottagningen vid Haartmanska sjukhuset har öppet vardagar kl. 14–21 och lör–sön kl. 8–21.
Tfn (09) 310 49999
Mun- och tandhälsovårdenfinska _ svenska
Privat tandvård
I Grankulla finns också privata tandläkare.
Om om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna, kan du gå till en privat tandläkare.
Privat tandvård är dyrare än offentlig tandvård.
Privat tandläkarefinska _ svenska
Läs mer: Tandvård
Mental hälsa
Om du behöver psykisk hjälp och psykiskt stöd kan du kontakta hälsostationen.
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
Tfn (09) 5056 600
Mental hälsafinska _ svenska
Esbo social- och krisjour vid Jorv sjukhus betjänar personer som bor i Grankulla.
I krissituationer kan du ringa eller åka till jouren.
Esbo social- och krisjour
Jorv sjukhus, Åbovägen 150, Esbo
Tfn (09) 816 42439
Vardagar kl. 15–08, fre–sön och helgdagar dygnet runt
Kristjänsterfinska _ svenska
Läs mer: Mental hälsa
Sexualhälsa
Vid mödra- och preventivrådgivningen får du hjälp med graviditetsprevention och familjeplanering.
Könssjukdomar behandlas på hälsostationen och på polikliniken för könssjukdomar i Helsingfors. .
Hälsostationenfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Polikliniken för könssjukdomarfinska _ svenska _ engelska
När du väntar barn
Vid mödrarådgivningen följs moderns, fostrets och hela familjens hälsotillstånd under graviditeten.
Kontakta rådgivningsbyrån när du upptäcker att du är gravid.
Tidsbokning vardagar kl. 12–13
Tfn (09) 8789 1344
Rådgivningsbyråerfinska _ svenska _ engelska
Det närmaste förlossningssjukhuset är Jorv sjukhus i Esbo.
Om du vill kan du även föda barnet på något annat sjukhus inom Helsingfors och Nylands sjukvårdsdistrikt (HNS).
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Val av förlossningssjukhusfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Läs mer: Förlossning
Handikappade personer
Grankulla stad erbjuder olika tjänster för handikappade, till exempel hjälpmedel och dagverksamhet.
Du kan fråga om tjänsterna för handikappade hos socialarbetaren för ditt område.
Tjänster inom handikappvårdenfinska _ svenska
Läs mer: Handikappade personer
Hälsovårdstjänsterna i Grankulla
Barns hälsa
Äldre människors hälsa
Tandvård
Mental hälsa
Sexualhälsa
När du väntar barn
Handikappade personer
Ring nödnumret 112 om det är fråga om en brådskande nödsituation.
Ring nödnumret till exempel vid en allvarlig olycka eller när någon drabbas av en sjukdomsattack.
Ring inte nödnumret om det inte är en nödsituation.
Om du har din hemkommun i Grankulla, kan du utnyttja de offentliga hälso- och sjukvårdstjänsterna.
Offentliga hälso- och sjukvårdstjänster tillhandahålls till exempel vid hälsostationer, tandkliniker, rådgivningsbyråer och sjukhus.
Om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna, kan du söka dig till en privat läkarstation.
På en privat läkarstation måste du betala samtliga kostnader själv.
Läs mer: Hälsa
Hälsovårdstjänsterna i Grankulla
I Grankulla tillhandahålls offentliga hälso- och sjukvårdstjänster på hälsostationen.
På hälsostationen finns läkarens, sjukskötarens och hälsovårdarens mottagningar.
Hälsostationen har öppet vardagar kl. 8.00–16.00.
Om du behöver vård under samma dag ska du kontakta hälsostationen direkt på morgonen när hälsostationen öppnar.
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
Tfn (09) 8789 1300
Hälsostationenfinska _ svenska
Privata hälsotjänster
Information om privata hälsotjänster hittar du på sidorna Hälsa i Esbo och Hälsa i Helsingfors.
Läkemedel
Du kan köpa läkemedel på apoteket.
Adressen till apoteket i Grankulla är Kyrkovägen 15, Grankulla.
Läs mer: Läkemedel.
Apotekfinska _ svenska
linkkiApotekareförbundet:
Hälsovård för papperslösa
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärvård.
Tfn 044 977 4547
Kontaktuppgifterfinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Läs mer: Hälsovårdstjänster i Finland
Kvällstid och under veckoslut har hälsostationen stängt.
Då vårdas akuta sjukdomar och olycksfall på jourmottagningen.
Den närmaste jourmottagningen finns vid Jorv sjukhus i Esbo.
Ring den kostnadsfria Jourhjälpen på tfn 116 117 innan du kommer till jourmottagningen.
Jouren vid Jorv sjukhus
Åbovägen 150
Tfn (09) 4711
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Jourfinska _ svenska _ engelska
Läs mer: Hälsovårdstjänster i Finland
Barns hälsa
I hälso- och sjukvården av barn under skolåldern får man hjälp av rådgivningens hälsovårdare och läkare.
Dem kan du fråga om råd och få stöd i föräldraskapet och fostran av barn.
På rådgivningsbyrån följs barnets hälsa och tillväxt.
Rådgivningsbyråerfinska _ svenska _ engelska
När barnet blir sjukt ska du vid behov kontakta Grankulla hälsostation.
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
Tfn (09) 8789 1300
Hälsostationenfinska _ svenska
Skolhälsovårdaren tar hand om skolbarns hälsa.
Skolhälsovårdenfinska _ svenska
Under kvällar och veckoslut finns jourmottagningen för barn under 16 år vid Jorv sjukhus i Esbo och på Barnkliniken i Helsingfors.
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Jourmottagning för barnfinska _ svenska _ engelska
Läs mer: Barns hälsa
Äldre människors hälsa
Om du är över 65 år kan du kontakta seniorrådgivningen vid Grankulla hälsostation.
Information om tjänster för äldrefinska _ svenska
Äldre människor
Tandvård
Tidsbeställningen till tandkliniken vid Grankulla hälsostation mån–fre:
Tfn (09) 505 6379
Jourmottagningen vid Haartmanska sjukhuset har öppet vardagar kl. 14–21 och lör–sön kl. 8–21.
Tfn (09) 310 49999
Mun- och tandhälsovårdenfinska _ svenska
Privat tandvård
I Grankulla finns också privata tandläkare.
Om om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna, kan du gå till en privat tandläkare.
Privat tandvård är dyrare än offentlig tandvård.
Privat tandläkarefinska _ svenska
Läs mer: Tandvård
Mental hälsa
Om du behöver psykisk hjälp och psykiskt stöd kan du kontakta hälsostationen.
Grankulla hälsostation
Stationsvägen 19
02700 Grankulla
Tfn (09) 5056 600
Mental hälsafinska _ svenska
Esbo social- och krisjour vid Jorv sjukhus betjänar personer som bor i Grankulla.
I krissituationer kan du ringa eller åka till jouren.
Esbo social- och krisjour
Jorv sjukhus, Åbovägen 150, Esbo
Tfn (09) 816 42439
Vardagar kl. 15–08, fre–sön och helgdagar dygnet runt
Kristjänsterfinska _ svenska
Läs mer: Mental hälsa
Sexualhälsa
Vid mödra- och preventivrådgivningen får du hjälp med graviditetsprevention och familjeplanering.
Könssjukdomar behandlas på hälsostationen och på polikliniken för könssjukdomar i Helsingfors. .
Hälsostationenfinska _ svenska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Polikliniken för könssjukdomarfinska _ svenska _ engelska
När du väntar barn
Vid mödrarådgivningen följs moderns, fostrets och hela familjens hälsotillstånd under graviditeten.
Kontakta rådgivningsbyrån när du upptäcker att du är gravid.
Tidsbokning vardagar kl. 12–13
Tfn (09) 8789 1344
Rådgivningsbyråerfinska _ svenska _ engelska
Det närmaste förlossningssjukhuset är Jorv sjukhus i Esbo.
Om du vill kan du även föda barnet på något annat sjukhus inom Helsingfors och Nylands sjukvårdsdistrikt (HNS).
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Val av förlossningssjukhusfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Läs mer: Förlossning
Handikappade personer
Grankulla stad erbjuder olika tjänster för handikappade, till exempel hjälpmedel och dagverksamhet.
Du kan fråga om tjänsterna för handikappade hos socialarbetaren för ditt område.
Tjänster inom handikappvårdenfinska _ svenska
Läs mer: Handikappade personer
Dagvård
Förskoleundervisning
Grundläggande utbildning
Yrkesutbildning
Gymnasium
Högskoleutbildning
Andra studiemöjligheter
Dagvård
I Grankulla finns stadens egna daghem, privata daghem och privata familjedagvårdare.
Dagvård fås på finska och på svenska.
I Grankulla finns också ett engelskspråkigt daghem.
Ansök om dagvårdsplats för ditt barn minst fyra månader innan barnet ska börja i dagvården.
Om du ansöker om dagvårdplats för första gången ska du använda den elektroniska ansökan.
Du kan också hämta ansökningsblanketten på daghemmet eller vid informationen i stadshuset.
Lämna in ansökan till daghemmet eller stadshuset.
Familjer som bor i Grankulla kan också söka dagvårdsplats till sitt barn i Esbo, Helsingfors eller Vanda.
Du ska ändå lämna in din ansökan i Grankulla.
Mer information finns på tjänsten HelsingforsRegionen.fi.
Läs mer: Dagvård
Dagvård och förskoleundervisningfinska _ svenska _ engelska
Ansökan om dagvårdsplatsfinska _ svenska
Engelsk-finskspråkigt daghemfinska _ engelska
Dagvårdens samanvändningsområdefinska _ svenska _ engelska
Förskoleundervisning
I Grankulla anordnas förskoleundervisningen i daghemmen.
Förskoleundervisningen börjar i augusti och ansökningstiden är i januari.
Läs mer: Förskoleundervisning
Information om förskoleundervisningenfinska _ svenska _ engelska
Grundläggande utbildning
I Grankulla finns både en finsk- och en svenskspråkig grundskola. Anmälan till grundskolan ska ske i början av året.
Om du har frågor om den grundläggande utbildningen kan du kontakta skolbyrån.
Skolbyrån
Grankulla stadshus
Grankullavägen 10
02700 Grankulla
Tfn (09) 50 561 (växel)
Grundläggande utbildning
Grundläggande utbildning och gymnasiumfinska _ svenska _ engelska
Internationella skolor i huvudstadsregionenfinska
linkkiExpatFinland.fi:
Internationella skolor i huvudstadsregionenengelska
Yrkesutbildning
De närmaste yrkesläroanstalterna finns i Esbo och Helsingfors.
Läs mer: Yrkesutbildning
Yrkesutbildningfinska _ engelska
Yrkesinriktad utbildningfinska
Gymnasium
I Grankulla finns två gymnasier, ett finskspråkigt och ett svenskspråkigt.
I Esbo finns ett vuxengymnasium där vuxna kan avlägga gymnasiet och studentexamen.
Läs mer: Gymnasium
Grundläggande utbildning och gymnasiumfinska _ svenska _ engelska
linkkiEsbo stad:
Vuxengymnasietfinska
Högskoleutbildning
I anslutning till folkhögskolan Työväen Akatemia i Grankulla finns en enhet för Humanistiska Yrkeshögskolan, där du kan avlägga yrkeshögskoleexamen för kulturproducenter.
Vid yrkeshögskolorna och universiteten i Esbo och Helsingfors kan du studera inom många områden.
Mer information om högskolorna i Esbo och Helsingfors hittar du på städernas webbplatser.
Läs mer: Högskoleutbildning
linkkiHumanistiska yrkeshögskolan:
Information om Humanistiska yrkeshögskolanfinska _ engelska
linkkiEsbo stad:
Högskolorfinska _ engelska
Högskolorfinska
Andra studiemöjligheter
Vid Grankulla medborgarinstitut kan du studera till exempel språk, handarbete och matlagning eller delta i ledd motion.
Medborgarinstitutetfinska _ svenska _ engelska
Vid Grankulla konstskola kan barn och unga studera bildkonst och vid Grankulla musikinstitut kan barn och vuxna studera musik.
Information om Konstskolanfinska _ svenska
Information om Musikinstitutetfinska _ svenska
I Grankulla ligger Finska Bibelinstitutet.
Vid institutet kan du avlägga enskilda kurser eller studera på någon av institutets studielinjer.
Studierna på studielinjerna pågår i 1–2 år.
Vid bibelinstitutet finns även en studielinje som är särskilt avsedd för invandrare.
Kristliga folkhögskolanfinska _ engelska
Folkhögskolan Työväen Akatemia tillhandahåller undervisning inom många akademiska discipliner samt träning för dem som vill läsa på universitet.
Information om Työväen Akatemiafinska _ engelska
Läs mer: Andra studiemöjligheter
Dagvård
Förskoleundervisning
Grundläggande utbildning
Yrkesutbildning
Gymnasium
Högskoleutbildning
Andra studiemöjligheter
Dagvård
I Grankulla finns stadens egna daghem, privata daghem och privata familjedagvårdare.
Dagvård fås på finska och på svenska.
I Grankulla finns också ett engelskspråkigt daghem.
Ansök om dagvårdsplats för ditt barn minst fyra månader innan barnet ska börja i dagvården.
Om du ansöker om dagvårdplats för första gången ska du använda den elektroniska ansökan.
Du kan också hämta ansökningsblanketten på daghemmet eller vid informationen i stadshuset.
Lämna in ansökan till daghemmet eller stadshuset.
Familjer som bor i Grankulla kan också söka dagvårdsplats till sitt barn i Esbo, Helsingfors eller Vanda.
Du ska ändå lämna in din ansökan i Grankulla.
Mer information finns på tjänsten HelsingforsRegionen.fi.
Läs mer: Dagvård
Dagvård och förskoleundervisningfinska _ svenska _ engelska
Ansökan om dagvårdsplatsfinska _ svenska
Engelsk-finskspråkigt daghemfinska _ engelska
Dagvårdens samanvändningsområdefinska _ svenska _ engelska
Förskoleundervisning
I Grankulla anordnas förskoleundervisningen i daghemmen.
Förskoleundervisningen börjar i augusti och ansökningstiden är i januari.
Läs mer: Förskoleundervisning
Information om förskoleundervisningenfinska _ svenska _ engelska
Grundläggande utbildning
I Grankulla finns både en finsk- och en svenskspråkig grundskola. Anmälan till grundskolan ska ske i början av året.
Om du har frågor om den grundläggande utbildningen kan du kontakta skolbyrån.
Skolbyrån
Grankulla stadshus
Grankullavägen 10
02700 Grankulla
Tfn (09) 50 561 (växel)
Grundläggande utbildning
Grundläggande utbildning och gymnasiumfinska _ svenska _ engelska
Internationella skolor i huvudstadsregionenfinska
linkkiExpatFinland.fi:
Internationella skolor i huvudstadsregionenengelska
Yrkesutbildning
De närmaste yrkesläroanstalterna finns i Esbo och Helsingfors.
Läs mer: Yrkesutbildning
Yrkesutbildningfinska _ engelska
Yrkesinriktad utbildningfinska
Gymnasium
I Grankulla finns två gymnasier, ett finskspråkigt och ett svenskspråkigt.
I Esbo finns ett vuxengymnasium där vuxna kan avlägga gymnasiet och studentexamen.
Läs mer: Gymnasium
Grundläggande utbildning och gymnasiumfinska _ svenska _ engelska
linkkiEsbo stad:
Vuxengymnasietfinska
Högskoleutbildning
I anslutning till folkhögskolan Työväen Akatemia i Grankulla finns en enhet för Humanistiska Yrkeshögskolan, där du kan avlägga yrkeshögskoleexamen för kulturproducenter.
Vid yrkeshögskolorna och universiteten i Esbo och Helsingfors kan du studera inom många områden.
Mer information om högskolorna i Esbo och Helsingfors hittar du på städernas webbplatser.
Läs mer: Högskoleutbildning
linkkiHumanistiska yrkeshögskolan:
Information om Humanistiska yrkeshögskolanfinska _ engelska
linkkiEsbo stad:
Högskolorfinska _ engelska
Högskolorfinska
Andra studiemöjligheter
Vid Grankulla medborgarinstitut kan du studera till exempel språk, handarbete och matlagning eller delta i ledd motion.
Medborgarinstitutetfinska _ svenska _ engelska
Vid Grankulla konstskola kan barn och unga studera bildkonst och vid Grankulla musikinstitut kan barn och vuxna studera musik.
Information om Konstskolanfinska _ svenska
Information om Musikinstitutetfinska _ svenska
I Grankulla ligger Finska Bibelinstitutet.
Vid institutet kan du avlägga enskilda kurser eller studera på någon av institutets studielinjer.
Studierna på studielinjerna pågår i 1–2 år.
Vid bibelinstitutet finns även en studielinje som är särskilt avsedd för invandrare.
Kristliga folkhögskolanfinska _ engelska
Folkhögskolan Työväen Akatemia tillhandahåller undervisning inom många akademiska discipliner samt träning för dem som vill läsa på universitet.
Information om Työväen Akatemiafinska _ engelska
Läs mer: Andra studiemöjligheter
Dagvård
Förskoleundervisning
Grundläggande utbildning
Yrkesutbildning
Gymnasium
Högskoleutbildning
Andra studiemöjligheter
Dagvård
I Grankulla finns stadens egna daghem, privata daghem och privata familjedagvårdare.
Dagvård fås på finska och på svenska.
I Grankulla finns också ett engelskspråkigt daghem.
Ansök om dagvårdsplats för ditt barn minst fyra månader innan barnet ska börja i dagvården.
Om du ansöker om dagvårdplats för första gången ska du använda den elektroniska ansökan.
Du kan också hämta ansökningsblanketten på daghemmet eller vid informationen i stadshuset.
Lämna in ansökan till daghemmet eller stadshuset.
Familjer som bor i Grankulla kan också söka dagvårdsplats till sitt barn i Esbo, Helsingfors eller Vanda.
Du ska ändå lämna in din ansökan i Grankulla.
Mer information finns på tjänsten HelsingforsRegionen.fi.
Läs mer: Dagvård
Dagvård och förskoleundervisningfinska _ svenska _ engelska
Ansökan om dagvårdsplatsfinska _ svenska
Engelsk-finskspråkigt daghemfinska _ engelska
Dagvårdens samanvändningsområdefinska _ svenska _ engelska
Förskoleundervisning
I Grankulla anordnas förskoleundervisningen i daghemmen.
Förskoleundervisningen börjar i augusti och ansökningstiden är i januari.
Läs mer: Förskoleundervisning
Information om förskoleundervisningenfinska _ svenska _ engelska
Grundläggande utbildning
I Grankulla finns både en finsk- och en svenskspråkig grundskola. Anmälan till grundskolan ska ske i början av året.
Om du har frågor om den grundläggande utbildningen kan du kontakta skolbyrån.
Skolbyrån
Grankulla stadshus
Grankullavägen 10
02700 Grankulla
Tfn (09) 50 561 (växel)
Grundläggande utbildning
Grundläggande utbildning och gymnasiumfinska _ svenska _ engelska
Internationella skolor i huvudstadsregionenfinska
linkkiExpatFinland.fi:
Internationella skolor i huvudstadsregionenengelska
Yrkesutbildning
De närmaste yrkesläroanstalterna finns i Esbo och Helsingfors.
Läs mer: Yrkesutbildning
Yrkesutbildningfinska _ engelska
Yrkesinriktad utbildningfinska
Gymnasium
I Grankulla finns två gymnasier, ett finskspråkigt och ett svenskspråkigt.
I Esbo finns ett vuxengymnasium där vuxna kan avlägga gymnasiet och studentexamen.
Läs mer: Gymnasium
Grundläggande utbildning och gymnasiumfinska _ svenska _ engelska
linkkiEsbo stad:
Vuxengymnasietfinska
Högskoleutbildning
I anslutning till folkhögskolan Työväen Akatemia i Grankulla finns en enhet för Humanistiska Yrkeshögskolan, där du kan avlägga yrkeshögskoleexamen för kulturproducenter.
Vid yrkeshögskolorna och universiteten i Esbo och Helsingfors kan du studera inom många områden.
Mer information om högskolorna i Esbo och Helsingfors hittar du på städernas webbplatser.
Läs mer: Högskoleutbildning
linkkiHumanistiska yrkeshögskolan:
Information om Humanistiska yrkeshögskolanfinska _ engelska
linkkiEsbo stad:
Högskolorfinska _ engelska
Högskolorfinska
Andra studiemöjligheter
Vid Grankulla medborgarinstitut kan du studera till exempel språk, handarbete och matlagning eller delta i ledd motion.
Medborgarinstitutetfinska _ svenska _ engelska
Vid Grankulla konstskola kan barn och unga studera bildkonst och vid Grankulla musikinstitut kan barn och vuxna studera musik.
Information om Konstskolanfinska _ svenska
Information om Musikinstitutetfinska _ svenska
I Grankulla ligger Finska Bibelinstitutet.
Vid institutet kan du avlägga enskilda kurser eller studera på någon av institutets studielinjer.
Studierna på studielinjerna pågår i 1–2 år.
Vid bibelinstitutet finns även en studielinje som är särskilt avsedd för invandrare.
Kristliga folkhögskolanfinska _ engelska
Folkhögskolan Työväen Akatemia tillhandahåller undervisning inom många akademiska discipliner samt träning för dem som vill läsa på universitet.
Information om Työväen Akatemiafinska _ engelska
Läs mer: Andra studiemöjligheter
Hyresbostad
Ägarbostad
Stöd- och serviceboende
Avfallshantering i bostaden
Hyresbostad
Hyresbostäderna är dyra i huvudstadsregionen.
Stadens hyresbostäder är förmånligare än bostäder som hyrs ut av företag och privatpersoner.
Privata hyresbostäder
Du hittar bostäder som hyrs ut av företag och privatpersoner via bostadssidor på internet.
Sökning av hyresbostäderfinska
Sökning av hyresbostäderfinska _ engelska
Stadens hyresbostäder
Om du vill söka en av stadens hyresbostäder ska du fylla i en ansökningsblankett för hyresbostäder.
Blanketten får du antingen vid informationen på Grankulla stadshus, på socialbyrån eller på Grankulla stads webbplats.
På stadens webbplats hittar du också anvisningar om hur du söker hyresbostad.
Skicka din ansökan till adressen:
PB 52
02701 Grankulla
Stadens hyresbostäderfinska _ svenska _ engelska
Om du är studerande kan du få en hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS.
linkkiHOAS:
Hyresbostäder för studerandefinska _ svenska _ engelska
Läs mer: Hyresbostad
Ägarbostad
På internet finns många annonser om bostäder som är till salu.
Bostäderna i Grankulla är tämligen dyra.
Information om köp av bostad hittar du på InfoFinlands sida Ägarbostad.
Om du blir bostadslös på grund av en kris eller en olycka, ska du kontakta socialbyrån.
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta ett skyddshem.
Steniusvägen 20
Du kan ringa skyddshemmet dygnet runt, telefonnumret är 09 4777 180.
Du behöver inte uppge ditt namn när du ringer.
Om du är ung och har problem hemma, kan du kontakta Finlands Röda Kors De ungas skyddshus.
Det närmaste skyddshuset finns i Esbo.
De ungas skyddshus
Tfn 09 819 55360
Hjälp till offer för familjevåldfinska
linkkiFörbundet för mödra- och skyddshem:
Information om skyddshem och mödrahemfinska
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Stöd- och serviceboende
Personer som har svårt att klara av de dagliga sysslorna utan hjälp, till exempel äldre eller personer med funktionsnedsättning, kan få ta del av hemvårdens stödtjänster.
En person som inte kan bo på egen hand kan bo på en anstalt.
På Grankulla socialbyrå kan du fråga mer om hemvårdens stödtjänster och boende på anstalt.
Grankulla socialbyrå
Köpcentret Grani
Grankullavägen 7 02700 Grankulla
Tfn 09 505 61
Läs mer: Stöd- och serviceboende
Information om hemvårdens stödtjänsterfinska _ svenska
Information om boende på anstaltfinska _ svenska
Avfallshantering och återvinning
På InfoFinlands sida Avfallshantering och återvinning hittar du information om sopsortering.
linkkiHelsingforsregionens miljötjänster:
Sopsorteringsanvisningarfinska _ svenska _ engelska
Avfallsinsamlingsstationerfinska
Hyresbostad
Ägarbostad
Stöd- och serviceboende
Avfallshantering i bostaden
Hyresbostad
Hyresbostäderna är dyra i huvudstadsregionen.
Stadens hyresbostäder är förmånligare än bostäder som hyrs ut av företag och privatpersoner.
Privata hyresbostäder
Du hittar bostäder som hyrs ut av företag och privatpersoner via bostadssidor på internet.
Sökning av hyresbostäderfinska
Sökning av hyresbostäderfinska _ engelska
Stadens hyresbostäder
Om du vill söka en av stadens hyresbostäder ska du fylla i en ansökningsblankett för hyresbostäder.
Blanketten får du antingen vid informationen på Grankulla stadshus, på socialbyrån eller på Grankulla stads webbplats.
På stadens webbplats hittar du också anvisningar om hur du söker hyresbostad.
Skicka din ansökan till adressen:
PB 52
02701 Grankulla
Stadens hyresbostäderfinska _ svenska _ engelska
Om du är studerande kan du få en hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS.
linkkiHOAS:
Hyresbostäder för studerandefinska _ svenska _ engelska
Läs mer: Hyresbostad
Ägarbostad
På internet finns många annonser om bostäder som är till salu.
Bostäderna i Grankulla är tämligen dyra.
Information om köp av bostad hittar du på InfoFinlands sida Ägarbostad.
Om du blir bostadslös på grund av en kris eller en olycka, ska du kontakta socialbyrån.
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta ett skyddshem.
Steniusvägen 20
Du kan ringa skyddshemmet dygnet runt, telefonnumret är 09 4777 180.
Du behöver inte uppge ditt namn när du ringer.
Om du är ung och har problem hemma, kan du kontakta Finlands Röda Kors De ungas skyddshus.
Det närmaste skyddshuset finns i Esbo.
De ungas skyddshus
Tfn 09 819 55360
Hjälp till offer för familjevåldfinska
linkkiFörbundet för mödra- och skyddshem:
Information om skyddshem och mödrahemfinska
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Stöd- och serviceboende
Personer som har svårt att klara av de dagliga sysslorna utan hjälp, till exempel äldre eller personer med funktionsnedsättning, kan få ta del av hemvårdens stödtjänster.
En person som inte kan bo på egen hand kan bo på en anstalt.
På Grankulla socialbyrå kan du fråga mer om hemvårdens stödtjänster och boende på anstalt.
Grankulla socialbyrå
Köpcentret Grani
Grankullavägen 7 02700 Grankulla
Tfn 09 505 61
Läs mer: Stöd- och serviceboende
Information om hemvårdens stödtjänsterfinska _ svenska
Information om boende på anstaltfinska _ svenska
Avfallshantering och återvinning
På InfoFinlands sida Avfallshantering och återvinning hittar du information om sopsortering.
linkkiHelsingforsregionens miljötjänster:
Sopsorteringsanvisningarfinska _ svenska _ engelska
Avfallsinsamlingsstationerfinska
Hyresbostad
Ägarbostad
Stöd- och serviceboende
Avfallshantering i bostaden
Hyresbostad
Hyresbostäderna är dyra i huvudstadsregionen.
Stadens hyresbostäder är förmånligare än bostäder som hyrs ut av företag och privatpersoner.
Privata hyresbostäder
Du hittar bostäder som hyrs ut av företag och privatpersoner via bostadssidor på internet.
Sökning av hyresbostäderfinska
Sökning av hyresbostäderfinska _ engelska
Stadens hyresbostäder
Om du vill söka en av stadens hyresbostäder ska du fylla i en ansökningsblankett för hyresbostäder.
Blanketten får du antingen vid informationen på Grankulla stadshus, på socialbyrån eller på Grankulla stads webbplats.
På stadens webbplats hittar du också anvisningar om hur du söker hyresbostad.
Skicka din ansökan till adressen:
PB 52
02701 Grankulla
Stadens hyresbostäderfinska _ svenska _ engelska
Om du är studerande kan du få en hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS.
linkkiHOAS:
Hyresbostäder för studerandefinska _ svenska _ engelska
Läs mer: Hyresbostad
Ägarbostad
På internet finns många annonser om bostäder som är till salu.
Bostäderna i Grankulla är tämligen dyra.
Information om köp av bostad hittar du på InfoFinlands sida Ägarbostad.
Om du blir bostadslös på grund av en kris eller en olycka, ska du kontakta socialbyrån.
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta ett skyddshem.
Steniusvägen 20
Du kan ringa skyddshemmet dygnet runt, telefonnumret är 09 4777 180.
Du behöver inte uppge ditt namn när du ringer.
Om du är ung och har problem hemma, kan du kontakta Finlands Röda Kors De ungas skyddshus.
Det närmaste skyddshuset finns i Esbo.
De ungas skyddshus
Tfn 09 819 55360
Hjälp till offer för familjevåldfinska
linkkiFörbundet för mödra- och skyddshem:
Information om skyddshem och mödrahemfinska
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Stöd- och serviceboende
Personer som har svårt att klara av de dagliga sysslorna utan hjälp, till exempel äldre eller personer med funktionsnedsättning, kan få ta del av hemvårdens stödtjänster.
En person som inte kan bo på egen hand kan bo på en anstalt.
På Grankulla socialbyrå kan du fråga mer om hemvårdens stödtjänster och boende på anstalt.
Grankulla socialbyrå
Köpcentret Grani
Grankullavägen 7 02700 Grankulla
Tfn 09 505 61
Läs mer: Stöd- och serviceboende
Information om hemvårdens stödtjänsterfinska _ svenska
Information om boende på anstaltfinska _ svenska
Avfallshantering och återvinning
På InfoFinlands sida Avfallshantering och återvinning hittar du information om sopsortering.
linkkiHelsingforsregionens miljötjänster:
Sopsorteringsanvisningarfinska _ svenska _ engelska
Avfallsinsamlingsstationerfinska
Språkkurser
Med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors, Vanda, Esbo eller Grankulla.
I tjänsten finns också information om kurser i svenska.
Kurser i finska och svenska språketfinska _ engelska _ ryska
I Grankulla ordnas kurser i finska och svenska av Grankulla medborgarinstitut.
Du kan anmäla dig till medborgarinstitutets kurser per telefon eller via internet.
Medborgarinstitutetfinska _ svenska _ engelska
Läs mer: Studier i finska och svenska
Svenska språket i Finland.
Diskutera på finska
Information om bibliotekens språkkaféer och andra finska samtalsgrupper hittar du på InfoFinlands sidor Finska och svenska språket i Esbo och Finska och svenska språket i Helsingfors.
Allmän språkexamen
Du kan avlägga allmän språkexamen i finska eller svenska till exempel i Esbo och Helsingfors.
På Utbildningsstyrelsens webbplats finns en sökmotor med vilken du kan kontrollera var och när du kan avlägga examen.
Läs mer: Officiellt intyg på språkkunskaper.
linkkiUtbildningsstyrelsen:
Allmänna språkexaminafinska _ svenska _ engelska
Språkkurser
Med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors, Vanda, Esbo eller Grankulla.
I tjänsten finns också information om kurser i svenska.
Kurser i finska och svenska språketfinska _ engelska _ ryska
I Grankulla ordnas kurser i finska och svenska av Grankulla medborgarinstitut.
Du kan anmäla dig till medborgarinstitutets kurser per telefon eller via internet.
Medborgarinstitutetfinska _ svenska _ engelska
Läs mer: Studier i finska och svenska
Svenska språket i Finland.
Diskutera på finska
Information om bibliotekens språkkaféer och andra finska samtalsgrupper hittar du på InfoFinlands sidor Finska och svenska språket i Esbo och Finska och svenska språket i Helsingfors.
Allmän språkexamen
Du kan avlägga allmän språkexamen i finska eller svenska till exempel i Esbo och Helsingfors.
På Utbildningsstyrelsens webbplats finns en sökmotor med vilken du kan kontrollera var och när du kan avlägga examen.
Läs mer: Officiellt intyg på språkkunskaper.
linkkiUtbildningsstyrelsen:
Allmänna språkexaminafinska _ svenska _ engelska
Språkkurser
Med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors, Vanda, Esbo eller Grankulla.
I tjänsten finns också information om kurser i svenska.
Kurser i finska och svenska språketfinska _ engelska _ ryska
I Grankulla ordnas kurser i finska och svenska av Grankulla medborgarinstitut.
Du kan anmäla dig till medborgarinstitutets kurser per telefon eller via internet.
Medborgarinstitutetfinska _ svenska _ engelska
Läs mer: Studier i finska och svenska
Svenska språket i Finland.
Diskutera på finska
Information om bibliotekens språkkaféer och andra finska samtalsgrupper hittar du på InfoFinlands sidor Finska och svenska språket i Esbo och Finska och svenska språket i Helsingfors.
Allmän språkexamen
Du kan avlägga allmän språkexamen i finska eller svenska till exempel i Esbo och Helsingfors.
På Utbildningsstyrelsens webbplats finns en sökmotor med vilken du kan kontrollera var och när du kan avlägga examen.
Läs mer: Officiellt intyg på språkkunskaper.
linkkiUtbildningsstyrelsen:
Allmänna språkexaminafinska _ svenska _ engelska
Var hittar jag jobb?
Att grunda ett företag
Beskattning
Var hittar jag jobb?
Nylands arbets- och näringsbyrå hjälper invånare i Grankulla att söka jobb.
Den närmaste byrån finns i Esbo.
Nylands arbets- och näringsbyrå, Esbo
Läs mer: Arbete och entreprenörskap i Esbo
Information om arbets- och näringsbyråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös.
Information om jobbsökning i Finland hittar du på InfoFinlands sida Var hittar jag jobb?
Seure erbjuder kortvariga jobb vid Helsingfors, Vanda, Esbo och Grankulla städer.
Jobben finns till exempel på skolor, daghem och sjukhus.
Arbetsplatser i kommunernafinska _ svenska
Lediga jobbfinska _ svenska _ engelska
Arbetslöshetsersättning
Information om att ansöka om arbetslöshetsersättning hittar du på InfoFinlands sida Arbetslöshetsförsäkring.
Att grunda ett företag
På InfoFinlands sida Att grunda ett företag hittar du information om hur man grundar ett företag i Finland.
Bekanta dig med de lokala tjänsterna på sidorna Arbete och entreprenörskap i Esbo och Arbete och entreprenörskap i Helsingfors.
Om du är företagare kan du bli medlem i företagarnas intressebevakningsorganisation Grankulla företagare rf som erbjuder sina medlemmar utbildning, nätverk och rådgivning.
Information för företagarefinska
Beskattning
Huvudstadsregionens skattebyrå ligger på Alexandersgatan 9 i Gloet i Helsingfors.
linkkiSkatteförvaltningen:
Kontaktuppgifter till skattebyråerfinska _ svenska _ engelska
Du kan även besöka servicestället In To Finland i Kampen i Helsingfors för att fråga om beskattningen.
Servicestället betjänar invandrare som kommer till Finland för att arbeta i ärenden som berör beskattning och social trygghet.
Albertsgatan 25
Lär mer Beskattning
Var hittar jag jobb?
Att grunda ett företag
Beskattning
Var hittar jag jobb?
Nylands arbets- och näringsbyrå hjälper invånare i Grankulla att söka jobb.
Den närmaste byrån finns i Esbo.
Nylands arbets- och näringsbyrå, Esbo
Läs mer: Arbete och entreprenörskap i Esbo
Information om arbets- och näringsbyråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös.
Information om jobbsökning i Finland hittar du på InfoFinlands sida Var hittar jag jobb?
Seure erbjuder kortvariga jobb vid Helsingfors, Vanda, Esbo och Grankulla städer.
Jobben finns till exempel på skolor, daghem och sjukhus.
Arbetsplatser i kommunernafinska _ svenska
Lediga jobbfinska _ svenska _ engelska
Arbetslöshetsersättning
Information om att ansöka om arbetslöshetsersättning hittar du på InfoFinlands sida Arbetslöshetsförsäkring.
Att grunda ett företag
På InfoFinlands sida Att grunda ett företag hittar du information om hur man grundar ett företag i Finland.
Bekanta dig med de lokala tjänsterna på sidorna Arbete och entreprenörskap i Esbo och Arbete och entreprenörskap i Helsingfors.
Om du är företagare kan du bli medlem i företagarnas intressebevakningsorganisation Grankulla företagare rf som erbjuder sina medlemmar utbildning, nätverk och rådgivning.
Information för företagarefinska
Beskattning
Huvudstadsregionens skattebyrå ligger på Alexandersgatan 9 i Gloet i Helsingfors.
linkkiSkatteförvaltningen:
Kontaktuppgifter till skattebyråerfinska _ svenska _ engelska
Invandrare kan även sköta ärenden vid servicestället International House Helsinki.
På servicestället hjälper FPA:s och Skatteförvaltningens experter invandrare som kommer till Finland för att arbeta i frågor som rör beskattning och social trygghet.
Lär mer Beskattning
Var hittar jag jobb?
Att grunda ett företag
Beskattning
Var hittar jag jobb?
Nylands arbets- och näringsbyrå hjälper invånare i Grankulla att söka jobb.
Den närmaste byrån finns i Esbo.
Nylands arbets- och näringsbyrå, Esbo
Läs mer: Arbete och entreprenörskap i Esbo
Information om arbets- och näringsbyråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös.
Information om jobbsökning i Finland hittar du på InfoFinlands sida Var hittar jag jobb?
Seure erbjuder kortvariga jobb vid Helsingfors, Vanda, Esbo och Grankulla städer.
Jobben finns till exempel på skolor, daghem och sjukhus.
Arbetsplatser i kommunernafinska _ svenska _ engelska
Lediga jobbfinska _ svenska _ engelska
Arbetslöshetsersättning
Information om att ansöka om arbetslöshetsersättning hittar du på InfoFinlands sida Arbetslöshetsförsäkring.
Att grunda ett företag
På InfoFinlands sida Att grunda ett företag hittar du information om hur man grundar ett företag i Finland.
Bekanta dig med de lokala tjänsterna på sidorna Arbete och entreprenörskap i Esbo och Arbete och entreprenörskap i Helsingfors.
Om du är företagare kan du bli medlem i företagarnas intressebevakningsorganisation Grankulla företagare rf som erbjuder sina medlemmar utbildning, nätverk och rådgivning.
Information för företagarefinska
Beskattning
Huvudstadsregionens skattebyrå ligger på Alexandersgatan 9 i Gloet i Helsingfors.
linkkiSkatteförvaltningen:
Kontaktuppgifter till skattebyråerfinska _ svenska _ engelska
Invandrare kan även sköta ärenden vid servicestället International House Helsinki.
På servicestället hjälper FPA:s och Skatteförvaltningens experter invandrare som kommer till Finland för att arbeta i frågor som rör beskattning och social trygghet.
IHH – serviceställe för dig som flyttar till Finland engelska
Lär mer Beskattning
Rådgivning för och integration av invandrare
Inledande kartläggning och integrationsplan
Behöver du en tolk?
Rådgivning för och integration av invandrare
Om du har frågor om tjänsterna vid Grankulla stad kan du kontakta stadens rådgivningstjänst via e-post på adressen neuvontapalvelu(at)kauniainen.fi.
Du kan skriva på finska, svenska eller engelska.
Helsingfors stads rådgivning för invandrare, Helsingfors-info, betjänar alla invandrare i huvudstadsregionen.
Helsingfors-infofinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
IHH – serviceställe för dig som flyttar till Finland engelska
Inledande kartläggning och integrationsplan
Tillsammans med en anställd vid arbets- och näringsbyrån (TE-byrån) gör du en inledande kartläggning och en integrationsplan i samband med att du registrerar dig som arbetssökande.
linkkiArbets- och näringsministeriet:
Arbets- och näringsbyråerna i Nylandfinska _ svenska
Om du inte är kund hos arbets- och näringsbyrån görs den inledande kartläggningen och integrationsplanen på socialbyrån.
Kontaktuppgifter till socialbyrån:
Köpcentret Grani
Grankullavägen 7
02700 Grankulla
Tfn (09) 50 561
Socialbyrånfinska _ svenska
Behöver du en tolk?
Om du inte kan finska eller svenska kan du anlita en tolk när du sköter ärenden med myndigheter.
Du kan anlita en tolk när som helst om du bokar tolken och betalar kostnaderna själv.
I vissa fall får du en tolk via myndigheten.
Då är tolkningen avgiftsfri för dig.
Läs mer: Behöver du en tolk?
linkkiFinlands översättar- och tolkförbund:
Sök tolk eller översättarefinska _ svenska _ engelska
Rådgivning för och integration av invandrare
Inledande kartläggning och integrationsplan
Behöver du en tolk?
Rådgivning för och integration av invandrare
Om du har frågor om tjänsterna vid Grankulla stad kan du kontakta stadens rådgivningstjänst via e-post på adressen neuvontapalvelu(at)kauniainen.fi.
Du kan skriva på finska, svenska eller engelska.
Helsingfors stads rådgivning för invandrare, Helsingfors-info, betjänar alla invandrare i huvudstadsregionen.
Helsingfors-infofinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
IHH – serviceställe för dig som flyttar till Finland engelska
Inledande kartläggning och integrationsplan
Tillsammans med en anställd vid arbets- och näringsbyrån (TE-byrån) gör du en inledande kartläggning och en integrationsplan i samband med att du registrerar dig som arbetssökande.
linkkiArbets- och näringsministeriet:
Arbets- och näringsbyråerna i Nylandfinska _ svenska
Om du inte är kund hos arbets- och näringsbyrån görs den inledande kartläggningen och integrationsplanen på socialbyrån.
Kontaktuppgifter till socialbyrån:
Köpcentret Grani
Grankullavägen 7
02700 Grankulla
Tfn (09) 50 561
Socialbyrånfinska _ svenska
Behöver du en tolk?
Om du inte kan finska eller svenska kan du anlita en tolk när du sköter ärenden med myndigheter.
Du kan anlita en tolk när som helst om du bokar tolken och betalar kostnaderna själv.
I vissa fall får du en tolk via myndigheten.
Då är tolkningen avgiftsfri för dig.
Läs mer: Behöver du en tolk?
linkkiFinlands översättar- och tolkförbund:
Sök tolk eller översättarefinska _ svenska _ engelska
Rådgivning för och integration av invandrare
Inledande kartläggning och integrationsplan
Behöver du en tolk?
Rådgivning för och integration av invandrare
Om du har frågor om tjänsterna vid Grankulla stad kan du kontakta stadens rådgivningstjänst via e-post på adressen neuvontapalvelu(at)kauniainen.fi.
Du kan skriva på finska, svenska eller engelska.
Helsingfors stads rådgivning för invandrare, Helsingfors-info, betjänar alla invandrare i huvudstadsregionen.
Helsingfors-infofinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
IHH – serviceställe för dig som flyttar till Finland engelska
Inledande kartläggning och integrationsplan
Tillsammans med en anställd vid arbets- och näringsbyrån (TE-byrån) gör du en inledande kartläggning och en integrationsplan i samband med att du registrerar dig som arbetssökande.
linkkiArbets- och näringsministeriet:
Arbets- och näringsbyråerna i Nylandfinska _ svenska
Om du inte är kund hos arbets- och näringsbyrån görs den inledande kartläggningen och integrationsplanen på socialbyrån.
Kontaktuppgifter till socialbyrån:
Köpcentret Grani
Grankullavägen 7
02700 Grankulla
Tfn (09) 50 561
Socialbyrånfinska _ svenska
Behöver du en tolk?
Om du inte kan finska eller svenska kan du anlita en tolk när du sköter ärenden med myndigheter.
Du kan anlita en tolk när som helst om du bokar tolken och betalar kostnaderna själv.
I vissa fall får du en tolk via myndigheten.
Då är tolkningen avgiftsfri för dig.
Läs mer: Behöver du en tolk?
linkkiFinlands översättar- och tolkförbund:
Sök tolk eller översättarefinska _ svenska _ engelska
Tillståndsärenden
På Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU-medborgarens uppehållsrätt.
Boka en tid i förväg.
Adress:
Göksgränd 3A
Elektronisk tidsbokningfinska _ svenska _ engelska
Du kan också ansöka om många slags uppehållstillstånd och EU-registrering på internet i tjänsten Enter Finland.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Läs mer: Flytta till Finland.
Registrering som invånare
Om du flyttar ditt stadigvarande boende till Grankulla, ska du registrera dig som invånare i kommunen.
Du kan registrera dig vid Helsingfors enhet vid magistraten i Nyland.
Helsingfors enhet
Albertsgatan 25
Tfn 029 55 39391
När du går till magistraten ska du ta med dig
legitimation (till exempel pass)
uppehållstillstånd och uppehållskort (om du behöver uppehållstillstånd i Finland)
registreringsintyget över uppehållsrätten (om du är EU-medborgare)
äktenskapsintyg
dina barns födelseattester.
Observera att utländska handlingar ska vara legaliserade samt översatta till finska eller svenska.
Läs mer: Registrering som invånare
Hemkommun i Finland
Registrering av utlänningarfinska _ svenska _ engelska
IHH – serviceställe för dig som flyttar till Finland engelska
Tillståndsärenden
På Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU-medborgarens uppehållsrätt.
Boka en tid i förväg.
Adress:
Göksgränd 3A
Elektronisk tidsbokningfinska _ svenska _ engelska
Du kan också ansöka om många slags uppehållstillstånd och EU-registrering på internet i tjänsten Enter Finland.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Läs mer: Flytta till Finland.
Registrering som invånare
Om du flyttar ditt stadigvarande boende till Grankulla, ska du registrera dig som invånare i kommunen.
Du kan registrera dig vid Helsingfors enhet vid magistraten i Nyland.
Helsingfors enhet
Tfn 029 55 39391
När du går till magistraten ska du ta med dig
legitimation (till exempel pass)
uppehållstillstånd och uppehållskort (om du behöver uppehållstillstånd i Finland)
registreringsintyget över uppehållsrätten (om du är EU-medborgare)
äktenskapsintyg
dina barns födelseattester.
Observera att utländska handlingar ska vara legaliserade samt översatta till finska eller svenska.
Läs mer: Registrering som invånare
Hemkommun i Finland
Registrering av utlänningarfinska _ svenska _ engelska
IHH – serviceställe för dig som flyttar till Finland engelska
Tillståndsärenden
På Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU-medborgarens uppehållsrätt.
Boka en tid i förväg.
Adress:
Göksgränd 3A
Elektronisk tidsbokningfinska _ svenska _ engelska
Du kan också ansöka om många slags uppehållstillstånd och EU-registrering på internet i tjänsten Enter Finland.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Läs mer: Flytta till Finland.
Registrering som invånare
Om du flyttar ditt stadigvarande boende till Grankulla, ska du registrera dig som invånare i kommunen.
Du kan registrera dig vid Helsingfors enhet vid magistraten i Nyland.
Helsingfors enhet
Tfn 029 55 39391
När du går till magistraten ska du ta med dig
legitimation (till exempel pass)
uppehållstillstånd och uppehållskort (om du behöver uppehållstillstånd i Finland)
registreringsintyget över uppehållsrätten (om du är EU-medborgare)
äktenskapsintyg
dina barns födelseattester.
Observera att utländska handlingar ska vara legaliserade samt översatta till finska eller svenska.
Läs mer: Registrering som invånare
Hemkommun i Finland
Registrering av utlänningarfinska _ svenska _ engelska
IHH – serviceställe för dig som flyttar till Finland engelska
Trafik
Beslutsfattande och påverkan
Religion
Grundläggande information
Historia
Trafik
Kollektivtrafiken
Vanda och hela huvudstadsregionen har goda kollektivtrafikförbindelser.
Längs stambanan och Mårtensdals bana finns flera tågstationer.
I staden finns flera busslinjer.
Vanda tillhör samkommunen Helsingforsregionens trafik (HRT) (Helsingin seudun liikenne -kuntayhtymä (HSL)), som ordnar kollektivtrafiken i huvudstadsregionen.
Mer information hittar du på HRT:s webbplats.
Du kan söka information om rutterna i Reseplaneraren (Reittiopas).
Tjänsten ger dig förslag på olika kollektivtrafikförbindelser från ett ställe till ett annat.
I kollektivtrafiken kan du betala med kontanter eller resekort.
I närtågen måste du köpa biljetten i förväg.
Du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat.
Reseplanerarefinska _ svenska _ engelska _ ryska
Resekort
Med ett resekort (matkakortti) reser du förmånligare än med kontanter.
Resekortet gäller i lokaltrafikens bussar, närtågen, metron, spårvagnarna och Sveaborgsfärjorna.
Det finns två slags resekort.
Det är det billigaste sättet att resa.
Ett innehavarkort (haltijakohtainen kortti) kan användas av flera personer.
Innan du skaffar dig ett personligt kort ska du registrera dig som invånare i någon av kommunerna inom HRT-området.
Du kan köpa resekort vid HRT:s försäljningsställen (myyntipiste) eller serviceställen (palvelupiste).
De finns runtom i huvudstadsregionen.
Personligt resekort kan du köpa vid serviceställena.
Ta med dig identitetsbevis om du ska köpa personligt resekort.
Om du har finska nätbankskoder kan du även köpa personligt resekort på HRT:s webbplats.
Du kan resa med resekortet när du laddar kortet med period (kausi) eller värde (arvo).
En period betyder tid: till exempel en månad.
Värde betyder pengar.
Om du använder kollektivtrafiken ofta tjänar du på att ladda kortet med period.
Du kan ladda resekortet på vilket serviceställe för resekort (matkakortin latauspiste) som helst.
Du hittar mer information på HRT:s webbplats.
Ansökan om försäljningsplatserfinska _ svenska _ engelska
Information och råd till resenärerfinska _ svenska _ engelska
Biljetter och priserfinska _ svenska _ engelska
Att gå och cykla
Om du vill gå eller cykla i Vanda kan du söka en lämplig rutt i reseplaneraren för cykling och gång.
En cykelkarta i pappersformat för Vanda kan du hämta i Vandainfo.
Cykelkartorna är kostnadsfria.
linkkiVanda stad:
Vandainfofinska _ svenska _ engelska
Bil och flyg
Helsingfors-Vanda internationella flygplats ligger i Vanda.
Flygplatsen har goda trafikförbindelser till exempel med bil, buss och tåg.
Du kan parkera bilen på många järnvägsstationer och fortsätta färden med kollektivtrafiken.
Tidtabellerna för bussar och tåg hittar du enkelt i reseplaneraren.
Läs mer: Trafik.
Flygplatsenfinska _ svenska _ engelska _ ryska _ kinesiska
Beslutsfattande och påverkan
I Vanda beslutas ärenden av stadsfullmäktige (kaupunginvaltuusto).
I stadsfullmäktige sitter 67 ledamöter som representerar olika politiska grupper.
Fullmäktige väljs var fjärde år genom kommunalval (kunnallisvaalit).
Invånarna i Vanda kan påverka beslutsfattandet och beredning av ärenden på många olika sätt.
På Vandakanalen kan du följa fullmäktiges sammanträden och få mer information om beslutsfattandet.
I Vanda finns en delegation för mångkulturella frågor (monikulttuurisuusasiain neuvottelukunta) som lägger fram propositioner i ärenden som rör invandrare.
Läs mer på Vanda stads webbplats.
I Vanda finns många politiska föreningar, invandrarföreningar och andra föreningar via vilka du också kan påverka beslutsfattandet.
Mer information om föreningarna hittar du på sidan Vantaalla.info.
linkkiVanda stad:
Beslutsfattandefinska _ svenska _ engelska
linkkiVanda stad:
Delta och påverkafinska
Stadsfullmäktiges sammanträden på Internetfinska
linkkiVanda stad:
Delegationen för mångkulturella frågorfinska
Religion
Många religiösa samfund är verksamma i Vanda och Helsingfors.
Via tjänsten Uskonnot Suomessa kan du söka information efter det religiösa samfundet och orten.
Den evangelisk-lutherska kyrkan har sex finskspråkiga församlingar och en svenskspråkig församling i Vanda.
Läs mer på Vanda kyrkliga samfällighets webbplats.
I Dickursby finns en ortodox kyrka.
Mer information om verksamheten vid den ortodoxa kyrkan i Vanda hittar du på Helsingfors ortodoxa församlings webbplats.
Läs mer: Kulturer och religioner i Finland.
linkkiVanda kyrkliga samfällighet:
Evangelisk-lutherska församlingarfinska
linkkiHelsingfors ortodoxa församling:
Ortodoxa församlingenfinska _ ryska
Religiösa samfundfinska _ engelska
Grundläggande information
Vanda är en av de fyra kommunerna i huvudstadsregionen.
Den ligger intill Esbo och Helsingfors.
Vanda centrum ligger i Dickursby.
Därtill finns det andra stora tätorter i Vanda, till exempel Korso, Björkby-Havukoski, Myrbacka, Mårtensdal, Håkansböle, Västerkulla och Backas.
Vanda har drygt 205 000 invånare.
Av dem är cirka 2,8 procent svenskspråkiga och 11 procent har något annat modersmål än finska eller svenska.
Arealen är cirka 240 km2, varav cirka 2 km2 består av vatten.
linkkiVanda stad:
Grundläggande informationfinska _ svenska _ engelska
Historia
Vanda område har varit bebott länge.
Man har hittat upp till 7 000 år gamla lämningar efter bosättning.
Nuvarande Vanda har uppstått på ett område som förr var Helsingfors socken.
Helsingfors sockens historia sträcker sig ända till 1300-talet.
Helsingfors socken blev först Helsingfors landskommun, sedan Vanda köping år 1972 och till slut Vanda stad år 1974.
Läget som granne till huvudstaden Helsingfors har varit viktigt för Vanda.
Viktiga vägar, såsom vägen från Åbo via Helsingfors till Viborg och senare järnvägen norrut från Helsingfors, har gått genom Vanda.
Längs med vägarna och järnvägen har det utvecklats industrier och bostadsområden.
Vanda är än idag en viktig trafikknutpunkt.
Till exempel ligger Helsingfors-Vanda flygplats i Vanda.
linkkiVanda stad:
Information om Vandafinska
linkkiVanda stad:
Stadsmuseetfinska _ svenska _ engelska
Trafik
Beslutsfattande och påverkan
Religion
Grundläggande information
Historia
Trafik
Kollektivtrafiken
Vanda och hela huvudstadsregionen har goda kollektivtrafikförbindelser.
Längs stambanan och Mårtensdals bana finns flera tågstationer.
I staden finns flera busslinjer.
Vanda tillhör samkommunen Helsingforsregionens trafik (HRT) (Helsingin seudun liikenne -kuntayhtymä (HSL)), som ordnar kollektivtrafiken i huvudstadsregionen.
Mer information hittar du på HRT:s webbplats.
Du kan söka information om rutterna i Reseplaneraren (Reittiopas).
Tjänsten ger dig förslag på olika kollektivtrafikförbindelser från ett ställe till ett annat.
I kollektivtrafiken kan du betala med kontanter eller resekort.
I närtågen måste du köpa biljetten i förväg.
Du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat.
Reseplanerarefinska _ svenska _ engelska _ ryska
Resekort
Med ett resekort (matkakortti) reser du förmånligare än med kontanter.
Resekortet gäller i lokaltrafikens bussar, närtågen, metron, spårvagnarna och Sveaborgsfärjorna.
Det finns två slags resekort.
Det är det billigaste sättet att resa.
Ett innehavarkort (haltijakohtainen kortti) kan användas av flera personer.
Innan du skaffar dig ett personligt kort ska du registrera dig som invånare i någon av kommunerna inom HRT-området.
Du kan köpa resekort vid HRT:s försäljningsställen (myyntipiste) eller serviceställen (palvelupiste).
De finns runtom i huvudstadsregionen.
Personligt resekort kan du köpa vid serviceställena.
Ta med dig identitetsbevis om du ska köpa personligt resekort.
Om du har finska nätbankskoder kan du även köpa personligt resekort på HRT:s webbplats.
Du kan resa med resekortet när du laddar kortet med period (kausi) eller värde (arvo).
En period betyder tid: till exempel en månad.
Värde betyder pengar.
Om du använder kollektivtrafiken ofta tjänar du på att ladda kortet med period.
Du kan ladda resekortet på vilket serviceställe för resekort (matkakortin latauspiste) som helst.
Du hittar mer information på HRT:s webbplats.
Ansökan om försäljningsplatserfinska _ svenska _ engelska
Information och råd till resenärerfinska _ svenska _ engelska
Biljetter och priserfinska _ svenska _ engelska
Att gå och cykla
Om du vill gå eller cykla i Vanda kan du söka en lämplig rutt i reseplaneraren för cykling och gång.
En cykelkarta i pappersformat för Vanda kan du hämta i Vandainfo.
Cykelkartorna är kostnadsfria.
linkkiVanda stad:
Vandainfofinska _ svenska _ engelska
Bil och flyg
Helsingfors-Vanda internationella flygplats ligger i Vanda.
Flygplatsen har goda trafikförbindelser till exempel med bil, buss och tåg.
Du kan parkera bilen på många järnvägsstationer och fortsätta färden med kollektivtrafiken.
Tidtabellerna för bussar och tåg hittar du enkelt i reseplaneraren.
Läs mer: Trafik.
Flygplatsenfinska _ svenska _ engelska _ ryska _ kinesiska
Beslutsfattande och påverkan
I Vanda beslutas ärenden av stadsfullmäktige (kaupunginvaltuusto).
I stadsfullmäktige sitter 67 ledamöter som representerar olika politiska grupper.
Fullmäktige väljs var fjärde år genom kommunalval (kunnallisvaalit).
Invånarna i Vanda kan påverka beslutsfattandet och beredning av ärenden på många olika sätt.
På Vandakanalen kan du följa fullmäktiges sammanträden och få mer information om beslutsfattandet.
I Vanda finns en delegation för mångkulturella frågor (monikulttuurisuusasiain neuvottelukunta) som lägger fram propositioner i ärenden som rör invandrare.
Läs mer på Vanda stads webbplats.
I Vanda finns många politiska föreningar, invandrarföreningar och andra föreningar via vilka du också kan påverka beslutsfattandet.
Mer information om föreningarna hittar du på sidan Vantaalla.info.
linkkiVanda stad:
Beslutsfattandefinska _ svenska _ engelska
linkkiVanda stad:
Delta och påverkafinska
Stadsfullmäktiges sammanträden på Internetfinska
linkkiVanda stad:
Delegationen för mångkulturella frågorfinska
Religion
Många religiösa samfund är verksamma i Vanda och Helsingfors.
Via tjänsten Uskonnot Suomessa kan du söka information efter det religiösa samfundet och orten.
Den evangelisk-lutherska kyrkan har sex finskspråkiga församlingar och en svenskspråkig församling i Vanda.
Läs mer på Vanda kyrkliga samfällighets webbplats.
I Dickursby finns en ortodox kyrka.
Mer information om verksamheten vid den ortodoxa kyrkan i Vanda hittar du på Helsingfors ortodoxa församlings webbplats.
Läs mer: Kulturer och religioner i Finland.
linkkiVanda kyrkliga samfällighet:
Evangelisk-lutherska församlingarfinska
linkkiHelsingfors ortodoxa församling:
Ortodoxa församlingenfinska _ ryska
Religiösa samfundfinska _ engelska
Grundläggande information
Vanda är en av de fyra kommunerna i huvudstadsregionen.
Den ligger intill Esbo och Helsingfors.
Vanda centrum ligger i Dickursby.
Därtill finns det andra stora tätorter i Vanda, till exempel Korso, Björkby-Havukoski, Myrbacka, Mårtensdal, Håkansböle, Västerkulla och Backas.
Vanda har drygt 205 000 invånare.
Av dem är cirka 2,8 procent svenskspråkiga och 11 procent har något annat modersmål än finska eller svenska.
Arealen är cirka 240 km2, varav cirka 2 km2 består av vatten.
linkkiVanda stad:
Grundläggande informationfinska _ svenska _ engelska
Historia
Vanda område har varit bebott länge.
Man har hittat upp till 7 000 år gamla lämningar efter bosättning.
Nuvarande Vanda har uppstått på ett område som förr var Helsingfors socken.
Helsingfors sockens historia sträcker sig ända till 1300-talet.
Helsingfors socken blev först Helsingfors landskommun, sedan Vanda köping år 1972 och till slut Vanda stad år 1974.
Läget som granne till huvudstaden Helsingfors har varit viktigt för Vanda.
Viktiga vägar, såsom vägen från Åbo via Helsingfors till Viborg och senare järnvägen norrut från Helsingfors, har gått genom Vanda.
Längs med vägarna och järnvägen har det utvecklats industrier och bostadsområden.
Vanda är än idag en viktig trafikknutpunkt.
Till exempel ligger Helsingfors-Vanda flygplats i Vanda.
linkkiVanda stad:
Information om Vandafinska
linkkiVanda stad:
Stadsmuseetfinska _ svenska _ engelska
Trafik
Beslutsfattande och påverkan
Religion
Grundläggande information
Historia
Trafik
Kollektivtrafiken
Vanda och hela huvudstadsregionen har goda kollektivtrafikförbindelser.
Längs stambanan och Mårtensdals bana finns flera tågstationer.
I staden finns flera busslinjer.
Vanda tillhör samkommunen Helsingforsregionens trafik (HRT) (Helsingin seudun liikenne -kuntayhtymä (HSL)), som ordnar kollektivtrafiken i huvudstadsregionen.
Mer information hittar du på HRT:s webbplats.
Du kan söka information om rutterna i Reseplaneraren (Reittiopas).
Tjänsten ger dig förslag på olika kollektivtrafikförbindelser från ett ställe till ett annat.
I kollektivtrafiken kan du betala med kontanter eller resekort.
I närtågen måste du köpa biljetten i förväg.
Du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat.
Reseplanerarefinska _ svenska _ engelska
Resekort
Med ett resekort (matkakortti) reser du förmånligare än med kontanter.
Resekortet gäller i lokaltrafikens bussar, närtågen, metron, spårvagnarna och Sveaborgsfärjorna.
Det finns två slags resekort.
Det är det billigaste sättet att resa.
Ett innehavarkort (haltijakohtainen kortti) kan användas av flera personer.
Innan du skaffar dig ett personligt kort ska du registrera dig som invånare i någon av kommunerna inom HRT-området.
Du kan köpa resekort vid HRT:s försäljningsställen (myyntipiste) eller serviceställen (palvelupiste).
De finns runtom i huvudstadsregionen.
Personligt resekort kan du köpa vid serviceställena.
Ta med dig identitetsbevis om du ska köpa personligt resekort.
Om du har finska nätbankskoder kan du även köpa personligt resekort på HRT:s webbplats.
Du kan resa med resekortet när du laddar kortet med period (kausi) eller värde (arvo).
En period betyder tid: till exempel en månad.
Värde betyder pengar.
Om du använder kollektivtrafiken ofta tjänar du på att ladda kortet med period.
Du kan ladda resekortet på vilket serviceställe för resekort (matkakortin latauspiste) som helst.
Du hittar mer information på HRT:s webbplats.
Ansökan om försäljningsplatserfinska _ svenska _ engelska
Information och råd till resenärerfinska _ svenska _ engelska
Biljetter och priserfinska _ svenska _ engelska
Att gå och cykla
Om du vill gå eller cykla i Vanda kan du söka en lämplig rutt i reseplaneraren för cykling och gång.
En cykelkarta i pappersformat för Vanda kan du hämta i Vandainfo.
Cykelkartorna är kostnadsfria.
linkkiVanda stad:
Vandainfofinska _ svenska _ engelska
Bil och flyg
Helsingfors-Vanda internationella flygplats ligger i Vanda.
Flygplatsen har goda trafikförbindelser till exempel med bil, buss och tåg.
Du kan parkera bilen på många järnvägsstationer och fortsätta färden med kollektivtrafiken.
Tidtabellerna för bussar och tåg hittar du enkelt i reseplaneraren.
Läs mer: Trafik.
Flygplatsenfinska _ svenska _ engelska _ ryska _ kinesiska
Beslutsfattande och påverkan
I Vanda beslutas ärenden av stadsfullmäktige (kaupunginvaltuusto).
I stadsfullmäktige sitter 67 ledamöter som representerar olika politiska grupper.
Fullmäktige väljs var fjärde år genom kommunalval (kunnallisvaalit).
Invånarna i Vanda kan påverka beslutsfattandet och beredning av ärenden på många olika sätt.
På Vandakanalen kan du följa fullmäktiges sammanträden och få mer information om beslutsfattandet.
I Vanda finns en delegation för mångkulturella frågor (monikulttuurisuusasiain neuvottelukunta) som lägger fram propositioner i ärenden som rör invandrare.
Läs mer på Vanda stads webbplats.
I Vanda finns många politiska föreningar, invandrarföreningar och andra föreningar via vilka du också kan påverka beslutsfattandet.
Mer information om föreningarna hittar du på sidan Vantaalla.info.
linkkiVanda stad:
Beslutsfattandefinska _ svenska _ engelska
linkkiVanda stad:
Delta och påverkafinska
Stadsfullmäktiges sammanträden på Internetfinska
linkkiVanda stad:
Delegationen för mångkulturella frågorfinska
Religion
Många religiösa samfund är verksamma i Vanda och Helsingfors.
Via tjänsten Uskonnot Suomessa kan du söka information efter det religiösa samfundet och orten.
Den evangelisk-lutherska kyrkan har sex finskspråkiga församlingar och en svenskspråkig församling i Vanda.
Läs mer på Vanda kyrkliga samfällighets webbplats.
I Dickursby finns en ortodox kyrka.
Mer information om verksamheten vid den ortodoxa kyrkan i Vanda hittar du på Helsingfors ortodoxa församlings webbplats.
Läs mer: Kulturer och religioner i Finland.
linkkiVanda kyrkliga samfällighet:
Evangelisk-lutherska församlingarfinska
linkkiHelsingfors ortodoxa församling:
Ortodoxa församlingenfinska _ ryska
Religiösa samfundfinska _ engelska
Grundläggande information
Vanda är en av de fyra kommunerna i huvudstadsregionen.
Den ligger intill Esbo och Helsingfors.
Vanda centrum ligger i Dickursby.
Därtill finns det andra stora tätorter i Vanda, till exempel Korso, Björkby-Havukoski, Myrbacka, Mårtensdal, Håkansböle, Västerkulla och Backas.
Vanda har drygt 205 000 invånare.
Av dem är cirka 2,8 procent svenskspråkiga och 11 procent har något annat modersmål än finska eller svenska.
Arealen är cirka 240 km2, varav cirka 2 km2 består av vatten.
linkkiVanda stad:
Grundläggande informationfinska _ svenska _ engelska
Historia
Vanda område har varit bebott länge.
Man har hittat upp till 7 000 år gamla lämningar efter bosättning.
Nuvarande Vanda har uppstått på ett område som förr var Helsingfors socken.
Helsingfors sockens historia sträcker sig ända till 1300-talet.
Helsingfors socken blev först Helsingfors landskommun, sedan Vanda köping år 1972 och till slut Vanda stad år 1974.
Läget som granne till huvudstaden Helsingfors har varit viktigt för Vanda.
Viktiga vägar, såsom vägen från Åbo via Helsingfors till Viborg och senare järnvägen norrut från Helsingfors, har gått genom Vanda.
Längs med vägarna och järnvägen har det utvecklats industrier och bostadsområden.
Vanda är än idag en viktig trafikknutpunkt.
Till exempel ligger Helsingfors-Vanda flygplats i Vanda.
linkkiVanda stad:
Information om Vandafinska
linkkiVanda stad:
Stadsmuseetfinska _ svenska _ engelska
Bibliotek
Motion
Att röra sig i naturen
Teater och film
Museer
Fritidsverksamhet för barn och unga
Fritidsverksamhet för seniorer
Föreningar
Vid Vanda vuxenutbildningsinstitut (Vantaan Aikuisopisto) kan man till exempel skapa konst, handarbeten, laga mat eller dansa.
Man kan även studera språk.
I Vanda finns två kulturhus: konserthuset Martinus och allaktivitetscentret Myrbackahuset.
Dessutom ordnar allaktivitetscentret LUMO många evenemang.
Kulturhuset för barn och unga Fernissan, Konsthuset Pessi och Konsthuset Totem ordnar kulturevenemang för barn.
Läs mer: Fritid.
linkkiVanda vuxenutbildningsinstitut:
Studiehandbokfinska
linkkiVanda stad:
Kulturevenemangfinska _ svenska _ engelska
Konserterfinska _ svenska _ engelska
Evenemangfinska _ engelska
linkkiKulturhuset för barn och unga Fernissan:
Kulturevenemang för barnfinska
Kulturevenemang för barnfinska
Kulturevenemang för barnfinska _ svenska
linkkiVanda stad:
Evenemang och festivalerfinska _ engelska
Bibliotek
I Vanda finns 10 bibliotek (kirjasto) och två bokbussar (kirjastoauto).
På biblioteket kan du låna böcker, tidningar, musik, filmer, spel och mycket annat.
Böcker och annat material finns på flera olika språk.
På biblioteket kan du också använda dator.
På vissa bibliotek ordnas även språkcaféer i det finska språket för invandrare.
Biblioteken i Vanda är med i huvudstadsregionens bibliotekstjänst HelMet.
Du kan alltså använda samma bibliotekskort på stadsbiblioteken i Vanda, Esbo, Grankulla och Helsingfors.
I Helsingfors huvudbibliotek i Böle finns Flerspråkigt bibliotek.
Där hittar man böcker på över 60 olika språk.
Om du har ett Helmet-lånekort, kan du också låna böcker i Flerspråkiga biblioteket.
Läs mer: Bibliotek
linkkiVanda stad:
Information om bibliotekenfinska _ svenska _ engelska
linkkiHelsingfors stadsbibliotek:
Flerspråkiga biblioteketfinska _ svenska _ engelska
Motion
I Vanda finns fem kommunala simhallar.
Simhallen i Korso har ett eget simpass för invandrarkvinnor och -flickor.
I Vanda finns flera idrottshallar, idrottsplaner och andra idrottsplatser för olika idrottsgrenar.
På motionsslingorna kan man springa på somrarna och åka skidor på vintrarna.
Läs mer: Motion.
linkkiVanda stad:
Simhallarnas kontaktuppgifterfinska _ svenska _ engelska
linkkiVanda stad:
Simpass för invandrarkvinnorfinska _ engelska
linkkiVanda stad:
Idrottsklubbarfinska
Att röra sig i naturen
I Vanda finns många motionsslingor och naturstigar.
Du kan även röra dig i naturen i Petikkos rekreationsområde.
Du kan fiska på Vanda stads fiskeområden i Vanda å, Kervo å och på Finska viken.
Läs mer: Att röra sig i naturen.
linkkiVanda stad:
Rekreations- och campingområdenfinska _ svenska
linkkiVanda stad:
Idrottsplatser och friluftsområdenfinska _ svenska
Friluftsområdenfinska
linkkiVanda stad:
Fiske och båtlivfinska
Teater och film
I Vanda finns flera yrkes- och amatörteatrar.
I Vanda finns fyra biografer.
Mer information om filmerna hittar du på biografernas webbplatser.
Därtill ordnar Vanda stad filmvisningar.
Läs mer: Teater och film.
linkkiVanda stad:
Film, dans och teaterfinska _ engelska
Museer
I Vanda finns flera museer.
På Vanda konstmuseum ordnas växlande utställningar med inhemsk och utländsk modern konst.
Om de övriga museerna hittar du information på Vanda stads webbplats.
Läs mer: Museer.
linkkiVanda stad:
Museerfinska _ engelska
linkkiVanda stad:
Stadsmuseetfinska _ svenska _ engelska
linkkiVanda stad:
Konstmuseetfinska _ svenska _ engelska
Fritidsverksamhet för barn och unga
I Vanda finns flera läroanstalter som ger grundundervisning i konst speciellt för barn och unga.
Olika konstarter är musik, bildkonst, dans, teater, cirkuskonst, ordkonst, handarbete och arkitektur.
Stadens ungdomsgårdar är öppna för alla ungdomar i åldrarna 10–17 år.
Projektet Sport för alla (Sporttia kaikille-hanke) ordnar idrottsklubbar, turneringar och läger för barn och ungdomar med invandrarbakgrund.
Också föreningar och idrottsklubbar ordnar mycket verksamhet för ungdomar.
Mer information hittar du på Vanda stads webbplats.
Läs mer: Fritidsverksamhet för barn och unga.
linkkiVanda stad:
Information om hobbymöjligheter för ungdomarfinska
linkkiVanda stad:
Kultur för barn och ungafinska _ svenska _ engelska
linkkiVanda stad:
Information om konstundervisningfinska _ engelska
Ungdomsgårdarfinska
Motionsmöjligheterfinska
Hobbysökningfinska
linkkiVanda stad:
Delta och påverkafinska _ svenska
Fritidsverksamhet för seniorer
Om du har fyllt 70 år och Vanda är din hemkommun kan du kostnadsfritt använda Vanda stads simhallar och gym. Du kommer gratis in till idrottsanläggningarna om du har ett Sportkort (Sporttikortti).
Du kan avhämta Sportkortet kostnadsfritt vid Vanda-informationspunkterna.
Ta med dig identitetsbevis och ett foto när du ansöker om kortet.
På Seniorrådgivningen (seniorineuvonta) får du information om hobbyer och tjänster för seniorer som olika organisationer, företag och staden erbjuder.
Seniorrådgivningen
Tfn: (09) 8392 4202
Motionsmöjligheterfinska _ svenska
Föreningar
I Vanda finns många olika föreningar, till exempel kulturföreningar och idrottsklubbar.
Mer information hittar du på Vanda stads webbplats.
Läs mer: Föreningar.
linkkiVanda stad:
Kulturföreningarfinska
linkkiVanda stad:
Idrottsklubbarfinska
Bibliotek
Motion
Att röra sig i naturen
Teater och film
Museer
Fritidsverksamhet för barn och unga
Fritidsverksamhet för seniorer
Föreningar
Vid Vanda vuxenutbildningsinstitut (Vantaan Aikuisopisto) kan man till exempel skapa konst, handarbeten, laga mat eller dansa.
Man kan även studera språk.
I Vanda finns två kulturhus: konserthuset Martinus och allaktivitetscentret Myrbackahuset.
Dessutom ordnar allaktivitetscentret LUMO många evenemang.
Kulturhuset för barn och unga Fernissan, Konsthuset Pessi och Konsthuset Totem ordnar kulturevenemang för barn.
Läs mer: Fritid.
linkkiVanda vuxenutbildningsinstitut:
Studiehandbokfinska
linkkiVanda stad:
Kulturevenemangfinska _ svenska _ engelska
Konserterfinska _ svenska _ engelska
Evenemangfinska _ engelska
linkkiKulturhuset för barn och unga Fernissan:
Kulturevenemang för barnfinska
Kulturevenemang för barnfinska
Kulturevenemang för barnfinska _ svenska
linkkiVanda stad:
Evenemang och festivalerfinska _ engelska
Bibliotek
I Vanda finns 10 bibliotek (kirjasto) och två bokbussar (kirjastoauto).
På biblioteket kan du låna böcker, tidningar, musik, filmer, spel och mycket annat.
Böcker och annat material finns på flera olika språk.
På biblioteket kan du också använda dator.
På vissa bibliotek ordnas även språkcaféer i det finska språket för invandrare.
Biblioteken i Vanda är med i huvudstadsregionens bibliotekstjänst HelMet.
Du kan alltså använda samma bibliotekskort på stadsbiblioteken i Vanda, Esbo, Grankulla och Helsingfors.
I Helsingfors huvudbibliotek i Böle finns Flerspråkigt bibliotek.
Där hittar man böcker på över 60 olika språk.
Om du har ett Helmet-lånekort, kan du också låna böcker i Flerspråkiga biblioteket.
Läs mer: Bibliotek
linkkiVanda stad:
Information om bibliotekenfinska _ svenska _ engelska
linkkiHelsingfors stadsbibliotek:
Flerspråkiga biblioteketfinska _ svenska _ engelska
Motion
I Vanda finns fem kommunala simhallar.
Simhallen i Korso har ett eget simpass för invandrarkvinnor och -flickor.
I Vanda finns flera idrottshallar, idrottsplaner och andra idrottsplatser för olika idrottsgrenar.
På motionsslingorna kan man springa på somrarna och åka skidor på vintrarna.
Läs mer: Motion.
linkkiVanda stad:
Simhallarnas kontaktuppgifterfinska _ svenska _ engelska
linkkiVanda stad:
Simpass för invandrarkvinnorfinska _ engelska
linkkiVanda stad:
Idrottsklubbarfinska
Att röra sig i naturen
I Vanda finns många motionsslingor och naturstigar.
Du kan även röra dig i naturen i Petikkos rekreationsområde.
Du kan fiska på Vanda stads fiskeområden i Vanda å, Kervo å och på Finska viken.
Läs mer: Att röra sig i naturen.
linkkiVanda stad:
Rekreations- och campingområdenfinska _ svenska
linkkiVanda stad:
Idrottsplatser och friluftsområdenfinska _ svenska
Friluftsområdenfinska
linkkiVanda stad:
Fiske och båtlivfinska
Teater och film
I Vanda finns flera yrkes- och amatörteatrar.
I Vanda finns fyra biografer.
Mer information om filmerna hittar du på biografernas webbplatser.
Därtill ordnar Vanda stad filmvisningar.
Läs mer: Teater och film.
linkkiVanda stad:
Film, dans och teaterfinska _ engelska
Museer
I Vanda finns flera museer.
På Vanda konstmuseum ordnas växlande utställningar med inhemsk och utländsk modern konst.
Om de övriga museerna hittar du information på Vanda stads webbplats.
Läs mer: Museer.
linkkiVanda stad:
Museerfinska _ engelska
linkkiVanda stad:
Stadsmuseetfinska _ svenska _ engelska
linkkiVanda stad:
Konstmuseetfinska _ svenska _ engelska
Fritidsverksamhet för barn och unga
I Vanda finns flera läroanstalter som ger grundundervisning i konst speciellt för barn och unga.
Olika konstarter är musik, bildkonst, dans, teater, cirkuskonst, ordkonst, handarbete och arkitektur.
Stadens ungdomsgårdar är öppna för alla ungdomar i åldrarna 10–17 år.
Projektet Sport för alla (Sporttia kaikille-hanke) ordnar idrottsklubbar, turneringar och läger för barn och ungdomar med invandrarbakgrund.
Också föreningar och idrottsklubbar ordnar mycket verksamhet för ungdomar.
Mer information hittar du på Vanda stads webbplats.
Läs mer: Fritidsverksamhet för barn och unga.
linkkiVanda stad:
Information om hobbymöjligheter för ungdomarfinska
linkkiVanda stad:
Kultur för barn och ungafinska _ svenska _ engelska
linkkiVanda stad:
Information om konstundervisningfinska _ engelska
Ungdomsgårdarfinska
Motionsmöjligheterfinska
Hobbysökningfinska
linkkiVanda stad:
Delta och påverkafinska _ svenska
Fritidsverksamhet för seniorer
Om du har fyllt 70 år och Vanda är din hemkommun kan du kostnadsfritt använda Vanda stads simhallar och gym. Du kommer gratis in till idrottsanläggningarna om du har ett Sportkort (Sporttikortti).
Du kan avhämta Sportkortet kostnadsfritt vid Vanda-informationspunkterna.
Ta med dig identitetsbevis och ett foto när du ansöker om kortet.
På Seniorrådgivningen (seniorineuvonta) får du information om hobbyer och tjänster för seniorer som olika organisationer, företag och staden erbjuder.
Seniorrådgivningen
Tfn: (09) 8392 4202
Motionsmöjligheterfinska _ svenska
Föreningar
I Vanda finns många olika föreningar, till exempel kulturföreningar och idrottsklubbar.
Mer information hittar du på Vanda stads webbplats.
Läs mer: Föreningar.
linkkiVanda stad:
Kulturföreningarfinska
linkkiVanda stad:
Idrottsklubbarfinska
Bibliotek
Motion
Att röra sig i naturen
Teater och film
Museer
Fritidsverksamhet för barn och unga
Fritidsverksamhet för seniorer
Föreningar
Vid Vanda vuxenutbildningsinstitut (Vantaan Aikuisopisto) kan man till exempel skapa konst, handarbeten, laga mat eller dansa.
Man kan även studera språk.
I Vanda finns två kulturhus: konserthuset Martinus och allaktivitetscentret Myrbackahuset.
Dessutom ordnar allaktivitetscentret LUMO många evenemang.
Kulturhuset för barn och unga Fernissan, Konsthuset Pessi och Konsthuset Totem ordnar kulturevenemang för barn.
Läs mer: Fritid.
linkkiVanda vuxenutbildningsinstitut:
Studiehandbokfinska
linkkiVanda stad:
Kulturevenemangfinska _ svenska _ engelska
Konserterfinska _ svenska _ engelska
Evenemangfinska _ engelska
linkkiKulturhuset för barn och unga Fernissan:
Kulturevenemang för barnfinska
Kulturevenemang för barnfinska
Kulturevenemang för barnfinska _ svenska
linkkiVanda stad:
Evenemang och festivalerfinska _ engelska
Bibliotek
I Vanda finns 10 bibliotek (kirjasto) och två bokbussar (kirjastoauto).
På biblioteket kan du låna böcker, tidningar, musik, filmer, spel och mycket annat.
Böcker och annat material finns på flera olika språk.
På biblioteket kan du också använda dator.
På vissa bibliotek ordnas även språkcaféer i det finska språket för invandrare.
Biblioteken i Vanda är med i huvudstadsregionens bibliotekstjänst HelMet.
Du kan alltså använda samma bibliotekskort på stadsbiblioteken i Vanda, Esbo, Grankulla och Helsingfors.
I Helsingfors huvudbibliotek i Böle finns Flerspråkigt bibliotek.
Där hittar man böcker på över 60 olika språk.
Om du har ett Helmet-lånekort, kan du också låna böcker i Flerspråkiga biblioteket.
Läs mer: Bibliotek
linkkiVanda stad:
Information om bibliotekenfinska _ svenska _ engelska
linkkiHelsingfors stadsbibliotek:
Flerspråkiga biblioteketfinska _ svenska _ engelska
Motion
I Vanda finns fem kommunala simhallar.
Simhallen i Korso har ett eget simpass för invandrarkvinnor och -flickor.
I Vanda finns flera idrottshallar, idrottsplaner och andra idrottsplatser för olika idrottsgrenar.
På motionsslingorna kan man springa på somrarna och åka skidor på vintrarna.
Läs mer: Motion.
linkkiVanda stad:
Simhallarnas kontaktuppgifterfinska _ svenska _ engelska
linkkiVanda stad:
Simpass för invandrarkvinnorfinska _ engelska
linkkiVanda stad:
Idrottsklubbarfinska
Att röra sig i naturen
I Vanda finns många motionsslingor och naturstigar.
Du kan även röra dig i naturen i Petikkos rekreationsområde.
Du kan fiska på Vanda stads fiskeområden i Vanda å, Kervo å och på Finska viken.
Läs mer: Att röra sig i naturen.
linkkiVanda stad:
Rekreations- och campingområdenfinska _ svenska
linkkiVanda stad:
Idrottsplatser och friluftsområdenfinska _ svenska
Friluftsområdenfinska
linkkiVanda stad:
Fiske och båtlivfinska
Teater och film
I Vanda finns flera yrkes- och amatörteatrar.
I Vanda finns fyra biografer.
Mer information om filmerna hittar du på biografernas webbplatser.
Därtill ordnar Vanda stad filmvisningar.
Läs mer: Teater och film.
linkkiVanda stad:
Film, dans och teaterfinska _ engelska
Museer
I Vanda finns flera museer.
På Vanda konstmuseum ordnas växlande utställningar med inhemsk och utländsk modern konst.
Om de övriga museerna hittar du information på Vanda stads webbplats.
Läs mer: Museer.
linkkiVanda stad:
Museerfinska _ engelska
linkkiVanda stad:
Stadsmuseetfinska _ svenska _ engelska
linkkiVanda stad:
Konstmuseetfinska _ svenska _ engelska
Fritidsverksamhet för barn och unga
I Vanda finns flera läroanstalter som ger grundundervisning i konst speciellt för barn och unga.
Olika konstarter är musik, bildkonst, dans, teater, cirkuskonst, ordkonst, handarbete och arkitektur.
Stadens ungdomsgårdar är öppna för alla ungdomar i åldrarna 10–17 år.
Projektet Sport för alla (Sporttia kaikille-hanke) ordnar idrottsklubbar, turneringar och läger för barn och ungdomar med invandrarbakgrund.
Också föreningar och idrottsklubbar ordnar mycket verksamhet för ungdomar.
Mer information hittar du på Vanda stads webbplats.
Läs mer: Fritidsverksamhet för barn och unga.
linkkiVanda stad:
Information om hobbymöjligheter för ungdomarfinska
linkkiVanda stad:
Kultur för barn och ungafinska _ svenska _ engelska
linkkiVanda stad:
Information om konstundervisningfinska _ engelska
Ungdomsgårdarfinska
Motionsmöjligheterfinska
Hobbysökningfinska
linkkiVanda stad:
Delta och påverkafinska _ svenska
Fritidsverksamhet för seniorer
Om du har fyllt 70 år och Vanda är din hemkommun kan du kostnadsfritt använda Vanda stads simhallar och gym. Du kommer gratis in till idrottsanläggningarna om du har ett Sportkort (Sporttikortti).
Du kan avhämta Sportkortet kostnadsfritt vid Vanda-informationspunkterna.
Ta med dig identitetsbevis och ett foto när du ansöker om kortet.
På Seniorrådgivningen (seniorineuvonta) får du information om hobbyer och tjänster för seniorer som olika organisationer, företag och staden erbjuder.
Seniorrådgivningen
Tfn: (09) 8392 4202
Motionsmöjligheterfinska _ svenska
Föreningar
I Vanda finns många olika föreningar, till exempel kulturföreningar och idrottsklubbar.
Mer information hittar du på Vanda stads webbplats.
Läs mer: Föreningar.
linkkiVanda stad:
Kulturföreningarfinska
linkkiVanda stad:
Idrottsklubbarfinska
Problem med uppehållstillståndet
Brott
Behöver du en jurist?
Våld
Missbruksproblem och spelberoende
Dödsfall
Om du behöver brådskande hjälp av polisen, brandkåren eller ambulansen, ring nödnumret 112.
Du får ringa nödnumret endast i brådskande nödfall där liv, hälsa, egendom eller miljö är i fara.
Om du drabbas av en akut krissituation, såsom att en närstående avlider eller på grund av familjevåld, kan du kontakta social- och krisjouren (sosiaali- ja kriisipäivystys).
Du kan också söka hjälp för en familjemedlem eller en vän.
Social- och krisjouren har öppet dygnet runt varje dag.
Social- och krisjouren
Tfn (09) 8392 4005
linkkiNödcentralsverket:
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
linkkiVanda stad:
Social- och krisjourenfinska _ svenska _ engelska
Problem med uppehållstillståndet
Om du har problem eller oklarheter med uppehållstillståndet, kontakta Migrationsverket.
Du kan även fråga om råd på rådgivningstjänsterna för invandrare.
Information om tjänsterna finns på sidan Som invandrare i Vanda.
Migrationsverkets närmaste tjänsteställe finns i Helsingfors:
Göksgränd 3A
Läs mer: Problem med uppehållstillståndet
Olika tillståndfinska _ svenska _ engelska
Hälsovård för papperslösa
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärhälsovård.
Tjänsterna vid Global Clinic är avgiftsfria för kunderna.
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter.
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
Telefonnumret till Global Clinic i Helsingfors är 044 977 4547.
Samtalet besvaras av en sjukskötare eller en läkare.
E-postadressen är globalclinic.finland(at)gmail.com.
Läs mer: Problem med uppehållstillstånd
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Brott
Brottsanmälan (rikosilmoitus) kan göras per telefon eller personligen på polisstationen.
Du kan också göra brottsanmälan på internet om brottet i fråga är ringa och du inte behöver omedelbar hjälp av polisen.
Konvaljvägen 21
Tfn 0295 430291
Läs mer: Brott.
Kontaktuppgifterfinska _ svenska
Elektronisk polisanmälanfinska _ svenska _ engelska
Behöver du en jurist?
Östra Nylands rättshjälpsbyrå (Itä-Uudenmaan oikeusaputoimisto) betjänar invånarna i Vanda.
Pyrolavägen 37
Tfn 029 5660 160
Du kan också söka information om privata jurister på till exempel Finlands Juristförbunds (Suomen Asianajajaliitto) webbplats.
Läs mer: Behöver du en jurist?
linkkiÖstra Nylands rättshjälpsbyrå:
Information om rättshjälpfinska _ svenska _ engelska
linkkiFinlands Advokatförbund:
Advokaterfinska _ svenska _ engelska
Våld
I nödsituationer ringer du nödnumret 112.
I krissituationer får man även hjälp vid Vanda stads social- och krisjour (sosiaali- ja kriisipäivystys), som har öppet dygnet runt.
Social- och krisjouren
Tfn (09) 8392 4005
linkkiNödcentralsverket:
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
Skyddshem
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta ett skyddshem (turvakoti).
Skyddshemmen har jourmottagning dygnet runt.
Skyddshemmet Mona (turvakoti Mona) är ett skyddshem avsett för invandrarkvinnor och deras barn.
Tfn 045 639 6274
linkkiTurvakoti Mona:
Skyddshemfinska
Du kan även gå till Vanda skyddshem (Vantaan turvakoti) eller huvudstadsregionens skyddshem (pääkaupunkiseudun turvakoti).
Puh. (09) 8392 0071
Skyddshemfinska _ engelska
Steniusvägen 20
Tfn (09) 4777 180
Hjälp till offer för familjevåldfinska
Hjälp för invandrarkvinnor
Föreningen Monika-Naiset liitto (Monika-Naiset Liitto) ger råd och stöd till invandrarkvinnor.
Föreningen har ett resurscenter (voimavarakeskus) i Vanda där man får stöd och råd.
Tfn (09) 839 35013
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Hjälp för män
Män som har utövat våld mot sina familjemedlemmar eller har själva blivit offer för våld i hemmet, kan få hjälp från Jussi-arbetet i Vanda (Vantaan Jussi-työ).
Hjälp för män att sluta med våldsamt beteendefinska
Miehen linja (Miehen linja) hjälper invandrarmän som har problem med våld.
Tfn (09) 276 62899
Hjälp för män för att sluta med våldsamt beteendefinska _ engelska
Hjälp för unga
Finlands Röda Kors De ungas skyddshus (Suomen Punaisen Ristin Nuorten turvatalo) ger stöd och hjälp i krissituationer för 12–19-åringar.
Skyddshuset har öppet kl. 17–10, telefonjouren betjänar dygnet runt.
Sjukhusgatan 3 (Räckhals gård)
Tfn (09) 871 4043
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Läs mer: Våld
Problem i äktenskap eller parförhållande
Par med barn under 13 år kan vid problem i äktenskap och parförhållande få hjälp vid familjerådgivningen (perheneuvola).
Kontaktuppgifterna hittar du på Vanda stads webbplats.
Familjerådgivningens tjänster är konfidentiella och avgiftsfria.
Vid akuta krissituationer inom familjen kan du kontakta social- och krisjouren (sosiaali- ja kriisipäivystys), som har öppet dygnet runt varje dag.
Social- och krisjouren
Tfn (09) 8392 4005
Vid problem i parförhållandet och familjen får man även hjälp av familjerådgivningen vid Vanda församlingar (Vantaan seurakunnan perheneuvonta).
Läs mer: Problem i äktenskap och parförhållande
linkkiVanda stad:
Familjerådgivningarfinska _ svenska
linkkiVanda kyrkliga samfällighet:
Familjerådgivningfinska _ engelska
Barnrådgivningsbyråerna (lastenneuvola) och familjerådgivningsbyråerna (perheneuvola) ger råd i frågor som rör barns hälsa, uppväxt och utveckling.
Vid problem hos barn i skolåldern får man hjälp hos skolhälsovårdarna (kouluterveydenhoitaja), skolkuratorerna (koulukuraattori) och socialhandledarna (sosiaaliohjaaja).
Mer information hittar du på Vanda stads webbplats.
Läs mer: Barns och ungas problem
linkkiVanda stad:
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad:
Familjerådgivningarfinska _ svenska
linkkiVanda stad:
Information om tjänster för barn, ungdomar och familjerfinska _ svenska _ engelska
I skolan får de unga hjälp av skol- och studenthälsovårdarna (koulu- ja opiskeluterveydenhoitajat), skolkuratorerna (koulukuraattorit) och skolpsykologerna (koulupsykologit).
linkkiVanda stad:
Information om skolhälsovårdenfinska _ svenska _ engelska
linkkiVanda stad:
Skolkuratorerfinska _ svenska
linkkiVanda stad:
Skolpsykologerfinska _ svenska
Nuppi
13–21-åriga barn och ungdomar samt deras familjer kan få hjälp hos ungdomscentralen (nuortenkeskus).
På Nuppi kan du till exempel få hjälp med mentala problem och missbruksproblem.
Hjälp för ungafinska _ svenska _ engelska
Om du är under 30 år, kan du få råd och handledning via tjänsten Navigatorn.
Personalen vid Navigatorn hjälper dig om du inte har något arbete eller en studieplats.
Du kan även be om råd gällande andra saker, till exempel boende och ekonomi.
De ungas skyddshus
Finlands Röda Kors De ungas skyddshus (Suomen Punaisen Ristin Nuorten turvatalo) ger stöd och hjälp i krissituationer för 12–19-åringar.
Skyddshuset har öppet kl. 17–10, telefonjouren betjänar dygnet runt.
Sjukhusgatan 3
Tfn (09) 871 4043
Läs mer: Barns och ungas problem
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Vägledning och stöd för ungafinska _ svenska
Socialrådgivningen (sosiaalineuvonta) ger information om utkomststöd (toimeentulotuki) och andra bidrag om du har ekonomiska problem.
Tfn (09) 83 911.
linkkiVanda stad:
Socialrådgivningenfinska _ svenska _ engelska
Utkomststöd
Utkomststödet (toimeentulotuki) är avsett som en sista utväg då du inte har några andra inkomster eller medel, eller om dina inkomster är mycket låga.
Utkomststöd kan du få om du inte lyckas få tillräckliga inkomster genom eget arbete, andras omsorg eller på något annat sätt.
Du kan be om råd gällande ansökan om utkomststöd via den centraliserade telefontjänsten tfn (09) 8392 1119.
linkkiVanda stad:
Information om utkomststödfinska _ svenska _ engelska
Ekonomi- och skuldrådgivning
Om du inte kan betala dina räkningar eller skulder då de förfaller, ska du kontakta skuldrådgivningen (velkaneuvonta).
Tfn (09) 8392 2120.
linkkiVanda ekonomi- och skuldrådgivning:
Ekonomi- och skuldrådgivningfinska _ svenska _ engelska
Social kreditgivning
Om du har låga inkomster och är medellös samt har svårt att få lån, kan du ansöka om lån via den sociala kreditgivningen (sosiaalinen luototus).
Telefonnumret till kundrådgivningen och tidsbokningen är (09) 8392 0173.
linkkiVanda stad:
Information om social kreditgivningfinska _ svenska _ engelska
Missbruksproblem och spelberoende
Itä-Vantaan A-klinikka
Konvaljvägen 20 C vån.
tfn (09) 8392 3415
Länsi-Vantaan A-klinikka
tfn (09) 8393 5534
H-klinikka
Eldstadsvägen 7 B, vån.
Tfn (09) 839 21064
H-kliniken har också verksamhetsställen på Dickursby och Myrbacka hälsostationer.
Om du har spelproblem kan du söka hjälp vid Spelkliniken (Peliklinikka), som finns i centrala Helsingfors.
Peliklinikka
tfn 040 152 3918.
Ungdomscentralen Nuppi (nuortenkeskus Nuppi) hjälper ungdomar med missbruksproblem, Internetberoende eller spelberoende.
Nuppi ger också stöd till ungdomar som oroar sig för rusmedelsbruket hos någon närstående person.
Läs mer: Missbruksproblem.
linkkiVanda stad:
Hjälp med missbruksproblemfinska _ svenska _ engelska
linkkiVanda stad:
Information om vård av drogproblemfinska _ svenska _ engelska
Hjälp med penningspelproblemfinska
Hjälp för ungafinska _ svenska _ engelska
Dödsfall
I Vanda finns fyra begravningsplatser som tillhör de evangelisk-lutherska församlingarna.
I Furumo i Vanda finns dessutom Vandas och Helsingfors gemensamma begravningsplats för avlidna personer som inte har varit medlemmar i något religionssamfund.
Information om begravning får du på Vanda församlingars gravkontor (Vantaan seurakuntien hautaustoimisto) och vid privata begravningsbyråer (hautaustoimisto).
Vanda församlingars gravkontor
Prästgårdsgränden 5
Tfn (09) 8306 220
Om din närstående avlider plötsligt, kan du få hjälp med att återhämta dig från den chockartade upplevelsen och stöd i att klara dig efter förlusten av Vandas social- och krisjour (sosiaali- ja kriisipäivystys).
Jouren har öppet varje dag dygnet runt.
Social- och krisjouren
Tfn (09) 8392 4005
Läs mer: Död
linkkiVanda kyrkliga samfällighet:
Begravningsplatserfinska
linkkiHelsingfors kyrkliga samfällighet:
Konfessionslös begravningsplatsfinska
linkkiFinlands Begravningbyråers Förbund:
Begravningsbyråerfinska _ svenska _ engelska
När en närstående har avliditfinska _ svenska _ engelska
linkkiVanda stad:
Social- och krisjourenfinska _ svenska _ engelska
Problem med uppehållstillståndet
Brott
Behöver du en jurist?
Våld
Missbruksproblem och spelberoende
Dödsfall
Om du behöver brådskande hjälp av polisen, brandkåren eller ambulansen, ring nödnumret 112.
Du får ringa nödnumret endast i brådskande nödfall där liv, hälsa, egendom eller miljö är i fara.
Om du drabbas av en akut krissituation, såsom att en närstående avlider eller på grund av familjevåld, kan du kontakta social- och krisjouren (sosiaali- ja kriisipäivystys).
Du kan också söka hjälp för en familjemedlem eller en vän.
Social- och krisjouren har öppet dygnet runt varje dag.
Social- och krisjouren
Tfn (09) 8392 4005
linkkiNödcentralsverket:
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
linkkiVanda stad:
Social- och krisjourenfinska _ svenska _ engelska
Problem med uppehållstillståndet
Om du har problem eller oklarheter med uppehållstillståndet, kontakta Migrationsverket.
Du kan även fråga om råd på rådgivningstjänsterna för invandrare.
Information om tjänsterna finns på sidan Som invandrare i Vanda.
Migrationsverkets närmaste tjänsteställe finns i Helsingfors:
Göksgränd 3A
Läs mer: Problem med uppehållstillståndet
Olika tillståndfinska _ svenska _ engelska
Hälsovård för papperslösa
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärhälsovård.
Tjänsterna vid Global Clinic är avgiftsfria för kunderna.
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter.
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
Telefonnumret till Global Clinic i Helsingfors är 044 977 4547.
Samtalet besvaras av en sjukskötare eller en läkare.
E-postadressen är globalclinic.finland(at)gmail.com.
Läs mer: Problem med uppehållstillstånd
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Brott
Brottsanmälan (rikosilmoitus) kan göras per telefon eller personligen på polisstationen.
Du kan också göra brottsanmälan på internet om brottet i fråga är ringa och du inte behöver omedelbar hjälp av polisen.
Konvaljvägen 21
Tfn 0295 430291
Läs mer: Brott.
Kontaktuppgifterfinska _ svenska
Elektronisk polisanmälanfinska _ svenska _ engelska
Behöver du en jurist?
Östra Nylands rättshjälpsbyrå (Itä-Uudenmaan oikeusaputoimisto) betjänar invånarna i Vanda.
Pyrolavägen 37
Tfn 029 5660 160
Du kan också söka information om privata jurister på till exempel Finlands Juristförbunds (Suomen Asianajajaliitto) webbplats.
Läs mer: Behöver du en jurist?
linkkiÖstra Nylands rättshjälpsbyrå:
Information om rättshjälpfinska _ svenska _ engelska
linkkiFinlands Advokatförbund:
Advokaterfinska _ svenska _ engelska
Våld
I nödsituationer ringer du nödnumret 112.
I krissituationer får man även hjälp vid Vanda stads social- och krisjour (sosiaali- ja kriisipäivystys), som har öppet dygnet runt.
Social- och krisjouren
Tfn (09) 8392 4005
linkkiNödcentralsverket:
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
Skyddshem
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta ett skyddshem (turvakoti).
Skyddshemmen har jourmottagning dygnet runt.
Skyddshemmet Mona (turvakoti Mona) är ett skyddshem avsett för invandrarkvinnor och deras barn.
Tfn 045 639 6274
linkkiTurvakoti Mona:
Skyddshemfinska
Du kan även gå till Vanda skyddshem (Vantaan turvakoti) eller huvudstadsregionens skyddshem (pääkaupunkiseudun turvakoti).
Puh. (09) 8392 0071
Skyddshemfinska _ engelska
Steniusvägen 20
Tfn (09) 4777 180
Hjälp till offer för familjevåldfinska
Hjälp för invandrarkvinnor
Föreningen Monika-Naiset liitto (Monika-Naiset Liitto) ger råd och stöd till invandrarkvinnor.
Föreningen har ett resurscenter (voimavarakeskus) i Vanda där man får stöd och råd.
Tfn (09) 839 35013
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Hjälp för män
Män som har utövat våld mot sina familjemedlemmar eller har själva blivit offer för våld i hemmet, kan få hjälp från Jussi-arbetet i Vanda (Vantaan Jussi-työ).
Hjälp för män att sluta med våldsamt beteendefinska
Miehen linja (Miehen linja) hjälper invandrarmän som har problem med våld.
Tfn (09) 276 62899
Hjälp för män för att sluta med våldsamt beteendefinska _ engelska
Hjälp för unga
Finlands Röda Kors De ungas skyddshus (Suomen Punaisen Ristin Nuorten turvatalo) ger stöd och hjälp i krissituationer för 12–19-åringar.
Skyddshuset har öppet kl. 17–10, telefonjouren betjänar dygnet runt.
Sjukhusgatan 3 (Räckhals gård)
Tfn (09) 871 4043
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Läs mer: Våld
Problem i äktenskap eller parförhållande
Par med barn under 13 år kan vid problem i äktenskap och parförhållande få hjälp vid familjerådgivningen (perheneuvola).
Kontaktuppgifterna hittar du på Vanda stads webbplats.
Familjerådgivningens tjänster är konfidentiella och avgiftsfria.
Vid akuta krissituationer inom familjen kan du kontakta social- och krisjouren (sosiaali- ja kriisipäivystys), som har öppet dygnet runt varje dag.
Social- och krisjouren
Tfn (09) 8392 4005
Vid problem i parförhållandet och familjen får man även hjälp av familjerådgivningen vid Vanda församlingar (Vantaan seurakunnan perheneuvonta).
Läs mer: Problem i äktenskap och parförhållande
linkkiVanda stad:
Familjerådgivningarfinska _ svenska
linkkiVanda kyrkliga samfällighet:
Familjerådgivningfinska _ engelska
Barnrådgivningsbyråerna (lastenneuvola) och familjerådgivningsbyråerna (perheneuvola) ger råd i frågor som rör barns hälsa, uppväxt och utveckling.
Vid problem hos barn i skolåldern får man hjälp hos skolhälsovårdarna (kouluterveydenhoitaja), skolkuratorerna (koulukuraattori) och socialhandledarna (sosiaaliohjaaja).
Mer information hittar du på Vanda stads webbplats.
Läs mer: Barns och ungas problem
linkkiVanda stad:
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad:
Familjerådgivningarfinska _ svenska
linkkiVanda stad:
Information om tjänster för barn, ungdomar och familjerfinska _ svenska _ engelska
I skolan får de unga hjälp av skol- och studenthälsovårdarna (koulu- ja opiskeluterveydenhoitajat), skolkuratorerna (koulukuraattorit) och skolpsykologerna (koulupsykologit).
linkkiVanda stad:
Information om skolhälsovårdenfinska _ svenska _ engelska
linkkiVanda stad:
Skolkuratorerfinska _ svenska
linkkiVanda stad:
Skolpsykologerfinska _ svenska
Nuppi
13–21-åriga barn och ungdomar samt deras familjer kan få hjälp hos ungdomscentralen (nuortenkeskus).
På Nuppi kan du till exempel få hjälp med mentala problem och missbruksproblem.
Hjälp för ungafinska _ svenska _ engelska
Om du är under 30 år, kan du få råd och handledning via tjänsten Navigatorn.
Personalen vid Navigatorn hjälper dig om du inte har något arbete eller en studieplats.
Du kan även be om råd gällande andra saker, till exempel boende och ekonomi.
De ungas skyddshus
Finlands Röda Kors De ungas skyddshus (Suomen Punaisen Ristin Nuorten turvatalo) ger stöd och hjälp i krissituationer för 12–19-åringar.
Skyddshuset har öppet kl. 17–10, telefonjouren betjänar dygnet runt.
Sjukhusgatan 3
Tfn (09) 871 4043
Läs mer: Barns och ungas problem
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Vägledning och stöd för ungafinska _ svenska
Socialrådgivningen (sosiaalineuvonta) ger information om utkomststöd (toimeentulotuki) och andra bidrag om du har ekonomiska problem.
Tfn (09) 83 911.
linkkiVanda stad:
Socialrådgivningenfinska _ svenska _ engelska
Utkomststöd
Utkomststödet (toimeentulotuki) är avsett som en sista utväg då du inte har några andra inkomster eller medel, eller om dina inkomster är mycket låga.
Utkomststöd kan du få om du inte lyckas få tillräckliga inkomster genom eget arbete, andras omsorg eller på något annat sätt.
Du kan be om råd gällande ansökan om utkomststöd via den centraliserade telefontjänsten tfn (09) 8392 1119.
linkkiVanda stad:
Information om utkomststödfinska _ svenska _ engelska
Ekonomi- och skuldrådgivning
Om du inte kan betala dina räkningar eller skulder då de förfaller, ska du kontakta skuldrådgivningen (velkaneuvonta).
Tfn (09) 8392 2120.
linkkiVanda ekonomi- och skuldrådgivning:
Ekonomi- och skuldrådgivningfinska _ svenska _ engelska
Social kreditgivning
Om du har låga inkomster och är medellös samt har svårt att få lån, kan du ansöka om lån via den sociala kreditgivningen (sosiaalinen luototus).
Telefonnumret till kundrådgivningen och tidsbokningen är (09) 8392 0173.
linkkiVanda stad:
Information om social kreditgivningfinska _ svenska _ engelska
Missbruksproblem och spelberoende
Itä-Vantaan A-klinikka
Konvaljvägen 20 C vån.
tfn (09) 8392 3415
Länsi-Vantaan A-klinikka
tfn (09) 8393 5534
H-klinikka
Eldstadsvägen 7 B, vån.
Tfn (09) 839 21064
H-kliniken har också verksamhetsställen på Dickursby och Myrbacka hälsostationer.
Om du har spelproblem kan du söka hjälp vid Spelkliniken (Peliklinikka), som finns i centrala Helsingfors.
Peliklinikka
tfn 040 152 3918.
Ungdomscentralen Nuppi (nuortenkeskus Nuppi) hjälper ungdomar med missbruksproblem, Internetberoende eller spelberoende.
Nuppi ger också stöd till ungdomar som oroar sig för rusmedelsbruket hos någon närstående person.
Läs mer: Missbruksproblem.
linkkiVanda stad:
Hjälp med missbruksproblemfinska _ svenska _ engelska
linkkiVanda stad:
Information om vård av drogproblemfinska _ svenska _ engelska
Hjälp med penningspelproblemfinska
Hjälp för ungafinska _ svenska _ engelska
Dödsfall
I Vanda finns fyra begravningsplatser som tillhör de evangelisk-lutherska församlingarna.
I Furumo i Vanda finns dessutom Vandas och Helsingfors gemensamma begravningsplats för avlidna personer som inte har varit medlemmar i något religionssamfund.
Information om begravning får du på Vanda församlingars gravkontor (Vantaan seurakuntien hautaustoimisto) och vid privata begravningsbyråer (hautaustoimisto).
Vanda församlingars gravkontor
Prästgårdsgränden 5
Tfn (09) 8306 220
Om din närstående avlider plötsligt, kan du få hjälp med att återhämta dig från den chockartade upplevelsen och stöd i att klara dig efter förlusten av Vandas social- och krisjour (sosiaali- ja kriisipäivystys).
Jouren har öppet varje dag dygnet runt.
Social- och krisjouren
Tfn (09) 8392 4005
Läs mer: Död
linkkiVanda kyrkliga samfällighet:
Begravningsplatserfinska
linkkiHelsingfors kyrkliga samfällighet:
Konfessionslös begravningsplatsfinska
linkkiFinlands Begravningbyråers Förbund:
Begravningsbyråerfinska
När en närstående har avliditfinska _ svenska _ engelska
linkkiVanda stad:
Social- och krisjourenfinska _ svenska _ engelska
Problem med uppehållstillståndet
Brott
Behöver du en jurist?
Våld
Missbruksproblem och spelberoende
Dödsfall
Om du behöver brådskande hjälp av polisen, brandkåren eller ambulansen, ring nödnumret 112.
Du får ringa nödnumret endast i brådskande nödfall där liv, hälsa, egendom eller miljö är i fara.
Om du drabbas av en akut krissituation, såsom att en närstående avlider eller på grund av familjevåld, kan du kontakta social- och krisjouren (sosiaali- ja kriisipäivystys).
Du kan också söka hjälp för en familjemedlem eller en vän.
Social- och krisjouren har öppet dygnet runt varje dag.
Social- och krisjouren
Tfn (09) 8392 4005
linkkiNödcentralsverket:
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
linkkiVanda stad:
Social- och krisjourenfinska _ svenska _ engelska
Problem med uppehållstillståndet
Om du har problem eller oklarheter med uppehållstillståndet, kontakta Migrationsverket.
Du kan även fråga om råd på rådgivningstjänsterna för invandrare.
Information om tjänsterna finns på sidan Som invandrare i Vanda.
Migrationsverkets närmaste tjänsteställe finns i Helsingfors:
Göksgränd 3A
Läs mer: Problem med uppehållstillståndet
Olika tillståndfinska _ svenska _ engelska
Hälsovård för papperslösa
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärhälsovård.
Tjänsterna vid Global Clinic är avgiftsfria för kunderna.
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter.
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
Telefonnumret till Global Clinic i Helsingfors är 044 977 4547.
Samtalet besvaras av en sjukskötare eller en läkare.
E-postadressen är globalclinic.finland(at)gmail.com.
Läs mer: Problem med uppehållstillstånd
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Brott
Brottsanmälan (rikosilmoitus) kan göras per telefon eller personligen på polisstationen.
Du kan också göra brottsanmälan på internet om brottet i fråga är ringa och du inte behöver omedelbar hjälp av polisen.
Konvaljvägen 21
Tfn 0295 430291
Läs mer: Brott.
Kontaktuppgifterfinska _ svenska
Elektronisk polisanmälanfinska _ svenska _ engelska
Behöver du en jurist?
Östra Nylands rättshjälpsbyrå (Itä-Uudenmaan oikeusaputoimisto) betjänar invånarna i Vanda.
Pyrolavägen 37
Tfn 029 5660 160
Du kan också söka information om privata jurister på till exempel Finlands Juristförbunds (Suomen Asianajajaliitto) webbplats.
Läs mer: Behöver du en jurist?
linkkiÖstra Nylands rättshjälpsbyrå:
Information om rättshjälpfinska _ svenska _ engelska
linkkiFinlands Advokatförbund:
Advokaterfinska _ svenska _ engelska
Våld
I nödsituationer ringer du nödnumret 112.
I krissituationer får man även hjälp vid Vanda stads social- och krisjour (sosiaali- ja kriisipäivystys), som har öppet dygnet runt.
Social- och krisjouren
Tfn (09) 8392 4005
linkkiNödcentralsverket:
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
Skyddshem
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta ett skyddshem (turvakoti).
Skyddshemmen har jourmottagning dygnet runt.
Skyddshemmet Mona (turvakoti Mona) är ett skyddshem avsett för invandrarkvinnor och deras barn.
Tfn 045 639 6274
linkkiTurvakoti Mona:
Skyddshemfinska
Du kan även gå till Vanda skyddshem (Vantaan turvakoti) eller huvudstadsregionens skyddshem (pääkaupunkiseudun turvakoti).
Puh. (09) 8392 0071
Skyddshemfinska _ engelska
Steniusvägen 20
Tfn (09) 4777 180
Hjälp till offer för familjevåldfinska
Hjälp för invandrarkvinnor
Föreningen Monika-Naiset liitto (Monika-Naiset Liitto) ger råd och stöd till invandrarkvinnor.
Föreningen har ett resurscenter (voimavarakeskus) i Vanda där man får stöd och råd.
Tfn (09) 839 35013
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Hjälp för män
Män som har utövat våld mot sina familjemedlemmar eller har själva blivit offer för våld i hemmet, kan få hjälp från Jussi-arbetet i Vanda (Vantaan Jussi-työ).
Hjälp för män att sluta med våldsamt beteendefinska
Miehen linja (Miehen linja) hjälper invandrarmän som har problem med våld.
Tfn (09) 276 62899
Hjälp för män för att sluta med våldsamt beteendefinska _ engelska
Hjälp för unga
Finlands Röda Kors De ungas skyddshus (Suomen Punaisen Ristin Nuorten turvatalo) ger stöd och hjälp i krissituationer för 12–19-åringar.
Skyddshuset har öppet kl. 17–10, telefonjouren betjänar dygnet runt.
Sjukhusgatan 3 (Räckhals gård)
Tfn (09) 871 4043
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Läs mer: Våld
Problem i äktenskap eller parförhållande
Par med barn under 13 år kan vid problem i äktenskap och parförhållande få hjälp vid familjerådgivningen (perheneuvola).
Kontaktuppgifterna hittar du på Vanda stads webbplats.
Familjerådgivningens tjänster är konfidentiella och avgiftsfria.
Vid akuta krissituationer inom familjen kan du kontakta social- och krisjouren (sosiaali- ja kriisipäivystys), som har öppet dygnet runt varje dag.
Social- och krisjouren
Tfn (09) 8392 4005
Vid problem i parförhållandet och familjen får man även hjälp av familjerådgivningen vid Vanda församlingar (Vantaan seurakunnan perheneuvonta).
Läs mer: Problem i äktenskap och parförhållande
linkkiVanda stad:
Familjerådgivningarfinska _ svenska
linkkiVanda kyrkliga samfällighet:
Familjerådgivningfinska _ engelska
Barnrådgivningsbyråerna (lastenneuvola) och familjerådgivningsbyråerna (perheneuvola) ger råd i frågor som rör barns hälsa, uppväxt och utveckling.
Vid problem hos barn i skolåldern får man hjälp hos skolhälsovårdarna (kouluterveydenhoitaja), skolkuratorerna (koulukuraattori) och socialhandledarna (sosiaaliohjaaja).
Mer information hittar du på Vanda stads webbplats.
Läs mer: Barns och ungas problem
linkkiVanda stad:
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad:
Familjerådgivningarfinska _ svenska
linkkiVanda stad:
Information om tjänster för barn, ungdomar och familjerfinska _ svenska _ engelska
I skolan får de unga hjälp av skol- och studenthälsovårdarna (koulu- ja opiskeluterveydenhoitajat), skolkuratorerna (koulukuraattorit) och skolpsykologerna (koulupsykologit).
linkkiVanda stad:
Information om skolhälsovårdenfinska _ svenska _ engelska
linkkiVanda stad:
Skolkuratorerfinska _ svenska
linkkiVanda stad:
Skolpsykologerfinska _ svenska
Nuppi
13–21-åriga barn och ungdomar samt deras familjer kan få hjälp hos ungdomscentralen (nuortenkeskus).
På Nuppi kan du till exempel få hjälp med mentala problem och missbruksproblem.
Hjälp för ungafinska _ svenska _ engelska
Om du är under 30 år, kan du få råd och handledning via tjänsten Navigatorn.
Personalen vid Navigatorn hjälper dig om du inte har något arbete eller en studieplats.
Du kan även be om råd gällande andra saker, till exempel boende och ekonomi.
De ungas skyddshus
Finlands Röda Kors De ungas skyddshus (Suomen Punaisen Ristin Nuorten turvatalo) ger stöd och hjälp i krissituationer för 12–19-åringar.
Skyddshuset har öppet kl. 17–10, telefonjouren betjänar dygnet runt.
Sjukhusgatan 3
Tfn (09) 871 4043
Läs mer: Barns och ungas problem
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Vägledning och stöd för ungafinska _ svenska
Socialrådgivningen (sosiaalineuvonta) ger information om utkomststöd (toimeentulotuki) och andra bidrag om du har ekonomiska problem.
Tfn (09) 83 911.
linkkiVanda stad:
Socialrådgivningenfinska _ svenska _ engelska
Utkomststöd
Utkomststödet (toimeentulotuki) är avsett som en sista utväg då du inte har några andra inkomster eller medel, eller om dina inkomster är mycket låga.
Utkomststöd kan du få om du inte lyckas få tillräckliga inkomster genom eget arbete, andras omsorg eller på något annat sätt.
Du kan be om råd gällande ansökan om utkomststöd via den centraliserade telefontjänsten tfn (09) 8392 1119.
linkkiVanda stad:
Information om utkomststödfinska _ svenska _ engelska
Ekonomi- och skuldrådgivning
Om du inte kan betala dina räkningar eller skulder då de förfaller, ska du kontakta skuldrådgivningen (velkaneuvonta).
Tfn 029 566 0175.
linkkiVanda ekonomi- och skuldrådgivning:
Ekonomi- och skuldrådgivningfinska _ svenska _ engelska
Social kreditgivning
Om du har låga inkomster och är medellös samt har svårt att få lån, kan du ansöka om lån via den sociala kreditgivningen (sosiaalinen luototus).
Telefonnumret till kundrådgivningen och tidsbokningen är (09) 8392 0173.
linkkiVanda stad:
Information om social kreditgivningfinska _ svenska _ engelska
Missbruksproblem och spelberoende
Itä-Vantaan A-klinikka
Konvaljvägen 20 C vån.
tfn (09) 8392 3415
Länsi-Vantaan A-klinikka
tfn (09) 8393 5534
H-klinikka
Eldstadsvägen 7 B, vån.
Tfn (09) 839 21064
H-kliniken har också verksamhetsställen på Dickursby och Myrbacka hälsostationer.
Om du har spelproblem kan du söka hjälp vid Spelkliniken (Peliklinikka), som finns i centrala Helsingfors.
Peliklinikka
tfn 040 152 3918.
Ungdomscentralen Nuppi (nuortenkeskus Nuppi) hjälper ungdomar med missbruksproblem, Internetberoende eller spelberoende.
Nuppi ger också stöd till ungdomar som oroar sig för rusmedelsbruket hos någon närstående person.
Läs mer: Missbruksproblem.
linkkiVanda stad:
Hjälp med missbruksproblemfinska _ svenska _ engelska
linkkiVanda stad:
Information om vård av drogproblemfinska _ svenska _ engelska
Hjälp med penningspelproblemfinska
Hjälp för ungafinska _ svenska _ engelska
Dödsfall
I Vanda finns fyra begravningsplatser som tillhör de evangelisk-lutherska församlingarna.
I Furumo i Vanda finns dessutom Vandas och Helsingfors gemensamma begravningsplats för avlidna personer som inte har varit medlemmar i något religionssamfund.
Information om begravning får du på Vanda församlingars gravkontor (Vantaan seurakuntien hautaustoimisto) och vid privata begravningsbyråer (hautaustoimisto).
Vanda församlingars gravkontor
Prästgårdsgränden 5
Tfn (09) 8306 220
Om din närstående avlider plötsligt, kan du få hjälp med att återhämta dig från den chockartade upplevelsen och stöd i att klara dig efter förlusten av Vandas social- och krisjour (sosiaali- ja kriisipäivystys).
Jouren har öppet varje dag dygnet runt.
Social- och krisjouren
Tfn (09) 8392 4005
Läs mer: Död
linkkiVanda kyrkliga samfällighet:
Begravningsplatserfinska
linkkiHelsingfors kyrkliga samfällighet:
Konfessionslös begravningsplatsfinska
linkkiFinlands Begravningbyråers Förbund:
Begravningsbyråerfinska
När en närstående har avliditfinska _ svenska _ engelska
linkkiVanda stad:
Social- och krisjourenfinska _ svenska _ engelska
Äktenskap
Skilsmässa
Barnets födelse
Vård av barn
Problem i familjen
Äktenskap
Före äktenskapet ska du skriftligt begära hindersprövning (avioliiton esteiden tutkiminen).
Hindersprövningen görs på magistraten (maistraatti).
Du kan begära hindersprövning på vilken magistrat som helst.
Mer information hittar du på magistratens webbplats.
Också borgerliga vigslar förrättas på magistraten.
Konvaljvägen 15, PB 112
01301 Vanda
Läs mer: Äktenskap.
Anhållan om prövning av hinder mot äktenskapfinska _ svenska
Ingående av äktenskapfinska _ svenska _ engelska
linkkiVanda församlingar:
Information om kyrklig vigselfinska _ svenska _ engelska
linkkiHelsingfors ortodoxa församling:
Information om ortodox vigselfinska _ ryska
Skilsmässa
Kvinnan eller mannen kan lämna in skilsmässoansökan i Vanda tingsrätts kansli.
Makarna kan ansöka om skilsmässa tillsammans eller också kan den ena maken göra det ensam.
Ansökan kan lämnas till tingsrättens kansli eller skickas dit per post, fax eller via e-post.
Tfn 029 56 45200
Läs mer: Skilsmässa.
linkkiVanda stad:
Information om skilsmässafinska _ engelska
Att ansöka om skilsmässafinska _ svenska _ engelska
Om du har barn och ska skilja dig tar du kontakt med barnatillsyningsmannen (lastenvalvoja) vid Vanda stad.
Socialväsendet bekräftar ett avtal om barnens boende, vårdnad, umgängesrätt och underhållsbidrag.
Barnatillsyningsmännen ger även råd till föräldrar som ska skiljas.
Kontaktuppgifterna till barnatillsyningsmannen hittar du på Vanda stads webbplats.
Läs mer:
Barn vid skilsmässa.
linkkiVanda stad:
Kontaktuppgifter till barnatillsyningsmännenfinska _ svenska _ engelska
Barnets födelse
Uppgifterna om barnets födelse skickas från sjukhuset till befolkningsdataregistret i Finland.
Du ska meddela barnets namn, modersmål och andra erforderliga uppgifter till magistraten (Maistraatti) med en separat blankett som skickas hem till dig.
Du kan läsa mer om registrering av barnets födelse, faderskapserkännande och vårdnaden om barnet på InfoFinlands sida: När ett barn föds i Finland.
Vård av barn
Dagvård
På InfoFinlands sida Utbildning i Vanda hittar du information om dagvård för barn i Vanda.
Hemvårdsstöd
Om du tar hand om ett under treårigt barn, kan du få hemvårdsstöd (kotihoidon tuki).
Du ansöker om hemvårdsstödet hos FPA.
Vanda stad betalar dessutom ett kommuntillägg till hemvårdsstödet för barn till de familjer som vårdar ett under 1 ½-årigt barn i hemmet.
Du behöver inte ansöka separat om stödet, utan FPA betalar ut Vandatillägget (Vantaa-lisä) med hemvårdsstödet.
Information om hemvårdsstödfinska _ svenska _ engelska
linkkiVanda stad:
Information om hemvårdsstödets kommuntilläggfinska _ svenska _ engelska
Öppna daghem och invånarparker
Öppna daghem (avoin päiväkoti) är avsedda för barn under skolåldern och de föräldrar och vårdare som tar hand om dem.
Invånarparker (asukaspuistot) är avsedda för barn i alla åldrar och deras föräldrar eller vårdare.
Små barn kan delta i verksamheten tillsammans med sin förälder eller vårdare.
Verksamheten i öppna daghem och invånarparker är kostnadsfri och du behöver inte anmäla dig på förhand.
I verksamheten ingår lek och ledda aktiviteter, till exempel musik, motion och utflykter.
linkkiVanda stad:
Parker för invånare och öppna daghemfinska _ svenska _ engelska
Klubbar
Vanda stad ordnar även klubbar (kerho) för 2,5–5-åriga barn som vårdas i hemmet.
Klubbarna är avgiftsfria.
I klubben lär sig barnet tala finska, fungera i en grupp och där kan barnet träffa andra barn.
Till klubben ansöker du om plats med samma ansökan om småbarnsfostran (varhaiskasvatushakemus), med vilken du även ansöker om dagvårdsplats.
linkkiVanda stad:
Klubbverksamhetfinska _ svenska _ engelska
Barnpassningsservice för barn
Om du vårdar ditt barn i hemmet och behöver tillfälligt en vårdplats för barnet, till exempel när du ska sköta ärenden, kan du kontakta barnpassningsservicen (hoitoapupalvelu).
Barnpassningen är avgiftsbelagd.
linkkiVanda stad:
Barnpassningsservice för barnfinska _ engelska
Tillfällig barnpassning
Om du behöver tillfällig barnpassning i hemmet, kan du kontakta Mannerheims Barnskyddsförbund eller Väestöliitto.
Den tillfälliga barnpassningshjälpen är avgiftsbelagd.
Läs mer: Vård av barnet
linkkiMannerheims barnskyddsförbund:
Barnvaktshjälpfinska _ engelska
linkkiVanda stad:
Hjälp i hemmet för barnfamiljer(pdf, 500 kb)finska _ engelska
Problem i familjen
Om du misstänker att ditt barn eller din ungdom behöver barnskyddets (lastensuojelu) hjälp, ska du kontakta en socialarbetare.
Tfn växeln 09 83 911
mån–fre kl. 8.15–16.00
Kvällar och helger
Social- och krisjouren
tfn 09 8392 4005
linkkiVanda stad:
Barnskyddsanmälanfinska _ engelska
På InfoFinlands sida Problematiska situationer i Vanda hittar du information om var någonstans i Vanda det finns hjälp att få till barns och ungas problem.
Information om barns och ungas problem finns även på InfoFinlands sidor Barns och ungas problem och Barnskydd.
På InfoFinlands sida Problem i äktenskap och parförhållande finns information om var man kan få hjälp med problem i parförhållanden.
Äktenskap
Skilsmässa
Barnets födelse
Vård av barn
Problem i familjen
Äldre människor
Äktenskap
Före äktenskapet ska du skriftligt begära hindersprövning (avioliiton esteiden tutkiminen).
Hindersprövningen görs på magistraten (maistraatti).
Du kan begära hindersprövning på vilken magistrat som helst.
Mer information hittar du på magistratens webbplats.
Också borgerliga vigslar förrättas på magistraten.
Konvaljvägen 15, PB 112
01301 Vanda
Läs mer: Äktenskap.
Anhållan om prövning av hinder mot äktenskapfinska _ svenska
Ingående av äktenskapfinska _ svenska _ engelska
linkkiVanda församlingar:
Information om kyrklig vigselfinska _ svenska _ engelska
linkkiHelsingfors ortodoxa församling:
Information om ortodox vigselfinska _ ryska
Skilsmässa
Kvinnan eller mannen kan lämna in skilsmässoansökan i Vanda tingsrätts kansli.
Makarna kan ansöka om skilsmässa tillsammans eller också kan den ena maken göra det ensam.
Ansökan kan lämnas till tingsrättens kansli eller skickas dit per post, fax eller via e-post.
Tfn 029 56 45200
Läs mer: Skilsmässa.
linkkiVanda stad:
Information om skilsmässafinska _ engelska
Att ansöka om skilsmässafinska _ svenska _ engelska
Om du har barn och ska skilja dig tar du kontakt med barnatillsyningsmannen (lastenvalvoja) vid Vanda stad.
Socialväsendet bekräftar ett avtal om barnens boende, vårdnad, umgängesrätt och underhållsbidrag.
Barnatillsyningsmännen ger även råd till föräldrar som ska skiljas.
Kontaktuppgifterna till barnatillsyningsmannen hittar du på Vanda stads webbplats.
Läs mer:
Barn vid skilsmässa.
linkkiVanda stad:
Kontaktuppgifter till barnatillsyningsmännenfinska _ svenska _ engelska
Barnets födelse
Uppgifterna om barnets födelse skickas från sjukhuset till befolkningsdataregistret i Finland.
Du ska meddela barnets namn, modersmål och andra erforderliga uppgifter till magistraten (Maistraatti) med en separat blankett som skickas hem till dig.
Du kan läsa mer om registrering av barnets födelse, faderskapserkännande och vårdnaden om barnet på InfoFinlands sida: När ett barn föds i Finland.
Vård av barn
Dagvård
På InfoFinlands sida Utbildning i Vanda hittar du information om dagvård för barn i Vanda.
Hemvårdsstöd
Om du tar hand om ett under treårigt barn, kan du få hemvårdsstöd (kotihoidon tuki).
Du ansöker om hemvårdsstödet hos FPA.
Vanda stad betalar dessutom ett kommuntillägg till hemvårdsstödet för barn till de familjer som vårdar ett under 1 ½-årigt barn i hemmet.
Du behöver inte ansöka separat om stödet, utan FPA betalar ut Vandatillägget (Vantaa-lisä) med hemvårdsstödet.
Information om hemvårdsstödfinska _ svenska _ engelska
linkkiVanda stad:
Information om hemvårdsstödets kommuntilläggfinska _ svenska _ engelska
Öppna daghem och invånarparker
Öppna daghem (avoin päiväkoti) är avsedda för barn under skolåldern och de föräldrar och vårdare som tar hand om dem.
Invånarparker (asukaspuistot) är avsedda för barn i alla åldrar och deras föräldrar eller vårdare.
Små barn kan delta i verksamheten tillsammans med sin förälder eller vårdare.
Verksamheten i öppna daghem och invånarparker är kostnadsfri och du behöver inte anmäla dig på förhand.
I verksamheten ingår lek och ledda aktiviteter, till exempel musik, motion och utflykter.
linkkiVanda stad:
Parker för invånare och öppna daghemfinska _ svenska _ engelska
Klubbar
Vanda stad ordnar även klubbar (kerho) för 2,5–5-åriga barn som vårdas i hemmet.
Klubbarna är avgiftsfria.
I klubben lär sig barnet tala finska, fungera i en grupp och där kan barnet träffa andra barn.
Till klubben ansöker du om plats med samma ansökan om småbarnsfostran (varhaiskasvatushakemus), med vilken du även ansöker om dagvårdsplats.
linkkiVanda stad:
Klubbverksamhetfinska _ svenska _ engelska
Barnpassningsservice för barn
Om du vårdar ditt barn i hemmet och behöver tillfälligt en vårdplats för barnet, till exempel när du ska sköta ärenden, kan du kontakta barnpassningsservicen (hoitoapupalvelu).
Barnpassningen är avgiftsbelagd.
linkkiVanda stad:
Barnpassningsservice för barnfinska _ engelska
Tillfällig barnpassning
Om du behöver tillfällig barnpassning i hemmet, kan du kontakta Mannerheims Barnskyddsförbund eller Väestöliitto.
Den tillfälliga barnpassningshjälpen är avgiftsbelagd.
Läs mer: Vård av barnet
linkkiMannerheims barnskyddsförbund:
Barnvaktshjälpfinska _ engelska
linkkiVanda stad:
Hjälp i hemmet för barnfamiljer(pdf, 500 kb)finska _ engelska
Problem i familjen
Om du misstänker att ditt barn eller din ungdom behöver barnskyddets (lastensuojelu) hjälp, ska du kontakta en socialarbetare.
Tfn växeln 09 83 911
mån–fre kl. 8.15–16.00
Kvällar och helger
Social- och krisjouren
tfn 09 8392 4005
linkkiVanda stad:
Barnskyddsanmälanfinska _ engelska
På InfoFinlands sida Problematiska situationer i Vanda hittar du information om var någonstans i Vanda det finns hjälp att få till barns och ungas problem.
Information om barns och ungas problem finns även på InfoFinlands sidor Barns och ungas problem och Barnskydd.
På InfoFinlands sida Problem i äktenskap och parförhållande finns information om var man kan få hjälp med problem i parförhållanden.
Äldre människor
I Vanda finns tjänster som är särskilt avsedda för äldre.
Du får information om dem vid seniorrådgivningen.
Seniorrådgivningen Tfn: 09 8392 4202
När du tar hand om en anhörig i hemmet
När en familjemedlem behöver kontinuerlig hjälp och vården är både bindande och krävande, finns det möjlighet att få stöd för närståendevård av kommunen.
Seniorrådgivningen bedömer behovet av anhörigvård för en äldre person.
Läs mer: Äldre människor.
linkkiVanda stad:
Seniorrådgivningenfinska _ svenska _ engelska
Äktenskap
Skilsmässa
Barnets födelse
Vård av barn
Problem i familjen
Äldre människor
Äktenskap
Före äktenskapet ska du skriftligt begära hindersprövning (avioliiton esteiden tutkiminen).
Hindersprövningen görs på magistraten (maistraatti).
Du kan begära hindersprövning på vilken magistrat som helst.
Mer information hittar du på magistratens webbplats.
Också borgerliga vigslar förrättas på magistraten.
Konvaljvägen 15, PB 112
01301 Vanda
Läs mer: Äktenskap.
Anhållan om prövning av hinder mot äktenskapfinska _ svenska _ engelska
Ingående av äktenskapfinska _ svenska _ engelska
linkkiVanda församlingar:
Information om kyrklig vigselfinska _ svenska _ engelska
linkkiHelsingfors ortodoxa församling:
Information om ortodox vigselfinska _ ryska
Skilsmässa
Kvinnan eller mannen kan lämna in skilsmässoansökan i Vanda tingsrätts kansli.
Makarna kan ansöka om skilsmässa tillsammans eller också kan den ena maken göra det ensam.
Ansökan kan lämnas till tingsrättens kansli eller skickas dit per post, fax eller via e-post.
Tfn 029 56 45200
Läs mer: Skilsmässa.
linkkiVanda stad:
Information om skilsmässafinska _ engelska
Att ansöka om skilsmässafinska _ svenska _ engelska
Om du har barn och ska skilja dig tar du kontakt med barnatillsyningsmannen (lastenvalvoja) vid Vanda stad.
Socialväsendet bekräftar ett avtal om barnens boende, vårdnad, umgängesrätt och underhållsbidrag.
Barnatillsyningsmännen ger även råd till föräldrar som ska skiljas.
Kontaktuppgifterna till barnatillsyningsmannen hittar du på Vanda stads webbplats.
Läs mer:
Barn vid skilsmässa.
linkkiVanda stad:
Kontaktuppgifter till barnatillsyningsmännenfinska _ svenska _ engelska
Barnets födelse
Uppgifterna om barnets födelse skickas från sjukhuset till befolkningsdataregistret i Finland.
Du ska meddela barnets namn, modersmål och andra erforderliga uppgifter till magistraten (Maistraatti) med en separat blankett som skickas hem till dig.
Du kan läsa mer om registrering av barnets födelse, faderskapserkännande och vårdnaden om barnet på InfoFinlands sida: När ett barn föds i Finland.
Vård av barn
Dagvård
På InfoFinlands sida Utbildning i Vanda hittar du information om dagvård för barn i Vanda.
Hemvårdsstöd
Om du tar hand om ett under treårigt barn, kan du få hemvårdsstöd (kotihoidon tuki).
Du ansöker om hemvårdsstödet hos FPA.
Vanda stad betalar dessutom ett kommuntillägg till hemvårdsstödet för barn till de familjer som vårdar ett under 1 ½-årigt barn i hemmet.
Du behöver inte ansöka separat om stödet, utan FPA betalar ut Vandatillägget (Vantaa-lisä) med hemvårdsstödet.
Information om hemvårdsstödfinska _ svenska _ engelska
linkkiVanda stad:
Information om hemvårdsstödets kommuntilläggfinska _ svenska _ engelska
Öppna daghem och invånarparker
Öppna daghem (avoin päiväkoti) är avsedda för barn under skolåldern och de föräldrar och vårdare som tar hand om dem.
Invånarparker (asukaspuistot) är avsedda för barn i alla åldrar och deras föräldrar eller vårdare.
Små barn kan delta i verksamheten tillsammans med sin förälder eller vårdare.
Verksamheten i öppna daghem och invånarparker är kostnadsfri och du behöver inte anmäla dig på förhand.
I verksamheten ingår lek och ledda aktiviteter, till exempel musik, motion och utflykter.
linkkiVanda stad:
Parker för invånare och öppna daghemfinska _ svenska _ engelska
Klubbar
Vanda stad ordnar även klubbar (kerho) för 2,5–5-åriga barn som vårdas i hemmet.
Klubbarna är avgiftsfria.
I klubben lär sig barnet tala finska, fungera i en grupp och där kan barnet träffa andra barn.
Till klubben ansöker du om plats med samma ansökan om småbarnsfostran (varhaiskasvatushakemus), med vilken du även ansöker om dagvårdsplats.
linkkiVanda stad:
Klubbverksamhetfinska _ svenska _ engelska
Barnpassningsservice för barn
Om du vårdar ditt barn i hemmet och behöver tillfälligt en vårdplats för barnet, till exempel när du ska sköta ärenden, kan du kontakta barnpassningsservicen (hoitoapupalvelu).
Barnpassningen är avgiftsbelagd.
linkkiVanda stad:
Barnpassningsservice för barnfinska _ engelska
Tillfällig barnpassning
Om du behöver tillfällig barnpassning i hemmet, kan du kontakta Mannerheims Barnskyddsförbund eller Väestöliitto.
Den tillfälliga barnpassningshjälpen är avgiftsbelagd.
Läs mer: Vård av barnet
linkkiMannerheims barnskyddsförbund:
Barnvaktshjälpfinska _ engelska
linkkiVanda stad:
Hjälp i hemmet för barnfamiljer(pdf, 500 kb)finska _ engelska
Problem i familjen
Om du misstänker att ditt barn eller din ungdom behöver barnskyddets (lastensuojelu) hjälp, ska du kontakta en socialarbetare.
Tfn växeln 09 83 911
mån–fre kl. 8.15–16.00
Kvällar och helger
Social- och krisjouren
tfn 09 8392 4005
linkkiVanda stad:
Barnskyddsanmälanfinska _ engelska
På InfoFinlands sida Problematiska situationer i Vanda hittar du information om var någonstans i Vanda det finns hjälp att få till barns och ungas problem.
Information om barns och ungas problem finns även på InfoFinlands sidor Barns och ungas problem och Barnskydd.
På InfoFinlands sida Problem i äktenskap och parförhållande finns information om var man kan få hjälp med problem i parförhållanden.
Äldre människor
I Vanda finns tjänster som är särskilt avsedda för äldre.
Du får information om dem vid seniorrådgivningen.
Seniorrådgivningen Tfn: 09 8392 4202
När du tar hand om en anhörig i hemmet
När en familjemedlem behöver kontinuerlig hjälp och vården är både bindande och krävande, finns det möjlighet att få stöd för närståendevård av kommunen.
Seniorrådgivningen bedömer behovet av anhörigvård för en äldre person.
Läs mer: Äldre människor.
linkkiVanda stad:
Seniorrådgivningenfinska _ svenska _ engelska
Hälsotjänster i Vanda
Privata hälsotjänster
Barns hälsa
Äldre människors hälsa
Tandvård
Mental hälsa
Sexuell hälsa
När du väntar barn
Handikappade
Hälsotjänsterna i Vanda
Om du behöver information om hälsotjänsterna, kan du ringa hälsorådgivningstelefonen: Tfn (09) 839 10023, mån-fre kl. 8–16.
Via tjänsten kan du också fråga om anvisningar för vård av sjukdomar.
Du kan tala finska, svenska eller engelska.
Läs mer: Hälsa.
linkkiVanda stad:
Information om hälsorådgivningfinska _ svenska _ engelska
Offentliga hälsovårdstjänster
Om du har din hemkommun i Vanda, kan du utnyttja de offentliga hälsovårdstjänsterna.
Offentliga hälsovårdstjänster tillhandahålls till exempel vid hälsostationer, tandkliniker, rådgivningsbyråer och sjukhus.
Om du insjuknar plötsligt eller om du råkar ut för en olycka, får du akut sjukvård även om din hemkommun inte är Vanda.
I Vanda finns sju hälsostationer (terveysasema) som tillhandahåller offentliga hälsovårdstjänster.
Hälsostationerna har öppet vardagar kl. 8.00–16.00.
Hälsostationerna når du genom att ringa till respektive hälsostations eget telefonnummer eller hälsorådgivningens telefonnummer (09) 839 10023 och väljer din hälsostation med hjälpa av knappsatsen.
Om du behöver akut vård samma dag, ska du ringa hälsostationen direkt då den öppnar.
Hälsostationernas adresser:
Håkansböle hälsostation, Galoppbrinken 4
Korso hälsostation, Fjällrävsstigen 6
Västerkulla hälsostation, Kägelgränden 1
Myrbacka hälsostation, Jönsasvägen 4
Dickursby hälsostation, Konvaljvägen 11
Närmare information hittar du på hälsostationernas egna webbplatser.
linkkiVanda stad:
Hälsostationernafinska _ svenska _ engelska
Privata hälsotjänster
I Vanda finns flera läkarstationer som erbjuder privata hälsovårdstjänster.
Du kan gå till en privat läkarstation även om du inte har rätt att använda den offentliga hälsovårdens tjänster i Finland.
På en privat läkarstation måste du betala samtliga kostnader själv.
I vissa fall ersätter Kela en liten del av kostnaderna för privat sjukvård.
Privat läkarstationfinska _ svenska _ engelska
Privat läkarstationfinska _ svenska _ engelska _ ryska
Privat läkarstationfinska _ svenska _ engelska
linkkiAava:
Privat läkarstationfinska _ svenska _ engelska
Läkemedel
Information om köp av läkemedel hittar du på InfoFinlands sida Läkemedel.
linkkiApotekareförbundet:
Apotekens kontaktuppgifterfinska
Hälsovård för papperslösa
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärhälsovård.
Tjänsterna vid Global Clinic är avgiftsfria för kunderna.
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter.
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
Telefonnumret till Helsingfors Global Clinicin är 044 948 1698.
En sjuksköterska eller läkare svarar i telefonen.
Läs mer: Hälsovårdstjänster i Finland.
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
På kvällar, helger och storhelger är hälsostationerna stängda.
Då vårdas akuta sjukfall och olycksfall på jourmottagningen (päivystys).
Jourmottagningen är öppen alla dagar dygnet runt
I Vanda finns jourmottagningen på Pejas sjukhus (Peijaksen sairaala).
Adress:
Sjukhusgatan 1
Tfn 116 117
Om du blir akut sjuk, kan du även besöka någon annan jourmottagning i huvudstadsregionen.
Mer information om jourmottagningarna hittar du på Vanda stads webbplats om hälsovårdstjänster.
I nödsituationer ringer du det allmänna nödnumret 112.
Läs mer: Hälsovårdstjänster i Finland.
linkkiVanda stad:
Jourmottagningarfinska _ svenska _ engelska
Barns hälsa
I hälsovården av barn under skolåldern får man hjälp av rådgivningsbyråerna (neuvola).
Där kan du fråga om råd och få stöd i föräldraskapet och fostran av barn.
På rådgivningsbyrån följs barnets hälsa, tillväxt och utveckling upp och där ges även vaccinationerna.
Kontaktuppgifterna till rådgivningsbyråerna hittar du på Vanda webbplats.
Via rådgivningsbyråernas telefontjänst kan du boka tid på rådgivningsbyrån och fråga hälsovårdaren om råd beträffande graviditet och barns hälsa.
Numret till telefontjänsten är (09) 8392 5900.
Den är öppen mån-tors kl. 8–15 och fre kl. 8–13.
Skolhälsovården har hand om skolbarns hälsa.
Mer information hittar du på Vanda stads webbplats.
Om ett barn blir akut sjukt, ska du ta kontakt med hälsostationen eller jourmottagningen.
I nödsituationer ringer du det allmänna nödnumret 112.
Läs mer: Barns hälsa.
linkkiVanda stad:
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad:
Tidsbokning och rådgivningfinska _ svenska _ engelska
linkkiVanda stad:
Information om skolhälsovårdenfinska _ svenska _ engelska
linkkiVanda stad:
Hälsostationernafinska _ svenska _ engelska
linkkiVanda stad:
Jourmottagningarfinska _ svenska _ engelska
Äldre människors hälsa
Äldre människor använder samma hälsovårdstjänster som alla andra.
Dessutom finns det i Vanda särskilda tjänster för äldre som du får information om via seniorrådgivningen (seniorineuvonta).
Tfn: (09) 8392 4202
Mer information om tjänsterna för äldre hittar du på Vanda stads webbplats.
Läs mer: Äldre människors hälsa och Äldre människor.
linkkiVanda stad:
Seniorrådgivningenfinska _ svenska _ engelska
linkkiVanda stad:
Information om tjänster för äldrefinska _ svenska _ engelska
linkkiVanda stad:
Serviceguide för seniorer(pdf, 1 MB)finska
När du tar hand om en anhörig i hemmet
När en familjemedlem behöver kontinuerlig hjälp och vården är både bindande och krävande, finns det möjlighet att få stöd för närståendevård av kommunen.
Behovet av närståendevård bedöms inom seniorrådgivningen.
Tfn: (09) 8392 4202
Behovet av närståendevård för personer under 65 år bedöms inom handikapprådgivningen.
Tfn: (09) 8392 4682
linkkiVanda stad:
Stöd för närståendevårdfinska _ svenska
Tandvård
Offentlig tandvård
Tidsbokningsnumret till Vanda tandvård (hammashoito) är (09) 8393 5300.
Tidsbokningen kan du ringa:
Mån-tors 7.30–15
Fredagar och storhelgsaftnar 7.30–14.
Om ditt ärende inte är brådskande, ring efter kl. 10.00.
Om tjänsten är hårt belastad, kan du lämna ett meddelande om att bli uppringd vid ett senare tillfälle.
Om du behöver akut tandvård på en vardag, ska du ringa tidsbokningen så fort den öppnar.
linkkiVanda stad:
Information om tandvårdenfinska _ svenska _ engelska
linkkiVanda stad:
Tandklinikerfinska _ svenska
Tandvårdens jourmottagning
Under kvällar och veckoslut finns tandvårdsjouren (hammashoidon päivystys) vid Haartmanska sjukhuset i Helsingfors.
Tfn (09) 310 49999.
Tandvårdens nattjour (hammashoidon yöpäivystys) finns på Tölö sjukhus olycksfallsstation.
Tölö sjukhus olycksfallsstation, Oral och käkkirurgisk jourmottagning
Tfn 040 621 5699
Tandvårdens jourmottagning kvällar och veckoslutfinska _ svenska _ engelska
Barns tandvård
Om tandvården för barn under skolåldern får du information på barnrådgivningen (lastenneuvola) och vid tandklinikerna (hammashoitola).
Barn under 17 år kallas till tandkliniken för undersökning med cirka två års mellanrum.
linkkiVanda stad:
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad:
Information om tandvården för skolbarnfinska
Privata tandvårdstjänster
I Vanda finns också privata tandläkare.
Om du inte har rätt att använda de offentliga hälsovårdstjänsterna, kan du söka dig till en privat tandläkare.
Hos en privat tandläkare måste du betala samtliga kostnader själv.
I vissa fall ersätter Kela en liten del av kostnaderna för privat tandvård.
Läs mer: Tandvård.
Sök tandläkarefinska
Mental hälsa
Om du behöver psykisk hjälp eller stöd, ska du kontakta din hälsostation (terveysasema).
På hälsostationen behandlas de vanligaste psykiska problemen.
Från hälsostationen kan du remitteras vidare exempelvis till depressionsskötare.
Om hälsostationen inte har öppet och situationen är akut, ska du kontakta samjouren vid Pejas sjukhus (Peijaksen sairaalan yhteispäivystys).
Sjukhusgatan 1
Tfn (09) 4716 7060
Om du behöver omedelbar krishjälp, kan du också ta kontakt med social- och krisjouren.
Den har öppet dygnet runt.
Social- och krisjouren
Tfn (09) 8392 4005
Läs mer: Mental hälsa.
linkkiVanda stad:
Information om mentalvårdstjänsternafinska _ svenska _ engelska
linkkiVanda stad:
Hälsostationernafinska _ svenska _ engelska
linkkiVanda stad:
Jourmottagningarfinska _ svenska _ engelska
linkkiVanda stad:
Social- och krisjourenfinska _ svenska _ engelska
Sexuell hälsa
Om du vill har information om graviditetsprevention, abort, sexuell hälsa och könssjukdomar, kan du kontakta preventivmedels- och familjeplaneringsrådgivningen (ehkäisy- ja perhesuunnitteluneuvola).
Preventivmedels- och familjeplaneringsrådgivningarna betjänar kvinnor och män i alla åldrar.
Du måste beställa tid vid rådgivningarna.
Besöken är avgiftsfria för kunderna.
Information om kontaktuppgifter finns på Vanda stads webbplats.
Boka en tid hos preventivmedelsrådgivningens läkare eller hälsovårdare om du behöver preventivmedel (raskauden ehkäisy) eller om du överväger abort (abortti).
Boka en tid hos hälsostationens allmänläkare om du till exempel har problem med blödningar eller smärtor i underlivet.
Vid hälsostationerna vårdas även könssjukdomar (sukupuolitauti).
Vandabor kan även besöka polikliniken för könssjukdomar i Helsingfors.
linkkiVanda stad:
Rådgivningarna för familjeplaneringfinska _ svenska.
linkkiVanda stad:
Hälsostationernafinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Polikliniken för könssjukdomarfinska _ svenska _ engelska
När du väntar barn
Vid mödrarådgivningen (äitiysneuvola) följs moderns, fostrets och hela familjens hälsotillstånd under graviditeten.
Kontakta rådgivningsbyrån (neuvola) när du upptäcker att du är gravid.
Rådgivningarnas telefontjänst
mån-tors kl. 8–15 och fre kl. 8–13
Via rådgivningsbyråernas telefontjänst kan du boka tid på rådgivningsbyrån och fråga hälsovårdaren om råd beträffande graviditet och förlossning.
Mer information om graviditet och förlossning hittar du på Vanda stads mödra- och barnrådgivning på Internet (Nettineuvola).
Läs mer: När du väntar barn.
linkkiVanda stad:
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad:
Rådgivningarna för familjeplaneringfinska _ svenska
linkkiVanda stad:
Förlossningen
Läs mer: Förlossning.
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Förlossningfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Handikappade
Du kan få tjänster för handikappade (vammaispalvelut) om du eller en närstående till dig har en invaliditet eller en sjukdom som orsakar långvariga, betydande svårigheter att klara sig hemma och i livet utanför hemmet.
Tjänster för handikappade är till exempel personlig assistans, serviceboende, färdtjänst och ombyggnadsarbeten i bostaden.
Ta kontakt med handikapprådgivningen som utreder ditt behov av stöd, handledning och tjänster utifrån din situation.
Mån.-fre. kl. 9–15
Tfn: (09) 8392 4682
Läs mer: Handikappade personer.
linkkiVanda stad:
Information om handikapptjänsternafinska _ svenska _ engelska
Hälsotjänster i Vanda
Barns hälsa
Tandvård
Mental hälsa
Sexuell hälsa och prevention
Graviditet och förlossning
Handikappade
Hälsotjänsterna i Vanda
Det allmänna nödnumret är 112.
Ring nödnumret endast om det handlar om ett nödfall, till exempel en akut sjukdomsattack.
Om din hemkommun är Vanda kan du använda kommunens offentliga hälsovårdstjänster.
Offentliga hälsovårdstjänster tillhandahålls till exempel vid hälsostationer, tandkliniker, rådgivningsbyråer och sjukhus.
Om du insjuknar akut eller råkar ut för en olycka får du akut sjukvård även om din hemkommun inte är Vanda.
Om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna, kan du boka tid på en privat läkarstation.
Läs mer: Hälsovårdstjänster i Finland.
Offentliga hälsovårdstjänster
Telefonnumret till den gemensamma telefontjänsten för hälsostationerna i Vanda är 09 839 50 000.
Du kan ringa detta nummer om du behöver rådgivning i behandlingen av en sjukdom eller vill boka eller avboka en läkartid.
Tjänsten har öppet måndag till fredag kl. 8–16.
I Vanda finns sju hälsostationer som tillhandahåller offentliga hälsovårdstjänster.
På hälsostationerna finns läkarens, sjukskötarens och hälsovårdarens mottagningar.
Om du insjuknar akut kan du gå direkt till vilken som helst hälsostation.
Det är bäst att gå till hälsostationen direkt på morgonen.
Hälsostationerna har öppet vardagar kl. 8.00–16.00.
linkkiVanda stad:
Information om hälsorådgivningfinska _ svenska _ engelska
linkkiVanda stad:
Hälsostationernafinska _ svenska _ engelska
Privata hälsotjänster
I Vanda finns flera läkarstationer som erbjuder privata hälsovårdstjänster.
Du kan gå till en privat läkarstation även om du inte har rätt att använda den offentliga hälsovårdens tjänster i Finland.
På en privat läkarstation måste du betala samtliga kostnader själv.
I vissa fall ersätter Kela en liten del av kostnaderna för privat sjukvård.
Läs mer: Hälsovårdstjänster i Finland.
Privat läkarstationfinska _ svenska _ engelska
Privat läkarstationfinska _ svenska _ engelska _ ryska
Privat läkarstationfinska _ svenska _ engelska
linkkiAava:
Privat läkarstationfinska _ svenska _ engelska
Läkemedel
Information om köp av läkemedel hittar du på InfoFinlands sida Läkemedel.
linkkiApotekareförbundet:
Apotekens kontaktuppgifterfinska
Hälsovård för papperslösa
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärhälsovård.
Tjänsterna vid Global Clinic är avgiftsfria för kunderna.
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter.
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
Telefonnumret till Helsingfors Global Clinicin är 044 948 1698.
En sjuksköterska eller läkare svarar i telefonen.
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
På kvällar, helger och storhelger är hälsostationerna stängda.
Om du insjuknar akut eller råkar ut för en olycka och inte kan vänta tills hälsostationen öppnar, kontakta jourmottagningen.
I Vanda finns jourmottagningen på Pejas sjukhus (Peijaksen sairaala).
Adress:
Sjukhusgatan 1
Tfn 116 117
Om du blir akut sjuk, kan du även besöka någon annan jourmottagning i huvudstadsregionen.
Mer information om jourmottagningarna hittar du på Vanda stads webbplats om hälsovårdstjänster.
linkkiVanda stad:
Jourmottagningarfinska _ svenska _ engelska
Barns hälsa
I hälsovården av barn under skolåldern får man hjälp av rådgivningsbyråerna (neuvola).
Telefonnumret till rådgivningsbyråerna i Vanda är 09 8392 5900.
Du kan boka en tid på rådgivningen eller fråga om råd om du har frågor kring barnets hälsa.
Skolhälsovården har hand om skolbarns hälsa.
Mer information hittar du på Vanda stads webbplats.
Om ett barn insjuknar akut, ska du kontakta hälsostationen.
Hälsostationerna har öppet måndag till fredag kl. 8–16.
När hälsostationen har stängt ska du kontakta jourmottagningen vid Barnsjukhuset.
Jourmottagningen tar endast hand om barn med brådskande hjälpbehov.
Telefonnumret till jourmottagningen är 116 117.
Adress:
Barnsjukhuset
Stenbäcksgatan 9
Du kan även ta barnet till en privat läkarstation.
I Vanda finns många privata läkarstationer som även tar hand om barn.
Läs mer: Barns hälsa.
linkkiVanda stad:
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad:
Tidsbokning och rådgivningfinska _ svenska _ engelska
linkkiVanda stad:
Information om skolhälsovårdenfinska _ svenska _ engelska
linkkiVanda stad:
Hälsostationernafinska _ svenska _ engelska
linkkiVanda stad:
Jourmottagningarfinska _ svenska _ engelska
Tandvård
Offentlig tandvård
Tidsbokningsnumret till Vanda tandvård (hammashoito) är (09) 8393 5300.
Om du inte behöver brådskande tandvård, ring efter kl. 10.00.
Om du behöver brådskande tandvård, ska du ringa tidsbokningen så fort den öppnar kl. 7.30.
Mottagningen för brådskande vård finns vid Dickursby hälsostation måndag till fredag kl. 8–14.
linkkiVanda stad:
Information om tandvårdenfinska _ svenska _ engelska
linkkiVanda stad:
Tandklinikerfinska _ svenska
Tandvårdens jourmottagning
Under kvällar och veckoslut finns tandvårdsjouren (hammashoidon päivystys) vid Haartmanska sjukhuset i Helsingfors.
Telefonnumret är 09 471 71110.
Tidsbokningen har öppet vardagar kl. 14–21 och på veckoslut kl. 8–21.
Tandvårdens nattjour (hammashoidon yöpäivystys) finns på Tölö sjukhus olycksfallsstation.
Tölö sjukhus olycksfallsstation, Oral och käkkirurgisk jourmottagning
Tfn 040 621 5699
Tandvårdens jourmottagning kvällar och veckoslutfinska _ svenska _ engelska
Barns tandvård
Om tandvården för barn under skolåldern får du information på barnrådgivningen (lastenneuvola) och vid tandklinikerna (hammashoitola).
Barn under 17 år kallas till tandkliniken för undersökning med cirka två års mellanrum.
linkkiVanda stad:
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad:
Information om tandvården för skolbarnfinska
Privata tandvårdstjänster
I Vanda finns också privata tandläkare.
Om du inte har rätt att använda de offentliga hälsovårdstjänsterna, kan du söka dig till en privat tandläkare.
Hos en privat tandläkare måste du betala samtliga kostnader själv.
I vissa fall ersätter Kela en liten del av kostnaderna för privat tandvård.
Läs mer: Tandvård.
Sök tandläkarefinska
Mental hälsa
Om du behöver psykisk hjälp eller stöd, ska du kontakta din hälsostation (terveysasema).
På hälsostationen behandlas de vanligaste psykiska problemen.
Från hälsostationen kan du remitteras vidare exempelvis till depressionsskötare.
Om hälsostationen inte har öppet och situationen är akut, ska du kontakta samjouren vid Pejas sjukhus (Peijaksen sairaalan yhteispäivystys).
Sjukhusgatan 1
Tfn 116 117
Om du behöver omedelbar krishjälp, kan du också ta kontakt med social- och krisjouren.
Den har öppet dygnet runt.
Social- och krisjouren
Tfn (09) 8392 4005
Läs mer: Mental hälsa.
linkkiVanda stad:
Information om mentalvårdstjänsternafinska _ svenska _ engelska
linkkiVanda stad:
Hälsostationernafinska _ svenska _ engelska
linkkiVanda stad:
Jourmottagningarfinska _ svenska _ engelska
linkkiVanda stad:
Social- och krisjourenfinska _ svenska _ engelska
Sexuell hälsa och prevention
Om du behöver preventivmedel eller abort eller misstänker att du har en könssjukdom, kan du kontakta preventivmedels- och familjeplaneringsrådgivningen.
Du kan boka tid per telefon.
Numret är 09 839 50030.
Om du har en könssjukdom kan du även besöka polikliniken för könssjukdomar i Helsingfors eller en hälsostation.
Vanda erbjuder ungdomar under 20 år gratis preventivmedel.
Även unga vuxna under 24 år kan få gratis preventivmedel om de använder långvariga preventivmedel såsom spiral eller p-stav.
Läs mer: Sexuell hälsa och prevention.
linkkiVanda stad:
Rådgivningarna för familjeplaneringfinska _ svenska.
linkkiVanda stad:
Hälsostationernafinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Polikliniken för könssjukdomarfinska _ svenska _ engelska
Graviditet och förlossning
Vid mödrarådgivningen (äitiysneuvola) följs moderns, fostrets och hela familjens hälsotillstånd under graviditeten.
Kontakta rådgivningsbyrån (neuvola) när du upptäcker att du är gravid.
Rådgivningarnas telefontjänst
Via rådgivningsbyråernas telefontjänst kan du boka tid på rådgivningsbyrån och fråga hälsovårdaren om råd beträffande graviditet och förlossning.
Läs mer: Graviditet och förlossning och När ett barn föds i Finland.
linkkiVanda stad:
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad:
Rådgivningarna för familjeplaneringfinska _ svenska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Förlossningfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Handikappade
Du kan få tjänster för handikappade (vammaispalvelut) om du eller en närstående till dig har en invaliditet eller en sjukdom som orsakar långvariga, betydande svårigheter att klara sig hemma och i livet utanför hemmet.
Tjänster för handikappade är till exempel personlig assistans, serviceboende, färdtjänst och ombyggnadsarbeten i bostaden.
Ta kontakt med handikapprådgivningen som utreder ditt behov av stöd, handledning och tjänster utifrån din situation.
Mån.-fre. kl. 9–15
Tfn: (09) 8392 4682
Läs mer: Handikappade personer.
linkkiVanda stad:
Information om handikapptjänsternafinska _ svenska _ engelska
Hälsotjänster i Vanda
Barns hälsa
Tandvård
Mental hälsa
Sexuell hälsa och prevention
Graviditet och förlossning
Handikappade
Hälsotjänsterna i Vanda
Det allmänna nödnumret är 112.
Ring nödnumret endast om det handlar om ett nödfall, till exempel en akut sjukdomsattack.
Om din hemkommun är Vanda kan du använda kommunens offentliga hälsovårdstjänster.
Offentliga hälsovårdstjänster tillhandahålls till exempel vid hälsostationer, tandkliniker, rådgivningsbyråer och sjukhus.
Om du insjuknar akut eller råkar ut för en olycka får du akut sjukvård även om din hemkommun inte är Vanda.
Om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna, kan du boka tid på en privat läkarstation.
Läs mer: Hälsovårdstjänster i Finland.
Offentliga hälsovårdstjänster
Telefonnumret till den gemensamma telefontjänsten för hälsostationerna i Vanda är 09 839 50 000.
Du kan ringa detta nummer om du behöver rådgivning i behandlingen av en sjukdom eller vill boka eller avboka en läkartid.
Tjänsten har öppet måndag till fredag kl. 8–16.
I Vanda finns sju hälsostationer som tillhandahåller offentliga hälsovårdstjänster.
På hälsostationerna finns läkarens, sjukskötarens och hälsovårdarens mottagningar.
Om du insjuknar akut kan du gå direkt till vilken som helst hälsostation.
Det är bäst att gå till hälsostationen direkt på morgonen.
Hälsostationerna har öppet vardagar kl. 8.00–16.00.
linkkiVanda stad:
Information om hälsorådgivningfinska _ svenska _ engelska
linkkiVanda stad:
Hälsostationernafinska _ svenska _ engelska
Privata hälsotjänster
I Vanda finns flera läkarstationer som erbjuder privata hälsovårdstjänster.
Du kan gå till en privat läkarstation även om du inte har rätt att använda den offentliga hälsovårdens tjänster i Finland.
På en privat läkarstation måste du betala samtliga kostnader själv.
I vissa fall ersätter Kela en liten del av kostnaderna för privat sjukvård.
Läs mer: Hälsovårdstjänster i Finland.
Privat läkarstationfinska _ svenska _ engelska
Privat läkarstationfinska _ svenska _ engelska _ ryska
Privat läkarstationfinska _ svenska _ engelska
linkkiAava:
Privat läkarstationfinska _ svenska _ engelska
Läkemedel
Information om köp av läkemedel hittar du på InfoFinlands sida Läkemedel.
linkkiApotekareförbundet:
Apotekens kontaktuppgifterfinska
Hälsovård för papperslösa
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärhälsovård.
Tjänsterna vid Global Clinic är avgiftsfria för kunderna.
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter.
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
Telefonnumret till Helsingfors Global Clinicin är 044 948 1698.
En sjuksköterska eller läkare svarar i telefonen.
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
På kvällar, helger och storhelger är hälsostationerna stängda.
Om du insjuknar akut eller råkar ut för en olycka och inte kan vänta tills hälsostationen öppnar, kontakta jourmottagningen.
I Vanda finns jourmottagningen på Pejas sjukhus (Peijaksen sairaala).
Adress:
Sjukhusgatan 1
Tfn 116 117
Om du blir akut sjuk, kan du även besöka någon annan jourmottagning i huvudstadsregionen.
Mer information om jourmottagningarna hittar du på Vanda stads webbplats om hälsovårdstjänster.
linkkiVanda stad:
Jourmottagningarfinska _ svenska _ engelska
Barns hälsa
I hälsovården av barn under skolåldern får man hjälp av rådgivningsbyråerna (neuvola).
Telefonnumret till rådgivningsbyråerna i Vanda är 09 8392 5900.
Du kan boka en tid på rådgivningen eller fråga om råd om du har frågor kring barnets hälsa.
Skolhälsovården har hand om skolbarns hälsa.
Mer information hittar du på Vanda stads webbplats.
Om ett barn insjuknar akut, ska du kontakta hälsostationen.
Hälsostationerna har öppet måndag till fredag kl. 8–16.
När hälsostationen har stängt ska du kontakta jourmottagningen vid Barnsjukhuset.
Jourmottagningen tar endast hand om barn med brådskande hjälpbehov.
Telefonnumret till jourmottagningen är 116 117.
Adress:
Barnsjukhuset
Stenbäcksgatan 9
Du kan även ta barnet till en privat läkarstation.
I Vanda finns många privata läkarstationer som även tar hand om barn.
Läs mer: Barns hälsa.
linkkiVanda stad:
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad:
Tidsbokning och rådgivningfinska _ svenska _ engelska
linkkiVanda stad:
Information om skolhälsovårdenfinska _ svenska _ engelska
linkkiVanda stad:
Hälsostationernafinska _ svenska _ engelska
linkkiVanda stad:
Jourmottagningarfinska _ svenska _ engelska
Tandvård
Offentlig tandvård
Tidsbokningsnumret till Vanda tandvård (hammashoito) är (09) 8393 5300.
Om du inte behöver brådskande tandvård, ring efter kl. 10.00.
Om du behöver brådskande tandvård, ska du ringa tidsbokningen så fort den öppnar kl. 7.30.
Mottagningen för brådskande vård finns vid Dickursby hälsostation måndag till fredag kl. 8–14.
linkkiVanda stad:
Information om tandvårdenfinska _ svenska _ engelska
linkkiVanda stad:
Tandklinikerfinska _ svenska
Tandvårdens jourmottagning
Under kvällar och veckoslut finns tandvårdsjouren (hammashoidon päivystys) vid Haartmanska sjukhuset i Helsingfors.
Telefonnumret är 09 471 71110.
Tidsbokningen har öppet vardagar kl. 14–21 och på veckoslut kl. 8–21.
Tandvårdens nattjour (hammashoidon yöpäivystys) finns på Tölö sjukhus olycksfallsstation.
Tölö sjukhus olycksfallsstation, Oral och käkkirurgisk jourmottagning
Tfn 040 621 5699
Tandvårdens jourmottagning kvällar och veckoslutfinska _ svenska _ engelska
Barns tandvård
Om tandvården för barn under skolåldern får du information på barnrådgivningen (lastenneuvola) och vid tandklinikerna (hammashoitola).
Barn under 17 år kallas till tandkliniken för undersökning med cirka två års mellanrum.
linkkiVanda stad:
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad:
Information om tandvården för skolbarnfinska
Privata tandvårdstjänster
I Vanda finns också privata tandläkare.
Om du inte har rätt att använda de offentliga hälsovårdstjänsterna, kan du söka dig till en privat tandläkare.
Hos en privat tandläkare måste du betala samtliga kostnader själv.
I vissa fall ersätter Kela en liten del av kostnaderna för privat tandvård.
Läs mer: Tandvård.
Sök tandläkarefinska
Mental hälsa
Om du behöver psykisk hjälp eller stöd, ska du kontakta din hälsostation (terveysasema).
På hälsostationen behandlas de vanligaste psykiska problemen.
Från hälsostationen kan du remitteras vidare exempelvis till depressionsskötare.
Om hälsostationen inte har öppet och situationen är akut, ska du kontakta samjouren vid Pejas sjukhus (Peijaksen sairaalan yhteispäivystys).
Sjukhusgatan 1
Tfn 116 117
Om du behöver omedelbar krishjälp, kan du också ta kontakt med social- och krisjouren.
Den har öppet dygnet runt.
Social- och krisjouren
Tfn (09) 8392 4005
Läs mer: Mental hälsa.
linkkiVanda stad:
Information om mentalvårdstjänsternafinska _ svenska _ engelska
linkkiVanda stad:
Hälsostationernafinska _ svenska _ engelska
linkkiVanda stad:
Jourmottagningarfinska _ svenska _ engelska
linkkiVanda stad:
Social- och krisjourenfinska _ svenska _ engelska
Sexuell hälsa och prevention
Om du behöver preventivmedel eller abort eller misstänker att du har en könssjukdom, kan du kontakta preventivmedels- och familjeplaneringsrådgivningen.
Du kan boka tid per telefon.
Numret är 09 839 50030.
Om du har en könssjukdom kan du även besöka polikliniken för könssjukdomar i Helsingfors eller en hälsostation.
Vanda erbjuder ungdomar under 20 år gratis preventivmedel.
Även unga vuxna under 24 år kan få gratis preventivmedel om de använder långvariga preventivmedel såsom spiral eller p-stav.
Läs mer: Sexuell hälsa och prevention.
linkkiVanda stad:
Rådgivningarna för familjeplaneringfinska _ svenska.
linkkiVanda stad:
Hälsostationernafinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Polikliniken för könssjukdomarfinska _ svenska _ engelska
Graviditet och förlossning
Vid mödrarådgivningen (äitiysneuvola) följs moderns, fostrets och hela familjens hälsotillstånd under graviditeten.
Kontakta rådgivningsbyrån (neuvola) när du upptäcker att du är gravid.
Rådgivningarnas telefontjänst
Via rådgivningsbyråernas telefontjänst kan du boka tid på rådgivningsbyrån och fråga hälsovårdaren om råd beträffande graviditet och förlossning.
Läs mer: Graviditet och förlossning och När ett barn föds i Finland.
linkkiVanda stad:
Rådgivningsbyråerfinska _ svenska _ engelska
linkkiVanda stad:
Rådgivningarna för familjeplaneringfinska _ svenska
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS:
Förlossningfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Handikappade
Du kan få tjänster för handikappade (vammaispalvelut) om du eller en närstående till dig har en invaliditet eller en sjukdom som orsakar långvariga, betydande svårigheter att klara sig hemma och i livet utanför hemmet.
Tjänster för handikappade är till exempel personlig assistans, serviceboende, färdtjänst och ombyggnadsarbeten i bostaden.
Ta kontakt med handikapprådgivningen som utreder ditt behov av stöd, handledning och tjänster utifrån din situation.
Mån.-fre. kl. 9–15
Tfn: (09) 8392 4682
Läs mer: Handikappade personer.
linkkiVanda stad:
Information om handikapptjänsternafinska _ svenska _ engelska
Dagvård
Förskoleundervisning
Grundläggande utbildning
Yrkesutbildning
Gymnasium
Stöd och handledning för unga
Högskoleutbildning
Övriga studiemöjligheter
Dagvård
I Vanda finns både kommunala och privata daghem.
Kommunen övervakar också den privata dagvården.
I Vanda ges dagvård på finska, svenska, ryska och engelska.
Inom dagvården ges även undervisning i finska som andra språk.
Dagvård ordnas också inom familjedagvården och i gruppfamiljedaghem.
Man ska ansöka om dagvårdsplats för sitt barn minst fyra månader innan barnet ska börja i dagvården.
Du kan ansöka om plats i den kommunala dagvården via Internet eller med en pappersblankett.
För en elektronisk ansökan behöver du egna nätbankskoder eller en elektronisk legitimation.
Pappersblanketter kan hämtas till exempel vid Vandainfo eller daghemmen.
Privata dagvårdsplatser söks direkt på daghemmet.
Frågor kring dagvård och ansökan om dagvårdsplats kan du ställa till daghemsföreståndaren eller skicka till adressen varhaiskasvatus(at)vantaa.fi.
Vanligtvis ansöker man om dagvårdsplats i den egna kommunen.
Om familjen bor nära gränsen till Helsingfors eller Esbo, kan du också söka dagvårdsplats i grannkommunen.
Du ska ändå lämna in din ansökan i den egna kommunen.
Mer information hittar du via tjänsten Helsingforsregionen.fi.
Läs mer: Dagvård
linkkiVanda stad:
Privat dagvårdfinska _ svenska _ engelska
linkkiVanda stad:
Privat dagvårdfinska
linkkiVanda stad:
Ansökan om dagvårdsplatsfinska _ svenska _ engelska
linkkiVanda stad:
Elektronisk ansökningsblankett för dagvårdenfinska _ svenska _ engelska
Information om dagvården finska _ svenska _ engelska
Förskoleundervisning
Förskoleundervisning (esiopetus) ordnas i både kommunala och privata daghem samt i förskoleenheter i skolornas lokaler.
I Vanda kan man få förskoleundervisning på finska, svenska och engelska.
Du måste ansöka om plats i förskoleundervisningen.
Ansökan kan göras elektroniskt via stadens webbplats eller med en pappersblankett.
Ansökningstiden är i januari, men ansökan kan även lämnas in övriga tider, om familjen till exempel flyttar till Vanda mitt under året.
Förberedande undervisning tillhandahålls för invandrarbarn som inte har tillräckliga kunskaper i finska för att klara sig i förskoleundervisningen.
Den förberedande undervisningen är avsedd för 6-åriga barn med invandrarbakgrund.
Den ordnas i daghemmens förskolegrupper.
Daghemmet anvisar barnet till den förberedande undervisningen i samband med ansökningen till förskoleundervisningen.
Du hittar mer information om förskoleundervisningen, ansökning till förskoleundervisningen och om undervisning som förbereder för förskoleundervisning på Vanda stads (Vantaan kaupunki) webbplats.
Du kan även fråga om mer information på daghemmen.
Läs mer: Förskoleundervisning
linkkiVanda stad:
Ansökan till förskoleundervisningfinska _ svenska _ engelska
linkkiVanda stad:
Information om den förberedande undervisningenfinska _ engelska
linkkiVanda stad:
Elektronisk ansökningsblankett för förskoleundervisningenfinska _ svenska _ engelska
linkkiVanda stad:
Daghem som ger förskoleundervisningfinska _ engelska
Grundläggande utbildning
I Vanda finns finskspråkiga och svenskspråkiga grundskolor (peruskoulu).
I Vanda finns även en internationell skola, där man kan avlägga grundskolan på engelska.
Mer information om skolorna i Vanda hittar du på Vanda stads (Vantaan kaupunki) webbplats.
Anmälan till grundskolan ska göras på förhand.
Anmälningstiden är vanligtvis i januari.
På stadens webbplats hittar du kontaktuppgifterna till skolorna och mer information om anmälan.
Läs mer: Grundläggande utbildning
linkkiVanda stad:
Anmälan till skolanfinska _ svenska _ engelska
linkkiVanda stad:
Skolornas kontaktuppgifterfinska
Eftermiddagsverksamhetfinska _ svenska
Förberedande utbildning inför grundskola
Om barnets kunskaper i det finska språket inte är tillräckligt bra för studier i den finskspråkiga grundskolan, kan barnet få förberedande utbildning (valmistava opetus).
I den förberedande utbildningen läser barnen det finska språket och grundskolans läroämnen.
Undervisningen pågår vanligtvis i ett år.
Om du har anlänt till Finland för en kort tid sedan och har barn under skolåldern ska du ta kontakt med områdeskoordinatorn för ditt bostadsområde (aluekoordinaattori).
Områdeskoordinatorn berättar om hur undervisningen ordnas och hjälper dig i frågor som rör barnets skolgång.
Information om den förberedande undervisningenfinska
linkkiVanda stad:
Områdeskoordinatorerfinska
Grundläggande utbildning för unga invandrare
Vid Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto) kan 17–24-åriga invandrarungdomar avlägga grundskolans avgångsbetyg.
Om man har hoppat av grundskolan, kan man avlägga grundskolans lärokurs också vid Eira vuxengymnasium (Eiran aikuislukio).
Grundläggande utbildning för invandrarefinska
linkkiEira vuxengymnasium:
Grundundervisning för vuxnafinska
Tionde klasserna
Du kan ansöka till den grundläggande utbildningens tilläggsundervisning, det vill säga till en tionde klass (kymppiluokka), om du fick grundskolans avgångsbetyg samma år eller året innan, men inte har fått en studieplats på andra stadiet.
På tionde klassen kan du höja dina betyg från grundskolan och du får en plan för fortsatta studier.
Tiondeklasserna i Vanda finns i östra och västra Vanda vid Varias verksamhetsställen och vid Lumo gymnasium (Lumon lukio).
linkkiVanda stad:
Tiondeklasserfinska _ svenska
Invandrare och grundläggande utbildning
I skolorna i Vanda ges hemspråksundervisning i flera olika språk.
I grundskolorna ges även utbildning i finska som andraspråk (suomi toisena kielenä) till elever som har ett annat modersmål än finska, svenska eller samiska, och vars kunskaper i det finska språket inte är i nivå med modersmålet.
När du anmäler dig till skolan, kan du samtidigt anmäla dig till hemspråksundervisning och undervisning i din egen religion.
Du kan även anmäla dig till undervisningen genom att fylla i en blankett, som du får från din egen skola.
Den ifyllda blanketten returneras till den egna skolan.
Undervisning i den egna religionen kan ordnas om gruppen består av minst tre elever.
Mer information om hemspråksundervisning och om undervisning i elevens egen religion hittar du på stadens webbplats och hos områdeskoordinatorerna (aluekoordinaattori).
linkkiVanda stad:
Information om hemspråksundervisningfinska
linkkiVanda stad:
Undervisning i den egna religionenfinska
Finska som andra språk i den grundläggande undervisningenfinska
linkkiVanda stad:
Områdeskoordinatorerfinska
Yrkesutbildning
I Vanda ordnas yrkesutbildning vid yrkesinstitutet Vantaan ammattiopisto Varia, handelsläroanstalten MERCURIA samt TTS Arbetseffektivitetsföreningen rf:s verksamhetsställe i Vanda.
I Varia ordnas även engelskspråkig undervisning samt finskspråkiga yrkesutbildningar särskilt avsedda för invandrare.
Edupoli ordnar yrkesutbildning för vuxna.
I Vanda finns även Finavia Avia College som ger utbildning för olika luftfartsyrken.
Läs mer: Yrkesutbildning.
linkkiVanda stad:
Yrkesutbildningfinska _ svenska
linkkiYrkesläroanstalten Varia i Vanda:
Yrkesutbildningfinska _ engelska
Yrkesutbildningfinska _ engelska
linkkiTTS Arbetseffektivitetsföreningen rf:s verksamhetsställe i Vanda:
Yrkesutbildningfinska
Utbildning som handleder för yrkesutbildning (VALMA)
Utbildning som handleder för grundläggande yrkesutbildning (Ammatilliseen peruskoulutukseen valmentava koulutus) d.v.s. VALMA är avsedd för dem som vill avlägga en grundläggande yrkesutbildning.
Under VALMA-utbildningen får du kunskap och färdigheter som hjälper dig i dina senare yrkesinriktade studier.
Du kan även förbättra din språkkunskap. Du kan också höja dina grundskolebetyg.
I Vanda ordnas VALMA-utbildning av Varia.
Läs mer om VALMA-utbildningen på InfoFinlands sida Utbildning som handleder för yrkesutbildning.
linkkiVanda stad:
Information om VALMA-utbildningarfinska
linkkiYrkesläroanstalten Varia i Vanda:
I Vanda kan du studera på gymnasiet (lukio) på finska, svenska eller engelska.
Undervisning på engelska erbjuds på IB-linjen vid gymnasieskolan Tikkurilan lukio.
I Vanda finns även ett vuxengymnasium.
Läs mer: Gymnasium.
linkkiVanda stad:
Information om gymnasieutbildningfinska _ svenska
linkkiVanda stad:
Gymnasierna och gymnasiernas hemsidorfinska
linkkiVanda stad:
Vuxengymnasiumfinska
linkkiVanda stad:
Distansgymnasiumfinska
linkkiVanda stad:
Steinergymnasietfinska
Förberedande gymnasieutbildning (LUVA)
Om du vill förbättra dina kunskaper i finska eller svenska innan du söker till ett gymnasium, kan du söka till en förberedande gymnasieutbildning.
Den är avsedd för invandrare.
I Vanda ordnas LUVA-utbildning av Lumon lukio.
Läs mer om LUVA-utbildningen på InfoFinlands sida Förberedande gymnasieutbildning.
linkkiVanda stad:
Förberedande gymnasieutbildningfinska
Stöd och handledning för unga
Om du är under 30 år gammal kan du få råd och handledning via Ohjaamo-tjänsten.
Ohjaamos personal hjälper dig om du inte har ett arbete eller en studieplats.
Du kan även fråga om andra saker, som till exempel boende eller ekonomiska frågor.
linkkiOhjaamo:
Stöd och handledning för ungafinska _ engelska
Vägledningscentret Kipinä
Om du är under 29 år gammal, bor i Vanda och inte har ett jobb eller en studieplats, kan du få råd och handledning i Kipinä.
Ring och boka en tid i förväg.
Utan tidsbokning kan du besöka Kipinä på tisdagar och onsdagar kl. 12.00–18.00.
Mer information hittar du på webbplatsen.
Kipinä
Banvägen 2, Dickursby
Tfn 050 312 4372
Vägledning och stöd för ungafinska _ svenska
Högskoleutbildning
I Vanda finns två yrkeshögskolor (ammattikorkeakoulu), Laurea och Metropolia.
De erbjuder utbildning inom många olika branscher.
Mer information om utbildningsprogram och om ansökan hittar du på läroanstalternas webbplats.
Också Helsingfors universitets öppna universitet (avoin yliopisto) har verksamhetsställen i Vanda. Där ges undervisning på högskolenivå och fortbildning.
Läs mer: Högskoleutbildning.
linkkiVanda stad:
Högskoleutbildningfinska
Yrkeshögskolafinska _ engelska
linkkiMetropolia:
Yrkeshögskolafinska _ engelska
Ubildning vid öppna universitetet i Vandafinska _ svenska _ engelska
Övriga studiemöjligheter
Vid Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto) kan du studera till exempel språk, handarbete och matlagning eller delta i ledd motion.
Kurserna är avgiftsbelagda och de ordnas både dag- och kvällstid.
Vuxenutbildningsinstitutet ordnar även kurser för invandrare.
Mer information hittar du på Vanda stads webbplats.
Läs mer: Andra studiemöjligheter.
linkkiVanda vuxenutbildningsinstitut:
Studiehandbokfinska
linkkiVanda vuxenutbildningsinstitut:
Kurser i finska och svenska språket för invandrarefinska
linkkiEdupoli:
Vuxenutbildningscenterfinska
Dagvård
Förskoleundervisning
Grundläggande utbildning
Yrkesutbildning
Gymnasium
Stöd och handledning för unga
Högskoleutbildning
Övriga studiemöjligheter
Dagvård
I Vanda finns både kommunala och privata daghem.
Kommunen övervakar också den privata dagvården.
I Vanda ges dagvård på finska, svenska, ryska och engelska.
Inom dagvården ges även undervisning i finska som andra språk.
Dagvård ordnas också inom familjedagvården och i gruppfamiljedaghem.
Man ska ansöka om dagvårdsplats för sitt barn minst fyra månader innan barnet ska börja i dagvården.
Du kan ansöka om plats i den kommunala dagvården via Internet eller med en pappersblankett.
För en elektronisk ansökan behöver du egna nätbankskoder eller en elektronisk legitimation.
Pappersblanketter kan hämtas till exempel vid Vandainfo eller daghemmen.
Privata dagvårdsplatser söks direkt på daghemmet.
Frågor kring dagvård och ansökan om dagvårdsplats kan du ställa till daghemsföreståndaren eller skicka till adressen varhaiskasvatus(at)vantaa.fi.
Vanligtvis ansöker man om dagvårdsplats i den egna kommunen.
Om familjen bor nära gränsen till Helsingfors eller Esbo, kan du också söka dagvårdsplats i grannkommunen.
Du ska ändå lämna in din ansökan i den egna kommunen.
Mer information hittar du via tjänsten Helsingforsregionen.fi.
Läs mer: Dagvård
linkkiVanda stad:
Privat dagvårdfinska _ svenska _ engelska
linkkiVanda stad:
Privat dagvårdfinska
linkkiVanda stad:
Ansökan om dagvårdsplatsfinska _ svenska _ engelska
linkkiVanda stad:
Elektronisk ansökningsblankett för dagvårdenfinska _ svenska _ engelska
Information om dagvården finska _ svenska _ engelska
Förskoleundervisning
Förskoleundervisning (esiopetus) ordnas i både kommunala och privata daghem samt i förskoleenheter i skolornas lokaler.
I Vanda kan man få förskoleundervisning på finska, svenska och engelska.
Du måste ansöka om plats i förskoleundervisningen.
Ansökan kan göras elektroniskt via stadens webbplats eller med en pappersblankett.
Ansökningstiden är i januari, men ansökan kan även lämnas in övriga tider, om familjen till exempel flyttar till Vanda mitt under året.
Förberedande undervisning tillhandahålls för invandrarbarn som inte har tillräckliga kunskaper i finska för att klara sig i förskoleundervisningen.
Den förberedande undervisningen är avsedd för 6-åriga barn med invandrarbakgrund.
Den ordnas i daghemmens förskolegrupper.
Daghemmet anvisar barnet till den förberedande undervisningen i samband med ansökningen till förskoleundervisningen.
Du hittar mer information om förskoleundervisningen, ansökning till förskoleundervisningen och om undervisning som förbereder för förskoleundervisning på Vanda stads (Vantaan kaupunki) webbplats.
Du kan även fråga om mer information på daghemmen.
Läs mer: Förskoleundervisning
linkkiVanda stad:
Ansökan till förskoleundervisningfinska _ svenska _ engelska
linkkiVanda stad:
Information om den förberedande undervisningenfinska _ engelska
linkkiVanda stad:
Elektronisk ansökningsblankett för förskoleundervisningenfinska _ svenska _ engelska
linkkiVanda stad:
Daghem som ger förskoleundervisningfinska _ engelska
Grundläggande utbildning
I Vanda finns finskspråkiga och svenskspråkiga grundskolor (peruskoulu).
I Vanda finns även en internationell skola, där man kan avlägga grundskolan på engelska.
Mer information om skolorna i Vanda hittar du på Vanda stads (Vantaan kaupunki) webbplats.
Anmälan till grundskolan ska göras på förhand.
Anmälningstiden är vanligtvis i januari.
På stadens webbplats hittar du kontaktuppgifterna till skolorna och mer information om anmälan.
Läs mer: Grundläggande utbildning
linkkiVanda stad:
Anmälan till skolanfinska _ svenska _ engelska
linkkiVanda stad:
Skolornas kontaktuppgifterfinska
Eftermiddagsverksamhetfinska _ svenska
Förberedande utbildning inför grundskola
Om barnets kunskaper i det finska språket inte är tillräckligt bra för studier i den finskspråkiga grundskolan, kan barnet få förberedande utbildning (valmistava opetus).
I den förberedande utbildningen läser barnen det finska språket och grundskolans läroämnen.
Undervisningen pågår vanligtvis i ett år.
Om du har anlänt till Finland för en kort tid sedan och har barn under skolåldern ska du ta kontakt med områdeskoordinatorn för ditt bostadsområde (aluekoordinaattori).
Områdeskoordinatorn berättar om hur undervisningen ordnas och hjälper dig i frågor som rör barnets skolgång.
Information om den förberedande undervisningenfinska
linkkiVanda stad:
Områdeskoordinatorerfinska
Grundläggande utbildning för unga invandrare
Vid Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto) kan 17–24-åriga invandrarungdomar avlägga grundskolans avgångsbetyg.
Om man har hoppat av grundskolan, kan man avlägga grundskolans lärokurs också vid Eira vuxengymnasium (Eiran aikuislukio).
Grundläggande utbildning för invandrarefinska
linkkiEira vuxengymnasium:
Grundundervisning för vuxnafinska
Tionde klasserna
Du kan ansöka till den grundläggande utbildningens tilläggsundervisning, det vill säga till en tionde klass (kymppiluokka), om du fick grundskolans avgångsbetyg samma år eller året innan, men inte har fått en studieplats på andra stadiet.
På tionde klassen kan du höja dina betyg från grundskolan och du får en plan för fortsatta studier.
Tiondeklasserna i Vanda finns i östra och västra Vanda vid Varias verksamhetsställen och vid Lumo gymnasium (Lumon lukio).
linkkiVanda stad:
Tiondeklasserfinska _ svenska
Invandrare och grundläggande utbildning
I skolorna i Vanda ges hemspråksundervisning i flera olika språk.
I grundskolorna ges även utbildning i finska som andraspråk (suomi toisena kielenä) till elever som har ett annat modersmål än finska, svenska eller samiska, och vars kunskaper i det finska språket inte är i nivå med modersmålet.
När du anmäler dig till skolan, kan du samtidigt anmäla dig till hemspråksundervisning och undervisning i din egen religion.
Du kan även anmäla dig till undervisningen genom att fylla i en blankett, som du får från din egen skola.
Den ifyllda blanketten returneras till den egna skolan.
Undervisning i den egna religionen kan ordnas om gruppen består av minst tre elever.
Mer information om hemspråksundervisning och om undervisning i elevens egen religion hittar du på stadens webbplats och hos områdeskoordinatorerna (aluekoordinaattori).
linkkiVanda stad:
Information om hemspråksundervisningfinska
linkkiVanda stad:
Undervisning i den egna religionenfinska
Finska som andra språk i den grundläggande undervisningenfinska
linkkiVanda stad:
Områdeskoordinatorerfinska
Yrkesutbildning
I Vanda ordnas yrkesutbildning vid yrkesinstitutet Vantaan ammattiopisto Varia, handelsläroanstalten MERCURIA samt TTS Arbetseffektivitetsföreningen rf:s verksamhetsställe i Vanda.
I Varia ordnas även engelskspråkig undervisning samt finskspråkiga yrkesutbildningar särskilt avsedda för invandrare.
Edupoli ordnar yrkesutbildning för vuxna.
I Vanda finns även Finavia Avia College som ger utbildning för olika luftfartsyrken.
Läs mer: Yrkesutbildning.
linkkiVanda stad:
Yrkesutbildningfinska _ svenska
linkkiYrkesläroanstalten Varia i Vanda:
Yrkesutbildningfinska _ engelska
Yrkesutbildningfinska _ engelska
linkkiTTS Arbetseffektivitetsföreningen rf:s verksamhetsställe i Vanda:
Yrkesutbildningfinska
Utbildning som handleder för yrkesutbildning (VALMA)
Utbildning som handleder för grundläggande yrkesutbildning (Ammatilliseen peruskoulutukseen valmentava koulutus) d.v.s. VALMA är avsedd för dem som vill avlägga en grundläggande yrkesutbildning.
Under VALMA-utbildningen får du kunskap och färdigheter som hjälper dig i dina senare yrkesinriktade studier.
Du kan även förbättra din språkkunskap. Du kan också höja dina grundskolebetyg.
I Vanda ordnas VALMA-utbildning av Varia.
Läs mer om VALMA-utbildningen på InfoFinlands sida Utbildning som handleder för yrkesutbildning.
linkkiVanda stad:
Information om VALMA-utbildningarfinska
linkkiYrkesläroanstalten Varia i Vanda:
I Vanda kan du studera på gymnasiet (lukio) på finska, svenska eller engelska.
Undervisning på engelska erbjuds på IB-linjen vid gymnasieskolan Tikkurilan lukio.
I Vanda finns även ett vuxengymnasium.
Läs mer: Gymnasium.
linkkiVanda stad:
Information om gymnasieutbildningfinska _ svenska
linkkiVanda stad:
Gymnasierna och gymnasiernas hemsidorfinska
linkkiVanda stad:
Vuxengymnasiumfinska
linkkiVanda stad:
Distansgymnasiumfinska
linkkiVanda stad:
Steinergymnasietfinska
Förberedande gymnasieutbildning (LUVA)
Om du vill förbättra dina kunskaper i finska eller svenska innan du söker till ett gymnasium, kan du söka till en förberedande gymnasieutbildning.
Den är avsedd för invandrare.
I Vanda ordnas LUVA-utbildning av Lumon lukio.
Läs mer om LUVA-utbildningen på InfoFinlands sida Förberedande gymnasieutbildning.
linkkiVanda stad:
Förberedande gymnasieutbildningfinska
Stöd och handledning för unga
Om du är under 30 år gammal kan du få råd och handledning via Ohjaamo-tjänsten.
Ohjaamos personal hjälper dig om du inte har ett arbete eller en studieplats.
Du kan även fråga om andra saker, som till exempel boende eller ekonomiska frågor.
linkkiOhjaamo:
Stöd och handledning för ungafinska _ engelska
Vägledningscentret Kipinä
Om du är under 29 år gammal, bor i Vanda och inte har ett jobb eller en studieplats, kan du få råd och handledning i Kipinä.
Ring och boka en tid i förväg.
Utan tidsbokning kan du besöka Kipinä på tisdagar och onsdagar kl. 12.00–18.00.
Mer information hittar du på webbplatsen.
Kipinä
Banvägen 2, Dickursby
Tfn 050 312 4372
Vägledning och stöd för ungafinska _ svenska
Högskoleutbildning
I Vanda finns två yrkeshögskolor (ammattikorkeakoulu), Laurea och Metropolia.
De erbjuder utbildning inom många olika branscher.
Mer information om utbildningsprogram och om ansökan hittar du på läroanstalternas webbplats.
Också Helsingfors universitets öppna universitet (avoin yliopisto) har verksamhetsställen i Vanda. Där ges undervisning på högskolenivå och fortbildning.
Läs mer: Högskoleutbildning.
linkkiVanda stad:
Högskoleutbildningfinska
Yrkeshögskolafinska _ engelska
linkkiMetropolia:
Yrkeshögskolafinska _ engelska
Ubildning vid öppna universitetet i Vandafinska _ svenska _ engelska
Övriga studiemöjligheter
Vid Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto) kan du studera till exempel språk, handarbete och matlagning eller delta i ledd motion.
Kurserna är avgiftsbelagda och de ordnas både dag- och kvällstid.
Vuxenutbildningsinstitutet ordnar även kurser för invandrare.
Mer information hittar du på Vanda stads webbplats.
Läs mer: Andra studiemöjligheter.
linkkiVanda vuxenutbildningsinstitut:
Studiehandbokfinska
linkkiVanda vuxenutbildningsinstitut:
Kurser i finska och svenska språket för invandrarefinska
linkkiEdupoli:
Vuxenutbildningscenterfinska
Dagvård
Förskoleundervisning
Grundläggande utbildning
Yrkesutbildning
Gymnasium
Stöd och handledning för unga
Högskoleutbildning
Övriga studiemöjligheter
Dagvård
I Vanda finns både kommunala och privata daghem.
Kommunen övervakar också den privata dagvården.
I Vanda ges dagvård på finska, svenska, ryska och engelska.
Inom dagvården ges även undervisning i finska som andra språk.
Dagvård ordnas också inom familjedagvården och i gruppfamiljedaghem.
Man ska ansöka om dagvårdsplats för sitt barn minst fyra månader innan barnet ska börja i dagvården.
Du kan ansöka om plats i den kommunala dagvården via Internet eller med en pappersblankett.
För en elektronisk ansökan behöver du egna nätbankskoder eller en elektronisk legitimation.
Pappersblanketter kan hämtas till exempel vid Vandainfo eller daghemmen.
Privata dagvårdsplatser söks direkt på daghemmet.
Frågor kring dagvård och ansökan om dagvårdsplats kan du ställa till daghemsföreståndaren eller skicka till adressen varhaiskasvatus(at)vantaa.fi.
Vanligtvis ansöker man om dagvårdsplats i den egna kommunen.
Om familjen bor nära gränsen till Helsingfors eller Esbo, kan du också söka dagvårdsplats i grannkommunen.
Du ska ändå lämna in din ansökan i den egna kommunen.
Mer information hittar du via tjänsten Helsingforsregionen.fi.
Läs mer: Dagvård
linkkiVanda stad:
Privat dagvårdfinska _ svenska _ engelska
linkkiVanda stad:
Privat dagvårdfinska
linkkiVanda stad:
Ansökan om dagvårdsplatsfinska _ svenska _ engelska
linkkiVanda stad:
Elektronisk ansökningsblankett för dagvårdenfinska _ svenska _ engelska
Information om dagvården finska _ svenska _ engelska
Förskoleundervisning
Förskoleundervisning (esiopetus) ordnas i både kommunala och privata daghem samt i förskoleenheter i skolornas lokaler.
I Vanda kan man få förskoleundervisning på finska, svenska och engelska.
Du måste ansöka om plats i förskoleundervisningen.
Ansökan kan göras elektroniskt via stadens webbplats eller med en pappersblankett.
Ansökningstiden är i januari, men ansökan kan även lämnas in övriga tider, om familjen till exempel flyttar till Vanda mitt under året.
Förberedande undervisning tillhandahålls för invandrarbarn som inte har tillräckliga kunskaper i finska för att klara sig i förskoleundervisningen.
Den förberedande undervisningen är avsedd för 6-åriga barn med invandrarbakgrund.
Den ordnas i daghemmens förskolegrupper.
Daghemmet anvisar barnet till den förberedande undervisningen i samband med ansökningen till förskoleundervisningen.
Du hittar mer information om förskoleundervisningen, ansökning till förskoleundervisningen och om undervisning som förbereder för förskoleundervisning på Vanda stads (Vantaan kaupunki) webbplats.
Du kan även fråga om mer information på daghemmen.
Läs mer: Förskoleundervisning
linkkiVanda stad:
Ansökan till förskoleundervisningfinska _ svenska _ engelska
linkkiVanda stad:
Information om den förberedande undervisningenfinska _ engelska
linkkiVanda stad:
Elektronisk ansökningsblankett för förskoleundervisningenfinska _ svenska _ engelska
linkkiVanda stad:
Daghem som ger förskoleundervisningfinska _ engelska
Grundläggande utbildning
I Vanda finns finskspråkiga och svenskspråkiga grundskolor (peruskoulu).
I Vanda finns även en internationell skola, där man kan avlägga grundskolan på engelska.
Mer information om skolorna i Vanda hittar du på Vanda stads (Vantaan kaupunki) webbplats.
Anmälan till grundskolan ska göras på förhand.
Anmälningstiden är vanligtvis i januari.
På stadens webbplats hittar du kontaktuppgifterna till skolorna och mer information om anmälan.
Läs mer: Grundläggande utbildning
linkkiVanda stad:
Anmälan till skolanfinska _ svenska _ engelska
linkkiVanda stad:
Skolornas kontaktuppgifterfinska
Eftermiddagsverksamhetfinska _ svenska
Förberedande utbildning inför grundskola
Om barnets kunskaper i det finska språket inte är tillräckligt bra för studier i den finskspråkiga grundskolan, kan barnet få förberedande utbildning (valmistava opetus).
I den förberedande utbildningen läser barnen det finska språket och grundskolans läroämnen.
Undervisningen pågår vanligtvis i ett år.
Om du har anlänt till Finland för en kort tid sedan och har barn under skolåldern ska du ta kontakt med områdeskoordinatorn för ditt bostadsområde (aluekoordinaattori).
Områdeskoordinatorn berättar om hur undervisningen ordnas och hjälper dig i frågor som rör barnets skolgång.
Information om den förberedande undervisningenfinska
linkkiVanda stad:
Områdeskoordinatorerfinska
Grundläggande utbildning för unga invandrare
Vid Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto) kan 17–24-åriga invandrarungdomar avlägga grundskolans avgångsbetyg.
Om man har hoppat av grundskolan, kan man avlägga grundskolans lärokurs också vid Eira vuxengymnasium (Eiran aikuislukio).
Grundläggande utbildning för invandrarefinska
linkkiEira vuxengymnasium:
Grundundervisning för vuxnafinska
Tionde klasserna
Du kan ansöka till den grundläggande utbildningens tilläggsundervisning, det vill säga till en tionde klass (kymppiluokka), om du fick grundskolans avgångsbetyg samma år eller året innan, men inte har fått en studieplats på andra stadiet.
På tionde klassen kan du höja dina betyg från grundskolan och du får en plan för fortsatta studier.
Tiondeklasserna i Vanda finns i östra och västra Vanda vid Varias verksamhetsställen och vid Lumo gymnasium (Lumon lukio).
linkkiVanda stad:
Tiondeklasserfinska _ svenska
Invandrare och grundläggande utbildning
I skolorna i Vanda ges hemspråksundervisning i flera olika språk.
I grundskolorna ges även utbildning i finska som andraspråk (suomi toisena kielenä) till elever som har ett annat modersmål än finska, svenska eller samiska, och vars kunskaper i det finska språket inte är i nivå med modersmålet.
När du anmäler dig till skolan, kan du samtidigt anmäla dig till hemspråksundervisning och undervisning i din egen religion.
Du kan även anmäla dig till undervisningen genom att fylla i en blankett, som du får från din egen skola.
Den ifyllda blanketten returneras till den egna skolan.
Undervisning i den egna religionen kan ordnas om gruppen består av minst tre elever.
Mer information om hemspråksundervisning och om undervisning i elevens egen religion hittar du på stadens webbplats och hos områdeskoordinatorerna (aluekoordinaattori).
linkkiVanda stad:
Information om hemspråksundervisningfinska
linkkiVanda stad:
Undervisning i den egna religionenfinska
Finska som andra språk i den grundläggande undervisningenfinska
linkkiVanda stad:
Områdeskoordinatorerfinska
Yrkesutbildning
I Vanda ordnas yrkesutbildning vid yrkesinstitutet Vantaan ammattiopisto Varia, handelsläroanstalten MERCURIA samt TTS Arbetseffektivitetsföreningen rf:s verksamhetsställe i Vanda.
I Varia ordnas även engelskspråkig undervisning samt finskspråkiga yrkesutbildningar särskilt avsedda för invandrare.
Edupoli ordnar yrkesutbildning för vuxna.
I Vanda finns även Finavia Avia College som ger utbildning för olika luftfartsyrken.
Läs mer: Yrkesutbildning.
linkkiVanda stad:
Yrkesutbildningfinska _ svenska
linkkiYrkesläroanstalten Varia i Vanda:
Yrkesutbildningfinska _ engelska
Yrkesutbildningfinska _ engelska
linkkiTTS Arbetseffektivitetsföreningen rf:s verksamhetsställe i Vanda:
Yrkesutbildningfinska
Utbildning som handleder för yrkesutbildning (VALMA)
Utbildning som handleder för grundläggande yrkesutbildning (Ammatilliseen peruskoulutukseen valmentava koulutus) d.v.s. VALMA är avsedd för dem som vill avlägga en grundläggande yrkesutbildning.
Under VALMA-utbildningen får du kunskap och färdigheter som hjälper dig i dina senare yrkesinriktade studier.
Du kan även förbättra din språkkunskap. Du kan också höja dina grundskolebetyg.
I Vanda ordnas VALMA-utbildning av Varia.
Läs mer om VALMA-utbildningen på InfoFinlands sida Utbildning som handleder för yrkesutbildning.
linkkiVanda stad:
Information om VALMA-utbildningarfinska
linkkiYrkesläroanstalten Varia i Vanda:
I Vanda kan du studera på gymnasiet (lukio) på finska, svenska eller engelska.
Undervisning på engelska erbjuds på IB-linjen vid gymnasieskolan Tikkurilan lukio.
I Vanda finns även ett vuxengymnasium.
Läs mer: Gymnasium.
linkkiVanda stad:
Information om gymnasieutbildningfinska _ svenska
linkkiVanda stad:
Gymnasierna och gymnasiernas hemsidorfinska
linkkiVanda stad:
Vuxengymnasiumfinska
linkkiVanda stad:
Distansgymnasiumfinska
linkkiVanda stad:
Steinergymnasietfinska
Förberedande gymnasieutbildning (LUVA)
Om du vill förbättra dina kunskaper i finska eller svenska innan du söker till ett gymnasium, kan du söka till en förberedande gymnasieutbildning.
Den är avsedd för invandrare.
I Vanda ordnas LUVA-utbildning av Lumon lukio.
Läs mer om LUVA-utbildningen på InfoFinlands sida Förberedande gymnasieutbildning.
linkkiVanda stad:
Förberedande gymnasieutbildningfinska
Stöd och handledning för unga
Om du är under 30 år gammal kan du få råd och handledning via Ohjaamo-tjänsten.
Ohjaamos personal hjälper dig om du inte har ett arbete eller en studieplats.
Du kan även fråga om andra saker, som till exempel boende eller ekonomiska frågor.
linkkiOhjaamo:
Stöd och handledning för ungafinska _ engelska
Vägledningscentret Kipinä
Om du är under 29 år gammal, bor i Vanda och inte har ett jobb eller en studieplats, kan du få råd och handledning i Kipinä.
Ring och boka en tid i förväg.
Utan tidsbokning kan du besöka Kipinä på tisdagar och onsdagar kl. 12.00–18.00.
Mer information hittar du på webbplatsen.
Kipinä
Banvägen 2, Dickursby
Tfn 050 312 4372
Vägledning och stöd för ungafinska _ svenska
Högskoleutbildning
I Vanda finns två yrkeshögskolor (ammattikorkeakoulu), Laurea och Metropolia.
De erbjuder utbildning inom många olika branscher.
Mer information om utbildningsprogram och om ansökan hittar du på läroanstalternas webbplats.
Också Helsingfors universitets öppna universitet (avoin yliopisto) har verksamhetsställen i Vanda. Där ges undervisning på högskolenivå och fortbildning.
Läs mer: Yrkeshögskolor, Universitet.
linkkiVanda stad:
Högskoleutbildningfinska
Yrkeshögskolafinska _ engelska
linkkiMetropolia:
Yrkeshögskolafinska _ engelska
Ubildning vid öppna universitetet i Vandafinska _ svenska _ engelska
Övriga studiemöjligheter
Vid Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto) kan du studera till exempel språk, handarbete och matlagning eller delta i ledd motion.
Kurserna är avgiftsbelagda och de ordnas både dag- och kvällstid.
Vuxenutbildningsinstitutet ordnar även kurser för invandrare.
Mer information hittar du på Vanda stads webbplats.
Läs mer: Studier som hobby.
linkkiVanda vuxenutbildningsinstitut:
Studiehandbokfinska
linkkiVanda vuxenutbildningsinstitut:
Kurser i finska och svenska språket för invandrarefinska
linkkiEdupoli:
Vuxenutbildningscenterfinska
Detta innehåll finns inte på det språk som du har valt.
Välj något annat språk.
Finska
Detta innehåll finns inte på det språk som du har valt.
Välj något annat språk.
Finska
Detta innehåll finns inte på det språk som du har valt.
Välj något annat språk.
Finska
Hyresbostad
Boende i en krissituation
Bostadslöshet
Stöd- och serviceboende
Bostadens avfallshantering
Hyresbostad
Hyresbostäderna är ofta dyra i huvudstadsregionen.
Du är själv ansvarig för att skaffa bostad åt dig själv.
Varken staden eller andra hyresvärdar har skyldighet att erbjuda dig bostad.
Läs mer: Hyresbostad.
Privata hyresbostäder
I Vanda finns också många andra hyresvärdar, varav de största är VVO, Sato och Avara.
Därtill ägs hyresbostäder i Vanda av många försäkringsbolag, Kuntien eläkevakuutus och Kunta-asunnot.
Det kan gå snabbt att få bostad via en privat hyresvärd.
Om du är studerande kan du ansöka om en hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS (Helsingin seudun Opiskelija-asuntosäätiö HOAS).
Om du är yngre än 30 år, kan du söka bostad hos Förbundet för ungdomsbostäder (Nuorisoasuntoliitto) och stiftelsen Nuorisosäätiö (Nuorisosäätiö).
linkkiSATO:
Hyresbostäderfinska _ engelska
linkkiAvara:
Hyresbostäderfinska
linkkiKommunbostäder:
Hyresbostäderfinska _ svenska _ engelska
linkkiFörbundet för ungdomsbostäder:
Hyresbostäder för personer under 30 årfinska _ engelska
Hyresbostäder för ungafinska _ engelska
linkkiHOAS:
Hyresbostäder för studerandefinska _ svenska _ engelska
Stadens hyresbostäder
Stadens hyresbostäder är vanligtvis förmånligare än de bostäder som hyrs ut av företag och privatpersoner.
Väntetiden för dessa bostäder kan dock vara lång och endast en liten del av de sökande får en bostad.
Vanda stads hyresbostäder ägs och hyrs ut av VAV Asunnot Oy.
Lokgränden 7
Tfn 010 235 1450 (kundtjänst)
Du kan göra en bostadsansökan på VAV Asunnot Oy:s webbplats.
Ansökan är giltig i fyra månader och måste sedan förnyas.
Vid val av invånare till stadens hyresbostäder prioriteras de sökande som har ett akut bostadsbehov.
Också sökandens inkomster beaktas, eftersom bostäderna främst är avsedda för personer med låga inkomster.
Information om stadens hyresbostäderfinska _ engelska
Ansökan om hyresbostad i stadenfinska _ engelska
Boende i en krissituation
Om din bostad har skadats till exempel till följd av brand eller vattenskada kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
Kontakta ditt försäkringsbolag direkt när skadan har inträffat.
I krissituationer får man även hjälp vid Vanda stads social- och krisjour (sosiaali- ja kriisipäivystys), som har öppet dygnet runt.
Telefonnumret till social- och krisjouren är (09) 8392 4005
linkkiVanda stad:
Social- och krisjourenfinska _ svenska _ engelska
Skyddshem
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta ett skyddshem (turvakoti).
Skyddshemmen har jourmottagning dygnet runt.
Skyddshemmet Mona är ett skyddshem avsett för invandrarkvinnor och deras barn.
Tfn 045 639 6274
Du kan även gå till Vanda skyddshem eller huvudstadsregionens skyddshem.
Tfn (09) 8392 0071
Steniusvägen 20
Tfn (09) 4777 180
linkkiTurvakoti Mona:
Skyddshemfinska
Skyddshemfinska _ engelska
Hjälp till offer för familjevåldfinska
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
De ungas skyddshus
Finlands Röda Kors De ungas skyddshus (Suomen Punaisen Ristin Nuorten turvatalo) ger stöd och hjälp i krissituationer för 12–19-åriga ungdomar.
Skyddshuset har öppet kl. 17–10, telefonjouren betjänar dygnet runt.
Sjukhusgatan 3 (Räckhals gård)
Tfn (09) 871 4043
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Bostadslöshet
Om du blir bostadslös ska du kontakta socialstationen (sosiaaliasema) för ditt eget område.
Kontaktuppgifterna hittar du på Vanda stads webbplats.
Om din hemkommun är Vanda, kan du få en bostad via Sininauha Oy eller Villenpirtti.
Läs mer: Bostadslöshet
linkkiVanda stad:
Socialtjänsterfinska _ svenska _ engelska
Bostäder för bostadslösafinska
Stödboende för personer med psykisk ohälsa och missbruksproblemfinska
Stöd- och serviceboende
Staden ordnar boendetjänster till exempel för åldringar och handikappade, som har svårt att klara av de dagliga sysslorna utan hjälp.
Åldringar och handikappade som inte klarar av att bo självständigt, kan bo i servicehus (palvelutalo) eller på en vårdinrättning (laitos).
Mer information om dessa tjänster får du från enheten för socialt arbete (sosiaalityön yksikkö) i ditt bostadsområde.
Läs mer: Stöd- och serviceboende.
linkkiVanda stad:
Information om hemvårdens stödtjänsterfinska
linkkiVanda stad:
Information om stadens servicebostäderfinska
linkkiVanda stad:
Privata servicehusfinska
linkkiVanda stad:
Socialtjänsterfinska _ svenska _ engelska
Bostadens avfallshantering
Information om var din närmaste återvinningsstation (kierrätyspiste) ligger hittar du på webbplatsen kierrätys.info.
Läs mer: Avfallshantering och återvinning.
linkkiAvfallsverksföreningen:
Återvinningsstationerfinska
linkkiHRM:
Återvinningsstationerfinska _ svenska _ engelska
Hyresbostad
Boende i en krissituation
Bostadslöshet
Stöd- och serviceboende
Bostadens avfallshantering
Hyresbostad
Hyresbostäderna är ofta dyra i huvudstadsregionen.
Du är själv ansvarig för att skaffa bostad åt dig själv.
Varken staden eller andra hyresvärdar har skyldighet att erbjuda dig bostad.
Läs mer: Hyresbostad.
Privata hyresbostäder
I Vanda finns också många andra hyresvärdar, varav de största är VVO, Sato och Avara.
Därtill ägs hyresbostäder i Vanda av många försäkringsbolag, Kuntien eläkevakuutus och Kunta-asunnot.
Det kan gå snabbt att få bostad via en privat hyresvärd.
Om du är studerande kan du ansöka om en hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS (Helsingin seudun Opiskelija-asuntosäätiö HOAS).
Om du är yngre än 30 år, kan du söka bostad hos Förbundet för ungdomsbostäder (Nuorisoasuntoliitto) och stiftelsen Nuorisosäätiö (Nuorisosäätiö).
linkkiSATO:
Hyresbostäderfinska _ engelska
linkkiAvara:
Hyresbostäderfinska
linkkiKommunbostäder:
Hyresbostäderfinska _ svenska _ engelska
linkkiFörbundet för ungdomsbostäder:
Hyresbostäder för personer under 30 årfinska _ engelska
Hyresbostäder för ungafinska _ engelska
linkkiHOAS:
Hyresbostäder för studerandefinska _ svenska _ engelska
Stadens hyresbostäder
Stadens hyresbostäder är vanligtvis förmånligare än de bostäder som hyrs ut av företag och privatpersoner.
Väntetiden för dessa bostäder kan dock vara lång och endast en liten del av de sökande får en bostad.
Vanda stads hyresbostäder ägs och hyrs ut av VAV Asunnot Oy.
Lokgränden 7
Tfn 010 235 1450 (kundtjänst)
Du kan göra en bostadsansökan på VAV Asunnot Oy:s webbplats.
Ansökan är giltig i fyra månader och måste sedan förnyas.
Vid val av invånare till stadens hyresbostäder prioriteras de sökande som har ett akut bostadsbehov.
Också sökandens inkomster beaktas, eftersom bostäderna främst är avsedda för personer med låga inkomster.
Information om stadens hyresbostäderfinska _ engelska
Ansökan om hyresbostad i stadenfinska _ engelska
Boende i en krissituation
Om din bostad har skadats till exempel till följd av brand eller vattenskada kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
Kontakta ditt försäkringsbolag direkt när skadan har inträffat.
I krissituationer får man även hjälp vid Vanda stads social- och krisjour (sosiaali- ja kriisipäivystys), som har öppet dygnet runt.
Telefonnumret till social- och krisjouren är (09) 8392 4005
linkkiVanda stad:
Social- och krisjourenfinska _ svenska _ engelska
Skyddshem
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta ett skyddshem (turvakoti).
Skyddshemmen har jourmottagning dygnet runt.
Skyddshemmet Mona är ett skyddshem avsett för invandrarkvinnor och deras barn.
Tfn 045 639 6274
Du kan även gå till Vanda skyddshem eller huvudstadsregionens skyddshem.
Tfn (09) 8392 0071
Steniusvägen 20
Tfn (09) 4777 180
linkkiTurvakoti Mona:
Skyddshemfinska
Skyddshemfinska _ engelska
Hjälp till offer för familjevåldfinska
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
De ungas skyddshus
Finlands Röda Kors De ungas skyddshus (Suomen Punaisen Ristin Nuorten turvatalo) ger stöd och hjälp i krissituationer för 12–19-åriga ungdomar.
Skyddshuset har öppet kl. 17–10, telefonjouren betjänar dygnet runt.
Sjukhusgatan 3 (Räckhals gård)
Tfn (09) 871 4043
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Bostadslöshet
Om du blir bostadslös ska du kontakta socialstationen (sosiaaliasema) för ditt eget område.
Kontaktuppgifterna hittar du på Vanda stads webbplats.
Om din hemkommun är Vanda, kan du få en bostad via Sininauha Oy eller Villenpirtti.
Läs mer: Bostadslöshet
linkkiVanda stad:
Socialtjänsterfinska _ svenska _ engelska
Bostäder för bostadslösafinska
Stödboende för personer med psykisk ohälsa och missbruksproblemfinska
Stöd- och serviceboende
Staden ordnar boendetjänster till exempel för åldringar och handikappade, som har svårt att klara av de dagliga sysslorna utan hjälp.
Åldringar och handikappade som inte klarar av att bo självständigt, kan bo i servicehus (palvelutalo) eller på en vårdinrättning (laitos).
Mer information om dessa tjänster får du från enheten för socialt arbete (sosiaalityön yksikkö) i ditt bostadsområde.
Läs mer: Stöd- och serviceboende.
linkkiVanda stad:
Information om hemvårdens stödtjänsterfinska
linkkiVanda stad:
Information om stadens servicebostäderfinska
linkkiVanda stad:
Privata servicehusfinska
linkkiVanda stad:
Socialtjänsterfinska _ svenska _ engelska
Bostadens avfallshantering
Information om var din närmaste återvinningsstation (kierrätyspiste) ligger hittar du på webbplatsen kierrätys.info.
Läs mer: Avfallshantering och återvinning.
linkkiAvfallsverksföreningen:
Återvinningsstationerfinska
linkkiHRM:
Återvinningsstationerfinska _ svenska _ engelska
Hyresbostad
Boende i en krissituation
Bostadslöshet
Stöd- och serviceboende
Bostadens avfallshantering
Hyresbostad
Hyresbostäderna är ofta dyra i huvudstadsregionen.
Du är själv ansvarig för att skaffa bostad åt dig själv.
Varken staden eller andra hyresvärdar har skyldighet att erbjuda dig bostad.
Läs mer: Hyresbostad.
Privata hyresbostäder
I Vanda finns också många andra hyresvärdar, varav de största är VVO, Sato och Avara.
Därtill ägs hyresbostäder i Vanda av många försäkringsbolag, Kuntien eläkevakuutus och Kunta-asunnot.
Det kan gå snabbt att få bostad via en privat hyresvärd.
Om du är studerande kan du ansöka om en hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS (Helsingin seudun Opiskelija-asuntosäätiö HOAS).
Om du är yngre än 30 år, kan du söka bostad hos Förbundet för ungdomsbostäder (Nuorisoasuntoliitto) och stiftelsen Nuorisosäätiö (Nuorisosäätiö).
linkkiSATO:
Hyresbostäderfinska _ engelska
linkkiAvara:
Hyresbostäderfinska
linkkiKommunbostäder:
Hyresbostäderfinska _ svenska _ engelska
linkkiFörbundet för ungdomsbostäder:
Hyresbostäder för personer under 30 årfinska _ engelska
Hyresbostäder för ungafinska _ engelska
linkkiHOAS:
Hyresbostäder för studerandefinska _ svenska _ engelska
Stadens hyresbostäder
Stadens hyresbostäder är vanligtvis förmånligare än de bostäder som hyrs ut av företag och privatpersoner.
Väntetiden för dessa bostäder kan dock vara lång och endast en liten del av de sökande får en bostad.
Vanda stads hyresbostäder ägs och hyrs ut av VAV Asunnot Oy.
Lokgränden 7
Tfn 010 235 1450 (kundtjänst)
Du kan göra en bostadsansökan på VAV Asunnot Oy:s webbplats.
Ansökan är giltig i fyra månader och måste sedan förnyas.
Vid val av invånare till stadens hyresbostäder prioriteras de sökande som har ett akut bostadsbehov.
Också sökandens inkomster beaktas, eftersom bostäderna främst är avsedda för personer med låga inkomster.
Information om stadens hyresbostäderfinska _ engelska
Ansökan om hyresbostad i stadenfinska _ engelska
Boende i en krissituation
Om din bostad har skadats till exempel till följd av brand eller vattenskada kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
Kontakta ditt försäkringsbolag direkt när skadan har inträffat.
I krissituationer får man även hjälp vid Vanda stads social- och krisjour (sosiaali- ja kriisipäivystys), som har öppet dygnet runt.
Telefonnumret till social- och krisjouren är (09) 8392 4005
linkkiVanda stad:
Social- och krisjourenfinska _ svenska _ engelska
Skyddshem
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta ett skyddshem (turvakoti).
Skyddshemmen har jourmottagning dygnet runt.
Skyddshemmet Mona är ett skyddshem avsett för invandrarkvinnor och deras barn.
Tfn 045 639 6274
Du kan även gå till Vanda skyddshem eller huvudstadsregionens skyddshem.
Tfn (09) 8392 0071
Steniusvägen 20
Tfn (09) 4777 180
linkkiTurvakoti Mona:
Skyddshemfinska
Skyddshemfinska _ engelska
Hjälp till offer för familjevåldfinska
Hjälp och stöd för invandrarkvinnorfinska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
De ungas skyddshus
Finlands Röda Kors De ungas skyddshus (Suomen Punaisen Ristin Nuorten turvatalo) ger stöd och hjälp i krissituationer för 12–19-åriga ungdomar.
Skyddshuset har öppet kl. 17–10, telefonjouren betjänar dygnet runt.
Sjukhusgatan 3 (Räckhals gård)
Tfn (09) 871 4043
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Bostadslöshet
Om du blir bostadslös ska du kontakta socialstationen (sosiaaliasema) för ditt eget område.
Kontaktuppgifterna hittar du på Vanda stads webbplats.
Om din hemkommun är Vanda, kan du få en bostad via Sininauha Oy eller Villenpirtti.
Läs mer: Bostadslöshet
linkkiVanda stad:
Socialtjänsterfinska _ svenska _ engelska
Bostäder för bostadslösafinska
Stödboende för personer med psykisk ohälsa och missbruksproblemfinska
Stöd- och serviceboende
Staden ordnar boendetjänster till exempel för åldringar och handikappade, som har svårt att klara av de dagliga sysslorna utan hjälp.
Åldringar och handikappade som inte klarar av att bo självständigt, kan bo i servicehus (palvelutalo) eller på en vårdinrättning (laitos).
Mer information om dessa tjänster får du från enheten för socialt arbete (sosiaalityön yksikkö) i ditt bostadsområde.
Läs mer: Stöd- och serviceboende.
linkkiVanda stad:
Information om hemvårdens stödtjänsterfinska
linkkiVanda stad:
Information om stadens servicebostäderfinska
linkkiVanda stad:
Privata servicehusfinska
linkkiVanda stad:
Socialtjänsterfinska _ svenska _ engelska
Bostadens avfallshantering
Information om var din närmaste återvinningsstation (kierrätyspiste) ligger hittar du på webbplatsen kierrätys.info.
Läs mer: Avfallshantering och återvinning.
linkkiAvfallsverksföreningen:
Återvinningsstationerfinska
linkkiHRM:
Återvinningsstationerfinska _ svenska _ engelska
Möjligheter att studera det finska eller svenska språket
Språkkurser
Med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors, Vanda, Esbo eller Grankulla.
Kurserna i svenska hittar du genom att klicka på länken på tjänstens startsida.
Kurserna i tjänsten finnishcourses.fi är öppna för alla.
Tjänsten omfattar inte arbets- och näringsbyråns kurser.
I Vanda anordnas kurser i finska och svenska språket för invandrare av Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto) Kurserna vid institutet är öppna för alla.
Vuxenutbildningsinstitutet ligger i Dickursby, men kurser ordnas runtom i Vanda.
Adress:
Näckrosvägen 5
Tfn (09) 8392 4342
Ytterligare information om kurser och anmälan hittar du på Vanda vuxenutbildningsinstituts webbplats och i studiehandboken.
Du får studiehandboken till exempel på bibliotek eller Vandainfo samt i elektroniskt format på Vanda stads webbplats.
Arbets- och näringsbyrån anvisar invandrare till kurser i finska språket som ingår i integrationsprocessen.
I samband med att en integrations- eller sysselsättningsplan upprättas för dig, kan du också få också en studieplats på en finskakurs reserverad eller också kan du ställas i kö för en studieplats.
Mer information hittar du vid arbets- och näringsbyrån.
Läs mer: Studier i finska och svenska
Kurser i finska och svenska språketfinska _ engelska _ ryska
linkkiVanda vuxenutbildningsinstitut:
Kurser i finska och svenska språket för invandrarefinska
linkkiArbets- och näringsministeriet:
Utbildning i finska och svenska språketfinska _ svenska _ engelska
linkkiVanda vuxenutbildningsinstitut:
Grundundervisning för vuxnafinska
Samtal på finska
På Vanda stadsbibliotek anordnas språkcaféer (kielikahvila), där man kan öva på att prata finska.
Alla som vill lära sig tala finska är välkomna till caféerna.
På språkcaféerna talar vi finska, så det är bra om du redan kan lite finska.
Språkcaféerna är avgiftsfria.
Mer information om språkcaféerna får du från biblioteken.
I Vanda anordnas samtalsklubbar på finska också på Silkesportens verksamhetscenter (Silkinportin toimintakeskus) och Kafnettis och Myyrinkis boendeträffpunkter (Kafnetin ja Myyringin asukastila).
Finskaklubbar avsedda för föräldrar som vårdar barn i hemmet anordnas i invånarparkerna (asukaspuisto) och i de öppna daghemmen (avoin päiväkoti).
Klubbarna för att lära sig tala finska är avgiftsfria.
Läsundervisning
Nätverket Vi läser tillsammans (Luetaan yhdessä-verkosto) erbjuder undervisning i läsning och det finska språket för invandrarkvinnor.
Flera olika Vi läser tillsammans-nätverk är verksamma på olika håll i Vanda.
Det är avgiftsfritt att delta i grupperna.
Språkkaféerfinska _ engelska _ ryska
linkkiVanda stad:
Invånarlokalfinska _ engelska
linkkiVanda stad:
Invånarlokalfinska _ engelska
linkkiVanda stad:
Parker för invånare och öppna daghemfinska _ svenska _ engelska
linkkiVi läser tillsammans-nätverket:
Vi läser tillsammans i Vandafinska _ svenska _ engelska
Allmän språkexamen
Du kan avlägga allmän språkexamen i finska eller svenska språket.
På utbildningsstyrelsens (Opetushallitus) webbplats finns en sökmotor med vilken du kan kontrollera var och när du kan avlägga examen.
I Vanda ordnas språkexamina till exempel vid Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto).
Läs mer: Officiellt intyg på språkkunskaper.
linkkiUtbildningsstyrelsen:
Att anmäla sig till en allmän språkexamen och examensavgifterfinska _ svenska _ engelska
linkkiVanda vuxenutbildningsinstitut:
Allmän språkexamenfinska
linkkiUtbildningsstyrelsen:
Examenssökningfinska
Möjligheter att studera det finska eller svenska språket
Språkkurser
Med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors, Vanda, Esbo eller Grankulla.
Kurserna i svenska hittar du genom att klicka på länken på tjänstens startsida.
Kurserna i tjänsten finnishcourses.fi är öppna för alla.
Tjänsten omfattar inte arbets- och näringsbyråns kurser.
I Vanda anordnas kurser i finska och svenska språket för invandrare av Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto) Kurserna vid institutet är öppna för alla.
Vuxenutbildningsinstitutet ligger i Dickursby, men kurser ordnas runtom i Vanda.
Adress:
Näckrosvägen 5
Tfn (09) 8392 4342
Ytterligare information om kurser och anmälan hittar du på Vanda vuxenutbildningsinstituts webbplats och i studiehandboken.
Du får studiehandboken till exempel på bibliotek eller Vandainfo samt i elektroniskt format på Vanda stads webbplats.
Arbets- och näringsbyrån anvisar invandrare till kurser i finska språket som ingår i integrationsprocessen.
I samband med att en integrations- eller sysselsättningsplan upprättas för dig, kan du också få också en studieplats på en finskakurs reserverad eller också kan du ställas i kö för en studieplats.
Mer information hittar du vid arbets- och näringsbyrån.
Läs mer: Studier i finska och svenska
Kurser i finska och svenska språketfinska _ engelska _ ryska
linkkiVanda vuxenutbildningsinstitut:
Kurser i finska och svenska språket för invandrarefinska
linkkiArbets- och näringsministeriet:
Utbildning i finska och svenska språketfinska _ svenska _ engelska
linkkiVanda vuxenutbildningsinstitut:
Grundundervisning för vuxnafinska
Samtal på finska
På Vanda stadsbibliotek anordnas språkcaféer (kielikahvila), där man kan öva på att prata finska.
Alla som vill lära sig tala finska är välkomna till caféerna.
På språkcaféerna talar vi finska, så det är bra om du redan kan lite finska.
Språkcaféerna är avgiftsfria.
Mer information om språkcaféerna får du från biblioteken.
I Vanda anordnas samtalsklubbar på finska också på Silkesportens verksamhetscenter (Silkinportin toimintakeskus) och Kafnettis och Myyrinkis boendeträffpunkter (Kafnetin ja Myyringin asukastila).
Finskaklubbar avsedda för föräldrar som vårdar barn i hemmet anordnas i invånarparkerna (asukaspuisto) och i de öppna daghemmen (avoin päiväkoti).
Klubbarna för att lära sig tala finska är avgiftsfria.
Läsundervisning
Nätverket Vi läser tillsammans (Luetaan yhdessä-verkosto) erbjuder undervisning i läsning och det finska språket för invandrarkvinnor.
Flera olika Vi läser tillsammans-nätverk är verksamma på olika håll i Vanda.
Det är avgiftsfritt att delta i grupperna.
Språkkaféerfinska _ engelska _ ryska
linkkiVanda stad:
Invånarlokalfinska _ engelska
linkkiVanda stad:
Invånarlokalfinska _ engelska
linkkiVanda stad:
Parker för invånare och öppna daghemfinska _ svenska _ engelska
linkkiVi läser tillsammans-nätverket:
Vi läser tillsammans i Vandafinska _ svenska _ engelska
Allmän språkexamen
Du kan avlägga allmän språkexamen i finska eller svenska språket.
På utbildningsstyrelsens (Opetushallitus) webbplats finns en sökmotor med vilken du kan kontrollera var och när du kan avlägga examen.
I Vanda ordnas språkexamina till exempel vid Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto).
Läs mer: Officiellt intyg på språkkunskaper.
linkkiUtbildningsstyrelsen:
Att anmäla sig till en allmän språkexamen och examensavgifterfinska _ svenska _ engelska
linkkiVanda vuxenutbildningsinstitut:
Allmän språkexamenfinska
linkkiUtbildningsstyrelsen:
Examenssökningfinska
Möjligheter att studera det finska eller svenska språket
Språkkurser
Med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors, Vanda, Esbo eller Grankulla.
Kurserna i svenska hittar du genom att klicka på länken på tjänstens startsida.
Kurserna i tjänsten finnishcourses.fi är öppna för alla.
Tjänsten omfattar inte arbets- och näringsbyråns kurser.
I Vanda anordnas kurser i finska och svenska språket för invandrare av Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto) Kurserna vid institutet är öppna för alla.
Vuxenutbildningsinstitutet ligger i Dickursby, men kurser ordnas runtom i Vanda.
Adress:
Näckrosvägen 5
Tfn (09) 8392 4342
Ytterligare information om kurser och anmälan hittar du på Vanda vuxenutbildningsinstituts webbplats och i studiehandboken.
Du får studiehandboken till exempel på bibliotek eller Vandainfo samt i elektroniskt format på Vanda stads webbplats.
Arbets- och näringsbyrån anvisar invandrare till kurser i finska språket som ingår i integrationsprocessen.
I samband med att en integrations- eller sysselsättningsplan upprättas för dig, kan du också få också en studieplats på en finskakurs reserverad eller också kan du ställas i kö för en studieplats.
Mer information hittar du vid arbets- och näringsbyrån.
Läs mer: Studier i finska och svenska
Kurser i finska och svenska språketfinska _ engelska _ ryska
linkkiVanda vuxenutbildningsinstitut:
Kurser i finska och svenska språket för invandrarefinska
linkkiArbets- och näringsministeriet:
Utbildning i finska och svenska språketfinska _ svenska _ engelska
linkkiVanda vuxenutbildningsinstitut:
Grundundervisning för vuxnafinska
Samtal på finska
På Vanda stadsbibliotek anordnas språkcaféer (kielikahvila), där man kan öva på att prata finska.
Alla som vill lära sig tala finska är välkomna till caféerna.
På språkcaféerna talar vi finska, så det är bra om du redan kan lite finska.
Språkcaféerna är avgiftsfria.
Mer information om språkcaféerna får du från biblioteken.
I Vanda anordnas samtalsklubbar på finska också på Silkesportens verksamhetscenter (Silkinportin toimintakeskus) och Kafnettis och Myyrinkis boendeträffpunkter (Kafnetin ja Myyringin asukastila).
Finskaklubbar avsedda för föräldrar som vårdar barn i hemmet anordnas i invånarparkerna (asukaspuisto) och i de öppna daghemmen (avoin päiväkoti).
Klubbarna för att lära sig tala finska är avgiftsfria.
Läsundervisning
Nätverket Vi läser tillsammans (Luetaan yhdessä-verkosto) erbjuder undervisning i läsning och det finska språket för invandrarkvinnor.
Flera olika Vi läser tillsammans-nätverk är verksamma på olika håll i Vanda.
Det är avgiftsfritt att delta i grupperna.
Språkkaféerfinska _ engelska _ ryska
linkkiVanda stad:
Invånarlokalfinska _ engelska
linkkiVanda stad:
Invånarlokalfinska _ engelska
linkkiVanda stad:
Parker för invånare och öppna daghemfinska _ svenska _ engelska
linkkiVi läser tillsammans-nätverket:
Vi läser tillsammans i Vandafinska _ svenska _ engelska
Allmän språkexamen
Du kan avlägga allmän språkexamen i finska eller svenska språket.
På utbildningsstyrelsens (Opetushallitus) webbplats finns en sökmotor med vilken du kan kontrollera var och när du kan avlägga examen.
I Vanda ordnas språkexamina till exempel vid Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto).
Läs mer: Officiellt intyg på språkkunskaper.
linkkiUtbildningsstyrelsen:
Att anmäla sig till en allmän språkexamen och examensavgifterfinska _ svenska _ engelska
linkkiVanda vuxenutbildningsinstitut:
Allmän språkexamenfinska
linkkiUtbildningsstyrelsen:
Examenssökningfinska
Var hittar jag jobb?
Hjälp med jobbsökningen
Att starta ett företag
Beskattning
Var hittar jag jobb?
TE-byrån (TE-toimisto) hjälper dig att söka arbete.
Om du är arbetslös och söker efter arbete, ska du anmäla dig som arbetssökande hos TE-byrån.
Du kan anmäla dig antingen via nättjänsten eller personligen hos TE-byrån.
Medborgare i EU-länderna, Island, Liechtenstein och Schweiz kan anmäla sig som arbetssökande via TE-byråns nättjänst.
Övriga länders medborgare måste anmäla sig personligen hos TE-byrån.
Ta med dig din legitimation och ditt uppehållstillstånd.
Kontaktuppgifter:
Information om TE-byråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös.
Information om att söka arbete i Finland hittar du på InfoFinlands sida: Var hittar jag jobb?
linkkiVanda arbets- och näringsbyrå:
Kontaktuppgifter och tjänsterfinska _ svenska
linkkiArbets- och näringsministeriet:
Lediga jobbfinska _ svenska
linkkiArbets- och näringsförvaltningen:
Länkar till jobbsajterfinska _ svenska _ engelska
linkkiVanda stad:
Stöd för att hitta sysselsättningfinska _ svenska _ engelska
Hjälp med jobbsökningen
Stadens tjänster för arbetssökande
Vanda stad tillhandahåller olika tjänster för arbetslösa som hjälper dem att få kontakt med arbetslivet och hitta jobb.
I Vanda ordnas även många rekryteringsevenemang där arbetsgivarna söker arbetstagare.
Du hittar mer information om stadens tjänster på Vanda stads webbplats.
linkkiVanda stad:
Stadens tjänster för arbetssökandefinska _ svenska _ engelska
Om du behöver hjälp med jobbsökningen eller med att hitta en studieplats kan du kontakta rådgivarna i Håkansböle internationella förenings Tsemppari-projekt.
Du hittar kontaktuppgifterna på Håkansböle internationella förenings webbplats.
Integrationscentret Kotoutumiskeskus Monika hjälper arbetslösa invandrarkvinnor att hitta jobb.
Du kan få hjälp med att skriva din CV eller en jobbansökan, studera vardagsfinska och digitala färdigheter.
Luckan integration
Luckan Integration är en rådgivningstjänst, som erbjuder personlig rådgivning för invandrare och anordnar bland annat evenemang och grupper relaterade till jobbsökning.
Språket som talas vid träffarna är engelska.
Råd om jobbsökningfinska _ svenska _ engelska _ spanska
Väestöliittos karriärmentorskap är avsett för utbildade invandrare.
Via programmet kan du få en mentor, som stödjer dig i sökningen efter arbete eller utbildningsplats eller i att starta eget företag.
Verksamheten sker på finska.
Mentorskap i fråga om arbetskarriärfinska _ engelska
Om du är under 30 år, kan du få råd och handledning via tjänsten Navigatorn.
Personalen vid Navigatorn hjälper dig om du inte har något arbete eller en studieplats.
Stödföreningen för unga invandrare R3 (R3 Maahanmuuttajanuorten tuki ry) hjälper ungdomar i frågor som rör utbildning och sysselsättning.
Mer information hittar du på föreningens webbplats.
Stöd för unga invandrarefinska
Att starta ett företag
Om du har ett företag i Vanda, kan du bli medlem i Vanda Företagare.
Vanda Företagare rf är företagarnas intressebevakningsorganisation som erbjuder sina medlemmar till exempel utbildning och rådgivning.
Mer information hittar du på föreningens webbplats.
NewCo Helsinki erbjuder rådgivning och hjälp med att starta eget företag på finska, svenska, engelska, ryska, arabiska, estniska, tyska och italienska.
Vid NewCo Helsinki ordnas informationsmöten om att starta eget för invandrare på finska, engelska, ryska, arabiska och estniska.
Infomötena är avgiftsfria.
NewCo Helsinki ordnar företagarutbildningar på finska, engelska och ryska.
En del av kurserna är avsedda för personer som ska starta eget företag och en del för dem som redan har eget företag.
Kurser hålls på finska, engelska och ryska.
Mer information och anmälan finns på NewCo Helsinki webbplats.
Nylands TE-byrå (TE-toimisto) erbjuder mångsidiga tjänster för personer som funderar på att starta eget och dem som är på väg att starta eget.
På Nylands TE-byrå kan du till exempel delta i företagarutbildning och söka startpeng för att starta eget företag.
Läs mer: Att grunda ett företag
Tjänster för företagare med invandrarbakgrundfinska _ engelska
linkkiFöretagsFinland:
Företagsrådgivningfinska _ svenska _ engelska
Företagsrådgivningfinska _ engelska
Företagarnas intressebevakningsorganisationfinska
Beskattning
Huvudstadsregionens skattebyrå betjänar kunderna i centrala Helsingfors.
Kontaktuppgifter:
Alexandersgatan 9 (Gloet)
Tfn: 029 512 000
Invandrare kan även sköta ärenden vid servicestället International House Helsinki.
På servicestället hjälper FPA:s och Skatteförvaltningens experter invandrare som kommer till Finland för att arbeta i frågor som rör beskattning och social trygghet
Kontaktuppgifter till servicestället International House Helsinki:
Albertinkatu 25
Läs mer: Beskattning
linkkiSkatteförvaltningen:
Kontaktuppgifterfinska _ svenska _ engelska
Rådgivning om social trygghet och beskattningfinska _ svenska _ engelska
IHH – serviceställe för dig som flyttar till Finland engelska
Var hittar jag jobb?
Hjälp med jobbsökningen
Att starta ett företag
Beskattning
Var hittar jag jobb?
TE-byrån (TE-toimisto) hjälper dig att söka arbete.
Om du är arbetslös och söker efter arbete, ska du anmäla dig som arbetssökande hos TE-byrån.
Du kan anmäla dig antingen via nättjänsten eller personligen hos TE-byrån.
Medborgare i EU-länderna, Island, Liechtenstein och Schweiz kan anmäla sig som arbetssökande via TE-byråns nättjänst.
Övriga länders medborgare måste anmäla sig personligen hos TE-byrån.
Ta med dig din legitimation och ditt uppehållstillstånd.
Kontaktuppgifter:
Information om TE-byråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös.
Information om att söka arbete i Finland hittar du på InfoFinlands sida: Var hittar jag jobb?
linkkiVanda arbets- och näringsbyrå:
Kontaktuppgifter och tjänsterfinska _ svenska
linkkiArbets- och näringsministeriet:
Lediga jobbfinska _ svenska
linkkiArbets- och näringsförvaltningen:
Länkar till jobbsajterfinska _ svenska _ engelska
linkkiVanda stad:
Stöd för att hitta sysselsättningfinska _ svenska _ engelska
Hjälp med jobbsökningen
Stadens tjänster för arbetssökande
Vanda stad tillhandahåller olika tjänster för arbetslösa som hjälper dem att få kontakt med arbetslivet och hitta jobb.
I Vanda ordnas även många rekryteringsevenemang där arbetsgivarna söker arbetstagare.
Du hittar mer information om stadens tjänster på Vanda stads webbplats.
linkkiVanda stad:
Stadens tjänster för arbetssökandefinska _ svenska _ engelska
Om du behöver hjälp med jobbsökningen eller med att hitta en studieplats kan du kontakta rådgivarna i Håkansböle internationella förenings Tsemppari-projekt.
Du hittar kontaktuppgifterna på Håkansböle internationella förenings webbplats.
Integrationscentret Kotoutumiskeskus Monika hjälper arbetslösa invandrarkvinnor att hitta jobb.
Du kan få hjälp med att skriva din CV eller en jobbansökan, studera vardagsfinska och digitala färdigheter.
Luckan integration
Luckan Integration är en rådgivningstjänst, som erbjuder personlig rådgivning för invandrare och anordnar bland annat evenemang och grupper relaterade till jobbsökning.
Språket som talas vid träffarna är engelska.
Råd om jobbsökningfinska _ svenska _ engelska _ spanska
Väestöliittos karriärmentorskap är avsett för utbildade invandrare.
Via programmet kan du få en mentor, som stödjer dig i sökningen efter arbete eller utbildningsplats eller i att starta eget företag.
Verksamheten sker på finska.
Mentorskap i fråga om arbetskarriärfinska _ engelska
Om du är under 30 år, kan du få råd och handledning via tjänsten Navigatorn.
Personalen vid Navigatorn hjälper dig om du inte har något arbete eller en studieplats.
Stödföreningen för unga invandrare R3 (R3 Maahanmuuttajanuorten tuki ry) hjälper ungdomar i frågor som rör utbildning och sysselsättning.
Mer information hittar du på föreningens webbplats.
Stöd för unga invandrarefinska
Att starta ett företag
Om du har ett företag i Vanda, kan du bli medlem i Vanda Företagare.
Vanda Företagare rf är företagarnas intressebevakningsorganisation som erbjuder sina medlemmar till exempel utbildning och rådgivning.
Mer information hittar du på föreningens webbplats.
NewCo Helsinki erbjuder rådgivning och hjälp med att starta eget företag på finska, svenska, engelska, ryska, arabiska, estniska, tyska och italienska.
Vid NewCo Helsinki ordnas informationsmöten om att starta eget för invandrare på finska, engelska, ryska, arabiska och estniska.
Infomötena är avgiftsfria.
NewCo Helsinki ordnar företagarutbildningar på finska, engelska och ryska.
En del av kurserna är avsedda för personer som ska starta eget företag och en del för dem som redan har eget företag.
Kurser hålls på finska, engelska och ryska.
Mer information och anmälan finns på NewCo Helsinki webbplats.
Nylands TE-byrå (TE-toimisto) erbjuder mångsidiga tjänster för personer som funderar på att starta eget och dem som är på väg att starta eget.
På Nylands TE-byrå kan du till exempel delta i företagarutbildning och söka startpeng för att starta eget företag.
Läs mer: Att grunda ett företag
Tjänster för företagare med invandrarbakgrundfinska _ engelska
linkkiFöretagsFinland:
Företagsrådgivningfinska _ svenska _ engelska
Företagsrådgivningfinska _ engelska
Företagarnas intressebevakningsorganisationfinska
Beskattning
Huvudstadsregionens skattebyrå betjänar kunderna i centrala Helsingfors.
Kontaktuppgifter:
Alexandersgatan 9 (Gloet)
Tfn: 029 512 000
Invandrare kan även sköta ärenden vid servicestället International House Helsinki.
På servicestället hjälper FPA:s och Skatteförvaltningens experter invandrare som kommer till Finland för att arbeta i frågor som rör beskattning och social trygghet
Kontaktuppgifter till servicestället International House Helsinki:
Albertinkatu 25
Läs mer: Beskattning
linkkiSkatteförvaltningen:
Kontaktuppgifterfinska _ svenska _ engelska
Rådgivning om social trygghet och beskattningfinska _ svenska _ engelska
IHH – serviceställe för dig som flyttar till Finland engelska
Var hittar jag jobb?
Hjälp med jobbsökningen
Att starta ett företag
Beskattning
Var hittar jag jobb?
TE-byrån (TE-toimisto) hjälper dig att söka arbete.
Om du är arbetslös och söker efter arbete, ska du anmäla dig som arbetssökande hos TE-byrån.
Du kan anmäla dig antingen via nättjänsten eller personligen hos TE-byrån.
Medborgare i EU-länderna, Island, Liechtenstein och Schweiz kan anmäla sig som arbetssökande via TE-byråns nättjänst.
Övriga länders medborgare måste anmäla sig personligen hos TE-byrån.
Ta med dig din legitimation och ditt uppehållstillstånd.
Kontaktuppgifter:
Information om TE-byråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös.
Information om att söka arbete i Finland hittar du på InfoFinlands sida: Var hittar jag jobb?
linkkiVanda arbets- och näringsbyrå:
Kontaktuppgifter och tjänsterfinska _ svenska
linkkiArbets- och näringsministeriet:
Lediga jobbfinska _ svenska
linkkiArbets- och näringsförvaltningen:
Länkar till jobbsajterfinska _ svenska _ engelska
linkkiVanda stad:
Stöd för att hitta sysselsättningfinska _ svenska _ engelska
Hjälp med jobbsökningen
Stadens tjänster för arbetssökande
Vanda stad tillhandahåller olika tjänster för arbetslösa som hjälper dem att få kontakt med arbetslivet och hitta jobb.
I Vanda ordnas även många rekryteringsevenemang där arbetsgivarna söker arbetstagare.
Du hittar mer information om stadens tjänster på Vanda stads webbplats.
linkkiVanda stad:
Stadens tjänster för arbetssökandefinska _ svenska _ engelska
Om du behöver hjälp med jobbsökningen eller med att hitta en studieplats kan du kontakta rådgivarna i Håkansböle internationella förenings Tsemppari-projekt.
Du hittar kontaktuppgifterna på Håkansböle internationella förenings webbplats.
Integrationscentret Kotoutumiskeskus Monika hjälper arbetslösa invandrarkvinnor att hitta jobb.
Du kan få hjälp med att skriva din CV eller en jobbansökan, studera vardagsfinska och digitala färdigheter.
Luckan integration
Luckan Integration är en rådgivningstjänst, som erbjuder personlig rådgivning för invandrare och anordnar bland annat evenemang och grupper relaterade till jobbsökning.
Språket som talas vid träffarna är engelska.
Råd om jobbsökningfinska _ svenska _ engelska _ spanska
Väestöliittos karriärmentorskap är avsett för utbildade invandrare.
Via programmet kan du få en mentor, som stödjer dig i sökningen efter arbete eller utbildningsplats eller i att starta eget företag.
Verksamheten sker på finska.
Mentorskap i fråga om arbetskarriärfinska _ engelska
Om du är under 30 år, kan du få råd och handledning via tjänsten Navigatorn.
Personalen vid Navigatorn hjälper dig om du inte har något arbete eller en studieplats.
Stödföreningen för unga invandrare R3 (R3 Maahanmuuttajanuorten tuki ry) hjälper ungdomar i frågor som rör utbildning och sysselsättning.
Mer information hittar du på föreningens webbplats.
Stöd för unga invandrarefinska
Att starta ett företag
Om du har ett företag i Vanda, kan du bli medlem i Vanda Företagare.
Vanda Företagare rf är företagarnas intressebevakningsorganisation som erbjuder sina medlemmar till exempel utbildning och rådgivning.
Mer information hittar du på föreningens webbplats.
NewCo Helsinki erbjuder rådgivning och hjälp med att starta eget företag på finska, svenska, engelska, ryska, arabiska, estniska, tyska och italienska.
Vid NewCo Helsinki ordnas informationsmöten om att starta eget för invandrare på finska, engelska, ryska, arabiska och estniska.
Infomötena är avgiftsfria.
NewCo Helsinki ordnar företagarutbildningar på finska, engelska och ryska.
En del av kurserna är avsedda för personer som ska starta eget företag och en del för dem som redan har eget företag.
Kurser hålls på finska, engelska och ryska.
Mer information och anmälan finns på NewCo Helsinki webbplats.
Nylands TE-byrå (TE-toimisto) erbjuder mångsidiga tjänster för personer som funderar på att starta eget och dem som är på väg att starta eget.
På Nylands TE-byrå kan du till exempel delta i företagarutbildning och söka startpeng för att starta eget företag.
Läs mer: Att grunda ett företag
Tjänster för företagare med invandrarbakgrundfinska _ engelska
linkkiFöretagsFinland:
Företagsrådgivningfinska _ svenska _ engelska
Företagsrådgivningfinska _ engelska
Företagarnas intressebevakningsorganisationfinska
Beskattning
Huvudstadsregionens skattebyrå betjänar kunderna i centrala Helsingfors.
Kontaktuppgifter:
Alexandersgatan 9 (Gloet)
Tfn: 029 512 000
Invandrare kan även sköta ärenden vid servicestället International House Helsinki.
På servicestället hjälper FPA:s och Skatteförvaltningens experter invandrare som kommer till Finland för att arbeta i frågor som rör beskattning och social trygghet
Kontaktuppgifter till servicestället International House Helsinki:
Albertinkatu 25
Läs mer: Beskattning
linkkiSkatteförvaltningen:
Kontaktuppgifterfinska _ svenska _ engelska
Rådgivning om social trygghet och beskattningfinska _ svenska _ engelska
IHH – serviceställe för dig som flyttar till Finland engelska
Rådgivning för och integration av invandrare
Inledande kartläggning
Behöver du en tolk?
Rådgivning för och integration av invandrare
Invandrartjänster
Vanda stads tjänster för invandrare omfattar
mottagningstjänster för invandrare
integrationstjänster
Vanda stads tjänster för invandrare (Vantaan maahanmuuttajapalvelut) ger dig information om integration, social- och hälsovårdstjänster och om stadens och olika organisationers tjänster.
Du kan bli klient om du flyttat till Finland på grund av familjeband, är flykting, offer för människohandel eller har rätt till en inledande kartläggning.
Tfn (09) 839 21074 och (09) 839 32042
linkkiVanda stad:
Invandrartjänsterfinska _ engelska
Verksamhetscentret Silkesporten (Silkinportin toimintakeskus) ger rådgivning för invandrare och där ordnas många slags aktiviteter.
dickursbyvägen 44 F, vån.
Tfn (09) 839 23651
linkkiSilkesportens verksamhetscenter:
Rådgivning och verksamhet för invandrarefinska _ engelska
Vandainfo ger dig information om såväl Vandas stads som statens tjänster.
Vandainfon finns i Dickursby, Korso och Myrbacka.
Adresserna är:
Dixi, Banvägen 11, 2:a vån.
tfn (09) 839 22133
Tfn (09) 839 22133
Tfn (09) 839 22133
Kontaktuppgifterna och öppettiderna hittar du på Vanda stads webbplats.
linkkiVanda stad:
Vandainfofinska _ svenska _ engelska
Den internationella föreningen i Håkansböle (Hakunilan kansainvälinen yhdistys) har en rådgivningspunkt som betjänar invandrare i Håkansböle, Björkby och andra områden i Vanda, som vill ha information om till exempel studier, språkkurser, arbete, hobbyverksamhet, krissituationer eller juridiska frågor.
Sporrgränden 2 A, vån. 3 (Håkansböle)
Tfn (09) 272 2775 och 040 501 3199.
linkkiInternationella föreningen i Håkansböle:
Rådgivning för invandrarefinska _ engelska _ ryska _ somaliska _ arabiska
På invandrarrådgivningen vid föreningen Vantaan Järjestörinki ry (Vantaan Järjestörinki ry:n Maahanmuuttajien neuvontapiste) kan du fråga om sådant som rör till exempel arbetslivet, social trygghet, hälsa, utbildning och uppehållstillstånd.
Adress:
Ranunkelvägen 22
Asukastila Myyrinki
Eldstadstorget 1 eller Kopparbergsvägen 10 B, vån.
Vanda Tfn (09) 839 35703 och 040 183 0930
Rautbergsgatan 3
Tfn 045 134 1711
Rådgivning för invandrarefinska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
IHH – serviceställe för dig som flyttar till Finland engelska
Inledande kartläggning
Den inledande kartläggningen (alkukartoitus) hjälper dig att hitta lämpliga tjänster i din hemstad.
Vanda stad eller Nylands TE-byrå ordnar en inledande kartläggning för varje ny invandrare i Vanda.
Du har rätt att få en inledande kartläggning om
din hemkommun är Vanda
du har flyttat till Vanda från ett annat land eller en annan ort i Finland
någon inledande kartläggning inte har gjorts för dig tidigare
du har haft hemkommun i Finland i högst tre år.
I den inledande kartläggningen får du information om utbildning i finska eller svenska, arbetssökning, utbildning och tjänster i Vanda.
Vid den inledande kartläggningen talas man vid med hjälp av tolk.
Den inledande kartläggningen är avgiftsfri.
Begäran om inledande kartläggning
Du kan begära en inledande kartläggning via e-post eller så kan du boka en tid per telefon.
Tfn 09 839 32622, 09 839 27525 eller 09 839 31766
Om du söker arbete, bör du anmäla dig till TE-byrån.
TE-byrån gör den inledande kartläggningen.
Läs mer om den inledande kartläggningen och integrationsplanen på InfoFinlands webbplats Integration i Finland
linkkiVanda stad:
Inledande kartläggningfinska _ engelska
Behöver du en tolk?
Om du måste sköta ärenden med myndigheter, men inte kan finska eller svenska och det inte heller finns något annat språk som både du och myndigheten talar, kan du använda en tolktjänst.
Meddela alltid myndigheten i förväg om du behöver en tolk.
Myndigheten bokar tolken och då får du tolkningstjänsten gratis.
Om du själv bokar tolken och betalar kostnaderna, kan du anlita en tolk när som helst.
Läs mer: Behöver du en tolk?
linkkiVanda stad:
Information om tolktjänsterfinska
linkkiFinlands översättar- och tolkförbund:
Sök tolk eller översättarefinska _ svenska _ engelska
Rådgivning för och integration av invandrare
Inledande kartläggning
Behöver du en tolk?
Rådgivning för och integration av invandrare
Invandrartjänster
Vanda stads tjänster för invandrare omfattar
mottagningstjänster för invandrare
integrationstjänster
Vanda stads tjänster för invandrare (Vantaan maahanmuuttajapalvelut) ger dig information om integration, social- och hälsovårdstjänster och om stadens och olika organisationers tjänster.
Du kan bli klient om du flyttat till Finland på grund av familjeband, är flykting, offer för människohandel eller har rätt till en inledande kartläggning.
Tfn (09) 839 21074 och (09) 839 32042
linkkiVanda stad:
Invandrartjänsterfinska _ engelska
Verksamhetscentret Silkesporten (Silkinportin toimintakeskus) ger rådgivning för invandrare och där ordnas många slags aktiviteter.
dickursbyvägen 44 F, vån.
Tfn (09) 839 23651
linkkiSilkesportens verksamhetscenter:
Rådgivning och verksamhet för invandrarefinska _ engelska
Vandainfo ger dig information om såväl Vandas stads som statens tjänster.
Vandainfon finns i Dickursby, Korso och Myrbacka.
Adresserna är:
Dixi, Banvägen 11, 2:a vån.
tfn (09) 839 22133
Tfn (09) 839 22133
Tfn (09) 839 22133
Kontaktuppgifterna och öppettiderna hittar du på Vanda stads webbplats.
linkkiVanda stad:
Vandainfofinska _ svenska _ engelska
Den internationella föreningen i Håkansböle (Hakunilan kansainvälinen yhdistys) har en rådgivningspunkt som betjänar invandrare i Håkansböle, Björkby och andra områden i Vanda, som vill ha information om till exempel studier, språkkurser, arbete, hobbyverksamhet, krissituationer eller juridiska frågor.
Sporrgränden 2 A, vån. 3 (Håkansböle)
Tfn (09) 272 2775 och 040 501 3199.
linkkiInternationella föreningen i Håkansböle:
Rådgivning för invandrarefinska _ engelska _ ryska _ somaliska _ arabiska
På invandrarrådgivningen vid föreningen Vantaan Järjestörinki ry (Vantaan Järjestörinki ry:n Maahanmuuttajien neuvontapiste) kan du fråga om sådant som rör till exempel arbetslivet, social trygghet, hälsa, utbildning och uppehållstillstånd.
Adress:
Ranunkelvägen 22
Asukastila Myyrinki
Eldstadstorget 1 eller Kopparbergsvägen 10 B, vån.
Vanda Tfn (09) 839 35703 och 040 183 0930
Rautbergsgatan 3
Tfn 045 134 1711
Rådgivning för invandrarefinska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
IHH – serviceställe för dig som flyttar till Finland engelska
Inledande kartläggning
Den inledande kartläggningen (alkukartoitus) hjälper dig att hitta lämpliga tjänster i din hemstad.
Vanda stad eller Nylands TE-byrå ordnar en inledande kartläggning för varje ny invandrare i Vanda.
Du har rätt att få en inledande kartläggning om
din hemkommun är Vanda
du har flyttat till Vanda från ett annat land eller en annan ort i Finland
någon inledande kartläggning inte har gjorts för dig tidigare
du har haft hemkommun i Finland i högst tre år.
I den inledande kartläggningen får du information om utbildning i finska eller svenska, arbetssökning, utbildning och tjänster i Vanda.
Vid den inledande kartläggningen talas man vid med hjälp av tolk.
Den inledande kartläggningen är avgiftsfri.
Begäran om inledande kartläggning
Du kan begära en inledande kartläggning via e-post eller så kan du boka en tid per telefon.
Tfn 09 839 32622, 09 839 27525 eller 09 839 31766
Om du söker arbete, bör du anmäla dig till TE-byrån.
TE-byrån gör den inledande kartläggningen.
Läs mer om den inledande kartläggningen och integrationsplanen på InfoFinlands webbplats Integration i Finland
linkkiVanda stad:
Inledande kartläggningfinska _ engelska
Behöver du en tolk?
Om du måste sköta ärenden med myndigheter, men inte kan finska eller svenska och det inte heller finns något annat språk som både du och myndigheten talar, kan du använda en tolktjänst.
Meddela alltid myndigheten i förväg om du behöver en tolk.
Myndigheten bokar tolken och då får du tolkningstjänsten gratis.
Om du själv bokar tolken och betalar kostnaderna, kan du anlita en tolk när som helst.
Läs mer: Behöver du en tolk?
linkkiVanda stad:
Information om tolktjänsterfinska
linkkiFinlands översättar- och tolkförbund:
Sök tolk eller översättarefinska _ svenska _ engelska
Rådgivning för och integration av invandrare
Inledande kartläggning
Behöver du en tolk?
Rådgivning för och integration av invandrare
Invandrartjänster
Vanda stads tjänster för invandrare omfattar
mottagningstjänster för invandrare
integrationstjänster
Vanda stads tjänster för invandrare (Vantaan maahanmuuttajapalvelut) ger dig information om integration, social- och hälsovårdstjänster och om stadens och olika organisationers tjänster.
Du kan bli klient om du flyttat till Finland på grund av familjeband, är flykting, offer för människohandel eller har rätt till en inledande kartläggning.
Tfn (09) 839 21074 och (09) 839 32042
linkkiVanda stad:
Invandrartjänsterfinska _ engelska
Vandainfo ger dig information om såväl Vandas stads som statens tjänster.
Vandainfon finns i Dickursby, Korso och Myrbacka.
Adresserna är:
Dixi, Banvägen 11, 2:a vån.
tfn (09) 839 22133
Tfn (09) 839 22133
Tfn (09) 839 22133
Kontaktuppgifterna och öppettiderna hittar du på Vanda stads webbplats.
linkkiVanda stad:
Vandainfofinska _ svenska _ engelska
Den internationella föreningen i Håkansböle (Hakunilan kansainvälinen yhdistys) har en rådgivningspunkt som betjänar invandrare i Håkansböle, Björkby och andra områden i Vanda, som vill ha information om till exempel studier, språkkurser, arbete, hobbyverksamhet, krissituationer eller juridiska frågor.
Sporrgränden 2 A, vån. 3 (Håkansböle)
Tfn (09) 272 2775 och 040 501 3199.
linkkiInternationella föreningen i Håkansböle:
Rådgivning för invandrarefinska _ engelska _ ryska _ somaliska _ arabiska
På invandrarrådgivningen vid föreningen Vantaan Järjestörinki ry (Vantaan Järjestörinki ry:n Maahanmuuttajien neuvontapiste) kan du fråga om sådant som rör till exempel arbetslivet, social trygghet, hälsa, utbildning och uppehållstillstånd.
Adress:
Ranunkelvägen 22
Asukastila Myyrinki
Eldstadstorget 1 eller Kopparbergsvägen 10 B, vån.
Vanda Tfn (09) 839 35703 och 040 183 0930
Rautbergsgatan 3
Tfn 045 134 1711
Rådgivning för invandrarefinska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
IHH – serviceställe för dig som flyttar till Finland engelska
Inledande kartläggning
Den inledande kartläggningen (alkukartoitus) hjälper dig att hitta lämpliga tjänster i din hemstad.
Vanda stad eller Nylands TE-byrå ordnar en inledande kartläggning för varje ny invandrare i Vanda.
Du har rätt att få en inledande kartläggning om
din hemkommun är Vanda
du har flyttat till Vanda från ett annat land eller en annan ort i Finland
någon inledande kartläggning inte har gjorts för dig tidigare
du har haft hemkommun i Finland i högst tre år.
I den inledande kartläggningen får du information om utbildning i finska eller svenska, arbetssökning, utbildning och tjänster i Vanda.
Vid den inledande kartläggningen talas man vid med hjälp av tolk.
Den inledande kartläggningen är avgiftsfri.
Begäran om inledande kartläggning
Du kan begära en inledande kartläggning via e-post eller så kan du boka en tid per telefon.
Tfn 09 839 32622, 09 839 27525 eller 09 839 31766
Om du söker arbete, bör du anmäla dig till TE-byrån.
TE-byrån gör den inledande kartläggningen.
Läs mer om den inledande kartläggningen och integrationsplanen på InfoFinlands webbplats Integration i Finland
linkkiVanda stad:
Inledande kartläggningfinska _ engelska
Behöver du en tolk?
Om du måste sköta ärenden med myndigheter, men inte kan finska eller svenska och det inte heller finns något annat språk som både du och myndigheten talar, kan du använda en tolktjänst.
Meddela alltid myndigheten i förväg om du behöver en tolk.
Myndigheten bokar tolken och då får du tolkningstjänsten gratis.
Om du själv bokar tolken och betalar kostnaderna, kan du anlita en tolk när som helst.
Läs mer: Behöver du en tolk?
linkkiVanda stad:
Information om tolktjänsterfinska
linkkiFinlands översättar- och tolkförbund:
Sök tolk eller översättarefinska _ svenska _ engelska
Tillståndsärenden
På Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU-medborgarens uppehållsrätt.
Migrationsverkets tjänsteställe i Helsingfors :
Göksgränd 3A
Du kan också ansöka om många slags uppehållstillstånd och EU-registrering på internet i tjänsten Enter Finland.
Om du inte är van vid att använda en dator, fyll i en ansökan på papper och lämna in den på Migrationsverkets tjänsteställe.
Dät är alltid bra att boka en tid i förväg på tjänstestället.
Du kan boka en tid på Migrationsverkets tidsbokningstjänst.
Observera att tjänstestället inte kan ge rådgivning om tillståndsärenden.
Läs mer: Flytta till Finland.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Registrering som invånare
Om du flyttar ditt stadigvarande boende till Vanda, ska du registrera dig som invånare i kommunen.
Du kan registrera dig vid magistraten.
Albertsgatan 25
Växel 029 55 39391
Registrering av utlänningar 029 55 36 300
När du går till magistraten ska du ta med dig
legitimation (till exempel pass)
uppehållstillstånd och uppehållskort (om du behöver uppehållstillstånd i Finland)
registreringsintyget över uppehållsrätten (oleskeluoikeuden rekisteröintitodistus) om du är EU-medborgare.
äktenskapsintyg
dina barns födelseattester.
Observera att utländska handlingar ska vara legaliserade.
Du får mer information om att legalisera officiella handlingar vid magistraten eller beskickningen för ditt eget land i Finland.
Läs mer: Registrering som invånare.
Registrering av utlänningarfinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
Du kan få:
kostnadsfri rådgivning och information kring att flytta på flera olika språk
en finländsk personbeteckning, registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1-intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
Adress
Albertsgatan 25
IHH – serviceställe för dig som flyttar till Finland engelska
Webbappen IHH Service Advisor App engelska
Tillståndsärenden
På Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU-medborgarens uppehållsrätt.
Migrationsverkets tjänsteställe i Helsingfors :
Göksgränd 3A
Du kan också ansöka om många slags uppehållstillstånd och EU-registrering på internet i tjänsten Enter Finland.
Om du inte är van vid att använda en dator, fyll i en ansökan på papper och lämna in den på Migrationsverkets tjänsteställe.
Dät är alltid bra att boka en tid i förväg på tjänstestället.
Du kan boka en tid på Migrationsverkets tidsbokningstjänst.
Observera att tjänstestället inte kan ge rådgivning om tillståndsärenden.
Läs mer: Flytta till Finland.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Registrering som invånare
Om du flyttar ditt stadigvarande boende till Vanda, ska du registrera dig som invånare i kommunen.
Du kan registrera dig vid magistraten.
Albertsgatan 25
Växel 029 55 39391
Registrering av utlänningar 029 55 36 300
När du går till magistraten ska du ta med dig
legitimation (till exempel pass)
uppehållstillstånd och uppehållskort (om du behöver uppehållstillstånd i Finland)
registreringsintyget över uppehållsrätten (oleskeluoikeuden rekisteröintitodistus) om du är EU-medborgare.
äktenskapsintyg
dina barns födelseattester.
Observera att utländska handlingar ska vara legaliserade.
Du får mer information om att legalisera officiella handlingar vid magistraten eller beskickningen för ditt eget land i Finland.
Läs mer: Registrering som invånare.
Registrering av utlänningarfinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
Du kan få:
kostnadsfri rådgivning och information kring att flytta på flera olika språk
en finländsk personbeteckning, registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1-intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
Adress
IHH – serviceställe för dig som flyttar till Finland engelska
Webbappen IHH Service Advisor App engelska
Tillståndsärenden
På Migrationsverkets tjänsteställe i Helsingfors kan du ansöka om uppehållstillstånd och registrera EU-medborgarens uppehållsrätt.
Migrationsverkets tjänsteställe i Helsingfors :
Göksgränd 3A
Du kan också ansöka om många slags uppehållstillstånd och EU-registrering på internet i tjänsten Enter Finland.
Om du inte är van vid att använda en dator, fyll i en ansökan på papper och lämna in den på Migrationsverkets tjänsteställe.
Dät är alltid bra att boka en tid i förväg på tjänstestället.
Du kan boka en tid på Migrationsverkets tidsbokningstjänst.
Observera att tjänstestället inte kan ge rådgivning om tillståndsärenden.
Läs mer: Flytta till Finland.
linkkiEnterfinland.fi:
Elektronisk ansökanfinska _ svenska _ engelska
Elektronisk tidsbokningfinska _ svenska _ engelska
Registrering som invånare
Om du flyttar ditt stadigvarande boende till Vanda, ska du registrera dig som invånare i kommunen.
Du kan registrera dig vid magistraten.
Albertsgatan 25
Växel 029 55 39391
Registrering av utlänningar 029 55 36 300
När du går till magistraten ska du ta med dig
legitimation (till exempel pass)
uppehållstillstånd och uppehållskort (om du behöver uppehållstillstånd i Finland)
registreringsintyget över uppehållsrätten (oleskeluoikeuden rekisteröintitodistus) om du är EU-medborgare.
äktenskapsintyg
dina barns födelseattester.
Observera att utländska handlingar ska vara legaliserade.
Du får mer information om att legalisera officiella handlingar vid magistraten eller beskickningen för ditt eget land i Finland.
Läs mer: Registrering som invånare.
Registrering av utlänningarfinska _ svenska _ engelska
Om du har flyttat till huvudstadsregionen nyligen, kan du vid International House Helsinki (IHH) få rådgivning och myndighetstjänster på ett och samma besök.
Du kan få:
kostnadsfri rådgivning och information kring att flytta på flera olika språk
en finländsk personbeteckning, registrera dig som invånare och anmäla din adress
skattekort och skattenummer samt rådgivning om beskattningen
information om den sociala tryggheten och sociala förmåner
rådgivning om arbets- och näringslivstjänsterna och om att komma igång med jobbsökningen
rådgivning om arbetspension och om A1-intyget
rådgivning om anställningar
rådgivning för företag och arbetsgivare.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
Adress
IHH – serviceställe för dig som flyttar till Finland engelska
Webbappen IHH Service Advisor App engelska
Trafik
Beslutsfattande och påverkan
Religion
Grundläggande information
Historia
Trafik
Kollektivtrafiken
Esbo och hela huvudstadsregionen har goda kollektivtrafikförbindelser.
I Esbo finns flera tåg- och metrostationer.
I staden finns flera busslinjer.
Information och råd till resenärerfinska _ svenska _ engelska
Esbo tillhör samkommunen Helsingforsregionens trafik HRT (HSL), som ordnar kollektivtrafiken i huvudstadsregionen.
Du kan söka information om rutterna i reseplanerartjänsten (Reittiopas).
Tjänsten ger dig råd om olika kollektivtrafikförbindelser från ett ställe till ett annat.
Reseplanerarefinska _ svenska _ engelska _ ryska
I kollektivtrafiken kan du betala med kontanter eller resekort.
I närtågen måste du köpa biljetten i förväg.
Mer information om resekorten och deras försäljningsställen i Esbo hittar du på HRT:s webbplats.
Du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat.
Biljetter och priserfinska _ svenska _ engelska
Att gå och cykla
Om du vill gå eller cykla i Esbo kan du söka en lämplig rutt i reseplaneraren för cykling och gång.
Resplan för cycling och gångfinska _ svenska _ engelska _ ryska
Cykelkartor för Helsingfors, Vanda och Esbo delas ut vid samservicekontoren och idrottsverkens serviceställen.
Cykelkartorna är kostnadsfria.
Friluftskartafinska
Bil och flyg
Du kan parkera bilen på många järnvägsstationer och fortsätta färden med kollektivtrafiken.
Helsingfors-Vanda flygplats ligger Esbos grannkommun Vanda.
Läs mer: Trafik.
linkkiEsbo stad:
Trafikfinska _ svenska _ engelska
linkkiEsbo stad:
Kartorfinska _ svenska _ engelska
Beslutsfattande och påverkan
I Esbo beslutas ärenden av stadsfullmäktige.
I stadsfullmäktige sitter 75 ledamöter som representerar olika politiska grupper.
Fullmäktige väljs var fjärde år genom kommunalval.
Invånarna i Esbo kan påverka beslutsfattandet och beredning av ärenden på många olika sätt.
Du kan ge respons till beslutsfattarna och tjänstemännen till exempel via det elektroniska responssystemet.
Du kan vara med i invånarverksamheten eller ta ett invånarinitiativ.
Läs mer om hur du kan påverka på Esbo stads webbplats.
I Esbo finns en delegation för mångkulturella frågor som utvecklar stadens mångkulturella politik.
I Esbo finns många politiska föreningar, invandrarföreningar och andra föreningar via vilka du också kan påverka beslutsfattandet.
Läs mer: Beslutsfattande och påverkan
linkkiEsbo stad:
Information om beslutsfattandefinska _ svenska _ engelska
linkkiEsbo stad:
Information om påverkanfinska _ svenska _ engelska
linkkiEsbo stad:
Elektroniskt responssystemfinska _ svenska _ engelska
linkkiEsbo stad:
Mångkulturella ärendenfinska _ svenska _ engelska
Religion
Många religiösa samfund är verksamma i Esbo och Helsingfors.
Via tjänsten Uskonnot Suomessa kan du söka information efter det religiösa samfundet och orten.
Läs mer: Kulturer och religioner i Finland.
Religiösa samfundfinska _ engelska
linkkiEsbo kyrkliga samfällighet:
Evangelisk-lutherska församlingarfinska _ svenska _ engelska
linkkiHelsingfors ortodoxa församling:
Ortodoxa församlingenfinska _ ryska
Grundläggande information
Esbo är en av huvudstadsregionens fyra kommuner.
Det ligger bredvid Helsingfors, väster om staden.
Utöver dessa finns det flera mindre tätorter, landsbygd och skogar i Esbo.
Esbo har cirka 280 000 invånare.
De flesta invånarna är finskspråkiga.
Ungefär 7 procent av invånarna är svenskspråkiga och 16 procent har andra modersmål.
Esbos areal är cirka 528 km2, varav cirka 216 km2 är vatten.
linkkiEsbo stad:
Information om Esbofinska _ svenska _ engelska
Historia
Esboområdet var bebott redan för ungefär 8 000 år sedan.
Då var södra Esbo fortfarande hav.
På 1200-talet flyttade många emigranter från Sverige till Esbo.
På 1400-talet blev Esbo en självständig socken med många byar.
I Esbo byggdes stora herrgårdar som hade stor betydelse för områdets utveckling.
När Finland blev en del av Ryssland blev Helsingfors huvudstad år 1812.
Även om Helsingfors växte snabbt, var Esbo ännu länge en fridfull landssocken.
Inflyttningen till Esbo blev livligare från och med 1940-talet.
År 1950 hade Esbo 25 000 invånare och 15 år senare redan 65 000 invånare.
Esbo blev en stad år 1972.
linkkiEsbo stad:
Historiafinska _ svenska
linkkiEsbo stad:
Museerfinska _ svenska _ engelska
Trafik
Beslutsfattande och påverkan
Religion
Grundläggande information
Historia
Trafik
Kollektivtrafiken
Esbo och hela huvudstadsregionen har goda kollektivtrafikförbindelser.
I Esbo finns flera tåg- och metrostationer.
I staden finns flera busslinjer.
Information och råd till resenärerfinska _ svenska _ engelska
Esbo tillhör samkommunen Helsingforsregionens trafik HRT (HSL), som ordnar kollektivtrafiken i huvudstadsregionen.
Du kan söka information om rutterna i reseplanerartjänsten (Reittiopas).
Tjänsten ger dig råd om olika kollektivtrafikförbindelser från ett ställe till ett annat.
Reseplanerarefinska _ svenska _ engelska _ ryska
I kollektivtrafiken kan du betala med kontanter eller resekort.
I närtågen måste du köpa biljetten i förväg.
Mer information om resekorten och deras försäljningsställen i Esbo hittar du på HRT:s webbplats.
Du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat.
Biljetter och priserfinska _ svenska _ engelska
Att gå och cykla
Om du vill gå eller cykla i Esbo kan du söka en lämplig rutt i reseplaneraren för cykling och gång.
Resplan för cycling och gångfinska _ svenska _ engelska _ ryska
Cykelkartor för Helsingfors, Vanda och Esbo delas ut vid samservicekontoren och idrottsverkens serviceställen.
Cykelkartorna är kostnadsfria.
Friluftskartafinska
Bil och flyg
Du kan parkera bilen på många järnvägsstationer och fortsätta färden med kollektivtrafiken.
Helsingfors-Vanda flygplats ligger Esbos grannkommun Vanda.
Läs mer: Trafik.
linkkiEsbo stad:
Trafikfinska _ svenska _ engelska
linkkiEsbo stad:
Kartorfinska _ svenska _ engelska
Beslutsfattande och påverkan
I Esbo beslutas ärenden av stadsfullmäktige.
I stadsfullmäktige sitter 75 ledamöter som representerar olika politiska grupper.
Fullmäktige väljs var fjärde år genom kommunalval.
Invånarna i Esbo kan påverka beslutsfattandet och beredning av ärenden på många olika sätt.
Du kan ge respons till beslutsfattarna och tjänstemännen till exempel via det elektroniska responssystemet.
Du kan vara med i invånarverksamheten eller ta ett invånarinitiativ.
Läs mer om hur du kan påverka på Esbo stads webbplats.
I Esbo finns en delegation för mångkulturella frågor som utvecklar stadens mångkulturella politik.
I Esbo finns många politiska föreningar, invandrarföreningar och andra föreningar via vilka du också kan påverka beslutsfattandet.
Läs mer: Beslutsfattande och påverkan
linkkiEsbo stad:
Information om beslutsfattandefinska _ svenska _ engelska
linkkiEsbo stad:
Information om påverkanfinska _ svenska _ engelska
linkkiEsbo stad:
Elektroniskt responssystemfinska _ svenska _ engelska
linkkiEsbo stad:
Mångkulturella ärendenfinska _ svenska _ engelska
Religion
Många religiösa samfund är verksamma i Esbo och Helsingfors.
Via tjänsten Uskonnot Suomessa kan du söka information efter det religiösa samfundet och orten.
Läs mer: Kulturer och religioner i Finland.
Religiösa samfundfinska _ engelska
linkkiEsbo kyrkliga samfällighet:
Evangelisk-lutherska församlingarfinska _ svenska _ engelska
linkkiHelsingfors ortodoxa församling:
Ortodoxa församlingenfinska _ ryska
Grundläggande information
Esbo är en av huvudstadsregionens fyra kommuner.
Det ligger bredvid Helsingfors, väster om staden.
Utöver dessa finns det flera mindre tätorter, landsbygd och skogar i Esbo.
Esbo har cirka 280 000 invånare.
De flesta invånarna är finskspråkiga.
Ungefär 7 procent av invånarna är svenskspråkiga och 16 procent har andra modersmål.
Esbos areal är cirka 528 km2, varav cirka 216 km2 är vatten.
linkkiEsbo stad:
Information om Esbofinska _ svenska _ engelska
Historia
Esboområdet var bebott redan för ungefär 8 000 år sedan.
Då var södra Esbo fortfarande hav.
På 1200-talet flyttade många emigranter från Sverige till Esbo.
På 1400-talet blev Esbo en självständig socken med många byar.
I Esbo byggdes stora herrgårdar som hade stor betydelse för områdets utveckling.
När Finland blev en del av Ryssland blev Helsingfors huvudstad år 1812.
Även om Helsingfors växte snabbt, var Esbo ännu länge en fridfull landssocken.
Inflyttningen till Esbo blev livligare från och med 1940-talet.
År 1950 hade Esbo 25 000 invånare och 15 år senare redan 65 000 invånare.
Esbo blev en stad år 1972.
linkkiEsbo stad:
Historiafinska _ svenska
linkkiEsbo stad:
Museerfinska _ svenska _ engelska
Trafik
Beslutsfattande och påverkan
Religion
Grundläggande information
Historia
Trafik
Kollektivtrafiken
Esbo och hela huvudstadsregionen har goda kollektivtrafikförbindelser.
I Esbo finns flera tåg- och metrostationer.
I staden finns flera busslinjer.
Information och råd till resenärerfinska _ svenska _ engelska
Esbo tillhör samkommunen Helsingforsregionens trafik HRT (HSL), som ordnar kollektivtrafiken i huvudstadsregionen.
Du kan söka information om rutterna i reseplanerartjänsten (Reittiopas).
Tjänsten ger dig råd om olika kollektivtrafikförbindelser från ett ställe till ett annat.
Reseplanerarefinska _ svenska _ engelska
I kollektivtrafiken kan du betala med kontanter eller resekort.
I närtågen måste du köpa biljetten i förväg.
Mer information om resekorten och deras försäljningsställen i Esbo hittar du på HRT:s webbplats.
Du kan även köpa en mobilbiljett med telefonen eller en enkelbiljett i en automat.
Biljetter och priserfinska _ svenska _ engelska
Att gå och cykla
Om du vill gå eller cykla i Esbo kan du söka en lämplig rutt i reseplaneraren för cykling och gång.
Resplan för cycling och gångfinska _ svenska _ engelska _ ryska
Bil och flyg
Du kan parkera bilen på många järnvägsstationer och fortsätta färden med kollektivtrafiken.
Helsingfors-Vanda flygplats ligger Esbos grannkommun Vanda.
Läs mer: Trafik.
linkkiEsbo stad:
Trafikfinska _ svenska _ engelska
linkkiEsbo stad:
Kartorfinska _ svenska _ engelska
Beslutsfattande och påverkan
I Esbo beslutas ärenden av stadsfullmäktige.
I stadsfullmäktige sitter 75 ledamöter som representerar olika politiska grupper.
Fullmäktige väljs var fjärde år genom kommunalval.
Invånarna i Esbo kan påverka beslutsfattandet och beredning av ärenden på många olika sätt.
Du kan ge respons till beslutsfattarna och tjänstemännen till exempel via det elektroniska responssystemet.
Du kan vara med i invånarverksamheten eller ta ett invånarinitiativ.
Läs mer om hur du kan påverka på Esbo stads webbplats.
I Esbo finns en delegation för mångkulturella frågor som utvecklar stadens mångkulturella politik.
I Esbo finns många politiska föreningar, invandrarföreningar och andra föreningar via vilka du också kan påverka beslutsfattandet.
Läs mer: Beslutsfattande och påverkan
linkkiEsbo stad:
Information om beslutsfattandefinska _ svenska _ engelska
linkkiEsbo stad:
Information om påverkanfinska _ svenska _ engelska
linkkiEsbo stad:
Elektroniskt responssystemfinska _ svenska _ engelska
linkkiEsbo stad:
Mångkulturella ärendenfinska _ svenska _ engelska
Religion
Många religiösa samfund är verksamma i Esbo och Helsingfors.
Via tjänsten Uskonnot Suomessa kan du söka information efter det religiösa samfundet och orten.
Läs mer: Kulturer och religioner i Finland.
Religiösa samfundfinska _ engelska
linkkiEsbo kyrkliga samfällighet:
Evangelisk-lutherska församlingarfinska _ svenska _ engelska
linkkiHelsingfors ortodoxa församling:
Ortodoxa församlingenfinska _ ryska
Grundläggande information
Esbo är en av huvudstadsregionens fyra kommuner.
Det ligger bredvid Helsingfors, väster om staden.
Utöver dessa finns det flera mindre tätorter, landsbygd och skogar i Esbo.
Esbo har cirka 280 000 invånare.
De flesta invånarna är finskspråkiga.
Ungefär 7 procent av invånarna är svenskspråkiga och 16 procent har andra modersmål.
Esbos areal är cirka 528 km2, varav cirka 216 km2 är vatten.
linkkiEsbo stad:
Information om Esbofinska _ svenska _ engelska
Historia
Esboområdet var bebott redan för ungefär 8 000 år sedan.
Då var södra Esbo fortfarande hav.
På 1200-talet flyttade många emigranter från Sverige till Esbo.
På 1400-talet blev Esbo en självständig socken med många byar.
I Esbo byggdes stora herrgårdar som hade stor betydelse för områdets utveckling.
När Finland blev en del av Ryssland blev Helsingfors huvudstad år 1812.
Även om Helsingfors växte snabbt, var Esbo ännu länge en fridfull landssocken.
Inflyttningen till Esbo blev livligare från och med 1940-talet.
År 1950 hade Esbo 25 000 invånare och 15 år senare redan 65 000 invånare.
Esbo blev en stad år 1972.
linkkiEsbo stad:
Historiafinska _ svenska
linkkiEsbo stad:
Museerfinska _ svenska _ engelska
Evenemang
Bibliotek
Motion
Att röra sig i naturen
Teater och film
Museer
Fritidsverksamhet för barn och unga
Föreningar
I Esbo finns många hobbymöjligheter.
Invånarhusen Kivenkolo och Kylämaja är öppna för alla.
I invånarhusen kan områdets invånare vistas och samlas samt få anvisningar och råd.
Invånarhuset Kivenkolo
Sjöstöveln 1 A
linkkiEsbo stad:
Kivenkolo invånarhusfinska _ svenska _ engelska
Invånarhuset Kylämaja
Mattsgatan 7
linkkiEsbo stad:
Invånarhus Kylämajafinska
Vid Esbo arbetarinstitut (Espoon työväenopisto) kan man till exempel skapa konst, handarbeten, laga mat, dansa eller idka motion.
Där kan man även studera finska och andra språk.
linkkiEsbo stad:
Arbetarinstitutetfinska _ svenska _ engelska
I Esbo finns flera läroanstalter som ger grundundervisning i konstämnen speciellt för barn och unga.
Olika konstarter är musik, bildkonst, dans, teater och cirkus.
linkkiEsbo stad:
Konstundervisningfinska _ engelska.
Konsthuset Lilla Aurora ordnar kulturevenemang för barn.
linkkiEsbo stad:
Kulturevenemang för barnfinska _ svenska _ engelska
Läs mer: Fritid.
Evenemang
Evenemangfinska _ svenska _ engelska _ ryska _ kinesiska
linkkiEsbo stad:
Evenemangfinska
Bibliotek
I Esbo finns flera bibliotek på olika håll i staden.
På biblioteket kan du låna böcker, tidningar, musik, filmer, spel och mycket annat.
Biblioteken har böcker och annat material på flera olika språk.
I biblioteket kan du också använda dator.
Ofta hålls också utställningar och evenemang på biblioteken.
linkkiEsbo stad:
Bibliotekfinska _ svenska _ engelska
Flerspråkiga biblioteket
Flerspråkiga biblioteket ligger i Böle i Helsingfors
Här finns böcker, musik, tidningar och tidskrifter samt ljudböcker på flera olika språk.
Du kan åka till Böle eller beställa material till ditt eget närbibliotek.
linkkiHelsingfors stadsbibliotek:
Flerspråkiga biblioteketfinska _ svenska _ engelska
Huvudstadsregionens gemensamma bibliotekstjänstfinska _ svenska _ engelska _ somaliska _ persiska _ arabiska
Läs mer: Bibliotek.
Motion
I Esbo finns simhallar, flera idrottshallar, idrottsplaner och andra idrottsplatser för olika idrottsgrenar.
På motionsslingorna kan man springa på somrarna och åka skidor på vintrarna.
Läs mer: Motion.
linkkiEsbo stad:
Information om motionstjänsternafinska _ svenska _ engelska
linkkiEsbo stad:
Idrottsklubbarfinska _ svenska
Att röra sig i naturen
I Esbo finns flera friluftsområden där man kan vandra i naturen.
Till exempel Noux nationalpark ligger delvis på Esbos område.
linkkiEsbo stad:
Naturobjekt i Esbofinska _ svenska _ engelska
Webbsidorfinska _ svenska _ engelska _ ryska _ kinesiska
Hemstadsstigarfinska _ svenska _ engelska
I naturhuset Villa Elfvik ordnas utflykter, evenemang och utställningar.
Naturhuset är öppet för alla och ligger vid sidan av Bredvikens naturskyddsområde.
linkkiVilla Elfvik:
Naturens husfinska _ svenska _ engelska
I Esbo finns motionsslingor och friluftsleder på olika håll i staden.
På vintern är många motionsslingor skidspår.
En del rutter är belysta.
linkkiEsbo stad:
Friluftslivfinska _ svenska _ engelska
linkkiEsbo stad:
Friluftsområdenfinska _ svenska _ engelska
Vid insjöarna och på havskusten finns många badstränder.
Alla Esbobor får fritt fiska med metspö och pimpla.
Om du använder andra fiskeredskap ska du ha ett fisketillstånd.
linkkiEsbo stad:
Fiske och jaktfinska _ svenska _ engelska
Läs mer: Att röra sig i naturen.
Teater och film
I Esbo finns flera yrkes- och amatörteatrar.
I Esbo finns tre biografer.
Mer information om filmerna hittar du på biografernas webbplatser.
Därtill ordnar Esbo stad filmvisningar.
Läs mer: Teater och film.
linkkiFinnkino:
Filmerfinska _ engelska
Filmerfinska
Filmerfinska _ svenska _ engelska
linkkiEsbo stad:
Teatrar i Esbofinska _ svenska _ engelska
Museer
I Esbo finns flera museer.
Esbo moderna konstmuseum EMMA är ett av Finlands största konstmuseer.
Läs mer: Museer.
linkkiEsbo stad:
Museerfinska _ svenska _ engelska
linkkiEsbo stad:
Stadsmuseetfinska _ svenska _ engelska
linkkiEsbo stad:
Museet för modern konst EMMAfinska _ svenska _ engelska _ ryska
Fritidsverksamhet för barn och unga
I Esbo finns flera läroanstalter som ger grundundervisning i konstämnen speciellt för barn och unga.
Olika konstarter är musik, bildkonst, dans, teater och cirkuskonst.
I Esbo finns ungdomsgårdar med utbildade ledare som övervakar verksamheten.
Ungdomsgårdarna är öppna för alla ungdomar i åldrarna 9–17.
På ungdomsgårdarna kan de unga vistas på fritiden.
Där bedrivs det även hobbyklubbar och ordnas kurser och evenemang.
Också föreningar och idrottsklubbar ordnar mycket verksamhet för ungdomar.
Läs mer: Fritidsverksamhet för barn och unga.
linkkiEsbo stad:
Verksamhet för ungafinska _ svenska _ engelska
linkkiEsbo stad:
Ungdomsgårdarfinska _ svenska _ engelska
linkkiEsbo stad:
Rådgivning för ungafinska _ svenska _ engelska
linkkiEsbo stad:
Idrottsklubbarfinska _ svenska
Hobbysökningfinska
Föreningar
I Esbo finns många olika föreningar, till exempel kulturföreningar och idrottsklubbar.
Läs mer: Föreningar.
linkkiEsbo stad:
Idrottsklubbarfinska _ svenska
Föreningsverksamhetfinska
linkkiEsbo stad:
Föreningar för seniorerfinska _ svenska
Evenemang
Bibliotek
Motion
Att röra sig i naturen
Teater och film
Museer
Fritidsverksamhet för barn och unga
Föreningar
I Esbo finns många hobbymöjligheter.
Invånarhusen Kivenkolo och Kylämaja är öppna för alla.
I invånarhusen kan områdets invånare vistas och samlas samt få anvisningar och råd.
Invånarhuset Kivenkolo
Sjöstöveln 1 A
linkkiEsbo stad:
Kivenkolo invånarhusfinska _ svenska _ engelska
Invånarhuset Kylämaja
Mattsgatan 7
linkkiEsbo stad:
Invånarhus Kylämajafinska
Vid Esbo arbetarinstitut (Espoon työväenopisto) kan man till exempel skapa konst, handarbeten, laga mat, dansa eller idka motion.
Där kan man även studera finska och andra språk.
linkkiEsbo stad:
Arbetarinstitutetfinska _ svenska _ engelska
I Esbo finns flera läroanstalter som ger grundundervisning i konstämnen speciellt för barn och unga.
Olika konstarter är musik, bildkonst, dans, teater och cirkus.
linkkiEsbo stad:
Konstundervisningfinska _ engelska.
Konsthuset Lilla Aurora ordnar kulturevenemang för barn.
linkkiEsbo stad:
Kulturevenemang för barnfinska _ svenska _ engelska
Läs mer: Fritid.
Evenemang
Evenemangfinska _ svenska _ engelska _ ryska
linkkiEsbo stad:
Evenemangfinska
Bibliotek
I Esbo finns flera bibliotek på olika håll i staden.
På biblioteket kan du låna böcker, tidningar, musik, filmer, spel och mycket annat.
Biblioteken har böcker och annat material på flera olika språk.
I biblioteket kan du också använda dator.
Ofta hålls också utställningar och evenemang på biblioteken.
linkkiEsbo stad:
Bibliotekfinska _ svenska _ engelska
Flerspråkiga biblioteket
Flerspråkiga biblioteket ligger i Böle i Helsingfors
Här finns böcker, musik, tidningar och tidskrifter samt ljudböcker på flera olika språk.
Du kan åka till Böle eller beställa material till ditt eget närbibliotek.
linkkiHelsingfors stadsbibliotek:
Flerspråkiga biblioteketfinska _ svenska _ engelska
Huvudstadsregionens gemensamma bibliotekstjänstfinska _ svenska _ engelska _ somaliska _ persiska _ arabiska
Läs mer: Bibliotek.
Motion
I Esbo finns simhallar, flera idrottshallar, idrottsplaner och andra idrottsplatser för olika idrottsgrenar.
På motionsslingorna kan man springa på somrarna och åka skidor på vintrarna.
Läs mer: Motion.
linkkiEsbo stad:
Information om motionstjänsternafinska _ svenska _ engelska
linkkiEsbo stad:
Idrottsklubbarfinska _ svenska
Att röra sig i naturen
I Esbo finns flera friluftsområden där man kan vandra i naturen.
Till exempel Noux nationalpark ligger delvis på Esbos område.
linkkiEsbo stad:
Naturobjekt i Esbofinska _ svenska _ engelska
Webbsidorfinska _ svenska _ engelska _ ryska _ kinesiska
Hemstadsstigarfinska _ svenska _ engelska
I naturhuset Villa Elfvik ordnas utflykter, evenemang och utställningar.
Naturhuset är öppet för alla och ligger vid sidan av Bredvikens naturskyddsområde.
linkkiVilla Elfvik:
Naturens husfinska _ svenska _ engelska
I Esbo finns motionsslingor och friluftsleder på olika håll i staden.
På vintern är många motionsslingor skidspår.
En del rutter är belysta.
linkkiEsbo stad:
Friluftslivfinska _ svenska _ engelska
linkkiEsbo stad:
Friluftsområdenfinska _ svenska _ engelska
Vid insjöarna och på havskusten finns många badstränder.
Alla Esbobor får fritt fiska med metspö och pimpla.
Om du använder andra fiskeredskap ska du ha ett fisketillstånd.
linkkiEsbo stad:
Fiske och jaktfinska _ svenska _ engelska
Läs mer: Att röra sig i naturen.
Teater och film
I Esbo finns flera yrkes- och amatörteatrar.
I Esbo finns tre biografer.
Mer information om filmerna hittar du på biografernas webbplatser.
Därtill ordnar Esbo stad filmvisningar.
Läs mer: Teater och film.
linkkiFinnkino:
Filmerfinska _ engelska
Filmerfinska
Filmerfinska _ svenska _ engelska
linkkiEsbo stad:
Teatrar i Esbofinska _ svenska _ engelska
Museer
I Esbo finns flera museer.
Esbo moderna konstmuseum EMMA är ett av Finlands största konstmuseer.
Läs mer: Museer.
linkkiEsbo stad:
Museerfinska _ svenska _ engelska
linkkiEsbo stad:
Stadsmuseetfinska _ svenska _ engelska
linkkiEsbo stad:
Museet för modern konst EMMAfinska _ svenska _ engelska _ ryska
Fritidsverksamhet för barn och unga
I Esbo finns flera läroanstalter som ger grundundervisning i konstämnen speciellt för barn och unga.
Olika konstarter är musik, bildkonst, dans, teater och cirkuskonst.
I Esbo finns ungdomsgårdar med utbildade ledare som övervakar verksamheten.
Ungdomsgårdarna är öppna för alla ungdomar i åldrarna 9–17.
På ungdomsgårdarna kan de unga vistas på fritiden.
Där bedrivs det även hobbyklubbar och ordnas kurser och evenemang.
Också föreningar och idrottsklubbar ordnar mycket verksamhet för ungdomar.
Läs mer: Fritidsverksamhet för barn och unga.
linkkiEsbo stad:
Verksamhet för ungafinska _ svenska _ engelska
linkkiEsbo stad:
Ungdomsgårdarfinska _ svenska _ engelska
linkkiEsbo stad:
Rådgivning för ungafinska _ svenska _ engelska
linkkiEsbo stad:
Idrottsklubbarfinska _ svenska
Hobbysökningfinska
Föreningar
I Esbo finns många olika föreningar, till exempel kulturföreningar och idrottsklubbar.
Läs mer: Föreningar.
linkkiEsbo stad:
Idrottsklubbarfinska _ svenska
Föreningsverksamhetfinska
linkkiEsbo stad:
Föreningar för seniorerfinska _ svenska
Evenemang
Bibliotek
Motion
Att röra sig i naturen
Teater och film
Museer
Fritidsverksamhet för barn och unga
Föreningar
I Esbo finns många hobbymöjligheter.
Invånarhusen Kivenkolo och Kylämaja är öppna för alla.
I invånarhusen kan områdets invånare vistas och samlas samt få anvisningar och råd.
Invånarhuset Kivenkolo
Sjöstöveln 1 A
linkkiEsbo stad:
Kivenkolo invånarhusfinska _ svenska _ engelska
Invånarhuset Kylämaja
Mattsgatan 7
linkkiEsbo stad:
Invånarhus Kylämajafinska
Vid Esbo arbetarinstitut (Espoon työväenopisto) kan man till exempel skapa konst, handarbeten, laga mat, dansa eller idka motion.
Där kan man även studera finska och andra språk.
linkkiEsbo stad:
Arbetarinstitutetfinska _ svenska _ engelska
I Esbo finns flera läroanstalter som ger grundundervisning i konstämnen speciellt för barn och unga.
Olika konstarter är musik, bildkonst, dans, teater och cirkus.
linkkiEsbo stad:
Konstundervisningfinska _ engelska.
Konsthuset Lilla Aurora ordnar kulturevenemang för barn.
linkkiEsbo stad:
Kulturevenemang för barnfinska _ svenska _ engelska
Läs mer: Fritid.
Evenemang
Evenemangfinska _ svenska _ engelska _ ryska
linkkiEsbo stad:
Evenemangfinska
Bibliotek
I Esbo finns flera bibliotek på olika håll i staden.
På biblioteket kan du låna böcker, tidningar, musik, filmer, spel och mycket annat.
Biblioteken har böcker och annat material på flera olika språk.
I biblioteket kan du också använda dator.
Ofta hålls också utställningar och evenemang på biblioteken.
linkkiEsbo stad:
Bibliotekfinska _ svenska _ engelska
Flerspråkiga biblioteket
Flerspråkiga biblioteket ligger i Böle i Helsingfors
Här finns böcker, musik, tidningar och tidskrifter samt ljudböcker på flera olika språk.
Du kan åka till Böle eller beställa material till ditt eget närbibliotek.
linkkiHelsingfors stadsbibliotek:
Flerspråkiga biblioteketfinska _ svenska _ engelska
Huvudstadsregionens gemensamma bibliotekstjänstfinska _ svenska _ engelska _ somaliska _ persiska _ arabiska
Läs mer: Bibliotek.
Motion
I Esbo finns simhallar, flera idrottshallar, idrottsplaner och andra idrottsplatser för olika idrottsgrenar.
På motionsslingorna kan man springa på somrarna och åka skidor på vintrarna.
Läs mer: Motion.
linkkiEsbo stad:
Information om motionstjänsternafinska _ svenska _ engelska
linkkiEsbo stad:
Idrottsklubbarfinska _ svenska
Att röra sig i naturen
I Esbo finns flera friluftsområden där man kan vandra i naturen.
Till exempel Noux nationalpark ligger delvis på Esbos område.
linkkiEsbo stad:
Naturobjekt i Esbofinska _ svenska _ engelska
Webbsidorfinska _ svenska _ engelska _ ryska _ kinesiska
Hemstadsstigarfinska _ svenska _ engelska
I naturhuset Villa Elfvik ordnas utflykter, evenemang och utställningar.
Naturhuset är öppet för alla och ligger vid sidan av Bredvikens naturskyddsområde.
linkkiVilla Elfvik:
Naturens husfinska _ svenska _ engelska
I Esbo finns motionsslingor och friluftsleder på olika håll i staden.
På vintern är många motionsslingor skidspår.
En del rutter är belysta.
linkkiEsbo stad:
Friluftslivfinska _ svenska _ engelska
linkkiEsbo stad:
Friluftsområdenfinska _ svenska _ engelska
Vid insjöarna och på havskusten finns många badstränder.
Alla Esbobor får fritt fiska med metspö och pimpla.
Om du använder andra fiskeredskap ska du ha ett fisketillstånd.
linkkiEsbo stad:
Fiske och jaktfinska _ svenska _ engelska
Läs mer: Att röra sig i naturen.
Teater och film
I Esbo finns flera yrkes- och amatörteatrar.
I Esbo finns tre biografer.
Mer information om filmerna hittar du på biografernas webbplatser.
Därtill ordnar Esbo stad filmvisningar.
Läs mer: Teater och film.
linkkiFinnkino:
Filmerfinska _ engelska
Filmerfinska
Filmerfinska _ svenska _ engelska
linkkiEsbo stad:
Teatrar i Esbofinska _ svenska _ engelska
Museer
I Esbo finns flera museer.
Esbo moderna konstmuseum EMMA är ett av Finlands största konstmuseer.
Läs mer: Museer.
linkkiEsbo stad:
Museerfinska _ svenska _ engelska
linkkiEsbo stad:
Stadsmuseetfinska _ svenska _ engelska
linkkiEsbo stad:
Museet för modern konst EMMAfinska _ svenska _ engelska _ ryska
Fritidsverksamhet för barn och unga
I Esbo finns flera läroanstalter som ger grundundervisning i konstämnen speciellt för barn och unga.
Olika konstarter är musik, bildkonst, dans, teater och cirkuskonst.
I Esbo finns ungdomsgårdar med utbildade ledare som övervakar verksamheten.
Ungdomsgårdarna är öppna för alla ungdomar i åldrarna 9–17.
På ungdomsgårdarna kan de unga vistas på fritiden.
Där bedrivs det även hobbyklubbar och ordnas kurser och evenemang.
Också föreningar och idrottsklubbar ordnar mycket verksamhet för ungdomar.
Läs mer: Fritidsverksamhet för barn och unga.
linkkiEsbo stad:
Verksamhet för ungafinska _ svenska _ engelska
linkkiEsbo stad:
Ungdomsgårdarfinska _ svenska _ engelska
linkkiEsbo stad:
Rådgivning för ungafinska _ svenska _ engelska
linkkiEsbo stad:
Idrottsklubbarfinska _ svenska
Hobbysökningfinska
Föreningar
I Esbo finns många olika föreningar, till exempel kulturföreningar och idrottsklubbar.
Läs mer: Föreningar.
linkkiEsbo stad:
Idrottsklubbarfinska _ svenska
Föreningsverksamhetfinska
linkkiEsbo stad:
Föreningar för seniorerfinska _ svenska
Problem med uppehållstillståndet
Brott
Behöver du en jurist?
Våld Problem i äktenskap eller parförhållande
Barns och ungas problem
Missbruksproblem
Dödsfall
Ring nödnumret 112 om det är fråga om en nödsituation.
Via nödnumret kan du tillkalla polis, ambulans eller brandkår.
Ring inte nödnumret om det inte är en nödsituation.
Läs mer:Nödsituationer
linkkiEsbo stad:
Jourmottagningarfinska _ svenska _ engelska
Social- och krisjouren
Social- och krisjouren (sosiaali- ja kriisipäivystys) hjälper dygnet runt om du eller din familj behöver hjälp i en akut krissituation.
Krisen kan till exempel ha med våld, parförhållandet eller barnens problem att göra.
Du kan även kontakta social- och krisjouren om du har problem med din mentala hälsa, missbruksproblem eller om du råkat ut för en traumatisk händelse i livet.
Social- och krisjouren
Jorvs sjukhus
Åbovägen 150
Tfn (09) 816 42439
Öppet varje dag dygnet runt.
linkkiEsbo stad:
Social- och krisjourenfinska _ svenska _ engelska
Föreningen för mental hälsa i Finland (Suomen Mielenterveysseura) har en krismottagning för invandrare.
Kontoret ligger i Böle i Helsingfors.
Krismottagningen ger dig hjälp och stöd i svåra situationer.
Boka en tid per telefon på numret (09) 4135 0501.
linkkiFöreningen för mental hälsa i Finland:
Krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Problem med uppehållstillståndet
Om du har problem eller oklarheter med uppehållstillståndet, ska du ta kontakt med migrationsverket.
Läs mer: Problem med uppehållstillstånd
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Om du är flykting, asylsökande eller vistas i Finland av någon annan anledning kan du be om juridisk hjälp och rådgivning vid Flyktingrådgivningen rf.
Kontoret ligger i Helsingfors.
Adress: Kaisaniemigatan 4 A
Tfn 09 2313 9325
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Brott
Om du blir utsatt för ett brott, gör en brottsanmälan hos polisen.
Du kan göra brottsanmälan på internet.
Du kan även fylla i en blankett och lämna den till Esbo huvudpolisstation.
Esbo huvudpolisstation
Knektbrogränden 4
Läs mer: Brott
Kontaktuppgifterfinska _ svenska _ engelska
Elektronisk polisanmälanfinska _ svenska _ engelska
Behöver du en jurist?
Om du behöver juridisk hjälp, kan du kontakta Västra Nylands rättshjälpsbyrå.
Biskopsbron 9 B
Tfn 029 56 61820
Läs mer: Behöver du en jurist?
linkkiVästra Nylands rättshjälpsbyrå:
Rättshjälpfinska
Våld
Omatila (Omatila) hjälper dig om du har blivit utsatt för närståendevåld eller våld inom familjen.
Omatila ordnar vid behov boende för dig och dina barn.
Du kan ringa Omatila-tjänsten dygnet runt. Du behöver inte uppge ditt namn när du ringer.
Du kan också komma utan tidsbokning för att prata om din situation, måndag till fredag kl. 9–11 och onsdagar kl. 16–20.
Omatila
Enheten för familjeärenden
Kamrersvägen 6 A
Tfn 043 825 0535
Läs mer: Våld
linkkiEsbo stad:
Hjälp till offer för familjevåldfinska _ svenska _ engelska
Miehen Linja (Miehen Linja) är en tjänst som hjälper män, som har utsatt sina familjemedlemmar för våld. Tjänsten är avsedd för invandrarmän.
Målargränden 3 B
Tfn (09) 276 62899
Hjälp för invandrarmänfinska _ engelska
Problem i äktenskap eller parförhållande
Om du har problem i ditt äktenskap eller parförhållande kan du kontakta familjerådgivningen.
Familjerådgivningsbyråerna är i synnerhet avsedda för familjer med barn.
linkkiEsbo stad:
Familjerådgivningarfinska _ svenska _ engelska
Väestöliitto erbjuder rådgivning och terapi för par på finska och engelska.
linkkiBefolkningsförbundet:
Rådgivning till invandrare telefonledes och via e-postfinska _ svenska _ engelska
Familia Clubs projekt Duo erbjuder relationsrådgivning för par från två kulturer på finska och engelska.
Rådgivningen är avgiftsbelagd.
Relationsrådgivning för par från två kulturerfinska _ engelska
Också kyrkans familjerådgivningscentral erbjuder familjerådgivning vid problem i parförhållandet.
Kyrkans familjerådgivningfinska _ svenska _ engelska
Läs mer: Problem i äktenskap och parförhållande
Barns och ungas problem
Hälsovårdaren vid barnrådgivningen ger råd i frågor som rör hälsan och utvecklingen av barn under skolåldern.
I Esbo finns flera rådgivningsbyråer runtom i staden.
Rådgivningsbyråernas tidsbokning och rådgivning
Tfn (09) 816 22800
linkkiEsbo stad:
Rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
Vid problem som berör barn i skolåldern hjälper till exempel skolans hälsovårdare.
linkkiEsbo stad:
Information om hälsovården för skolbarnfinska _ svenska _ engelska
Om du behöver råd i frågor kring barns psykiska utveckling, kan du boka en tid hos familjerådgivningen.
linkkiEsbo stad:
Familjerådgivningarfinska _ svenska _ engelska
Väestöliitto ger råd till invandrarfamiljer i frågor rörande barnfostran och familjens välmående.
Rådgivningen på olika språk:
Tfn 050 325 7173 (ryska, engelska)
Unga kan prata om sina problem med hälsovårdaren på den egna skolan eller läroanstalten.
Det finns även andra ställen där man kan få hjälp.
En ung i åldern 13–22 år kan få hjälp vid Ungdomspolikliniken Nupoli om hen har problem till exempel med den mentala hälsan, rusmedelsbruk, spelande eller fritidsaktiviteterna.
Man kan ringa eller besöka Nupoli.
Besök på Nupoli är kostnadsfria och konfidentiella.
Tfn 09 816 31300
linkkiEsbo stad:
Nupoli - hjälp för ungafinska _ svenska
Om den unga inte är trygg i sitt eget hem, kan hen kontakta Finlands Röda Kors De ungas skyddshus.
Skyddshuset finns i Alberga.
De ungas skyddshus
Tfn (09) 8195 5360
linkkiFinlands Röda Kors:
De ungas skyddshusfinska
Läs mer: Barns och ungas problem
Om du har ekonomiska problem kan du fråga om råd hos kommunens socialarbetare.
Om du eller din familj inte har tillräckliga inkomster eller tillgångar för den nödvändiga dagliga försörjningen kan du söka grundläggande utkomststöd hos FPA.
Information om utkomststödfinska _ svenska _ engelska _ ryska _ estniska
Om du har problem med skulder, kontakta rättshjälpsbyråns ekonomi- och skuldrådgivning.
Tjänsten är kostnadsfri.
linkkiRättshjälpsbyrå:
Ekonomi- och skuldrådgivningfinska _ svenska _ engelska
Missbruksproblem
Kliniken för mental- och missbruksvård erbjuder vuxna Esbobor hjälp och vård vid problem med den mentala hälsan och missbruk.
Köpcentret Iso Omena
Telefon: 09 816 31300
linkkiEsbo stad:
Information om mentalvårdstjänsternafinska _ svenska _ engelska
Unga i åldern 13-22 med missbruksproblem kan få hjälp vid Ungdomspolikliniken Nupoli.
Tfn 09 816 31300
linkkiEsbo stad:
Nupoli - hjälp för ungafinska _ svenska
Läs mer: Missbruksproblem
Dödsfall
Begravningsbyråer hjälper med de praktiska arrangemangen vid en begravning.
Du kan söka begravningsbyråer till exempel på Finlands begravningsbyråers förbunds webbplats.
linkkiFinlands Begravningbyråers Förbund:
Begravningsbyråerfinska _ svenska _ engelska
I Esbo finns fem kristna begravningsplatser.
På Klockarmalmens begravningsplats finns ett gravområde för konfessionslösa.
Där kan de avlidna begravas som hade en annan religionstillhörighet eller inte hörde till något religionssamfund.
linkkiEsbo församlingar:
Begravningsplatserfinska _ svenska _ engelska
Om en närstående dör oväntat och du behöver stöd kan du kontakta social- och krisjouren i Esbo, telefon (09) 816 42439.
Läs mer: Dödsfall
Problem med uppehållstillståndet
Brott
Behöver du en jurist?
Våld Problem i äktenskap eller parförhållande
Barns och ungas problem
Missbruksproblem
Dödsfall
Ring nödnumret 112 om det är fråga om en nödsituation.
Via nödnumret kan du tillkalla polis, ambulans eller brandkår.
Ring inte nödnumret om det inte är en nödsituation.
Läs mer:Nödsituationer
linkkiEsbo stad:
Jourmottagningarfinska _ svenska _ engelska
Social- och krisjouren
Social- och krisjouren (sosiaali- ja kriisipäivystys) hjälper dygnet runt om du eller din familj behöver hjälp i en akut krissituation.
Krisen kan till exempel ha med våld, parförhållandet eller barnens problem att göra.
Du kan även kontakta social- och krisjouren om du har problem med din mentala hälsa, missbruksproblem eller om du råkat ut för en traumatisk händelse i livet.
Social- och krisjouren
Jorvs sjukhus
Åbovägen 150
Tfn (09) 816 42439
Öppet varje dag dygnet runt.
linkkiEsbo stad:
Social- och krisjourenfinska _ svenska _ engelska
Föreningen för mental hälsa i Finland (Suomen Mielenterveysseura) har en krismottagning för invandrare.
Kontoret ligger i Böle i Helsingfors.
Krismottagningen ger dig hjälp och stöd i svåra situationer.
Boka en tid per telefon på numret (09) 4135 0501.
linkkiFöreningen för mental hälsa i Finland:
Krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Problem med uppehållstillståndet
Om du har problem eller oklarheter med uppehållstillståndet, ska du ta kontakt med migrationsverket.
Läs mer: Problem med uppehållstillstånd
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Om du är flykting, asylsökande eller vistas i Finland av någon annan anledning kan du be om juridisk hjälp och rådgivning vid Flyktingrådgivningen rf.
Kontoret ligger i Helsingfors.
Adress: Kaisaniemigatan 4 A
Tfn 09 2313 9325
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Brott
Om du blir utsatt för ett brott, gör en brottsanmälan hos polisen.
Du kan göra brottsanmälan på internet.
Du kan även fylla i en blankett och lämna den till Esbo huvudpolisstation.
Esbo huvudpolisstation
Knektbrogränden 4
Läs mer: Brott
Kontaktuppgifterfinska _ svenska _ engelska
Elektronisk polisanmälanfinska _ svenska _ engelska
Behöver du en jurist?
Om du behöver juridisk hjälp, kan du kontakta Västra Nylands rättshjälpsbyrå.
Biskopsbron 9 B
Tfn 029 56 61820
Läs mer: Behöver du en jurist?
linkkiVästra Nylands rättshjälpsbyrå:
Rättshjälpfinska
Våld
Omatila (Omatila) hjälper dig om du har blivit utsatt för närståendevåld eller våld inom familjen.
Omatila ordnar vid behov boende för dig och dina barn.
Du kan ringa Omatila-tjänsten dygnet runt. Du behöver inte uppge ditt namn när du ringer.
Du kan också komma utan tidsbokning för att prata om din situation, måndag till fredag kl. 9–11 och onsdagar kl. 16–20.
Omatila
Enheten för familjeärenden
Kamrersvägen 6 A
Tfn 043 825 0535
Läs mer: Våld
linkkiEsbo stad:
Hjälp till offer för familjevåldfinska _ svenska _ engelska
Miehen Linja (Miehen Linja) är en tjänst som hjälper män, som har utsatt sina familjemedlemmar för våld. Tjänsten är avsedd för invandrarmän.
Målargränden 3 B
Tfn (09) 276 62899
Hjälp för invandrarmänfinska _ engelska
Problem i äktenskap eller parförhållande
Om du har problem i ditt äktenskap eller parförhållande kan du kontakta familjerådgivningen.
Familjerådgivningsbyråerna är i synnerhet avsedda för familjer med barn.
linkkiEsbo stad:
Familjerådgivningarfinska _ svenska _ engelska
Väestöliitto erbjuder rådgivning och terapi för par på finska och engelska.
linkkiBefolkningsförbundet:
Rådgivning till invandrare telefonledes och via e-postfinska _ svenska _ engelska
Familia Clubs projekt Duo erbjuder relationsrådgivning för par från två kulturer på finska och engelska.
Rådgivningen är avgiftsbelagd.
Relationsrådgivning för par från två kulturerfinska _ engelska
Också kyrkans familjerådgivningscentral erbjuder familjerådgivning vid problem i parförhållandet.
Kyrkans familjerådgivningfinska _ svenska _ engelska
Läs mer: Problem i äktenskap och parförhållande
Barns och ungas problem
Hälsovårdaren vid barnrådgivningen ger råd i frågor som rör hälsan och utvecklingen av barn under skolåldern.
I Esbo finns flera rådgivningsbyråer runtom i staden.
Rådgivningsbyråernas tidsbokning och rådgivning
Tfn (09) 816 22800
linkkiEsbo stad:
Rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
Vid problem som berör barn i skolåldern hjälper till exempel skolans hälsovårdare.
linkkiEsbo stad:
Information om hälsovården för skolbarnfinska _ svenska _ engelska
Om du behöver råd i frågor kring barns psykiska utveckling, kan du boka en tid hos familjerådgivningen.
linkkiEsbo stad:
Familjerådgivningarfinska _ svenska _ engelska
Väestöliitto ger råd till invandrarfamiljer i frågor rörande barnfostran och familjens välmående.
Rådgivningen på olika språk:
Tfn 050 325 7173 (ryska, engelska)
Unga kan prata om sina problem med hälsovårdaren på den egna skolan eller läroanstalten.
Det finns även andra ställen där man kan få hjälp.
En ung i åldern 13–22 år kan få hjälp vid Ungdomspolikliniken Nupoli om hen har problem till exempel med den mentala hälsan, rusmedelsbruk, spelande eller fritidsaktiviteterna.
Man kan ringa eller besöka Nupoli.
Besök på Nupoli är kostnadsfria och konfidentiella.
Tfn 09 816 31300
linkkiEsbo stad:
Nupoli - hjälp för ungafinska _ svenska
Om den unga inte är trygg i sitt eget hem, kan hen kontakta Finlands Röda Kors De ungas skyddshus.
Skyddshuset finns i Alberga.
De ungas skyddshus
Tfn (09) 8195 5360
linkkiFinlands Röda Kors:
De ungas skyddshusfinska
Läs mer: Barns och ungas problem
Om du har ekonomiska problem kan du fråga om råd hos kommunens socialarbetare.
Om du eller din familj inte har tillräckliga inkomster eller tillgångar för den nödvändiga dagliga försörjningen kan du söka grundläggande utkomststöd hos FPA.
Information om utkomststödfinska _ svenska _ engelska _ ryska _ estniska
Om du har problem med skulder, kontakta rättshjälpsbyråns ekonomi- och skuldrådgivning.
Tjänsten är kostnadsfri.
linkkiRättshjälpsbyrå:
Ekonomi- och skuldrådgivningfinska _ svenska _ engelska
Missbruksproblem
Kliniken för mental- och missbruksvård erbjuder vuxna Esbobor hjälp och vård vid problem med den mentala hälsan och missbruk.
Köpcentret Iso Omena
Telefon: 09 816 31300
linkkiEsbo stad:
Information om mentalvårdstjänsternafinska _ svenska _ engelska
Unga i åldern 13-22 med missbruksproblem kan få hjälp vid Ungdomspolikliniken Nupoli.
Tfn 09 816 31300
linkkiEsbo stad:
Nupoli - hjälp för ungafinska _ svenska
Läs mer: Missbruksproblem
Dödsfall
Begravningsbyråer hjälper med de praktiska arrangemangen vid en begravning.
Du kan söka begravningsbyråer till exempel på Finlands begravningsbyråers förbunds webbplats.
linkkiFinlands Begravningbyråers Förbund:
Begravningsbyråerfinska
I Esbo finns fem kristna begravningsplatser.
På Klockarmalmens begravningsplats finns ett gravområde för konfessionslösa.
Där kan de avlidna begravas som hade en annan religionstillhörighet eller inte hörde till något religionssamfund.
linkkiEsbo församlingar:
Begravningsplatserfinska _ svenska _ engelska
Om en närstående dör oväntat och du behöver stöd kan du kontakta social- och krisjouren i Esbo, telefon (09) 816 42439.
Läs mer: Dödsfall
Problem med uppehållstillståndet
Brott
Behöver du en jurist?
Våld Problem i äktenskap eller parförhållande
Barns och ungas problem
Missbruksproblem
Dödsfall
Ring nödnumret 112 om det är fråga om en nödsituation.
Via nödnumret kan du tillkalla polis, ambulans eller brandkår.
Ring inte nödnumret om det inte är en nödsituation.
Läs mer:Nödsituationer
linkkiEsbo stad:
Jourmottagningarfinska _ svenska _ engelska
Social- och krisjouren
Social- och krisjouren (sosiaali- ja kriisipäivystys) hjälper dygnet runt om du eller din familj behöver hjälp i en akut krissituation.
Krisen kan till exempel ha med våld, parförhållandet eller barnens problem att göra.
Du kan även kontakta social- och krisjouren om du har problem med din mentala hälsa, missbruksproblem eller om du råkat ut för en traumatisk händelse i livet.
Social- och krisjouren
Jorvs sjukhus
Åbovägen 150
Tfn (09) 816 42439
Öppet varje dag dygnet runt.
linkkiEsbo stad:
Social- och krisjourenfinska _ svenska _ engelska
Föreningen för mental hälsa i Finland (Suomen Mielenterveysseura) har en krismottagning för invandrare.
Kontoret ligger i Böle i Helsingfors.
Krismottagningen ger dig hjälp och stöd i svåra situationer.
Boka en tid per telefon på numret (09) 4135 0501.
linkkiFöreningen för mental hälsa i Finland:
Krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Problem med uppehållstillståndet
Om du har problem eller oklarheter med uppehållstillståndet, ska du ta kontakt med migrationsverket.
Läs mer: Problem med uppehållstillstånd
Migrationsverkets tjänsteställenfinska _ svenska _ engelska
Om du är flykting, asylsökande eller vistas i Finland av någon annan anledning kan du be om juridisk hjälp och rådgivning vid Flyktingrådgivningen rf.
Kontoret ligger i Helsingfors.
Adress: Kaisaniemigatan 4 A
Tfn 09 2313 9325
linkkiFlyktingrådgivningen r.f.:
Rättshjälp till flyktingarfinska _ svenska _ engelska
Brott
Om du blir utsatt för ett brott, gör en brottsanmälan hos polisen.
Du kan göra brottsanmälan på internet.
Du kan även fylla i en blankett och lämna den till Esbo huvudpolisstation.
Esbo huvudpolisstation
Knektbrogränden 4
Läs mer: Brott
Kontaktuppgifterfinska _ svenska _ engelska
Elektronisk polisanmälanfinska _ svenska _ engelska
Behöver du en jurist?
Om du behöver juridisk hjälp, kan du kontakta Västra Nylands rättshjälpsbyrå.
Biskopsbron 9 B
Tfn 029 56 61820
Läs mer: Behöver du en jurist?
linkkiVästra Nylands rättshjälpsbyrå:
Rättshjälpfinska
Våld
Omatila (Omatila) hjälper dig om du har blivit utsatt för närståendevåld eller våld inom familjen.
Omatila ordnar vid behov boende för dig och dina barn.
Du kan ringa Omatila-tjänsten dygnet runt. Du behöver inte uppge ditt namn när du ringer.
Du kan också komma utan tidsbokning för att prata om din situation, måndag till fredag kl. 9–11 och onsdagar kl. 16–20.
Omatila
Enheten för familjeärenden
Kamrersvägen 6 A
Tfn 043 825 0535
Läs mer: Våld
linkkiEsbo stad:
Hjälp till offer för familjevåldfinska _ svenska _ engelska
Miehen Linja (Miehen Linja) är en tjänst som hjälper män, som har utsatt sina familjemedlemmar för våld. Tjänsten är avsedd för invandrarmän.
Målargränden 3 B
Tfn (09) 276 62899
Hjälp för invandrarmänfinska _ engelska
Problem i äktenskap eller parförhållande
Om du har problem i ditt äktenskap eller parförhållande kan du kontakta familjerådgivningen.
Familjerådgivningsbyråerna är i synnerhet avsedda för familjer med barn.
linkkiEsbo stad:
Familjerådgivningarfinska _ svenska _ engelska
Väestöliitto erbjuder rådgivning och terapi för par på finska och engelska.
linkkiBefolkningsförbundet:
Rådgivning till invandrare telefonledes och via e-postfinska _ svenska _ engelska
Familia Clubs projekt Duo erbjuder relationsrådgivning för par från två kulturer på finska och engelska.
Rådgivningen är avgiftsbelagd.
Relationsrådgivning för par från två kulturerfinska _ engelska
Också kyrkans familjerådgivningscentral erbjuder familjerådgivning vid problem i parförhållandet.
Kyrkans familjerådgivningfinska _ svenska _ engelska
Läs mer: Problem i äktenskap och parförhållande
Barns och ungas problem
Hälsovårdaren vid barnrådgivningen ger råd i frågor som rör hälsan och utvecklingen av barn under skolåldern.
I Esbo finns flera rådgivningsbyråer runtom i staden.
Rådgivningsbyråernas tidsbokning och rådgivning
Tfn (09) 816 22800
linkkiEsbo stad:
Rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
Vid problem som berör barn i skolåldern hjälper till exempel skolans hälsovårdare.
linkkiEsbo stad:
Information om hälsovården för skolbarnfinska _ svenska _ engelska
Om du behöver råd i frågor kring barns psykiska utveckling, kan du boka en tid hos familjerådgivningen.
linkkiEsbo stad:
Familjerådgivningarfinska _ svenska _ engelska
Väestöliitto ger råd till invandrarfamiljer i frågor rörande barnfostran och familjens välmående.
Rådgivningen på olika språk:
Tfn 050 325 7173 (ryska, engelska)
Unga kan prata om sina problem med hälsovårdaren på den egna skolan eller läroanstalten.
Det finns även andra ställen där man kan få hjälp.
En ung i åldern 13–22 år kan få hjälp vid Ungdomspolikliniken Nupoli om hen har problem till exempel med den mentala hälsan, rusmedelsbruk, spelande eller fritidsaktiviteterna.
Man kan ringa eller besöka Nupoli.
Besök på Nupoli är kostnadsfria och konfidentiella.
Tfn 09 816 31300
linkkiEsbo stad:
Nupoli - hjälp för ungafinska _ svenska
Om den unga inte är trygg i sitt eget hem, kan hen kontakta Finlands Röda Kors De ungas skyddshus.
Skyddshuset finns i Alberga.
De ungas skyddshus
Tfn (09) 8195 5360
linkkiFinlands Röda Kors:
De ungas skyddshusfinska
Läs mer: Barns och ungas problem
Om du har ekonomiska problem kan du fråga om råd hos kommunens socialarbetare.
Om du eller din familj inte har tillräckliga inkomster eller tillgångar för den nödvändiga dagliga försörjningen kan du söka grundläggande utkomststöd hos FPA.
Information om utkomststödfinska _ svenska _ engelska _ ryska _ estniska
Om du har problem med skulder, kontakta rättshjälpsbyråns ekonomi- och skuldrådgivning.
Tjänsten är kostnadsfri.
linkkiRättshjälpsbyrå:
Ekonomi- och skuldrådgivningfinska _ svenska _ engelska
Missbruksproblem
Kliniken för mental- och missbruksvård erbjuder vuxna Esbobor hjälp och vård vid problem med den mentala hälsan och missbruk.
Köpcentret Iso Omena
Telefon: 09 816 31300
linkkiEsbo stad:
Information om mentalvårdstjänsternafinska _ svenska _ engelska
Unga i åldern 13-22 med missbruksproblem kan få hjälp vid Ungdomspolikliniken Nupoli.
Tfn 09 816 31300
linkkiEsbo stad:
Nupoli - hjälp för ungafinska _ svenska
Läs mer: Missbruksproblem
Dödsfall
Begravningsbyråer hjälper med de praktiska arrangemangen vid en begravning.
Du kan söka begravningsbyråer till exempel på Finlands begravningsbyråers förbunds webbplats.
linkkiFinlands Begravningbyråers Förbund:
Begravningsbyråerfinska
I Esbo finns fem kristna begravningsplatser.
På Klockarmalmens begravningsplats finns ett gravområde för konfessionslösa.
Där kan de avlidna begravas som hade en annan religionstillhörighet eller inte hörde till något religionssamfund.
linkkiEsbo församlingar:
Begravningsplatserfinska _ svenska _ engelska
Om en närstående dör oväntat och du behöver stöd kan du kontakta social- och krisjouren i Esbo, telefon (09) 816 42439.
Läs mer: Dödsfall
Äktenskap
Skilsmässa
Registrerat parförhållande
Vård av barn Invånarparker och klubbar
Problem i familjen
Äktenskap
Före äktenskapet ska du skriftligt begära hindersprövning (avioliiton esteiden tutkiminen).
Hindersprövningen görs på magistraten (maistraatti).
Du kan begära hindersprövning på vilken magistrat som helst.
Magistraten i Nyland, Esbo enhet
Miestentie 3
Tfn 029 553 9391
Läs mer: Äktenskap.
Vigselfinska _ svenska _ engelska
Anhållan om prövning av hinder mot äktenskapfinska _ svenska
Skilsmässa
Kvinnan eller mannen kan lämna in skilsmässoansökan i Västra Nylands tingsrätts kansli.
Du kan också söka skilsmässa ensam, utan din makes eller makas samtycke.
Du kan skicka in ansökan till tingsrättens kansli per post, fax eller via e-post.
Tfn 029 564 4000
Läs mer: Skilsmässa.
linkkiVästra Nylands tingsrätt:
Kontaktuppgifterfinska _ svenska
Barn vid skilsmässa
Om du har barn under 13 år och överväger att skilja dig, ta kontakt med familjerådgivningen (perheneuvola).
På familjerådgivningen kan du diskutera familjens situation med de anställda.
Familjerådgivningarnas kontaktuppgifter finns på Esbo stads webbplats.
Om du planerar skilsmässa kan du också ta kontakt med barnatillsyningsmannen (lastenvalvoja) vid enheten för familjeärenden.
Med barnatillsyningsmannen kan du diskutera skilsmässan och barnens framtid.
Makarna ska ingå ett avtal om barnens boende, umgängesrätt och underhållsbidrag.
Barnatillsyningsmännen bekräftar avtalet.
Kontaktuppgifterna till barnatillsyningsmännen finns på Esbo stads webbplats.
Esbo stad har en rådgivningstelefon där man kan fråga om råd i frågor rörande barnen när föräldrarna skiljer sig.
Tfn 046 877 3267
Läs mer: Barn vid skilsmässa.
linkkiEsbo stad:
Kontaktuppgifter till barnatillsyningsmännenfinska _ svenska
linkkiEsbo stad:
Skilsmässa i en barnfamiljfinska _ svenska
Vård av barn
Information om dagvård av barn i Esbo finns på InfoFinlands sida Utbildning i Esbo.
Tillfällig vård av barn
Du kan föra barnet till en parktant för tillfällig vård.
Det innebär kortvarig (2–3 tim. per gång) vård av småbarn ute i en lekpark.
Du får närmare uppgifter av parktanterna per telefon.
Du hittar telefonnumren på Esbo stads webbplats.
linkkiEsbo stad:
Parktanterfinska
Om du behöver en tillfällig barnskötare hem, kan du kontakta Mannerheims Barnskyddsförbund eller Väestöliitto.
Barnavård och hemhjälpfinska
linkkiMannerheims Barnskyddsförbund:
Barnavårdfinska _ svenska _ engelska
Läs mer: Dagvård.
Hemvårdsstöd
Om familjens yngsta barn är under tre år, kan barnets förälder få hemvårdsstöd (kotihoidon tuki) när han eller hon vårdar barnet i hemmet.
Om du har rätt till hemvårdsstödet kan du ansöka om det hos FPA.
Du kan fylla i ansökan på Internet eller posta den till FPA.
Du kan också besöka FPA:s kontor.
Esbo stad betalar ett kommuntillägg till de familjer som vårdar ett under treårigt barn i hemmet.
Man kan ansöka om Esbotillägget om en förälder tar hand om familjens alla barn under skolåldern i hemmet.
linkkiEsbo stad:
Vård av barn i hemmetfinska _ svenska _ engelska
Information om hemvårdsstödfinska _ svenska _ engelska
Sköta ärenden på Internetfinska _ svenska _ engelska
Kontaktuppgifter till FPAfinska _ svenska _ engelska
Invånarparker och klubbar
Esbo stad ordnar mycket verksamhet för de föräldrar som vårdar barn i hemmet. Det finns till exempel invånarparker, öppna daghem och klubbar.
Läs mer: Stöd för vård av barn i hemmet
linkkiEsbo stad:
Invånarparker och klubbarfinska _ engelska
Problem i familjen
På InfoFinlands sida Problematiska situationer i Esbo hittar du uppgifter om vart du kan vända dig i Esbo för att få hjälp vid barns och ungas problem och problem i familjen.
Du hittar uppgifter om barns och ungas problem också på InfoFinlands sida Barns och ungas problem och Var hittar jag hjälp när barn eller unga har problem?
På InfoFinlands sida Problem i äktenskap och parförhållande finns uppgifter om vart du kan vända dig för att få hjälp vid problem i parförhållandet.
Äktenskap
Skilsmässa
Registrerat parförhållande
Vård av barn Invånarparker och klubbar
Problem i familjen
Äktenskap
Före äktenskapet ska du skriftligt begära hindersprövning (avioliiton esteiden tutkiminen).
Hindersprövningen görs på magistraten (maistraatti).
Du kan begära hindersprövning på vilken magistrat som helst.
Magistraten i Nyland, Esbo enhet
Miestentie 3
Tfn 029 553 9391
Läs mer: Äktenskap.
Vigselfinska _ svenska _ engelska
Anhållan om prövning av hinder mot äktenskapfinska _ svenska
Skilsmässa
Kvinnan eller mannen kan lämna in skilsmässoansökan i Västra Nylands tingsrätts kansli.
Du kan också söka skilsmässa ensam, utan din makes eller makas samtycke.
Du kan skicka in ansökan till tingsrättens kansli per post, fax eller via e-post.
Tfn 029 564 4000
Läs mer: Skilsmässa.
linkkiVästra Nylands tingsrätt:
Kontaktuppgifterfinska _ svenska
Barn vid skilsmässa
Om du har barn under 13 år och överväger att skilja dig, ta kontakt med familjerådgivningen (perheneuvola).
På familjerådgivningen kan du diskutera familjens situation med de anställda.
Familjerådgivningarnas kontaktuppgifter finns på Esbo stads webbplats.
Om du planerar skilsmässa kan du också ta kontakt med barnatillsyningsmannen (lastenvalvoja) vid enheten för familjeärenden.
Med barnatillsyningsmannen kan du diskutera skilsmässan och barnens framtid.
Makarna ska ingå ett avtal om barnens boende, umgängesrätt och underhållsbidrag.
Barnatillsyningsmännen bekräftar avtalet.
Kontaktuppgifterna till barnatillsyningsmännen finns på Esbo stads webbplats.
Esbo stad har en rådgivningstelefon där man kan fråga om råd i frågor rörande barnen när föräldrarna skiljer sig.
Tfn 046 877 3267
Läs mer: Barn vid skilsmässa.
linkkiEsbo stad:
Kontaktuppgifter till barnatillsyningsmännenfinska _ svenska
linkkiEsbo stad:
Skilsmässa i en barnfamiljfinska _ svenska
Vård av barn
Information om dagvård av barn i Esbo finns på InfoFinlands sida Utbildning i Esbo.
Tillfällig vård av barn
Du kan föra barnet till en parktant för tillfällig vård.
Det innebär kortvarig (2–3 tim. per gång) vård av småbarn ute i en lekpark.
Du får närmare uppgifter av parktanterna per telefon.
Du hittar telefonnumren på Esbo stads webbplats.
linkkiEsbo stad:
Parktanterfinska
Om du behöver en tillfällig barnskötare hem, kan du kontakta Mannerheims Barnskyddsförbund eller Väestöliitto.
Barnavård och hemhjälpfinska
linkkiMannerheims Barnskyddsförbund:
Barnavårdfinska _ svenska _ engelska
Läs mer: Dagvård.
Hemvårdsstöd
Om familjens yngsta barn är under tre år, kan barnets förälder få hemvårdsstöd (kotihoidon tuki) när han eller hon vårdar barnet i hemmet.
Om du har rätt till hemvårdsstödet kan du ansöka om det hos FPA.
Du kan fylla i ansökan på Internet eller posta den till FPA.
Du kan också besöka FPA:s kontor.
Esbo stad betalar ett kommuntillägg till de familjer som vårdar ett under treårigt barn i hemmet.
Man kan ansöka om Esbotillägget om en förälder tar hand om familjens alla barn under skolåldern i hemmet.
linkkiEsbo stad:
Vård av barn i hemmetfinska _ svenska _ engelska
Information om hemvårdsstödfinska _ svenska _ engelska
Sköta ärenden på Internetfinska _ svenska _ engelska
Kontaktuppgifter till FPAfinska _ svenska _ engelska
Invånarparker och klubbar
Esbo stad ordnar mycket verksamhet för de föräldrar som vårdar barn i hemmet. Det finns till exempel invånarparker, öppna daghem och klubbar.
Läs mer: Stöd för vård av barn i hemmet
linkkiEsbo stad:
Invånarparker och klubbarfinska _ engelska
Äldre människor
Åldringar kan använda tjänsterna vid de vanliga hälsostationerna.
Dessutom erbjuds åldringar i Esbo egna tjänster, till exempel hemvårdens tjänster.
Om du vill ha mer information om tjänster för äldre kan du kontakta seniorrådgivningen (seniorineuvonta).
tfn (09) 816 33333
linkkiEsbo stad:
Seniorrådgivningenfinska _ svenska _ engelska
När du tar hand om en anhörig i hemmet
Om du tar hand om en äldre, sjuk eller handikappad anhörig hemma så att hen ska kunna bo hemma, kan du ha rätt till stöd för närståendevård.
linkkiEsbo stad:
Stöd för närståendevårdfinska _ svenska
Äldre människor
Problem i familjen
På InfoFinlands sida Problematiska situationer i Esbo hittar du uppgifter om vart du kan vända dig i Esbo för att få hjälp vid barns och ungas problem och problem i familjen.
Du hittar uppgifter om barns och ungas problem också på InfoFinlands sida Barns och ungas problem och Var hittar jag hjälp när barn eller unga har problem?
På InfoFinlands sida Problem i äktenskap och parförhållande finns uppgifter om vart du kan vända dig för att få hjälp vid problem i parförhållandet.
Äktenskap
Skilsmässa
Registrerat parförhållande
Vård av barn Invånarparker och klubbar
Problem i familjen
Äktenskap
Före äktenskapet ska du skriftligt begära hindersprövning (avioliiton esteiden tutkiminen).
Hindersprövningen görs på magistraten (maistraatti).
Du kan begära hindersprövning på vilken magistrat som helst.
Magistraten i Nyland, Esbo enhet
Miestentie 3
Tfn 029 553 9391
Läs mer: Äktenskap.
Vigselfinska _ svenska _ engelska
Anhållan om prövning av hinder mot äktenskapfinska _ svenska
Skilsmässa
Kvinnan eller mannen kan lämna in skilsmässoansökan i Västra Nylands tingsrätts kansli.
Du kan också söka skilsmässa ensam, utan din makes eller makas samtycke.
Du kan skicka in ansökan till tingsrättens kansli per post, fax eller via e-post.
Tfn 029 564 4000
Läs mer: Skilsmässa.
linkkiVästra Nylands tingsrätt:
Kontaktuppgifterfinska _ svenska
Barn vid skilsmässa
Om du har barn under 13 år och överväger att skilja dig, ta kontakt med familjerådgivningen (perheneuvola).
På familjerådgivningen kan du diskutera familjens situation med de anställda.
Familjerådgivningarnas kontaktuppgifter finns på Esbo stads webbplats.
Om du planerar skilsmässa kan du också ta kontakt med barnatillsyningsmannen (lastenvalvoja) vid enheten för familjeärenden.
Med barnatillsyningsmannen kan du diskutera skilsmässan och barnens framtid.
Makarna ska ingå ett avtal om barnens boende, umgängesrätt och underhållsbidrag.
Barnatillsyningsmännen bekräftar avtalet.
Kontaktuppgifterna till barnatillsyningsmännen finns på Esbo stads webbplats.
Esbo stad har en rådgivningstelefon där man kan fråga om råd i frågor rörande barnen när föräldrarna skiljer sig.
Tfn 046 877 3267
Läs mer: Barn vid skilsmässa.
linkkiEsbo stad:
Kontaktuppgifter till barnatillsyningsmännenfinska _ svenska
linkkiEsbo stad:
Skilsmässa i en barnfamiljfinska _ svenska
Vård av barn
Information om dagvård av barn i Esbo finns på InfoFinlands sida Utbildning i Esbo.
Tillfällig vård av barn
Du kan föra barnet till en parktant för tillfällig vård.
Det innebär kortvarig (2–3 tim. per gång) vård av småbarn ute i en lekpark.
Du får närmare uppgifter av parktanterna per telefon.
Du hittar telefonnumren på Esbo stads webbplats.
linkkiEsbo stad:
Parktanterfinska _ svenska
Om du behöver en tillfällig barnskötare hem, kan du kontakta Mannerheims Barnskyddsförbund eller Väestöliitto.
Barnavård och hemhjälpfinska
linkkiMannerheims Barnskyddsförbund:
Barnavårdfinska _ svenska _ engelska
Läs mer: Dagvård.
Hemvårdsstöd
Om familjens yngsta barn är under tre år, kan barnets förälder få hemvårdsstöd (kotihoidon tuki) när han eller hon vårdar barnet i hemmet.
Om du har rätt till hemvårdsstödet kan du ansöka om det hos FPA.
Du kan fylla i ansökan på Internet eller posta den till FPA.
Du kan också besöka FPA:s kontor.
Esbo stad betalar ett kommuntillägg till de familjer som vårdar ett under treårigt barn i hemmet.
Man kan ansöka om Esbotillägget om en förälder tar hand om familjens alla barn under skolåldern i hemmet.
linkkiEsbo stad:
Vård av barn i hemmetfinska _ svenska _ engelska
Information om hemvårdsstödfinska _ svenska _ engelska
Sköta ärenden på Internetfinska _ svenska _ engelska
Kontaktuppgifter till FPAfinska _ svenska _ engelska
Invånarparker och klubbar
Esbo stad ordnar mycket verksamhet för de föräldrar som vårdar barn i hemmet. Det finns till exempel invånarparker, öppna daghem och klubbar.
Läs mer: Stöd för vård av barn i hemmet
linkkiEsbo stad:
Invånarparker och klubbarfinska _ engelska
Äldre människor
Åldringar kan använda tjänsterna vid de vanliga hälsostationerna.
Dessutom erbjuds åldringar i Esbo egna tjänster, till exempel hemvårdens tjänster.
Om du vill ha mer information om tjänster för äldre kan du kontakta seniorrådgivningen (seniorineuvonta).
tfn (09) 816 33333
linkkiEsbo stad:
Seniorrådgivningenfinska _ svenska _ engelska
När du tar hand om en anhörig i hemmet
Om du tar hand om en äldre, sjuk eller handikappad anhörig hemma så att hen ska kunna bo hemma, kan du ha rätt till stöd för närståendevård.
linkkiEsbo stad:
Stöd för närståendevårdfinska _ svenska
Äldre människor
Problem i familjen
På InfoFinlands sida Problematiska situationer i Esbo hittar du uppgifter om vart du kan vända dig i Esbo för att få hjälp vid barns och ungas problem och problem i familjen.
Du hittar uppgifter om barns och ungas problem också på InfoFinlands sida Barns och ungas problem och Var hittar jag hjälp när barn eller unga har problem?
På InfoFinlands sida Problem i äktenskap och parförhållande finns uppgifter om vart du kan vända dig för att få hjälp vid problem i parförhållandet.
Hälsovårdstjänsterna i Esbo
Äldre människors hälsa
Tandvården
Mental hälsa
Sexuell hälsa
När du väntar barn
Handikappade personer
Ring nödnumret 112 om det är fråga om en brådskande nödsituation.
Ring nödnumret till exempel vid en allvarlig olycka eller när någon drabbas av en sjukdomsattack.
Ring inte nödnumret om det inte är en nödsituation.
Om du har din hemkommun i Esbo kan du utnyttja de offentliga hälsovårdstjänsterna.
Offentliga hälsovårdstjänster tillhandahålls vid hälsostationer, tandkliniker, rådgivningsbyråer och sjukhus.
Om du inte har rätt till de offentliga hälsovårdstjänsterna, kan du söka hjälp på en privat läkarstation.
På en privat läkarstation måste du betala samtliga kostnader själv.
Läs mer: Hälsa.
Hälsovårdstjänsterna i Esbo
Offentliga hälsovårdstjänster tillhandahålls av hälsostationerna (terveysasema).
Hälsostationerna har öppet vardagar klockan 8–16.
På hälsostationerna finns vanligtvis läkarens, sjukskötarens och hälsovårdarens mottagningar.
Du kan boka tid på hälsostationen per telefon.
På Esbo stads webbplats finns kontaktuppgifterna och telefonnumren till hälsostationerna.
När du ringer hälsostationen, besvaras ditt samtal inte nödvändigtvis omedelbart.
Ditt nummer sparas dock i en automat och du blir uppringd.
Kom i tid till mottagningen.
Om du inte kan komma till mottagningen, kom ihåg att avboka din tid senast föregående vardag före klockan 14.
Om du behöver första hjälpen snabbt, kan du komma till hälsostationen utan tidsbeställning.
linkkiEsbo stad:
Hälsostationernafinska _ svenska _ engelska
linkkiEsbo stad:
Hälsovårdscentralsavgifterfinska _ svenska
Privata hälsovårdstjänster
Vem som helst kan gå till en privat hälsostation.
Också de personer som inte har rätt till den offentliga hälsovården i Finland kan besöka privata hälsostationer.
På en privat hälsostation måste kunden själv betala samtliga kostnader.
I Esbo finns flera privata läkarstationer.
Kontaktuppgifter till privata läkare hittar du till exempel på Internet.
linkkietsilaakari.fi:
Privata hälsovårdstjänsterfinska
Privat läkarstationfinska _ svenska _ engelska
Privat läkarstationfinska _ svenska _ engelska
Läkemedel
Information om köp av läkemedel hittar du på InfoFinlands sida Läkemedel.
Hälsovård för papperslösa
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärhälsovård.
Tjänsterna vid Global Clinic är avgiftsfria för kunderna.
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter.
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
Telefonnumret till Global Clinic i Helsingfors är 044 977 4547.
Samtalet besvaras av en sjukskötare eller en läkare.
Hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Läs mer: Hälsovårdstjänster i Finland
Kvällstid och under veckoslut har hälsostationen stängt.
Då vårdas akuta sjukfall och olycksfall på jourmottagningen (päivystys).
Den närmaste jourmottagningen för vuxna finns vid Jorv sjukhus.
Ring den kostnadsfria Jourhjälpen på tfn 116 117 innan du kommer till jourmottagningen.
Jourmottagningen vid Jorv sjukhus
Åbovägen 150
Tfn (09) 4711
Jourmottagningar för barn under 16 år finns i Jorv och på Barnkliniken i Helsingfors.
Du behöver inte boka tid på jourmottagningen.
linkkiEsbo stad:
Jourmottagningarfinska _ svenska _ engelska
Läs mer: Hälsovårdstjänster i Finland
Barns hälsa
I hälsovården av 1–6-åriga barn får man hjälp av rådgivningsbyråns (neuvola) hälsovårdare och läkare.
Dem kan du fråga om råd och få hjälp med fostran av barn.
På rådgivningsbyrån följs att barnet är friskt och växer som det ska.
I Esbo finns flera rådgivningsbyråer på olika håll i staden.
Rådgivningsbyråernas kontaktuppgifter finns på Esbo stads webbplats.
Du kan boka tid vid alla rådgivningsbyråer på samma nummer.
Om ett barn blir sjukt och behöver snabbt vård, ta kontakt med hälsostationen (terveysasema).
Skolhälsovårdaren har hand om skolbarns hälsa.
Under kvällar och veckoslut finns jourmottagningen för barn under 16 år vid Jorv sjukhus och på Barnkliniken i Helsingfors.
Du kan också ta ditt barn till en privat läkarstation.
Läs mer: Barns hälsa.
linkkiEsbo stad:
Barnrådgivningsbyråernas tjänsterfinska _ svenska _ engelska
linkkiEsbo stad:
Rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
linkkiEsbo stad:
Hälsostationernafinska _ svenska _ engelska
linkkiEsbo stad:
Information om hälsovården för skolbarnfinska _ svenska _ engelska
linkkiEsbo stad:
Jourmottagningarfinska _ svenska _ engelska
Äldre människors hälsa
Åldringar kan använda tjänsterna vid de vanliga hälsostationerna.
Dessutom erbjuds åldringar i Esbo egna tjänster, till exempel hemvårdens tjänster.
Om du vill ha mer information om tjänster för äldre kan du kontakta seniorrådgivningen (seniorineuvonta).
tfn (09) 816 33333
linkkiEsbo stad:
Seniorrådgivningenfinska _ svenska
När du tar hand om en anhörig i hemmet
Om du tar hand om en äldre, sjuk eller handikappad anhörig hemma så att hen ska kunna bo hemma, kan du ha rätt till stöd för närståendevård.
linkkiEsbo stad:
Stöd för närståendevårdfinska _ svenska
Äldre människors hälsa, Äldre människor
Tandvården
