����      ]�(�numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i4�����R�(K�<�NNNJ����J����K t�b�C8"   6  (      �	  \        �      0   �         �t�bhhK ��h��R�(KK��h�CX   E       �        �t�bhhK ��h��R�(KK��h�C0           I         $     �        �t�bhhK ��h��R�(KK	��h�C$   ?   #   !   
      F         �t�bhhK ��h��R�(KK��h�C�      a     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C  �        �   r      �t�bhhK ��h��R�(KK��h�C|
   3   6      w     @   (      !      �      @   2      0   <      �     �  m         "   m      �         �t�bhhK ��h��R�(KK��h�Cp   Y        S   X  i   ,            �  �  �     T        �  P        �                �t�bhhK ��h��R�(KK��h�C@�        �
        F     �         �  9  7         �t�bhhK ��h��R�(KK��h�CT   ,   �         �   f              9   q   L         �      �        �t�bhhK ��h��R�(KK��h�Ch�  �     =  �  (                                 A   :      a  �         	        �t�bhhK ��h��R�(KK��h�C4
         2   �        \   #  &   �        �t�bhhK ��h��R�(KK#��h�C�         �           .      0      n	  �  g	     &      �        $                       \      �  $            �t�bhhK ��h��R�(KK��h�C@   �      .        '   )   
               K         �t�bhhK ��h��R�(KK��h�C,�     �     �        e           �t�bhhK ��h��R�(KK��h�Ch	       p      u      �t�bhhK ��h��R�(KK
��h�C(   ^  v       �     �        �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   6                  �t�bhhK ��h��R�(KK��h�Cp            �   �     �      F        b  h      7      �   L   
        G      �   

        �t�bhhK ��h��R�(KK��h�CP              �     �   �   S     U   q   �  �    �  O        �t�bhhK ��h��R�(KK!��h�C�   �     8              )               
   $   �  �  N         I        R  D         M   �               �t�bhhK ��h��R�(KK��h�CD"   �             �           �    h  9   �        �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C      &     $   �         �t�bhhK ��h��R�(KK��h�Ch         �           �      �   9               ;      �  �   �     (      "        �t�bhhK ��h��R�(KK��h�C�  5	  	         �t�bhhK ��h��R�(KK	��h�C$)   �   Y           �         �t�bhhK ��h��R�(KK��h�C,      �
  `            �           �t�bhhK ��h��R�(KK	��h�C$X      �  T     [  
        �t�bhhK ��h��R�(KK��h�C@   �   �     Y      O               Y      O         �t�bhhK ��h��R�(KK��h�Cd      �  +      .         F	  �           
   $   �        `   �      `   �        �t�bhhK ��h��R�(KK��h�C<         $   k      e         ,  %   �           �t�bhhK ��h��R�(KK��h�C8   �        .               >      �        �t�bhhK ��h��R�(KK
��h�C(  �  )   [     C  �           �t�bhhK ��h��R�(KK��h�C)     $   �     �t�bhhK ��h��R�(KK��h�C�      V     �t�bhhK ��h��R�(KK��h�C0      A     �  Y     	      	         �t�bhhK ��h��R�(KK	��h�C$T   >   �  (       |        �t�bhhK ��h��R�(KK
��h�C(      )   6        �            �t�bhhK ��h��R�(KK��h�C      �     �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C,�  �     C      �  �  �           �t�bhhK ��h��R�(KK��h�C*      �  /      �t�bhhK ��h��R�(KK	��h�C$�      ^        $           �t�bhhK ��h��R�(KK��h�C<            G  >      �                       �t�bhhK ��h��R�(KK��h�C0      �        �   f                 �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C                �t�bhhK ��h��R�(KK��h�C �   �   �     �  �        �t�bhhK ��h��R�(KK��h�CH*                   (         w     �  �              �t�bhhK ��h��R�(KK��h�C\   H   7              �t�bhhK ��h��R�(KK��h�C   �  )         �t�bhhK ��h��R�(KK��h�C8  R   8   �  �  h    
   �     8   E        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C�  �      �t�bhhK ��h��R�(KK	��h�C$-   �        m              �t�bhhK ��h��R�(KK��h�C�	  �	     �t�bhhK ��h��R�(KK��h�C\
           �   �     -           T         �           �  
   �        �t�bhhK ��h��R�(KK��h�C�  
   a        �t�bhhK ��h��R�(KK��h�C<      )   �                        V  �         �t�bhhK ��h��R�(KK��h�C   e   '   �   �        �t�bhhK ��h��R�(KK��h�C0n     �     Y        	      	         �t�bhhK ��h��R�(KK��h�C8!      |      <  R      u   ,   	      	         �t�bhhK ��h��R�(KK��h�CT*   �   _  C   &   %   �              D   �      �  J                 �t�bhhK ��h��R�(KK��h�Cd   8                             &      �   �     b                  �        �t�bhhK ��h��R�(KK,��h�C�               n               *  
   �      �     $   k      x        w         $   k               �   D  �           .   �   �     �        �t�bhhK ��h��R�(KK��h�Cx      �      -  �      �t�bhhK ��h��R�(KK��h�C  0  �     `     �t�bhhK ��h��R�(KK��h�Cp   f   �         -   0            .         :  
      �     "            ~   
   B           �t�bhhK ��h��R�(KK��h�C  >     �  !         �t�bhhK ��h��R�(KK��h�C8   �           c  �   (      �  G   �         �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C1     �        �t�bhhK ��h��R�(KK��h�C4   >   v   �          �      �  4         �t�bhhK ��h��R�(KK��h�CD        `      �  �      �     A        �  �        �t�bhhK ��h��R�(KK��h�CLg      �  a  c   &         �   =            h         7         �t�bhhK ��h��R�(KK
��h�C(  
   �  �  W  
   �           �t�bhhK ��h��R�(KK��h�C8
   f     �   )            ,   �      u         �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�CX�     N     �     �                *     �   Y     �     �        �t�bhhK ��h��R�(KK��h�C0            \         +               �t�bhhK ��h��R�(KK��h�C   @   '   H            �t�bhhK ��h��R�(KK��h�CP         �     �     %   �   �     $     �        �   �        �t�bhhK ��h��R�(KK��h�CH      0   <      $         .   "   �                       �t�bhhK ��h��R�(KK��h�C8   
      {            �      �  $   
        �t�bhhK ��h��R�(KK��h�CP      -   =      H   �  4      Y      n  
        �   �           �t�bhhK ��h��R�(KK	��h�C$   e   '   �                  �t�bhhK ��h��R�(KK��h�C�   p      �t�bhhK ��h��R�(KK��h�CD   >   2     w        �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C8         �t�bhhK ��h��R�(KK��h�C<�   �  �     .   "   �     �	     +     y        �t�bhhK ��h��R�(KK��h�C,�      (  d            R        �t�bhhK ��h��R�(KK	��h�C$t     �      n     k         �t�bhhK ��h��R�(KK��h�C    @     �              �t�bhhK ��h��R�(KK��h�CD   �     y  �  4     P     �                       �t�bhhK ��h��R�(KK	��h�C$         I     "            �t�bhhK ��h��R�(KK��h�CL      5             9   �           U   Q  �     @         �t�bhhK ��h��R�(KK��h�C@      �                �     %                 �t�bhhK ��h��R�(KK��h�CD
        �     (      !        �     5               �t�bhhK ��h��R�(KK��h�C@   D         �   O   >   �   �   �   a   4               �t�bhhK ��h��R�(KK��h�CZ         �t�bhhK ��h��R�(KK��h�C4a  7  
   �      %   }                    �t�bhhK ��h��R�(KK��h�C   �         �        �t�bhhK ��h��R�(KK��h�C'  �        �t�bhhK ��h��R�(KK��h�C,�  �      �      /      �           �t�bhhK ��h��R�(KK��h�C4   @   '   )         5  O        �         �t�bhhK ��h��R�(KK��h�C  �
       �        �t�bhhK ��h��R�(KK	��h�C$   =         	      	         �t�bhhK ��h��R�(KK��h�C�  �  "        �t�bhhK ��h��R�(KK��h�C �        K              �t�bhhK ��h��R�(KK��h�C,      )   �            �   S        �t�bhhK ��h��R�(KK��h�CPE          <      �         �      S   :   �  �	     :            �t�bhhK ��h��R�(KK��h�CD   �  l  g      �	              �   �   �     [         �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C<   '            X        �   ^                 �t�bhhK ��h��R�(KK��h�C  
   �     �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6            �t�bhhK ��h��R�(KK��h�C�  R         	         �t�bhhK ��h��R�(KK��h�CP         9     7      B        2
     �   
   |         F         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C0     �	     2  *      �  (   �        �t�bhhK ��h��R�(KK��h�C,   �   )   x      8     &   �        �t�bhhK ��h��R�(KK	��h�C$      $  V                 �t�bhhK ��h��R�(KK��h�C�       �t�bhhK ��h��R�(KK��h�C8b      �  
      *   $   r  �     L  L        �t�bhhK ��h��R�(KK��h�C,b   "   �     	       $   x        �t�bhhK ��h��R�(KK
��h�C('  �  �         	      	         �t�bhhK ��h��R�(KK��h�Cd      '  �           �	     �  t     $   k   v   [                    +         �t�bhhK ��h��R�(KK��h�C,   �     u  Y        �  R         �t�bhhK ��h��R�(KK��h�Cl   �               �      &     ]                 A  �   �   �              �  �     �t�bhhK ��h��R�(KK��h�C,      �         �   �     J         �t�bhhK ��h��R�(KK��h�C    &   a   �   �  |        �t�bhhK ��h��R�(KK��h�C<      �  �	  �         
        J     �        �t�bhhK ��h��R�(KK��h�C�  k         �t�bhhK ��h��R�(KK��h�CL   Y      O         =      �  "      �        �              �t�bhhK ��h��R�(KK��h�C4      �           �                    �t�bhhK ��h��R�(KK��h�C@6  J     	      	      	   K   	     	   �  	   �      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C\   X   '              �                     ^        �      -  u         �t�bhhK ��h��R�(KK��h�C            	         �t�bhhK ��h��R�(KK
��h�C(4   
      d     	      	         �t�bhhK ��h��R�(KK��h�CH          &     �t�bhhK ��h��R�(KK��h�CL   $   �  {           =      �  �              "   �        �t�bhhK ��h��R�(KK��h�CD      0      :               T         +      f        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK
��h�C(     �      D   �  �   �        �t�bhhK ��h��R�(KK��h�C<�   L        G   t      �     \  L   �            �t�bhhK ��h��R�(KK'��h�C�      =      m                �   �                             S   �     Q     Q      x           _  �      "           �t�bhhK ��h��R�(KK
��h�C(   �        g   �   �            �t�bhhK ��h��R�(KK&��h�C�   n        t        Y      O   v  -         �         l           �  �        �  C   w      �   t     &   4              �t�bhhK ��h��R�(KK��h�CX         &   D  0      k         >      4        N   �   l              �t�bhhK ��h��R�(KK	��h�C$f     g  /  	      	         �t�bhhK ��h��R�(KK��h�C   k         �t�bhhK ��h��R�(KK��h�C{      s     �t�bhhK ��h��R�(KK
��h�C(�           d                  �t�bhhK ��h��R�(KK��h�C\        r      �t�bhhK ��h��R�(KK��h�CX         i     0     M   T   )     
        �  �     #  %   �        �t�bhhK ��h��R�(KK��h�CT      J   =         +     �        �     +  
   �  �  /  F         �t�bhhK ��h��R�(KK��h�C�      J  /         �t�bhhK ��h��R�(KK��h�C`@        0               0   �  b  �   �   {      �  }     
   �   S           �t�bhhK ��h��R�(KK��h�C<      =                 E         �           �t�bhhK ��h��R�(KK��h�CT�           ;     v  l      5      <   �            >              �t�bhhK ��h��R�(KK��h�C4        �        8   S     �  �        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C8            B  �      *         �   �         �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK	��h�C$0     0   �  "      �        �t�bhhK ��h��R�(KK��h�C@#   !   (         .   
   �	  F           @  �
        �t�bhhK ��h��R�(KK��h�C�   `     �t�bhhK ��h��R�(KK��h�CL
   �   F   '   )      �              !      �                  �t�bhhK ��h��R�(KK
��h�C(      )   
  �  ^   &  �         �t�bhhK ��h��R�(KK��h�C08      \     %  }        0           �t�bhhK ��h��R�(KK��h�C g	  &   5  M     �        �t�bhhK ��h��R�(KK��h�C         M     �t�bhhK ��h��R�(KK	��h�C$�	     �     	      	         �t�bhhK ��h��R�(KK��h�C1   #       �     �t�bhhK ��h��R�(KK��h�C,*      J   4  5         J  �         �t�bhhK ��h��R�(KK��h�CH      -   �         �  �   �      �   
   ,      
            �t�bhhK ��h��R�(KK��h�Cq        �t�bhhK ��h��R�(KK��h�C �  &   �  j
              �t�bhhK ��h��R�(KK
��h�C(m     Y      �   $  �  �        �t�bhhK ��h��R�(KK��h�C         .   �        �t�bhhK ��h��R�(KK��h�C      �  -            �t�bhhK ��h��R�(KK��h�CX   2   �     %        v     �         2   -   �   +     -	              �t�bhhK ��h��R�(KK	��h�C$      �          �        �t�bhhK ��h��R�(KK��h�C               �t�bhhK ��h��R�(KK��h�C,X        k         �  �            �t�bhhK ��h��R�(KK��h�C �        	      	         �t�bhhK ��h��R�(KK��h�CZ         Z         �t�bhhK ��h��R�(KK��h�C \   �   2         �  r      �t�bhhK ��h��R�(KK��h�CL         8   �   �      e      &      F  +           <        �t�bhhK ��h��R�(KK��h�C�  �  u        �t�bhhK ��h��R�(KK��h�C1   #            �t�bhhK ��h��R�(KK
��h�C(         �  �   �      D         �t�bhhK ��h��R�(KK	��h�C$�      �        �           �t�bhhK ��h��R�(KK��h�C\   $   �      z        $   �  �         �           �                    �t�bhhK ��h��R�(KK��h�C<j
     ;      �   ]         �  f
     o	  ]         �t�bhhK ��h��R�(KK��h�C\#   !                  �     >        �   �        �   '   
   �   F         �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�C�      R        �t�bhhK ��h��R�(KK%��h�C�         O      �      %     z        Y      Q         Q     Q         x     �               �      5      7  4         �t�bhhK ��h��R�(KK��h�C1   #       x     e      �t�bhhK ��h��R�(KK��h�C0      �   f    �   �  H   �  �        �t�bhhK ��h��R�(KK��h�C      0  c     N
     �t�bhhK ��h��R�(KK
��h�C(      �  c   I  
   �  F         �t�bhhK ��h��R�(KK��h�CD      /   �     :     &      M   �           �        �t�bhhK ��h��R�(KK	��h�C$�  �     �     ,            �t�bhhK ��h��R�(KK��h�C!     	      	         �t�bhhK ��h��R�(KK��h�CD%   �        
   ,            �      '   )   A   #         �t�bhhK ��h��R�(KK��h�C8   �   �  �      m  >   �     m     ]         �t�bhhK ��h��R�(KK	��h�C$      '   H   j     u         �t�bhhK ��h��R�(KK��h�C@@      q   b  E      V      q         V   '            �t�bhhK ��h��R�(KK��h�C<)      @           �   e   �  �                 �t�bhhK ��h��R�(KK��h�C$  �     �t�bhhK ��h��R�(KK��h�CT*      �  8   o           &      }        �     �  �      5        �t�bhhK ��h��R�(KK��h�C4   e   '   H   B      V   2      �   �        �t�bhhK ��h��R�(KK��h�C\   �        �          u            �   �      �     �                  �t�bhhK ��h��R�(KK��h�CH      P      1     .   
   q      F      ^   �               �t�bhhK ��h��R�(KK��h�C�     b        �t�bhhK ��h��R�(KK��h�CL      -   �           +      z     �        �  9   �        �t�bhhK ��h��R�(KK	��h�C$      �        (            �t�bhhK ��h��R�(KK��h�CX)         d  j  
      �     C      +         �   �  )   6  +   ,         �t�bhhK ��h��R�(KK��h�C,   �      %   �     "              �t�bhhK ��h��R�(KK��h�CL      �     u   �  {      Q       u               �        �t�bhhK ��h��R�(KK
��h�C("   6    %  �  �   D   5         �t�bhhK ��h��R�(KK��h�C@         .   M        �  <           �  3        �t�bhhK ��h��R�(KK��h�C,      ;      �   �      �  R         �t�bhhK ��h��R�(KK��h�C       )   \  �   c	        �t�bhhK ��h��R�(KK��h�C4#   !   ?      
   3   6   �        �         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CX�  �         .                                                      �t�bhhK ��h��R�(KK��h�C�   �     �t�bhhK ��h��R�(KK��h�C0�   l  w     7   T   D   �  #  7         �t�bhhK ��h��R�(KK��h�C,d   l    /  -      .   �   �        �t�bhhK ��h��R�(KK��h�C8        �   O      �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C      0          �t�bhhK ��h��R�(KK��h�CL      J   �  ,            1   #   
   3   6   �        �         �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C|                  �        �  a	  �   h     L   >   %   �  �     a	     0   �   
      S   �        �t�bhhK ��h��R�(KK��h�C,�  &   �   �     t      �           �t�bhhK ��h��R�(KK��h�Cp      �   :      S   Y      Q            f   �   ,  %                     A   Y      ?        �t�bhhK ��h��R�(KK��h�C<      (   #     i   #              $            �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�CD9        �  7         s         @   �
  �              �t�bhhK ��h��R�(KK	��h�C$�     ^        �   �         �t�bhhK ��h��R�(KK��h�C`N  �           �        �     ,   	      	      	   K   	   �   	   �   	   )     �t�bhhK ��h��R�(KK��h�C   �  �     �t�bhhK ��h��R�(KK��h�C48        �      
  X  �	  	      	         �t�bhhK ��h��R�(KK��h�CD   /         9     7         W     $   8     �   �     �t�bhhK ��h��R�(KK��h�C �     �  �      (	  r      �t�bhhK ��h��R�(KK��h�CH]   P        
   c  �            �  �  k  "     �        �t�bhhK ��h��R�(KK��h�CC  �  k             �t�bhhK ��h��R�(KK(��h�C�      J   =      o  �                  �
           �  �     ,         �      �            8  M        �  �  �   
   �  �        �t�bhhK ��h��R�(KK��h�C�	        �     �t�bhhK ��h��R�(KK��h�C0%   l  g      �  �      �     �        �t�bhhK ��h��R�(KK��h�C0�      �            �  +      S         �t�bhhK ��h��R�(KK��h�C�  	      	         �t�bhhK ��h��R�(KK��h�C   �                  �t�bhhK ��h��R�(KK��h�CH�      -   J     A   u      5   !  �            -  �        �t�bhhK ��h��R�(KK
��h�C(!      �         	      	         �t�bhhK ��h��R�(KK
��h�C(�   &   8   /   a      o  ~        �t�bhhK ��h��R�(KK��h�C8      �	  A  W  �          A     �        �t�bhhK ��h��R�(KK��h�C@b   $   �         �   �         ,   �   
   $   �        �t�bhhK ��h��R�(KK��h�C      a     �t�bhhK ��h��R�(KK	��h�C$"         �     �  z         �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C@�    �   �      
   $                    \        �t�bhhK ��h��R�(KK
��h�C(I   ?           �              �t�bhhK ��h��R�(KK��h�C�        �   ~        �t�bhhK ��h��R�(KK��h�CD#   !         i     �   n   (      
   P     G            �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C4   �   �      w            \              �t�bhhK ��h��R�(KK��h�C-   @   (              �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C<"   �   ,   9  M  �      ,      �     u   u         �t�bhhK ��h��R�(KK	��h�C$�  �      �     9  j   �     �t�bhhK ��h��R�(KK��h�C        �         �t�bhhK ��h��R�(KK��h�C    �      �              �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C@�      #  I           V           �     �        �t�bhhK ��h��R�(KK	��h�C$�   0  �   �  �               �t�bhhK ��h��R�(KK	��h�C$V     �  �  &   N            �t�bhhK ��h��R�(KK��h�C    �   )   �      u         �t�bhhK ��h��R�(KK��h�C,a  �  �  h      �  :   $            �t�bhhK ��h��R�(KK��h�CD�   �        E      +                �   
   y        �t�bhhK ��h��R�(KK��h�C  g   �     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK
��h�C(f      �     a     
   �
        �t�bhhK ��h��R�(KK��h�Cd         .      1
  L   G      �     �        �  �           
   �     L         �t�bhhK ��h��R�(KK��h�C<�        �           �     �                �t�bhhK ��h��R�(KK	��h�C$�      ,   �   
   4  	         �t�bhhK ��h��R�(KK	��h�C$p  L  
   t      �           �t�bhhK ��h��R�(KK(��h�C�)            �  ~           $   �     u  �        .         Z  �     u  �        R     4         8   L     4      a  c         �t�bhhK ��h��R�(KK��h�Cd   .   &   �  V   2   �                    �   k	  G   Q     y      �     �
        �t�bhhK ��h��R�(KK��h�CX         .         %  �        F     �  L         �   �              �t�bhhK ��h��R�(KK��h�CHD      0   �   W    �     �     #      �   ,              �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�CE           �t�bhhK ��h��R�(KK��h�Cy     �t�bhhK ��h��R�(KK��h�C�  �	         �t�bhhK ��h��R�(KK��h�C/  ^            �t�bhhK ��h��R�(KK��h�CH�  (   �        .   
   _           }     d     �        �t�bhhK ��h��R�(KK��h�C    '   B   %              �t�bhhK ��h��R�(KK��h�C8]        �             h      f  y        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C4      P   !      l                       �t�bhhK ��h��R�(KK��h�C8     6  I                   c            �t�bhhK ��h��R�(KK��h�C<9        �  :  D         �   ,      �  �        �t�bhhK ��h��R�(KK��h�CH     G  9            �   7           �                 �t�bhhK ��h��R�(KK#��h�C�      N      �     �                �           �        �           �
     �      "   k  �     %   6        �t�bhhK ��h��R�(KK��h�C      x  B            �t�bhhK ��h��R�(KK
��h�C(�     �   .  "   %   �  K        �t�bhhK ��h��R�(KK��h�C4         /   ;      �  �     �  }        �t�bhhK ��h��R�(KK��h�CP"   m      $   �  �   &           �   U   $   �   N     �          �t�bhhK ��h��R�(KK��h�CT   8   Q            &      K        �            g     $   �	        �t�bhhK ��h��R�(KK��h�C �   ?            +        �t�bhhK ��h��R�(KK��h�Cd      /            �              ,   	      	   K   	     	   �  	   �  	         �t�bhhK ��h��R�(KK��h�C@         �t�bhhK ��h��R�(KK��h�CL*      J   �     o   &      d  S  
               �            �t�bhhK ��h��R�(KK��h�CL         �           �        H    �                    �t�bhhK ��h��R�(KK
��h�C(`                              �t�bhhK ��h��R�(KK��h�C�            �t�bhhK ��h��R�(KK��h�C@)        8   /      �     8   E     D   �           �t�bhhK ��h��R�(KK
��h�C(1   #      �  
   3   6            �t�bhhK ��h��R�(KK��h�C      *  <         �t�bhhK ��h��R�(KK��h�CD   �
     �  �   &   �  �  �	           I               �t�bhhK ��h��R�(KK	��h�C$      -   N   $   �  �        �t�bhhK ��h��R�(KK��h�C\               
  �	        `            %                     �	        �t�bhhK ��h��R�(KK��h�C@�                             q   �              �t�bhhK ��h��R�(KK	��h�C$W  �     	  )               �t�bhhK ��h��R�(KK%��h�C��      v                  �  �     �           �  �   �        �  (   2   ;      �  �   �                     �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CK            �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C0E     )   U   e   �                     �t�bhhK ��h��R�(KK��h�C4�      e   (   )   <            e   �        �t�bhhK ��h��R�(KK��h�C      '               �t�bhhK ��h��R�(KK��h�CL*               �      �  :   c  �           �   ~  �         �t�bhhK ��h��R�(KK��h�C4f      �        )   %  +      
           �t�bhhK ��h��R�(KK��h�CH     �  1     x         �   �  �                       �t�bhhK ��h��R�(KK��h�C`         �              O        �   �        �  
      :                  �t�bhhK ��h��R�(KK��h�C0Z     )         o           >        �t�bhhK ��h��R�(KK	��h�C$   �  -      .               �t�bhhK ��h��R�(KK
��h�C(H  [        (   4               �t�bhhK ��h��R�(KK��h�C|         $   �              �              �           �        <   "               G   �        �t�bhhK ��h��R�(KK��h�CxF     -            �        .   s                                   �   %         �           �t�bhhK ��h��R�(KK��h�C1   #       �      �     �t�bhhK ��h��R�(KK��h�CL      H      	      	   K   	   �   	   I  	   U  	   /  	   s     �t�bhhK ��h��R�(KK��h�CG     �t�bhhK ��h��R�(KK��h�C,1           	   K   	     	   �      �t�bhhK ��h��R�(KK��h�C8
      �  ?      #   !      _     -  5        �t�bhhK ��h��R�(KK��h�C0v          .                        �t�bhhK ��h��R�(KK��h�CB        8   �	        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C<�     �  4   =     �   �        
   �  �        �t�bhhK ��h��R�(KK
��h�C(�  [     �    �              �t�bhhK ��h��R�(KK
��h�C(t   �  `   3        ,           �t�bhhK ��h��R�(KK��h�C,D      �   3  �   *   �   _  C         �t�bhhK ��h��R�(KK	��h�C$l     7   T   D   �  �  7      �t�bhhK ��h��R�(KK	��h�C$�     �      m     >	        �t�bhhK ��h��R�(KK��h�C<   �  t	           %   H   u        �   (         �t�bhhK ��h��R�(KK��h�C   �  �         �t�bhhK ��h��R�(KK��h�C,   5      �      `   8              �t�bhhK ��h��R�(KK��h�C,   �   �  *      �  �   $   �        �t�bhhK ��h��R�(KK��h�C8   '         
      i        :   �   E        �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C  N     �t�bhhK ��h��R�(KK��h�C0        Z     L        .   N          �t�bhhK ��h��R�(KK��h�C0>     �     %   �   �                �t�bhhK ��h��R�(KK��h�C0�        �	           �               �t�bhhK ��h��R�(KK��h�CF     	      	         �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C|�     �  
   >        .            �           �                 �  �                           �t�bhhK ��h��R�(KK
��h�C(�     4	  �  �     �  P        �t�bhhK ��h��R�(KK	��h�C$2     �
     8   �   ~  �     �t�bhhK ��h��R�(KK	��h�C$T                           �t�bhhK ��h��R�(KK��h�CD!      |      <  R   ?      
   3   6   �     �   f        �t�bhhK ��h��R�(KK	��h�C$�  1  '   
   e   �   F         �t�bhhK ��h��R�(KK��h�CP      
   _      �     \        �         0   �                 �t�bhhK ��h��R�(KK��h�C0                  �  �              �t�bhhK ��h��R�(KK��h�C0*         |  �	        �  �  C         �t�bhhK ��h��R�(KK��h�C,*           t   &      M      +      �t�bhhK ��h��R�(KK��h�C4      	  2   �
  3  i      H   A   ?        �t�bhhK ��h��R�(KK��h�C             �t�bhhK ��h��R�(KK��h�C                �t�bhhK ��h��R�(KK	��h�C$�              �  M        �t�bhhK ��h��R�(KK��h�CD
   H               $   G            x     �	        �t�bhhK ��h��R�(KK	��h�C$         �      �     �     �t�bhhK ��h��R�(KK��h�C8#   !      P  (      
   u          F         �t�bhhK ��h��R�(KK
��h�C(   =      �  )  	      	         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CP!     ~   �                  �    7      ;      �             �t�bhhK ��h��R�(KK��h�C �        	      	         �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C�                   �t�bhhK ��h��R�(KK��h�C8
         2      
         �     
            �t�bhhK ��h��R�(KK��h�CX      P      �   �        C  E   y              J  E      A   F        �t�bhhK ��h��R�(KK��h�C4"   >                      �  3        �t�bhhK ��h��R�(KK��h�C0      @  �     I   `   b     6
        �t�bhhK ��h��R�(KK��h�C4   R      �     l         k               �t�bhhK ��h��R�(KK��h�C   �      i     �     �t�bhhK ��h��R�(KK��h�C   �            �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C81   #      Y           )  �  
      F         �t�bhhK ��h��R�(KK��h�CP"           D     �      l   �     7            q              �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C<!      q      	   K   	   �   	   I  	   /  	   s     �t�bhhK ��h��R�(KK��h�C3        .   �        �t�bhhK ��h��R�(KK��h�CL   (         .   
           �      =  �
  
   X   �   F         �t�bhhK ��h��R�(KK��h�Cl   �      �  )   �                       b                  �   P  �     �        �t�bhhK ��h��R�(KK��h�C�      *            �t�bhhK ��h��R�(KK
��h�C(   &   P         �  E            �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CH   �   �   	  �   �  �        z        �	     �            �t�bhhK ��h��R�(KK��h�C    B      �  
   c        �t�bhhK ��h��R�(KK��h�C<#   !           �     u   (         �            �t�bhhK ��h��R�(KK��h�C4         �      
         H   A   }         �t�bhhK ��h��R�(KK��h�C04      �   R  A     s   7      �        �t�bhhK ��h��R�(KK��h�CH      �  �  +      �        3     +      �   `            �t�bhhK ��h��R�(KK��h�C�  �      �t�bhhK ��h��R�(KK��h�C82      �  n  �   �           W	              �t�bhhK ��h��R�(KK��h�C�     �  m      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C   �   �     s  r      �t�bhhK ��h��R�(KK��h�C%        	         �t�bhhK ��h��R�(KK��h�CPC        �  9   �  "         g   d   t  G   |          <        �t�bhhK ��h��R�(KK��h�C 1   #       �              �t�bhhK ��h��R�(KK��h�CPE     �  �   A   !     P   <      x      �   �  �  G   �  �        �t�bhhK ��h��R�(KK��h�CH*        H  C  H             0   4   
   �   �   _         �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�CXB  �           8   S                       c   b  :      
            �t�bhhK ��h��R�(KK��h�Cd      �     ~       F  8   �  �         W  t      �        2     �           �t�bhhK ��h��R�(KK��h�CtT      �      �  &      �         �      �     W     h  Z  �     �      J     �               �t�bhhK ��h��R�(KK	��h�C$#   !   (      ^   �            �t�bhhK ��h��R�(KK��h�C,w  l     E     �        �        �t�bhhK ��h��R�(KK��h�C*           �t�bhhK ��h��R�(KK��h�C!      �           �t�bhhK ��h��R�(KK��h�Cd         (   <      $      &      M   �      Y	  �              Z	                 �t�bhhK ��h��R�(KK��h�CD               �  �     9   �  T      ~      �         �t�bhhK ��h��R�(KK��h�CT*   2          �  2   �              :   %  �        �	           �t�bhhK ��h��R�(KK��h�C@%         c        j   C    m  ^   �     �        �t�bhhK ��h��R�(KK��h�C@  T  
   t         �t�bhhK ��h��R�(KK��h�CL   ?   !      x       �        
   3   6   x       �        �t�bhhK ��h��R�(KK
��h�C(�   �   )   �            �         �t�bhhK ��h��R�(KK��h�Cf   �  �           �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C<         k            ;      0   �   5           �t�bhhK ��h��R�(KK��h�C8      =      [        G   �     $   k         �t�bhhK ��h��R�(KK��h�C\           d   �      �     *   D         A   �  &      �  ]               �t�bhhK ��h��R�(KK��h�C,         �t�bhhK ��h��R�(KK��h�C8V                 �     $  �              �t�bhhK ��h��R�(KK��h�C8#   !        ?      
   3   6         8        �t�bhhK ��h��R�(KK
��h�C(X  O  �        	      	         �t�bhhK ��h��R�(KK��h�CT      �   �     C      =            T   �   �      �  i   A   =        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C<      �  )	  h   �   &      U   �     $   k         �t�bhhK ��h��R�(KK
��h�C(   �     �	           $   �      �t�bhhK ��h��R�(KK��h�C�         �       �t�bhhK ��h��R�(KK	��h�C$�  �     �   �     @         �t�bhhK ��h��R�(KK��h�C0                 f                  �t�bhhK ��h��R�(KK��h�C�  E      �   �        �t�bhhK ��h��R�(KK
��h�C(*  �     n                    �t�bhhK ��h��R�(KK��h�C,
   �	  F   ?      !      B   �        �t�bhhK ��h��R�(KK��h�C0�     B           �  �     :        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C8   �  u         �     �            �        �t�bhhK ��h��R�(KK��h�C8   ?         }      �            
   T        �t�bhhK ��h��R�(KK��h�CP      �   �   E      �      �     $   �      $   /	  �   �  k         �t�bhhK ��h��R�(KK��h�C1   #          �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C�
     A         �t�bhhK ��h��R�(KK��h�C\   �   �   r      �t�bhhK ��h��R�(KK��h�C@�     R     e	          �        H   !  �         �t�bhhK ��h��R�(KK��h�C8   &   \    h   �   �   g      a   �  E         �t�bhhK ��h��R�(KK��h�C8=  �     J         )   �  `   �     �        �t�bhhK ��h��R�(KK��h�C8�   &      a   k               �  �   n        �t�bhhK ��h��R�(KK#��h�C�            O      �      6              Q     Q         x     J   �     o            5         4      �         �t�bhhK ��h��R�(KK��h�C4      &   �  �        5                  �t�bhhK ��h��R�(KK��h�C  ^     ^  k     �t�bhhK ��h��R�(KK��h�C1   #       /   "   �      �t�bhhK ��h��R�(KK��h�CT   (   #   !            l  �  "   t      �     8   �   Q               �t�bhhK ��h��R�(KK��h�CD�        i  �  �   �         �   0        $   �         �t�bhhK ��h��R�(KK��h�C�     0      �  r      �t�bhhK ��h��R�(KK��h�C!      �           �t�bhhK ��h��R�(KK
��h�C(.  M     `  
   j             �t�bhhK ��h��R�(KK��h�C      ~        �t�bhhK ��h��R�(KK��h�Cx            ]        $   n   �         .   "              H        �     U   T   �  8   �        �t�bhhK ��h��R�(KK��h�C@'        1     �  
   3   6         b      x         �t�bhhK ��h��R�(KK!��h�C�      N  4  �   :         s   7         .   
   _      {      �            =   G   H        8   4      �        �t�bhhK ��h��R�(KK��h�C0]   >      �  �   �           �        �t�bhhK ��h��R�(KK��h�C/  ^            �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C\g   O     �          g              �  
   A   F                       �t�bhhK ��h��R�(KK��h�CZ      �            �t�be.