��      ]�(�numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i4�����R�(K�<�NNNJ����J����K t�b�C[         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK
��h�C(#         t   �  �  �  �        �t�bhhK ��h��R�(KK��h�C,#         �  �     �  �   �        �t�bhhK ��h��R�(KK��h�C �  �   �  H   )   �        �t�bhhK ��h��R�(KK��h�C4   #   I           �  �  �  �  �        �t�bhhK ��h��R�(KK��h�C �     U   �     Z        �t�bhhK ��h��R�(KK��h�C,&   �  J  �     �  �     �        �t�bhhK ��h��R�(KK��h�C,:   �     �     U   �     Z        �t�bhhK ��h��R�(KK��h�C0#         �     [      �     �        �t�bhhK ��h��R�(KK��h�C@#   �  �      �  �              �   �  �  �        �t�bhhK ��h��R�(KK��h�C,�     �     #      &   ~  �        �t�bhhK ��h��R�(KK��h�C@   #      &   �  �     �     �     �  .  K        �t�bhhK ��h��R�(KK��h�C #      -      �  �        �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C8  ?   �  �  .   �  	   �     �     #         �t�bhhK ��h��R�(KK��h�C,�  "   �     �  �     �          �t�bhhK ��h��R�(KK��h�CH&   "   �  �     �  �     �   e   �  �     �     �        �t�bhhK ��h��R�(KK��h�CT�  �  �     �  �  �     �  	   �  	   L     �  u   -   �  �        �t�bhhK ��h��R�(KK��h�CP�     �  	      �   [  K     �    	   �       �     Z        �t�bhhK ��h��R�(KK��h�Ch&   �  �  �  �  �  �  �  �  �     �     �  &   �  �     �     �  �              �t�bhhK ��h��R�(KK��h�C<�  �  u   �      �  �     �  a   �     �        �t�bhhK ��h��R�(KK��h�C8�  5  �  �   #      K        �     �        �t�bhhK ��h��R�(KK��h�C0�  �  �   e      �  	   �     �        �t�bhhK ��h��R�(KK��h�CP�  �  B   x           �  	     #      �     4   �            �t�bhhK ��h��R�(KK��h�C`I       �     	     �          	   �  M  N  &            	  �        �t�bhhK ��h��R�(KK��h�CX#   �   s     
        �          Z  M  N    �     �             �t�bhhK ��h��R�(KK��h�CPH       �            &   	   O                          �t�bhhK ��h��R�(KK	��h�C$#     u   ?     �   P        �t�bhhK ��h��R�(KK��h�Cd&     Q  �                 Z  	   5           �       M  N          �t�bhhK ��h��R�(KK��h�C4#   �      K    �  M  N               �t�bhhK ��h��R�(KK��h�C�                   �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C#   "   R          �t�bhhK ��h��R�(KK	��h�C$M   #      !  �     r        �t�bhhK ��h��R�(KK��h�C"        H   I        �t�bhhK ��h��R�(KK��h�C,#     �     9        �   �        �t�bhhK ��h��R�(KK��h�C8        �     x  �  $  %  U   #   I        �t�bhhK ��h��R�(KK��h�CH&    -   '   '  	   �  	   (     )  �     &   *  	        �t�bhhK ��h��R�(KK��h�C,#   "   +         �  ,     -        �t�bhhK ��h��R�(KK��h�C,.  /  :   >   0     �      \        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C1     
           �t�bhhK ��h��R�(KK��h�C2           �t�bhhK ��h��R�(KK��h�C3        �t�bhhK ��h��R�(KK��h�C 4                 E      �t�bhhK ��h��R�(KK��h�C5                 �t�bhhK ��h��R�(KK��h�C,�  U   #      �  6                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK	��h�C$   #      ^   >     S        �t�bhhK ��h��R�(KK��h�CH   q   �  �     7     1            
     S  6          �t�bhhK ��h��R�(KK��h�CD&   �      �   �  "   �   �  �        �  �     #         �t�bhhK ��h��R�(KK	��h�C$         #   �   �  2         �t�bhhK ��h��R�(KK��h�C    #         �  �        �t�bhhK ��h��R�(KK��h�CD      
   &   �   8  +     #         �  �   �  2         �t�bhhK ��h��R�(KK
��h�C(         T     �     1         �t�bhhK ��h��R�(KK��h�CU  �   �        �t�bhhK ��h��R�(KK��h�C #   �   �                 �t�bhhK ��h��R�(KK��h�C9  �   �        �t�bhhK ��h��R�(KK��h�C �  �   :           E      �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C0&   ;    <     #      =     �        �t�bhhK ��h��R�(KK��h�C0>     �  ?  �     �  �  �  I         �t�bhhK ��h��R�(KK��h�C0   H   2         
   �     �  �        �t�bhhK ��h��R�(KK��h�C,     �  H       �   �  @        �t�bhhK ��h��R�(KK��h�C8   
   >   �      �      �        H   2         �t�bhhK ��h��R�(KK��h�CPt  |   "   6  A  �       �   �   B     ]     �      V  �  +        �t�bhhK ��h��R�(KK��h�C@   #      C  	   D     E  \   '   f      F  G        �t�bhhK ��h��R�(KK��h�C0         �   H  	        I     1      �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK
��h�C(#         t   �  �  �  �        �t�bhhK ��h��R�(KK��h�C,#         �  �     �  �   �        �t�bhhK ��h��R�(KK��h�C �  �   �  H   )   �        �t�bhhK ��h��R�(KK��h�C4   #   I           �  �  �  �  �        �t�bhhK ��h��R�(KK��h�C �     U   �     Z        �t�bhhK ��h��R�(KK��h�C,&   �  J  �     �  �     �        �t�bhhK ��h��R�(KK��h�C,:   �     �     U   �     Z        �t�bhhK ��h��R�(KK��h�C0#         �     [      �     �        �t�bhhK ��h��R�(KK��h�C@#   �  �      �  �              �   �  �  �        �t�bhhK ��h��R�(KK��h�C,�     �     #      &   ~  �        �t�bhhK ��h��R�(KK��h�C@   #      &   �  �     �     �     �  .  K        �t�bhhK ��h��R�(KK��h�C #      -      �  �        �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C8  ?   �  �  .   �  	   �     �     #         �t�bhhK ��h��R�(KK��h�C,�  "   �     �  �     �          �t�bhhK ��h��R�(KK��h�CH&   "   �  �     �  �     �   e   �  �     �     �        �t�bhhK ��h��R�(KK��h�CT�  �  �     �  �  �     �  	   �  	   L     �  u   -   �  �        �t�bhhK ��h��R�(KK��h�CP�     �  	      �   [  K     �    	   �       �     Z        �t�bhhK ��h��R�(KK��h�Ch&   �  �  �  �  �  �  �  �  �     �     �  &   �  �     �     �  �              �t�bhhK ��h��R�(KK��h�C<�  �  u   �      �  �     �  a   �     �        �t�bhhK ��h��R�(KK��h�C8�  5  �  �   #      K        �     �        �t�bhhK ��h��R�(KK��h�C0�  �  �   e      �  	   �     �        �t�bhhK ��h��R�(KK��h�CP�  �  B   x           �  	     #      �     4   �            �t�bhhK ��h��R�(KK��h�C`I       �     	     �          	   �  M  N  &            	  �        �t�bhhK ��h��R�(KK��h�CX#   �   s     
        �          Z  M  N    �     �             �t�bhhK ��h��R�(KK��h�CPH       �            &   	   O                          �t�bhhK ��h��R�(KK	��h�C$#     u   ?     �   P        �t�bhhK ��h��R�(KK��h�Cd&     Q  �                 Z  	   5           �       M  N          �t�bhhK ��h��R�(KK��h�C4#   �      K    �  M  N               �t�bhhK ��h��R�(KK��h�C�                   �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C#   "   R          �t�bhhK ��h��R�(KK	��h�C$M   #      !  �     r        �t�bhhK ��h��R�(KK��h�C"        H   I        �t�bhhK ��h��R�(KK��h�C,#     �     9        �   �        �t�bhhK ��h��R�(KK��h�C8        �     x  �  $  %  U   #   I        �t�bhhK ��h��R�(KK��h�CH&    -   '   '  	   �  	   (     )  �     &   *  	        �t�bhhK ��h��R�(KK��h�C,#   "   +         �  ,     -        �t�bhhK ��h��R�(KK��h�C,.  /  :   >   0     �      \        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C1     
           �t�bhhK ��h��R�(KK��h�C2           �t�bhhK ��h��R�(KK��h�C3        �t�bhhK ��h��R�(KK��h�C 4                 E      �t�bhhK ��h��R�(KK��h�C5                 �t�bhhK ��h��R�(KK��h�C,�  U   #      �  6                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK	��h�C$   #      ^   >     S        �t�bhhK ��h��R�(KK��h�CH   q   �  �     7     1            
     S  6          �t�bhhK ��h��R�(KK��h�CD&   �      �   �  "   �   �  �        �  �     #         �t�bhhK ��h��R�(KK	��h�C$         #   �   �  2         �t�bhhK ��h��R�(KK��h�C    #         �  �        �t�bhhK ��h��R�(KK��h�CD      
   &   �   8  +     #         �  �   �  2         �t�bhhK ��h��R�(KK
��h�C(         T     �     1         �t�bhhK ��h��R�(KK��h�CU  �   �        �t�bhhK ��h��R�(KK��h�C #   �   �                 �t�bhhK ��h��R�(KK��h�C9  �   �        �t�bhhK ��h��R�(KK��h�C �  �   :           E      �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C0&   ;    <     #      =     �        �t�bhhK ��h��R�(KK��h�C0>     �  ?  �     �  �  �  I         �t�bhhK ��h��R�(KK��h�C0   H   2         
   �     �  �        �t�bhhK ��h��R�(KK��h�C,     �  H       �   �  @        �t�bhhK ��h��R�(KK��h�C8   
   >   �      �      �        H   2         �t�bhhK ��h��R�(KK��h�CPt  |   "   6  A  �       �   �   B     ]     �      V  �  +        �t�bhhK ��h��R�(KK��h�C@   #      C  	   D     E  \   '   f      F  G        �t�bhhK ��h��R�(KK��h�C0         �   H  	        I     1      �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C[         �t�bhhK ��h��R�(KK
��h�C(#         t   �  �  �  �        �t�bhhK ��h��R�(KK��h�C,#         �  �     �  �   �        �t�bhhK ��h��R�(KK��h�C �  �   �  H   )   �        �t�bhhK ��h��R�(KK��h�C4   #   I           �  �  �  �  �        �t�bhhK ��h��R�(KK��h�C �     U   �     Z        �t�bhhK ��h��R�(KK��h�C,&   �  J  �     �  �     �        �t�bhhK ��h��R�(KK��h�C,:   �     �     U   �     Z        �t�bhhK ��h��R�(KK��h�C0#         �     [      �     �        �t�bhhK ��h��R�(KK��h�C@#   �  �      �  �              �   �  �  �        �t�bhhK ��h��R�(KK��h�C,�     �     #      &   ~  �        �t�bhhK ��h��R�(KK��h�C@   #      &   �  �     �     �     �  .  K        �t�bhhK ��h��R�(KK��h�C #      -      �  �        �t�bhhK ��h��R�(KK��h�C    
   �                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C8  ?   �  �  .   �  	   �     �     #         �t�bhhK ��h��R�(KK��h�C,�  "   �     �  �     �          �t�bhhK ��h��R�(KK��h�CH&   "   �  �     �  �     �   e   �  �     �     �        �t�bhhK ��h��R�(KK��h�CT�  �  �     �  �  �     �  	   �  	   L     �  u   -   �  �        �t�bhhK ��h��R�(KK��h�CP�     �  	      �   [  K     �    	   �       �     Z        �t�bhhK ��h��R�(KK��h�Ch&   �  �  �  �  �  �  �  �  �     �     �  &   �  �     �     �  �              �t�bhhK ��h��R�(KK��h�C<�  �  u   �      �  �     �  a   �     �        �t�bhhK ��h��R�(KK��h�C8�  5  �  �   #      K        �     �        �t�bhhK ��h��R�(KK��h�C0�  �  �   e      �  	   �     �        �t�bhhK ��h��R�(KK��h�CP�  �  B   x           �  	     #      �     4   �            �t�bhhK ��h��R�(KK��h�C`I       �     	     �          	   �  M  N  &            	  �        �t�bhhK ��h��R�(KK��h�CX#   �   s     
        �          Z  M  N    �     �             �t�bhhK ��h��R�(KK��h�CPH       �            &   	   O                          �t�bhhK ��h��R�(KK	��h�C$#     u   ?     �   P        �t�bhhK ��h��R�(KK��h�Cd&     Q  �                 Z  	   5           �       M  N          �t�bhhK ��h��R�(KK��h�C4#   �      K    �  M  N               �t�bhhK ��h��R�(KK��h�C�                   �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C#   "   R          �t�bhhK ��h��R�(KK	��h�C$M   #      !  �     r        �t�bhhK ��h��R�(KK��h�C"        H   I        �t�bhhK ��h��R�(KK��h�C,#     �     9        �   �        �t�bhhK ��h��R�(KK��h�C8        �     x  �  $  %  U   #   I        �t�bhhK ��h��R�(KK��h�CH&    -   '   '  	   �  	   (     )  �     &   *  	        �t�bhhK ��h��R�(KK��h�C,#   "   +         �  ,     -        �t�bhhK ��h��R�(KK��h�C,.  /  :   >   0     �      \        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C1     
           �t�bhhK ��h��R�(KK��h�C2           �t�bhhK ��h��R�(KK��h�C3        �t�bhhK ��h��R�(KK��h�C 4                 E      �t�bhhK ��h��R�(KK��h�C5                 �t�bhhK ��h��R�(KK��h�C,�  U   #      �  6                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK	��h�C$   #      ^   >     S        �t�bhhK ��h��R�(KK��h�CH   q   �  �     7     1            
     S  6          �t�bhhK ��h��R�(KK��h�CD&   �      �   �  "   �   �  �        �  �     #         �t�bhhK ��h��R�(KK	��h�C$         #   �   �  2         �t�bhhK ��h��R�(KK��h�C    #         �  �        �t�bhhK ��h��R�(KK��h�CD      
   &   �   8  +     #         �  �   �  2         �t�bhhK ��h��R�(KK
��h�C(         T     �     1         �t�bhhK ��h��R�(KK��h�CU  �   �        �t�bhhK ��h��R�(KK��h�C #   �   �                 �t�bhhK ��h��R�(KK��h�C9  �   �        �t�bhhK ��h��R�(KK��h�C �  �   :           E      �t�bhhK ��h��R�(KK��h�C     Y     �t�bhhK ��h��R�(KK��h�C0&   ;    <     #      =     �        �t�bhhK ��h��R�(KK��h�C0>     �  ?  �     �  �  �  I         �t�bhhK ��h��R�(KK��h�C0   H   2         
   �     �  �        �t�bhhK ��h��R�(KK��h�C,     �  H       �   �  @        �t�bhhK ��h��R�(KK��h�C8   
   >   �      �      �        H   2         �t�bhhK ��h��R�(KK��h�CPt  |   "   6  A  �       �   �   B     ]     �      V  �  +        �t�bhhK ��h��R�(KK��h�C@   #      C  	   D     E  \   '   f      F  G        �t�bhhK ��h��R�(KK��h�C0         �   H  	        I     1      �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C4�  �     4      .   k         "           �t�bhhK ��h��R�(KK��h�C  �   e   k         �t�bhhK ��h��R�(KK��h�C)      �t�bhhK ��h��R�(KK��h�C4�  �     4      .   k         "           �t�bhhK ��h��R�(KK��h�C  �   e   k         �t�bhhK ��h��R�(KK��h�C)      �t�bhhK ��h��R�(KK��h�C4�  �     4      .   k         "           �t�bhhK ��h��R�(KK��h�C  �   e   k         �t�bhhK ��h��R�(KK��h�C)      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C    �   a      �      �t�bhhK ��h��R�(KK��h�C�      7     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�     $      L      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C<#         �  J     T   �  �     K             �t�bhhK ��h��R�(KK��h�C\Y   L       �  �     
   �  ?   M  �    �   a      �   �     �          �t�bhhK ��h��R�(KK��h�C,^   �       �  �  �     �        �t�bhhK ��h��R�(KK��h�CT�      �  \   N     �  W  T   �      �     �  \   �  k      �        �t�bhhK ��h��R�(KK��h�C@   O     P        H     Q    �     �  �        �t�bhhK ��h��R�(KK#��h�C�R  �      #      �   e   S  T     �     �  	   �  U     V  	   W  #   X  	   �  Y  \   Z     #      [  #   \        �t�bhhK ��h��R�(KK��h�C4      
   ]     #         #   Q   2         �t�bhhK ��h��R�(KK��h�CL   H   2      -           ^     _     
   H   �     `        �t�bhhK ��h��R�(KK��h�C         X        �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C #   �        H   I        �t�bhhK ��h��R�(KK��h�C<a        b  	   8  	   �  \   Y  c     d        �t�bhhK ��h��R�(KK��h�C0   
     �     ;         �  2         �t�bhhK ��h��R�(KK��h�C     -              �t�bhhK ��h��R�(KK��h�Ctv      Q  e         	   f  Z  	   g  �  �  	   �  h     [       9  ?      \     �         �t�bhhK ��h��R�(KK��h�CPM  N  .   i  j     1      k     �  l         m     #         �t�bhhK ��h��R�(KK��h�C#   �  �  n     �t�bhhK ��h��R�(KK��h�Co  :  	   �   #      �t�bhhK ��h��R�(KK��h�C]      p  	   q     �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�Cr                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK	��h�C$   #      �    �  �         �t�bhhK ��h��R�(KK��h�C,�   �    �     s  t     u        �t�bhhK ��h��R�(KK
��h�C(�      .   �     ^   >   �        �t�bhhK ��h��R�(KK��h�C4�  v     �         w  x     y          �t�bhhK ��h��R�(KK��h�CT�   z  {  	     	   |  	     	     	   }     ~  \                �t�bhhK ��h��R�(KK��h�C0   �   �           
   ]  �  �        �t�bhhK ��h��R�(KK��h�CH   #      �     �  �     >   �  \   �      !  �  �         �t�bhhK ��h��R�(KK��h�C4      
        #         #   Q   2         �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�     "     �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�C    �   a      �      �t�bhhK ��h��R�(KK��h�CP    �   a      �         �     �  �     �     #  ?      �        �t�bhhK ��h��R�(KK��h�Cl   1      B      V      �  �  �     �     �     �   a      �  	      �     �  �        �t�bhhK ��h��R�(KK��h�C0.      4   �      �  �  �  �   �        �t�bhhK ��h��R�(KK��h�C4   L  �  �  	      $     �     �        �t�bhhK ��h��R�(KK��h�C-   �  �  �        �t�bhhK ��h��R�(KK"��h�C��  p   4   �       �  �     �   	   %  �     �  	   �     %  �     �  	   �  �  �   �  >     &  �  �  �        �t�bhhK ��h��R�(KK��h�C\      
   �  	   �  	   �     L     �  \   �  �     #         H   2         �t�bhhK ��h��R�(KK��h�CT�     �  	   �  	   �  	   �       '     #         (             �t�bhhK ��h��R�(KK��h�C0   (  �  -   u   P  )     �           �t�bhhK ��h��R�(KK��h�CD      �   �  ;  #   d   #   �     �  �  	   �   #         �t�bhhK ��h��R�(KK
��h�C(             �   a      �         �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C �                 E      �t�bhhK ��h��R�(KK��h�C�  ;  �           �t�bhhK ��h��R�(KK��h�C     �           �t�bhhK ��h��R�(KK��h�C�      7     �t�bhhK ��h��R�(KK��h�CX#         �     �  �  	      T   �     �  *  �     �  +     �        �t�bhhK ��h��R�(KK��h�C4#   �        .   �  �     ,  �           �t�bhhK ��h��R�(KK��h�C<      �     
   �  +     �  2         �        �t�bhhK ��h��R�(KK��h�CH   #      �  -  .  	   �  <  �  �  �     �     /        �t�bhhK ��h��R�(KK
��h�C(-  .  �     ?   0  �  �        �t�bhhK ��h��R�(KK��h�C          �      7        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C1     �t�bhhK ��h��R�(KK
��h�C(�      �     �                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C@   �     �   	      .   �  �  �  	      �  �        �t�bhhK ��h��R�(KK��h�CT#      �  �  �  2  U      �     �  �  �  �     �     �           �t�bhhK ��h��R�(KK��h�CL   �     3  �     4  ^  U   �     �  �        �  5        �t�bhhK ��h��R�(KK��h�CH-      �    �     �  
   H   �     �     �     ^        �t�bhhK ��h��R�(KK��h�CD   �  �  2            
   �  ;   	   �  \   6  +        �t�bhhK ��h��R�(KK$��h�C�7  �  �  8  .   a       �   .   �  �  �     �     �  z  ^     �     �     \   :   Z   �       :   �  �     9        �t�bhhK ��h��R�(KK��h�C8�     �     �     �  �  �  �  �  �        �t�bhhK ��h��R�(KK��h�CD   8  	   �  =  �  :  U   #   	      �  �     �        �t�bhhK ��h��R�(KK��h�C0      
   �  �      ?   ;  �  �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C �      �                 �t�bhhK ��h��R�(KK��h�C0�  3  �  �   t   3   �                 �t�bhhK ��h��R�(KK
��h�C(�  	   #   �  �                 �t�bhhK ��h��R�(KK��h�C�  �     �        �t�bhhK ��h��R�(KK
��h�C(�  �     �  )                  �t�bhhK ��h��R�(KK��h�C^  �     �t�bhhK ��h��R�(KK��h�C�     $      L      �t�bhhK ��h��R�(KK��h�C,^   �       �  �  �     �        �t�bhhK ��h��R�(KK��h�CT^   >   �   \   �  W  p   L   �      �   �     �  \   �  k      �        �t�bhhK ��h��R�(KK��h�CH$      L      �      [   s      �   	   �  	   �     �        �t�bhhK ��h��R�(KK��h�C �   T   H   <     �        �t�bhhK ��h��R�(KK��h�C,H   <  =  >  �  �   
      #         �t�bhhK ��h��R�(KK��h�Cx:   �     �  �  T   �  +     $      �  :     �     L      �  r     _  I      >   ?     #         �t�bhhK ��h��R�(KK��h�C4   
   �     $      L         H   2         �t�bhhK ��h��R�(KK��h�CXL     �  @  p   6     
   �  �  	   R  	    	  	   G   	   �     �         �t�bhhK ��h��R�(KK��h�CH�   W  T   $      L   >   �     �  	   �     �     �         �t�bhhK ��h��R�(KK��h�C,�  _  �         �     ]  	        �t�bhhK ��h��R�(KK��h�C\#   �      �   �  T   -   �     $      L   	   �  	  	   �  	   	     A        �t�bhhK ��h��R�(KK��h�C,      
   �        #   �  2         �t�bhhK ��h��R�(KK��h�C�  @     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK
��h�C(         �     $      L         �t�bhhK ��h��R�(KK��h�C�  s      �           �t�bhhK ��h��R�(KK��h�C	                 �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�CU  �   �        �t�bhhK ��h��R�(KK��h�C #   �   �                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8#   "   '   	     	  	     |         �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C    �   a      �      �t�bhhK ��h��R�(KK��h�C�      7     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�     $      L      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C<#         �  J     T   �  �     K             �t�bhhK ��h��R�(KK��h�C\Y   L       �  �     
   �  ?   M  �    �   a      �   �     �          �t�bhhK ��h��R�(KK��h�C,^   �       �  �  �     �        �t�bhhK ��h��R�(KK��h�CT�      �  \   N     �  W  T   �      �     �  \   �  k      �        �t�bhhK ��h��R�(KK��h�C@   O     P        H     Q    �     �  �        �t�bhhK ��h��R�(KK#��h�C�R  �      #      �   e   S  T     �     �  	   �  U     V  	   W  #   X  	   �  Y  \   Z     #      [  #   \        �t�bhhK ��h��R�(KK��h�C4      
   ]     #         #   Q   2         �t�bhhK ��h��R�(KK��h�CL   H   2      -           ^     _     
   H   �     `        �t�bhhK ��h��R�(KK��h�C         X        �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C #   �        H   I        �t�bhhK ��h��R�(KK��h�C<a        b  	   8  	   �  \   Y  c     d        �t�bhhK ��h��R�(KK��h�C0   
     �     ;         �  2         �t�bhhK ��h��R�(KK��h�C     -              �t�bhhK ��h��R�(KK��h�Ctv      Q  e         	   f  Z  	   g  �  �  	   �  h     [       9  ?      \     �         �t�bhhK ��h��R�(KK��h�CPM  N  .   i  j     1      k     �  l         m     #         �t�bhhK ��h��R�(KK��h�C#   �  �  n     �t�bhhK ��h��R�(KK��h�Co  :  	   �   #      �t�bhhK ��h��R�(KK��h�C]      p  	   q     �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�Cr                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK	��h�C$   #      �    �  �         �t�bhhK ��h��R�(KK��h�C,�   �    �     s  t     u        �t�bhhK ��h��R�(KK
��h�C(�      .   �     ^   >   �        �t�bhhK ��h��R�(KK��h�C4�  v     �         w  x     y          �t�bhhK ��h��R�(KK��h�CT�   z  {  	     	   |  	     	     	   }     ~  \                �t�bhhK ��h��R�(KK��h�C0   �   �           
   ]  �  �        �t�bhhK ��h��R�(KK��h�CH   #      �     �  �     >   �  \   �      !  �  �         �t�bhhK ��h��R�(KK��h�C4      
        #         #   Q   2         �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�     "     �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�C    �   a      �      �t�bhhK ��h��R�(KK��h�CP    �   a      �         �     �  �     �     #  ?      �        �t�bhhK ��h��R�(KK��h�Cl   1      B      V      �  �  �     �     �     �   a      �  	      �     �  �        �t�bhhK ��h��R�(KK��h�C0.      4   �      �  �  �  �   �        �t�bhhK ��h��R�(KK��h�C4   L  �  �  	      $     �     �        �t�bhhK ��h��R�(KK��h�C-   �  �  �        �t�bhhK ��h��R�(KK"��h�C��  p   4   �       �  �     �   	   %  �     �  	   �     %  �     �  	   �  �  �   �  >     &  �  �  �        �t�bhhK ��h��R�(KK��h�C\      
   �  	   �  	   �     L     �  \   �  �     #         H   2         �t�bhhK ��h��R�(KK��h�CT�     �  	   �  	   �  	   �       '     #         (             �t�bhhK ��h��R�(KK��h�C0   (  �  -   u   P  )     �           �t�bhhK ��h��R�(KK��h�CD      �   �  ;  #   d   #   �     �  �  	   �   #         �t�bhhK ��h��R�(KK
��h�C(             �   a      �         �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C �                 E      �t�bhhK ��h��R�(KK��h�C�  ;  �           �t�bhhK ��h��R�(KK��h�C     �           �t�bhhK ��h��R�(KK��h�C�      7     �t�bhhK ��h��R�(KK��h�CX#         �     �  �  	      T   �     �  *  �     �  +     �        �t�bhhK ��h��R�(KK��h�C4#   �        .   �  �     ,  �           �t�bhhK ��h��R�(KK��h�C<      �     
   �  +     �  2         �        �t�bhhK ��h��R�(KK��h�CH   #      �  -  .  	   �  <  �  �  �     �     /        �t�bhhK ��h��R�(KK
��h�C(-  .  �     ?   0  �  �        �t�bhhK ��h��R�(KK��h�C          �      7        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C1     �t�bhhK ��h��R�(KK
��h�C(�      �     �                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C@   �     �   	      .   �  �  �  	      �  �        �t�bhhK ��h��R�(KK��h�CT#      �  �  �  2  U      �     �  �  �  �     �     �           �t�bhhK ��h��R�(KK��h�CL   �     3  �     4  ^  U   �     �  �        �  5        �t�bhhK ��h��R�(KK��h�CH-      �    �     �  
   H   �     �     �     ^        �t�bhhK ��h��R�(KK��h�CD   �  �  2            
   �  ;   	   �  \   6  +        �t�bhhK ��h��R�(KK$��h�C�7  �  �  8  .   a       �   .   �  �  �     �     �  z  ^     �     �     \   :   Z   �       :   �  �     9        �t�bhhK ��h��R�(KK��h�C8�     �     �     �  �  �  �  �  �        �t�bhhK ��h��R�(KK��h�CD   8  	   �  =  �  :  U   #   	      �  �     �        �t�bhhK ��h��R�(KK��h�C0      
   �  �      ?   ;  �  �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C �      �                 �t�bhhK ��h��R�(KK��h�C0�  3  �  �   t   3   �                 �t�bhhK ��h��R�(KK
��h�C(�  	   #   �  �                 �t�bhhK ��h��R�(KK��h�C�  �     �        �t�bhhK ��h��R�(KK
��h�C(�  �     �  )                  �t�bhhK ��h��R�(KK��h�C^  �     �t�bhhK ��h��R�(KK��h�C�     $      L      �t�bhhK ��h��R�(KK��h�C,^   �       �  �  �     �        �t�bhhK ��h��R�(KK��h�CT^   >   �   \   �  W  p   L   �      �   �     �  \   �  k      �        �t�bhhK ��h��R�(KK��h�CH$      L      �      [   s      �   	   �  	   �     �        �t�bhhK ��h��R�(KK��h�C �   T   H   <     �        �t�bhhK ��h��R�(KK��h�C,H   <  =  >  �  �   
      #         �t�bhhK ��h��R�(KK��h�Cx:   �     �  �  T   �  +     $      �  :     �     L      �  r     _  I      >   ?     #         �t�bhhK ��h��R�(KK��h�C4   
   �     $      L         H   2         �t�bhhK ��h��R�(KK��h�CXL     �  @  p   6     
   �  �  	   R  	    	  	   G   	   �     �         �t�bhhK ��h��R�(KK��h�CH�   W  T   $      L   >   �     �  	   �     �     �         �t�bhhK ��h��R�(KK��h�C,�  _  �         �     ]  	        �t�bhhK ��h��R�(KK��h�C\#   �      �   �  T   -   �     $      L   	   �  	  	   �  	   	     A        �t�bhhK ��h��R�(KK��h�C,      
   �        #   �  2         �t�bhhK ��h��R�(KK��h�C�  @     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK
��h�C(         �     $      L         �t�bhhK ��h��R�(KK��h�C�  s      �           �t�bhhK ��h��R�(KK��h�C	                 �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�CU  �   �        �t�bhhK ��h��R�(KK��h�C #   �   �                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8#   "   '   	     	  	     |         �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C    �   a      �      �t�bhhK ��h��R�(KK��h�C�      7     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C�     $      L      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C<#         �  J     T   �  �     K             �t�bhhK ��h��R�(KK��h�C\Y   L       �  �     
   �  ?   M  �    �   a      �   �     �          �t�bhhK ��h��R�(KK��h�C,^   �       �  �  �     �        �t�bhhK ��h��R�(KK��h�CT�      �  \   N     �  W  T   �      �     �  \   �  k      �        �t�bhhK ��h��R�(KK��h�C@   O     P        H     Q    �     �  �        �t�bhhK ��h��R�(KK#��h�C�R  �      #      �   e   S  T     �     �  	   �  U     V  	   W  #   X  	   �  Y  \   Z     #      [  #   \        �t�bhhK ��h��R�(KK��h�C4      
   ]     #         #   Q   2         �t�bhhK ��h��R�(KK��h�CL   H   2      -           ^     _     
   H   �     `        �t�bhhK ��h��R�(KK��h�C         X        �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C                 �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C #   �        H   I        �t�bhhK ��h��R�(KK��h�C<a        b  	   8  	   �  \   Y  c     d        �t�bhhK ��h��R�(KK��h�C0   
     �     ;         �  2         �t�bhhK ��h��R�(KK��h�C     -              �t�bhhK ��h��R�(KK��h�Ctv      Q  e         	   f  Z  	   g  �  �  	   �  h     [       9  ?      \     �         �t�bhhK ��h��R�(KK��h�CPM  N  .   i  j     1      k     �  l         m     #         �t�bhhK ��h��R�(KK��h�C#   �  �  n     �t�bhhK ��h��R�(KK��h�Co  :  	   �   #      �t�bhhK ��h��R�(KK��h�C]      p  	   q     �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�Cr                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK	��h�C$   #      �    �  �         �t�bhhK ��h��R�(KK��h�C,�   �    �     s  t     u        �t�bhhK ��h��R�(KK
��h�C(�      .   �     ^   >   �        �t�bhhK ��h��R�(KK��h�C4�  v     �         w  x     y          �t�bhhK ��h��R�(KK��h�CT�   z  {  	     	   |  	     	     	   }     ~  \                �t�bhhK ��h��R�(KK��h�C0   �   �           
   ]  �  �        �t�bhhK ��h��R�(KK��h�CH   #      �     �  �     >   �  \   �      !  �  �         �t�bhhK ��h��R�(KK��h�C4      
        #         #   Q   2         �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C�         �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C�     "     �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�C    �   a      �      �t�bhhK ��h��R�(KK��h�CP    �   a      �         �     �  �     �     #  ?      �        �t�bhhK ��h��R�(KK��h�Cl   1      B      V      �  �  �     �     �     �   a      �  	      �     �  �        �t�bhhK ��h��R�(KK��h�C0.      4   �      �  �  �  �   �        �t�bhhK ��h��R�(KK��h�C4   L  �  �  	      $     �     �        �t�bhhK ��h��R�(KK��h�C-   �  �  �        �t�bhhK ��h��R�(KK"��h�C��  p   4   �       �  �     �   	   %  �     �  	   �     %  �     �  	   �  �  �   �  >     &  �  �  �        �t�bhhK ��h��R�(KK��h�C\      
   �  	   �  	   �     L     �  \   �  �     #         H   2         �t�bhhK ��h��R�(KK��h�CT�     �  	   �  	   �  	   �       '     #         (             �t�bhhK ��h��R�(KK��h�C0   (  �  -   u   P  )     �           �t�bhhK ��h��R�(KK��h�CD      �   �  ;  #   d   #   �     �  �  	   �   #         �t�bhhK ��h��R�(KK
��h�C(             �   a      �         �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C �                 E      �t�bhhK ��h��R�(KK��h�C�  ;  �           �t�bhhK ��h��R�(KK��h�C     �           �t�bhhK ��h��R�(KK��h�C�      7     �t�bhhK ��h��R�(KK��h�CX#         �     �  �  	      T   �     �  *  �     �  +     �        �t�bhhK ��h��R�(KK��h�C4#   �        .   �  �     ,  �           �t�bhhK ��h��R�(KK��h�C<      �     
   �  +     �  2         �        �t�bhhK ��h��R�(KK��h�CH   #      �  -  .  	   �  <  �  �  �     �     /        �t�bhhK ��h��R�(KK
��h�C(-  .  �     ?   0  �  �        �t�bhhK ��h��R�(KK��h�C          �      7        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C1     �t�bhhK ��h��R�(KK
��h�C(�      �     �                 �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C@   �     �   	      .   �  �  �  	      �  �        �t�bhhK ��h��R�(KK��h�CT#      �  �  �  2  U      �     �  �  �  �     �     �           �t�bhhK ��h��R�(KK��h�CL   �     3  �     4  ^  U   �     �  �        �  5        �t�bhhK ��h��R�(KK��h�CH-      �    �     �  
   H   �     �     �     ^        �t�bhhK ��h��R�(KK��h�CD   �  �  2            
   �  ;   	   �  \   6  +        �t�bhhK ��h��R�(KK$��h�C�7  �  �  8  .   a       �   .   �  �  �     �     �  z  ^     �     �     \   :   Z   �       :   �  �     9        �t�bhhK ��h��R�(KK��h�C8�     �     �     �  �  �  �  �  �        �t�bhhK ��h��R�(KK��h�CD   8  	   �  =  �  :  U   #   	      �  �     �        �t�bhhK ��h��R�(KK��h�C0      
   �  �      ?   ;  �  �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C �      �                 �t�bhhK ��h��R�(KK��h�C0�  3  �  �   t   3   �                 �t�bhhK ��h��R�(KK
��h�C(�  	   #   �  �                 �t�bhhK ��h��R�(KK��h�C�  �     �        �t�bhhK ��h��R�(KK
��h�C(�  �     �  )                  �t�bhhK ��h��R�(KK��h�C^  �     �t�bhhK ��h��R�(KK��h�C�     $      L      �t�bhhK ��h��R�(KK��h�C,^   �       �  �  �     �        �t�bhhK ��h��R�(KK��h�CT^   >   �   \   �  W  p   L   �      �   �     �  \   �  k      �        �t�bhhK ��h��R�(KK��h�CH$      L      �      [   s      �   	   �  	   �     �        �t�bhhK ��h��R�(KK��h�C �   T   H   <     �        �t�bhhK ��h��R�(KK��h�C,H   <  =  >  �  �   
      #         �t�bhhK ��h��R�(KK��h�Cx:   �     �  �  T   �  +     $      �  :     �     L      �  r     _  I      >   ?     #         �t�bhhK ��h��R�(KK��h�C4   
   �     $      L         H   2         �t�bhhK ��h��R�(KK��h�CXL     �  @  p   6     
   �  �  	   R  	    	  	   G   	   �     �         �t�bhhK ��h��R�(KK��h�CH�   W  T   $      L   >   �     �  	   �     �     �         �t�bhhK ��h��R�(KK��h�C,�  _  �         �     ]  	        �t�bhhK ��h��R�(KK��h�C\#   �      �   �  T   -   �     $      L   	   �  	  	   �  	   	     A        �t�bhhK ��h��R�(KK��h�C,      
   �        #   �  2         �t�bhhK ��h��R�(KK��h�C�  @     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK
��h�C(         �     $      L         �t�bhhK ��h��R�(KK��h�C�  s      �           �t�bhhK ��h��R�(KK��h�C	                 �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�CU  �   �        �t�bhhK ��h��R�(KK��h�C #   �   �                 �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C8#   "   '   	     	  	     |         �        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C,      {      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�C`     �     �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C,      &   `  a     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C0      �        �   B     �  �         �t�bhhK ��h��R�(KK
��h�C(:   	     �  /   ^     		        �t�bhhK ��h��R�(KK��h�CP   6   x  �   B     �   �  	   v   C  	   D     
	        E        �t�bhhK ��h��R�(KK��h�C,      {      �t�bhhK ��h��R�(KK��h�C<
      "   ,      �     r   {         =   �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CF  G     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C          ,      {         �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CD
      �   5   +      H        M  6      �   �   �         �t�bhhK ��h��R�(KK��h�C4�   4   �   
   .   4      �   
      M        �t�bhhK ��h��R�(KK	��h�C$      �      I             �t�bhhK ��h��R�(KK��h�C             	  2         �t�bhhK ��h��R�(KK��h�C@      -   �  �   	          �   �   &      �        �t�bhhK ��h��R�(KK��h�C#   	     �t�bhhK ��h��R�(KK��h�C�  	     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C	                 �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�CD
      �   5   +      H        M  6      �   �   �         �t�bhhK ��h��R�(KK��h�C         l         �t�bhhK ��h��R�(KK��h�C`     �     �t�bhhK ��h��R�(KK��h�Cl
      u         �  b     `  �      	  �         J  6      �  w   y  �     J   �        �t�bhhK ��h��R�(KK��h�CP
   	  4      	     J  6      =   	     �     �      �  1         �t�bhhK ��h��R�(KK��h�Cc        �t�bhhK ��h��R�(KK��h�C�     �      �  1      �t�bhhK ��h��R�(KK��h�C	  K     �t�bhhK ��h��R�(KK��h�C	  �     �t�bhhK ��h��R�(KK��h�C]      	     �t�bhhK ��h��R�(KK��h�C8
      	     `        >  
   +      	        �t�bhhK ��h��R�(KK��h�CP
      	  �     '   	  	  �         �      I          �        �t�bhhK ��h��R�(KK��h�C          `     �        �t�bhhK ��h��R�(KK��h�C 	     �      �  1         �t�bhhK ��h��R�(KK��h�C,�     �      �  �                 �t�bhhK ��h��R�(KK'��h�C�+            Y      	     	  	                 E      s     �      �      /     v     �     �      �     �     �     L     �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�ChM  ;      �  5  
      "   �      	  �  	         @   !	     N  �  �  U   �          �t�bhhK ��h��R�(KK��h�Ct   3      3        �t�bhhK ��h��R�(KK��h�C#   �     �t�bhhK ��h��R�(KK
��h�C(c     "	  	   ,  #	  	   �   #      �t�bhhK ��h��R�(KK��h�C]      O     �t�bhhK ��h��R�(KK��h�C4   
   P  Q     �   e      �   $	  2         �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�C�   %	        �t�bhhK ��h��R�(KK��h�C�   &	                 �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C4&   �      �   �  �  �  '	     �  �        �t�bhhK ��h��R�(KK��h�C4v      -   �     4      �     �  R        �t�bhhK ��h��R�(KK��h�C,:      �  N        |      �         �t�bhhK ��h��R�(KK
��h�C(            #   �   �  2         �t�bhhK ��h��R�(KK��h�Cd
      �  �  S        g   �     J   �   �   	      T  (	     U     t   3   V        �t�bhhK ��h��R�(KK��h�C0:   �      �   W     �  T   -   )	        �t�bhhK ��h��R�(KK	��h�C$-   *	  +	  T   X     ,	        �t�bhhK ��h��R�(KK��h�C         �        �t�bhhK ��h��R�(KK��h�CU  �   �        �t�bhhK ��h��R�(KK��h�C #   �   �                 �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Ct           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK��h�Ct   ,      m      �   O      +      t   3   Y     -	     #   �   �     t   3   0      K   �  �        �t�bhhK ��h��R�(KK��h�C.	     �t�bhhK ��h��R�(KK��h�C]      /	        �t�bhhK ��h��R�(KK��h�C#   �     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C�     Z     �t�bhhK ��h��R�(KK
��h�C(         ,      m      �         �t�bhhK ��h��R�(KK��h�CP   3   0	        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C<b      [     d  	      e        \  �  ?        �t�bhhK ��h��R�(KK��h�C B   �   
   b      ]        �t�bhhK ��h��R�(KK
��h�C(       f     �     ^  g        �t�bhhK ��h��R�(KK��h�C3   h  #   �     �t�bhhK ��h��R�(KK��h�C c     �  i  	   �   #      �t�bhhK ��h��R�(KK��h�C]      _     �t�bhhK ��h��R�(KK��h�C         b         �t�bhhK ��h��R�(KK��h�CH?     �  p   f      �      V  �  n   G   	   �     �        �t�bhhK ��h��R�(KK��h�C0�  p      
        T   +      �        �t�bhhK ��h��R�(KK��h�C8   ,   d   L      �   x   �  j  0     1	        �t�bhhK ��h��R�(KK	��h�C$         n      _   ,         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C`           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Ca           �t�bhhK ��h��R�(KK��h�CD      w   y  ,      ?     @     2	     �      �        �t�bhhK ��h��R�(KK��h�C4            t   3   0      K   �  2         �t�bhhK ��h��R�(KK	��h�C$�     L   �     =   �         �t�bhhK ��h��R�(KK��h�C4v      B   �  
   ,      @   +      V         �t�bhhK ��h��R�(KK��h�C4            t   3   0      K   �  2         �t�bhhK ��h��R�(KK��h�Cb  w     Z        �t�bhhK ��h��R�(KK	��h�C$         n      _   ,         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C3	           �t�bhhK ��h��R�(KK��h�C�     4	  )            �t�bhhK ��h��R�(KK��h�C,      &   `  a     �t�bhhK ��h��R�(KK��h�CL
      5   +      V      J   `  G         �      {     �         �t�bhhK ��h��R�(KK��h�Cc  |  d        �t�bhhK ��h��R�(KK��h�C,   �  e  c     5	     6	  7	        �t�bhhK ��h��R�(KK��h�C         �   G         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C8	           �t�bhhK ��h��R�(KK ��h�C�
      "   Q  ,         >  
   f   d   t   3   0      K   �  9	     :	     �  	   (   ;	     <	  	   (   f        �t�bhhK ��h��R�(KK��h�C,
      "   ,      �  	   =   =	        �t�bhhK ��h��R�(KK��h�C4      �  ,     a    >	     J   S        �t�bhhK ��h��R�(KK��h�Ct   3      3        �t�bhhK ��h��R�(KK��h�C#   �     �t�bhhK ��h��R�(KK��h�C]      O     �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C?	           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK ��h�C�
      "   ,      @	  	   A	  	   -     B	        @   o      g     C	  	   t   3   0      K   �  D	     �         �t�bhhK ��h��R�(KK��h�Cx      w   y  E	     +  �   �     F	  	         G	  /   ^     H	  	      .  =   �  I	  	   (   J	        �t�bhhK ��h��R�(KK��h�CH   K	     L	  M	     N	  O	  -      P	  	   x  g     �        �t�bhhK ��h��R�(KK��h�C4-   #   �      �   �  Q	  T   X     �         �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CR	  1     �t�bhhK ��h��R�(KK��h�C�  #      �t�bhhK ��h��R�(KK��h�C]      S	     �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�     h           �t�bhhK ��h��R�(KK��h�CU  �      �   i        �t�bhhK ��h��R�(KK��h�C,#   �      �   �  �   �   h           �t�bhhK ��h��R�(KK��h�C,      {      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�C`     �     �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C,      &   `  a     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C0      �        �   B     �  �         �t�bhhK ��h��R�(KK
��h�C(:   	     �  /   ^     		        �t�bhhK ��h��R�(KK��h�CP   6   x  �   B     �   �  	   v   C  	   D     
	        E        �t�bhhK ��h��R�(KK��h�C,      {      �t�bhhK ��h��R�(KK��h�C<
      "   ,      �     r   {         =   �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CF  G     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C          ,      {         �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CD
      �   5   +      H        M  6      �   �   �         �t�bhhK ��h��R�(KK��h�C4�   4   �   
   .   4      �   
      M        �t�bhhK ��h��R�(KK	��h�C$      �      I             �t�bhhK ��h��R�(KK��h�C             	  2         �t�bhhK ��h��R�(KK��h�C@      -   �  �   	          �   �   &      �        �t�bhhK ��h��R�(KK��h�C#   	     �t�bhhK ��h��R�(KK��h�C�  	     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C	                 �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�CD
      �   5   +      H        M  6      �   �   �         �t�bhhK ��h��R�(KK��h�C         l         �t�bhhK ��h��R�(KK��h�C`     �     �t�bhhK ��h��R�(KK��h�Cl
      u         �  b     `  �      	  �         J  6      �  w   y  �     J   �        �t�bhhK ��h��R�(KK��h�CP
   	  4      	     J  6      =   	     �     �      �  1         �t�bhhK ��h��R�(KK��h�Cc        �t�bhhK ��h��R�(KK��h�C�     �      �  1      �t�bhhK ��h��R�(KK��h�C	  K     �t�bhhK ��h��R�(KK��h�C	  �     �t�bhhK ��h��R�(KK��h�C]      	     �t�bhhK ��h��R�(KK��h�C8
      	     `        >  
   +      	        �t�bhhK ��h��R�(KK��h�CP
      	  �     '   	  	  �         �      I          �        �t�bhhK ��h��R�(KK��h�C          `     �        �t�bhhK ��h��R�(KK��h�C 	     �      �  1         �t�bhhK ��h��R�(KK��h�C,�     �      �  �                 �t�bhhK ��h��R�(KK'��h�C�+            Y      	     	  	                 E      s     �      �      /     v     �     �      �     �     �     L     �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�ChM  ;      �  5  
      "   �      	  �  	         @   !	     N  �  �  U   �          �t�bhhK ��h��R�(KK��h�Ct   3      3        �t�bhhK ��h��R�(KK��h�C#   �     �t�bhhK ��h��R�(KK
��h�C(c     "	  	   ,  #	  	   �   #      �t�bhhK ��h��R�(KK��h�C]      O     �t�bhhK ��h��R�(KK��h�C4   
   P  Q     �   e      �   $	  2         �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�C�   %	        �t�bhhK ��h��R�(KK��h�C�   &	                 �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C4&   �      �   �  �  �  '	     �  �        �t�bhhK ��h��R�(KK��h�C4v      -   �     4      �     �  R        �t�bhhK ��h��R�(KK��h�C,:      �  N        |      �         �t�bhhK ��h��R�(KK
��h�C(            #   �   �  2         �t�bhhK ��h��R�(KK��h�Cd
      �  �  S        g   �     J   �   �   	      T  (	     U     t   3   V        �t�bhhK ��h��R�(KK��h�C0:   �      �   W     �  T   -   )	        �t�bhhK ��h��R�(KK	��h�C$-   *	  +	  T   X     ,	        �t�bhhK ��h��R�(KK��h�C         �        �t�bhhK ��h��R�(KK��h�CU  �   �        �t�bhhK ��h��R�(KK��h�C #   �   �                 �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Ct           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK��h�Ct   ,      m      �   O      +      t   3   Y     -	     #   �   �     t   3   0      K   �  �        �t�bhhK ��h��R�(KK��h�C.	     �t�bhhK ��h��R�(KK��h�C]      /	        �t�bhhK ��h��R�(KK��h�C#   �     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C�     Z     �t�bhhK ��h��R�(KK
��h�C(         ,      m      �         �t�bhhK ��h��R�(KK��h�CP   3   0	        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C<b      [     d  	      e        \  �  ?        �t�bhhK ��h��R�(KK��h�C B   �   
   b      ]        �t�bhhK ��h��R�(KK
��h�C(       f     �     ^  g        �t�bhhK ��h��R�(KK��h�C3   h  #   �     �t�bhhK ��h��R�(KK��h�C c     �  i  	   �   #      �t�bhhK ��h��R�(KK��h�C]      _     �t�bhhK ��h��R�(KK��h�C         b         �t�bhhK ��h��R�(KK��h�CH?     �  p   f      �      V  �  n   G   	   �     �        �t�bhhK ��h��R�(KK��h�C0�  p      
        T   +      �        �t�bhhK ��h��R�(KK��h�C8   ,   d   L      �   x   �  j  0     1	        �t�bhhK ��h��R�(KK	��h�C$         n      _   ,         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C`           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Ca           �t�bhhK ��h��R�(KK��h�CD      w   y  ,      ?     @     2	     �      �        �t�bhhK ��h��R�(KK��h�C4            t   3   0      K   �  2         �t�bhhK ��h��R�(KK	��h�C$�     L   �     =   �         �t�bhhK ��h��R�(KK��h�C4v      B   �  
   ,      @   +      V         �t�bhhK ��h��R�(KK��h�C4            t   3   0      K   �  2         �t�bhhK ��h��R�(KK��h�Cb  w     Z        �t�bhhK ��h��R�(KK	��h�C$         n      _   ,         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C3	           �t�bhhK ��h��R�(KK��h�C�     4	  )            �t�bhhK ��h��R�(KK��h�C,      &   `  a     �t�bhhK ��h��R�(KK��h�CL
      5   +      V      J   `  G         �      {     �         �t�bhhK ��h��R�(KK��h�Cc  |  d        �t�bhhK ��h��R�(KK��h�C,   �  e  c     5	     6	  7	        �t�bhhK ��h��R�(KK��h�C         �   G         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C8	           �t�bhhK ��h��R�(KK ��h�C�
      "   Q  ,         >  
   f   d   t   3   0      K   �  9	     :	     �  	   (   ;	     <	  	   (   f        �t�bhhK ��h��R�(KK��h�C,
      "   ,      �  	   =   =	        �t�bhhK ��h��R�(KK��h�C4      �  ,     a    >	     J   S        �t�bhhK ��h��R�(KK��h�Ct   3      3        �t�bhhK ��h��R�(KK��h�C#   �     �t�bhhK ��h��R�(KK��h�C]      O     �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C?	           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK ��h�C�
      "   ,      @	  	   A	  	   -     B	        @   o      g     C	  	   t   3   0      K   �  D	     �         �t�bhhK ��h��R�(KK��h�Cx      w   y  E	     +  �   �     F	  	         G	  /   ^     H	  	      .  =   �  I	  	   (   J	        �t�bhhK ��h��R�(KK��h�CH   K	     L	  M	     N	  O	  -      P	  	   x  g     �        �t�bhhK ��h��R�(KK��h�C4-   #   �      �   �  Q	  T   X     �         �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CR	  1     �t�bhhK ��h��R�(KK��h�C�  #      �t�bhhK ��h��R�(KK��h�C]      S	     �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�     h           �t�bhhK ��h��R�(KK��h�CU  �      �   i        �t�bhhK ��h��R�(KK��h�C,#   �      �   �  �   �   h           �t�bhhK ��h��R�(KK��h�C,      {      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�C`     �     �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C,      &   `  a     �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C0      �        �   B     �  �         �t�bhhK ��h��R�(KK
��h�C(:   	     �  /   ^     		        �t�bhhK ��h��R�(KK��h�CP   6   x  �   B     �   �  	   v   C  	   D     
	        E        �t�bhhK ��h��R�(KK��h�C,      {      �t�bhhK ��h��R�(KK��h�C<
      "   ,      �     r   {         =   �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CF  G     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C          ,      {         �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�CD
      �   5   +      H        M  6      �   �   �         �t�bhhK ��h��R�(KK��h�C4�   4   �   
   .   4      �   
      M        �t�bhhK ��h��R�(KK	��h�C$      �      I             �t�bhhK ��h��R�(KK��h�C             	  2         �t�bhhK ��h��R�(KK��h�C@      -   �  �   	          �   �   &      �        �t�bhhK ��h��R�(KK��h�C#   	     �t�bhhK ��h��R�(KK��h�C�  	     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�C�                 �t�bhhK ��h��R�(KK��h�C	                 �t�bhhK ��h��R�(KK��h�Cl      �t�bhhK ��h��R�(KK��h�CD
      �   5   +      H        M  6      �   �   �         �t�bhhK ��h��R�(KK��h�C         l         �t�bhhK ��h��R�(KK��h�C`     �     �t�bhhK ��h��R�(KK��h�Cl
      u         �  b     `  �      	  �         J  6      �  w   y  �     J   �        �t�bhhK ��h��R�(KK��h�CP
   	  4      	     J  6      =   	     �     �      �  1         �t�bhhK ��h��R�(KK��h�Cc        �t�bhhK ��h��R�(KK��h�C�     �      �  1      �t�bhhK ��h��R�(KK��h�C	  K     �t�bhhK ��h��R�(KK��h�C	  �     �t�bhhK ��h��R�(KK��h�C]      	     �t�bhhK ��h��R�(KK��h�C8
      	     `        >  
   +      	        �t�bhhK ��h��R�(KK��h�CP
      	  �     '   	  	  �         �      I          �        �t�bhhK ��h��R�(KK��h�C          `     �        �t�bhhK ��h��R�(KK��h�C 	     �      �  1         �t�bhhK ��h��R�(KK��h�C,�     �      �  �                 �t�bhhK ��h��R�(KK'��h�C�+            Y      	     	  	                 E      s     �      �      /     v     �     �      �     �     �     L     �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�ChM  ;      �  5  
      "   �      	  �  	         @   !	     N  �  �  U   �          �t�bhhK ��h��R�(KK��h�Ct   3      3        �t�bhhK ��h��R�(KK��h�C#   �     �t�bhhK ��h��R�(KK
��h�C(c     "	  	   ,  #	  	   �   #      �t�bhhK ��h��R�(KK��h�C]      O     �t�bhhK ��h��R�(KK��h�C4   
   P  Q     �   e      �   $	  2         �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C5           h      �t�bhhK ��h��R�(KK��h�C�   %	        �t�bhhK ��h��R�(KK��h�C�   &	                 �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C4&   �      �   �  �  �  '	     �  �        �t�bhhK ��h��R�(KK��h�C4v      -   �     4      �     �  R        �t�bhhK ��h��R�(KK��h�C,:      �  N        |      �         �t�bhhK ��h��R�(KK
���      h�C(            #   �   �  2         �t�bhhK ��h��R�(KK��h�Cd
      �  �  S        g   �     J   �   �   	      T  (	     U     t   3   V        �t�bhhK ��h��R�(KK��h�C0:   �      �   W     �  T   -   )	        �t�bhhK ��h��R�(KK	��h�C$-   *	  +	  T   X     ,	        �t�bhhK ��h��R�(KK��h�C         �        �t�bhhK ��h��R�(KK��h�CU  �   �        �t�bhhK ��h��R�(KK��h�C #   �   �                 �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Ct           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C,      m      �      �t�bhhK ��h��R�(KK��h�Ct   ,      m      �   O      +      t   3   Y     -	     #   �   �     t   3   0      K   �  �        �t�bhhK ��h��R�(KK��h�C.	     �t�bhhK ��h��R�(KK��h�C]      /	        �t�bhhK ��h��R�(KK��h�C#   �     �t�bhhK ��h��R�(KK��h�C�   #      �t�bhhK ��h��R�(KK��h�C�     Z     �t�bhhK ��h��R�(KK
��h�C(         ,      m      �         �t�bhhK ��h��R�(KK��h�CP   3   0	        �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�Cb      �t�bhhK ��h��R�(KK��h�C<b      [     d  	      e        \  �  ?        �t�bhhK ��h��R�(KK��h�C B   �   
   b      ]        �t�bhhK ��h��R�(KK
��h�C(       f     �     ^  g        �t�bhhK ��h��R�(KK��h�C3   h  #   �     �t�bhhK ��h��R�(KK��h�C c     �  i  	   �   #      �t�bhhK ��h��R�(KK��h�C]      _     �t�bhhK ��h��R�(KK��h�C         b         �t�bhhK ��h��R�(KK��h�CH?     �  p   f      �      V  �  n   G   	   �     �        �t�bhhK ��h��R�(KK��h�C0�  p      
        T   +      �        �t�bhhK ��h��R�(KK��h�C8   ,   d   L      �   x   �  j  0     1	        �t�bhhK ��h��R�(KK	��h�C$         n      _   ,         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C`           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�Ca           �t�bhhK ��h��R�(KK��h�CD      w   y  ,      ?     @     2	     �      �        �t�bhhK ��h��R�(KK��h�C4            t   3   0      K   �  2         �t�bhhK ��h��R�(KK	��h�C$�     L   �     =   �         �t�bhhK ��h��R�(KK��h�C4v      B   �  
   ,      @   +      V         �t�bhhK ��h��R�(KK��h�C4            t   3   0      K   �  2         �t�bhhK ��h��R�(KK��h�Cb  w     Z        �t�bhhK ��h��R�(KK	��h�C$         n      _   ,         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C3	           �t�bhhK ��h��R�(KK��h�C�     4	  )            �t�bhhK ��h��R�(KK��h�C,      &   `  a     �t�bhhK ��h��R�(KK��h�CL
      5   +      V      J   `  G         �      {     �         �t�bhhK ��h��R�(KK��h�Cc  |  d        �t�bhhK ��h��R�(KK��h�C,   �  e  c     5	     6	  7	        �t�bhhK ��h��R�(KK��h�C         �   G         �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C8	           �t�bhhK ��h��R�(KK ��h�C�
      "   Q  ,         >  
   f   d   t   3   0      K   �  9	     :	     �  	   (   ;	     <	  	   (   f        �t�bhhK ��h��R�(KK��h�C,
      "   ,      �  	   =   =	        �t�bhhK ��h��R�(KK��h�C4      �  ,     a    >	     J   S        �t�bhhK ��h��R�(KK��h�Ct   3      3        �t�bhhK ��h��R�(KK��h�C#   �     �t�bhhK ��h��R�(KK��h�C]      O     �t�bhhK ��h��R�(KK��h�C P   3   0      K   R         �t�bhhK ��h��R�(KK��h�C?	           �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK ��h�C�
      "   ,      @	  	   A	  	   -     B	        @   o      g     C	  	   t   3   0      K   �  D	     �         �t�bhhK ��h��R�(KK��h�Cx      w   y  E	     +  �   �     F	  	         G	  /   ^     H	  	      .  =   �  I	  	   (   J	        �t�bhhK ��h��R�(KK��h�CH   K	     L	  M	     N	  O	  -      P	  	   x  g     �        �t�bhhK ��h��R�(KK��h�C4-   #   �      �   �  Q	  T   X     �         �t�bhhK ��h��R�(KK��h�C�      �t�be.