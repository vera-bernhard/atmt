����      ]�(�numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i4�����R�(K�<�NNNJ����J����K t�b�C8�      \   �   7   C     �                    �t�bhhK ��h��R�(KK��h�C0E  H      �                           �t�bhhK ��h��R�(KK��h�C0�  
            S                     �t�bhhK ��h��R�(KK��h�C               �t�bhhK ��h��R�(KK��h�C4�   ,   m     �      e            4        �t�bhhK ��h��R�(KK��h�CP               x      	   w   C      X        .   K   �   F         �t�bhhK ��h��R�(KK��h�C0   �  �       )                     �t�bhhK ��h��R�(KK%��h�C��         �  �   
   �  [     I   	   �	     	   �      e   .        
            	                                       �t�bhhK ��h��R�(KK��h�CX            j   D     	   �                    p     )    �         �t�bhhK ��h��R�(KK(��h�C�9         9   D   �  1         `    &        0   %      �        �              0      �     �      M     	        �           �t�bhhK ��h��R�(KK��h�C,                  d     �         �t�bhhK ��h��R�(KK
��h�C(   1      "      '              �t�bhhK ��h��R�(KK��h�C87  
   �   �  D   
      =   �  #     1         �t�bhhK ��h��R�(KK��h�CP   �      �   �        �   �  �        �     �                  �t�bhhK ��h��R�(KK��h�Ch      
   L   �   c      
   �         �	                 9      D         3            �t�bhhK ��h��R�(KK	��h�C$"                 �         �t�bhhK ��h��R�(KK��h�C �  �  �        ^        �t�bhhK ��h��R�(KK��h�C4   m  Y        s   �            "         �t�bhhK ��h��R�(KK&��h�C�'   �   (      &   ^   �         o     L                            �      �        �   #        T              �        �t�bhhK ��h��R�(KK��h�CL�         �   ,   M               ^  �  l      
              �t�bhhK ��h��R�(KK��h�C�  g  &            �t�bhhK ��h��R�(KK-��h�C�
   �        m                     <         	      I      �     	   /      �  8      �      .   �        5   �         �  �      �   ,   /   N        �t�bhhK ��h��R�(KK��h�Cxv     O           �   b   �     �     `   �         	           U  ~        	        E         �t�bhhK ��h��R�(KK
��h�C(   R      	        �            �t�bhhK ��h��R�(KK��h�Cd'   >   (   �  
   �      �  �   B   �     C      T      L   �   "            Q         �t�bhhK ��h��R�(KK)��h�C�      h   |     �                  �        �               l   S  )   \                  \           B  -   �     �           �t�bhhK ��h��R�(KK��h�C4   _   
         =         
   6   �        �t�bhhK ��h��R�(KK��h�C0            Y     K     Y  u        �t�bhhK ��h��R�(KK ��h�C�
   �             s           �     a   �     "   )  �               `        �          /         �t�bhhK ��h��R�(KK��h�Cd         �       �   %  �  -      a            +         �      =  	   D        �t�bhhK ��h��R�(KK��h�C|               
      4               
      �                �        ^  V                     �t�bhhK ��h��R�(KK��h�CX
   L   �   �      �      R     *      �      u   �   [         �   �        �t�bhhK ��h��R�(KK��h�CD   s   �   �           L   9   �   �   	     �             �t�bhhK ��h��R�(KK��h�CH*   X  a         }                 Q    �  *   &        �t�bhhK ��h��R�(KK��h�C`   Q         	   8     �           |  H      �               r   �   T        �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�CHA  �        9         �
        )   �  V
  8      c         �t�bhhK ��h��R�(KK��h�CH*  &      �   3         <     �         �  �  �   �         �t�bhhK ��h��R�(KK��h�C\         T  !         3         3      �   3   |  	   k   �   )      �        �t�bhhK ��h��R�(KK/��h�C�
   �   :      �     ;        �   Q   i   F      i   �        �      _      9      M   "           /   �         �  �  0                                    �t�bhhK ��h��R�(KK��h�C|'   >   (   g     %   �      �   �     }   �  [         	   Y  2	        �        �   �  �      f	        �t�bhhK ��h��R�(KK��h�CX            n              w   �   +   T
  	      ,      J               �t�bhhK ��h��R�(KK��h�CT�      �           �        �              �  �      b            �t�bhhK ��h��R�(KK��h�CL            �      !            j      2   �  �               �t�bhhK ��h��R�(KK
��h�C(   a  N	        J  N	           �t�bhhK ��h��R�(KK��h�C8   B   �        $      h     �               �t�bhhK ��h��R�(KK��h�Cx      E   �
           �                 c   q               �  �  	   0  8  [      2   �        �t�bhhK ��h��R�(KK��h�C0U        '  @   !                    �t�bhhK ��h��R�(KK��h�CD      `   �        �           |                    �t�bhhK ��h��R�(KK��h�CT�     ,      �     \   �     w     $               l     =         �t�bhhK ��h��R�(KK��h�CD   	      z   	         /    <   �     k              �t�bhhK ��h��R�(KK��h�C0              ;  )      �            �t�bhhK ��h��R�(KK��h�C<*   4      <                        B           �t�bhhK ��h��R�(KK	��h�C$   G   R                     �t�bhhK ��h��R�(KK��h�C0        �    $   ^    �  �         �t�bhhK ��h��R�(KK#��h�C�        �        �   /   6         �            �   k      �  �
           �     t        m     �
              �t�bhhK ��h��R�(KK	��h�C$�         m     �   (        �t�bhhK ��h��R�(KK��h�C    
   R  9   ~           �t�bhhK ��h��R�(KK/��h�C�   �         	      �  
        8   �   *         �                        l     �           �   d      E   (  	      M     ,      M                 �t�bhhK ��h��R�(KK��h�CdG   Q         �  N     �   j        �        �  &         t                    �t�bhhK ��h��R�(KK2��h�C�
               �     
   �   �
  ?   	     �   o   	      �  �     �        $   �  �           
                    2      2      �           �   ?               �t�bhhK ��h��R�(KK��h�Cx                  B         =            
   Y  #      E   	   
   D   6         E      �  �        �t�bhhK ��h��R�(KK��h�C4"   /   ?   E      �                       �t�bhhK ��h��R�(KK��h�C    �   �   ~      �        �t�bhhK ��h��R�(KK��h�C0e      �      [     	   /   �            �t�bhhK ��h��R�(KK"��h�C�      �  K      }   �           	   Q  %   �            [	        !     �   q      �  K   �            q         �t�bhhK ��h��R�(KK��h�CP   �  @   g   �	     T      T      X         9                    �t�bhhK ��h��R�(KK��h�C`!         �  -   W            0      b                  O      e      (        �t�bhhK ��h��R�(KK��h�CP   �   5   �   �   V                    �         �              �t�bhhK ��h��R�(KK��h�C<      j      �           \   �     �           �t�bhhK ��h��R�(KK��h�CX        %   Q               �                                       �t�bhhK ��h��R�(KK��h�C      J  ^   s        �t�bhhK ��h��R�(KK��h�C47     �   �  J         �  E   �  @         �t�bhhK ��h��R�(KK	��h�C$         <   A      �         �t�bhhK ��h��R�(KK��h�C8K   �   �      �   �      �   ~      }   �        �t�bhhK ��h��R�(KK��h�C`      �   �  P         =     �     U   ~     �        �   B   .   %   �        �t�bhhK ��h��R�(KK��h�C      c            �t�bhhK ��h��R�(KK��h�C8
               �      S      l     �        �t�bhhK ��h��R�(KK��h�CL   7         ~  	      6   2       	         F   _   �          �t�bhhK ��h��R�(KK��h�C .   J      S   �             �t�bhhK ��h��R�(KK��h�C   �  	               �t�bhhK ��h��R�(KK��h�Cd   &      Z   
            &         �     �      r   E            }     M        �t�bhhK ��h��R�(KK��h�C,	      0      	   �  �  �             �t�bhhK ��h��R�(KK��h�C,         �   �        �   >        �t�bhhK ��h��R�(KK��h�C,u           	   C   1   0  �         �t�bhhK ��h��R�(KK��h�C�      <      �        �t�bhhK ��h��R�(KK��h�Cd
   �        ]   �   t  ,     t  \      !      �             .   1      �        �t�bhhK ��h��R�(KK��h�C        �           �t�bhhK ��h��R�(KK
��h�C(      �            #        �t�bhhK ��h��R�(KK��h�CDy   �     k      t                          �        �t�bhhK ��h��R�(KK��h�C,   E   �   �     �  	               �t�bhhK ��h��R�(KK��h�Cp?   ~   �  H   {      $      �     P  �              U   >     �   6   �  �   �   �  ~         �t�bhhK ��h��R�(KK
��h�C(1         a     �      �        �t�bhhK ��h��R�(KK��h�CL         7           &           �     +      B   &        �t�bhhK ��h��R�(KK��h�C8   R        ,      "   j   �     8   �         �t�bhhK ��h��R�(KK��h�Ct   �  �         �                 *   �  #      �        G  	   *   �      �   0               �t�bhhK ��h��R�(KK
��h�C(\        J   2      2   J         �t�bhhK ��h��R�(KK��h�C`     �           �  ,      :                    d   	            M         �t�bhhK ��h��R�(KK��h�C4   7   �   	         �            �        �t�bhhK ��h��R�(KK��h�C         F           �t�bhhK ��h��R�(KK��h�CX         �   @   �   	   
   �   �   
  4  �  [                           �t�bhhK ��h��R�(KK��h�C,         #   �      �               �t�bhhK ��h��R�(KK
��h�C(      K  g      �   �   \        �t�bhhK ��h��R�(KK
��h�C(                  B   &        �t�bhhK ��h��R�(KK1��h�C��   G        8      	   E   �     c     }   �   �      8         a                  J  �      �   �      .      R   �  j   -                B        �           �t�bhhK ��h��R�(KK��h�C<U        ?   	  i           _                 �t�bhhK ��h��R�(KK%��h�C�   �  .      �  �   �        �  .      �      �                          �            H   Y   �            H   P         �t�bhhK ��h��R�(KK��h�C   �   O   �        �t�bhhK ��h��R�(KK��h�C\   
   
  F            L  k  �   
   ]   a   �              b   @   g         �t�bhhK ��h��R�(KK��h�C4�    l   �    �      %                  �t�bhhK ��h��R�(KK��h�C .   �  f     �             �t�bhhK ��h��R�(KK��h�C,*   �   }   �        :  @   g         �t�bhhK ��h��R�(KK��h�CX                  �  c  �   5      .      �   r
     -      j   ~         �t�bhhK ��h��R�(KK8��h�C�'      (               J   �  �  �     c                 �  "      E  ,   �                                 �   �  2   %           E         "       	     "           3         �t�bhhK ��h��R�(KK	��h�C$      A  6                  �t�bhhK ��h��R�(KK<��h�C�         	                    �  �         1      :      .            =  �  ;         :   	      ;   �  	              �  1   �  c                        �            W   �   
                 �t�bhhK ��h��R�(KK
��h�C([  @   m   `         *            �t�bhhK ��h��R�(KK��h�C   
      �        �t�bhhK ��h��R�(KK��h�C0        �      *         G
           �t�bhhK ��h��R�(KK��h�C@               d   
      �   �  W      u   �         �t�bhhK ��h��R�(KK��h�C   &   y     �t�bhhK ��h��R�(KK��h�C\   
   �      �         �     u   �  &                  
   s   o  �         �t�bhhK ��h��R�(KK��h�C|!      �  H   3      ]  "            �      �  I            &      
         �      Y      �            �t�bhhK ��h��R�(KK��h�Cd   !   K   ;  H      !   K              �  @   �     �  
   V   �      =           �t�bhhK ��h��R�(KK��h�Ch   �   m         �   F      r                 �
        �     �   	   �  �   �        �t�bhhK ��h��R�(KK
��h�C(
   �              @   �         �t�bhhK ��h��R�(KK��h�Cl   �   �   �           �     *   p         b  �       0      �  {   	     $   .          �t�bhhK ��h��R�(KK��h�C@   
   �   �     "   m  �     '     |  �   @         �t�bhhK ��h��R�(KK��h�Cx	   J   B   �  
   <   �            W   .   >           a   E      �           �                     �t�bhhK ��h��R�(KK3��h�C�   !        ]        V                       c  �                                 �         *  !   %   �            �   7   D  1  0   �                           �t�bhhK ��h��R�(KK��h�C,i  r  X     �     <  �   K        �t�bhhK ��h��R�(KK��h�CP'   >   (   '   �   (   	  9           t     +                     �t�bhhK ��h��R�(KK��h�CP      j   �                   �         	         �            �t�bhhK ��h��R�(KK��h�CL	   �                 4  y           	   R  ,   8   1         �t�bhhK ��h��R�(KK��h�C�              �t�bhhK ��h��R�(KK��h�C@   Q      g  �                   �  �  %        �t�bhhK ��h��R�(KK��h�C<
      "
        �  .            �  ^            �t�bhhK ��h��R�(KK��h�C`!   *   C                       �         	            �     �   �           �t�bhhK ��h��R�(KK��h�C       �        4        �t�bhhK ��h��R�(KK��h�CD   7   B   	   �   �  <  !      )   V      %   Q            �t�bhhK ��h��R�(KK
��h�C(               :  @   �          �t�bhhK ��h��R�(KK��h�C,n   D   �   �   d      �   �  Q        �t�bhhK ��h��R�(KK%��h�C�s  z
     Q  �   �         e   Q        	     �   &   �  �   �
  M     �      k           2  	            "      �        �t�bhhK ��h��R�(KK��h�Ch!        P  Y           ,   .      M        g        ,   �   �        �            �t�bhhK ��h��R�(KK��h�C f         �   �   �        �t�bhhK ��h��R�(KK%��h�C�v  �   �   �                3      ,            1   	         �                  `   �  
            	   D   �           �t�bhhK ��h��R�(KK��h�CLK   5   �  �      K            �        K                     �t�bhhK ��h��R�(KK��h�CL           +      �           �           8   P   �        �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK"��h�C�
      �     }     5   �  	            �          C     �                 
   �   �  �           #        �t�bhhK ��h��R�(KK��h�C<�  )         -  Y   $           8      �        �t�bhhK ��h��R�(KK��h�C@   
   �   S      1            �         $            �t�bhhK ��h��R�(KK7��h�C�   
   e     
   �   3               )      a            �   �   
   3   R
     
   )   �      �  3         z                  �   �   �      �         �        s   �     �   d            �t�bhhK ��h��R�(KK/��h�C�   �  	      ;      1         _  2   F  ;         �  	      �   .              �        4           �   \           	   9   Q            f     !        �t�bhhK ��h��R�(KK	��h�C$      �   �                  �t�bhhK ��h��R�(KK��h�Cx      �           	            /
                    $            ?   �     	         �        �t�bhhK ��h��R�(KK��h�C4   �                 �                 �t�bhhK ��h��R�(KK��h�C4      �     �           �  �  j
        �t�bhhK ��h��R�(KK/��h�C�B      
   V      �     u   �   y   �           u   �         g         @  <  /   ?         2         u   �         �  �  �  
   �        "  V   �         �t�bhhK ��h��R�(KK��h�C<
   �        B	     �	     �  �                �t�bhhK ��h��R�(KK	��h�C$9   �   /            �        �t�bhhK ��h��R�(KK��h�CH!   V  �      �           I   	         5   U   �   s        �t�bhhK ��h��R�(KK	��h�C$%                           �t�bhhK ��h��R�(KK��h�C8�   ,      �   )        x   �                 �t�bhhK ��h��R�(KK��h�C`      �   �      �   �           �   �      �               �  �  2   �	        �t�bhhK ��h��R�(KK��h�C  �         x        �t�bhhK ��h��R�(KK��h�C`        �         �         �        )   n   C     l  A   �         �        �t�bhhK ��h��R�(KK��h�CH               G      �              �   �  N            �t�bhhK ��h��R�(KK2��h�C�   |                   2   �       �        !   
   �  0   a              0      	        �  �  �            	              Y  �      �  a                 �t�bhhK ��h��R�(KK��h�Cx   �      C                          �
  2                       q           �  s	  i        �t�bhhK ��h��R�(KK��h�C4   K   :   &   ;         I   =  7            �t�bhhK ��h��R�(KK��h�CT   y              B     	   �   �     +      2      F               �t�bhhK ��h��R�(KK!��h�C�K   r           �           �     3      K                     �     �   �   ^     K            3         �t�bhhK ��h��R�(KK	��h�C$   )   h         q   d        �t�bhhK ��h��R�(KK��h�C0*      Y   	      +   _   1   �           �t�bhhK ��h��R�(KK��h�CT         �     �            �   .  +         �     ~              �t�bhhK ��h��R�(KK��h�Cx         �   5   %   �            !   %   �     }         }              !   %   �     }   �        �t�bhhK ��h��R�(KK��h�Cp   9   /   C   �   G      S            �     8                     %   �            �         �t�bhhK ��h��R�(KK��h�C   t   �     X        �t�bhhK ��h��R�(KK��h�CL   �  3   	   )           t   �           ,   \   �  �        �t�bhhK ��h��R�(KK��h�C0                     M              �t�bhhK ��h��R�(KK'��h�C�	   �     �   
               �   w      r                     �   F         	      �   -   �	        	   D            �  k         �t�bhhK ��h��R�(KK��h�C,   �      �     �        �        �t�bhhK ��h��R�(KK��h�Ct
   �                                               %                        �   �
        �t�bhhK ��h��R�(KK��h�CP%   s                  M         P  �     �           F        �t�bhhK ��h��R�(KK
��h�C(H
     �     �  "              �t�bhhK ��h��R�(KK��h�C<      #   v   
   �   M
     =        �  G         �t�bhhK ��h��R�(KK��h�C@         p  @   g   �  
   #         �              �t�bhhK ��h��R�(KK��h�C\*   �     �     �   �        a   P  Y           g   �   -      a   ^        �t�bhhK ��h��R�(KK��h�C   
            �t�bhhK ��h��R�(KK��h�C   �   9         �      �t�bhhK ��h��R�(KK��h�CP
   4         �         �              �   	   b   E      6         �t�bhhK ��h��R�(KK��h�C`   ^   ?     )         U   #     �  X
  	      t  i      "      G   N            �t�bhhK ��h��R�(KK��h�C\      q     h  !   �        $            !         \   �  l      w	        �t�bhhK ��h��R�(KK��h�C0t         �         8   /   ?   d        �t�bhhK ��h��R�(KK
��h�C(  f      "   Z                   �t�bhhK ��h��R�(KK��h�C@K  �   |   =   �      y                     d	        �t�bhhK ��h��R�(KK��h�C`        <      �
        B     h   &        /      q         N   D   q         �t�bhhK ��h��R�(KK
��h�C(
   L      .      X              �t�bhhK ��h��R�(KK	��h�C$            �  P            �t�bhhK ��h��R�(KK��h�C8      j          \      	         �        �t�bhhK ��h��R�(KK��h�Cx   	   7      �        �  $   �   �   ?     	   C               �   0           -   V               �t�bhhK ��h��R�(KK��h�C`   �   �  r     �  P
  G                  �   �        	      �      �        �t�bhhK ��h��R�(KK��h�C1      +   �
        �t�bhhK ��h��R�(KK��h�CL      �   ,   [         B   E         $      "         8         �t�bhhK ��h��R�(KK��h�C\   6        	   �   7        �                 0         	              �t�bhhK ��h��R�(KK��h�CD
      �     �                 
                   �t�bhhK ��h��R�(KK��h�CX                 J        v           �     �        �   c         �t�bhhK ��h��R�(KK��h�Ch�      U         	               �     %              o     ?        2   y         �t�bhhK ��h��R�(KK��h�C4      P     G          �     #         �t�bhhK ��h��R�(KK��h�C|
            P   !      p      
   �   5   �        i     �           ]   �   �   3      =     '        �t�bhhK ��h��R�(KK$��h�C�'     (      �  �  2      ^	  9      �           P     �   5   9   U   �                  r      S   5   U              �t�bhhK ��h��R�(KK��h�CT        #  �  J   A  .     �  ~            �   �  &   �  �	        �t�bhhK ��h��R�(KK��h�CL
   N  K     �        ?  @                     r   �        �t�bhhK ��h��R�(KK��h�Ch   
   Z               �           �  +      v  !      �                           �t�bhhK ��h��R�(KK��h�CX         �              =   �     �   	               Q     �	        �t�bhhK ��h��R�(KK��h�C\                           	   K  �                 	   K  �            �t�bhhK ��h��R�(KK��h�C,   H  ,   .   %   �   R              �t�bhhK ��h��R�(KK��h�C8  �      �   i         �t�bhhK ��h��R�(KK��h�Cp        �           %   z
     �  $      �    �  @         �     �  %   V   �   /         �t�bhhK ��h��R�(KK	��h�C$      ~        Z  ~        �t�bhhK ��h��R�(KK��h�C`   �  3     �  �  $   �      A        D  �
  6     !      �         -        �t�bhhK ��h��R�(KK%��h�C�
      �      W        
   Z         
               ,  �   =   D        R    e   ,         �     	      5     D         �t�bhhK ��h��R�(KK��h�C          :   �           �t�bhhK ��h��R�(KK��h�C   
   f          �t�bhhK ��h��R�(KK��h�C          8  ^   �         �t�bhhK ��h��R�(KK��h�CR      6   �	         �t�bhhK ��h��R�(KK+��h�C�            %   �   �  �     �   @   G         "  .                  �  .      �      	     4  �      .      C   ,               A            �t�bhhK ��h��R�(KK��h�C`                          1                                 �        �t�bhhK ��h��R�(KK��h�C8   �         s   �           �     C         �t�bhhK ��h��R�(KK��h�C         (         �t�bhhK ��h��R�(KK��h�C<   ^            �     �   �      I   �        �t�bhhK ��h��R�(KK��h�C
         T  )        �t�bhhK ��h��R�(KK��h�C      �  +   3         �t�bhhK ��h��R�(KK��h�C@      r         �  
  	   T     +   �  �            �t�bhhK ��h��R�(KK��h�C,.   �        ;            E          �t�bhhK ��h��R�(KK
��h�C(      b   T                    �t�bhhK ��h��R�(KK ��h�C�            �        ]  �     �   \         	      �        �              	      �   	               �t�bhhK ��h��R�(KK��h�CtJ      ,   �   [   �      S  8   �   
     _      C   �          2     �     }  $   I   �         �t�bhhK ��h��R�(KK��h�C4'   �   (   �         }  g   
      ~         �t�bhhK ��h��R�(KK��h�C@      <   >     R              8   =               �t�bhhK ��h��R�(KK ��h�C�            �      �  	   |                      8   3   �     c      �            >  �   �  v        �t�bhhK ��h��R�(KK)��h�C�   �                  2      2      �      y
           �        o           �   �        J        o        m   t   �     A        �t�bhhK ��h��R�(KK��h�C\   
   N   �      �     	      =   �           �      
   ]   e      #         �t�bhhK ��h��R�(KK��h�CDt                       E     x           3         �t�bhhK ��h��R�(KK!��h�C�   
   �              h               $   I   =        g   8           �           F                    �t�bhhK ��h��R�(KK��h�C@�        n   �         �     G  �      �           �t�bhhK ��h��R�(KK��h�CT'   >   (   -              8   �        �      s  �  ,   �   �         �t�bhhK ��h��R�(KK��h�C   �      �t�bhhK ��h��R�(KK
��h�C(!      �   �   O	  
   F   V        �t�bhhK ��h��R�(KK.��h�C�!   1   �  ;   
   �     $  ;   
   )   �            �                 
   C            g        !      �   `               �          [  �  J        �t�bhhK ��h��R�(KK��h�Ch      S  x   �        Z     J         f   z               $      2                  �t�bhhK ��h��R�(KK��h�C          1   	   �        �t�bhhK ��h��R�(KK��h�CL      3  +      4  �	     U   �  v         \   �     �        �t�bhhK ��h��R�(KK��h�CT        /      	      �        �        �  �   Q                 �t�bhhK ��h��R�(KK��h�C4   )         v     '        2           �t�bhhK ��h��R�(KK��h�Cp      7              	         G     N                 q      �                       �t�bhhK ��h��R�(KK��h�Cty   �   j  /            	      +  t                 �        �   �  �   3      �  t   �        �t�bhhK ��h��R�(KK��h�C   f             �t�bhhK ��h��R�(KK��h�C8^      �  �      E     �        	            �t�bhhK ��h��R�(KK��h�C,�   
   �         �  �     D        �t�bhhK ��h��R�(KK&��h�C�   1         �              <               5           7   I   �  �         +   B   �       	      k         B   E         �t�bhhK ��h��R�(KK��h�C4�  @   !        �   $  &                 �t�bhhK ��h��R�(KK��h�CT7  z            ~      E        Y     �      Q   F      1   o          �t�bhhK ��h��R�(KK��h�C@   C   1   [      �   3  �  7     �  ,               �t�bhhK ��h��R�(KK��h�CD0      �               b     �     ^   c     Q        �t�bhhK ��h��R�(KK��h�C         "                �t�bhhK ��h��R�(KK��h�C@'   >   (   G     
   �      G  �   ]   
   �           �t�bhhK ��h��R�(KK*��h�C�                  �         �  )         d              �     �     �              j                 J      	      E  �  �         �t�bhhK ��h��R�(KK��h�C\'   L  (   �        e   �     n  N  
      �  �                   C     �t�bhhK ��h��R�(KK��h�C �   �   
     C   �        �t�bhhK ��h��R�(KK��h�CH
   L    [      8  �  �             +                 �t�bhhK ��h��R�(KK��h�Cb  H            �t�bhhK ��h��R�(KK ��h�C�
         #      �   o   ;   	         	      ;         #      �
  /            
         .   
      �        �t�bhhK ��h��R�(KK
��h�C(                     �        �t�bhhK ��h��R�(KK��h�CT=                        �  �  �                    �  7        �t�bhhK ��h��R�(KK!��h�C�   !   
   �      T   �           �   6                  �         �   T       �      �            �        �t�bhhK ��h��R�(KK$��h�C�      �     �  
   F         �     �  r      3            .  4     �            �	        
   9     
   O   �        �t�bhhK ��h��R�(KK��h�C@   T
        �         m      {  T
  	               �t�bhhK ��h��R�(KK��h�C,   O         =  �   	      M	        �t�bhhK ��h��R�(KK��h�C,K      �     E   	   w   �            �t�bhhK ��h��R�(KK��h�CL   4              s       �              `   �  ;        �t�bhhK ��h��R�(KK	��h�C$               �  N         �t�bhhK ��h��R�(KK��h�CH!      �  �   �           �             f              �t�bhhK ��h��R�(KK&��h�C�   �   
      �     �     
   D      e            
   D   :   M   f     ;   :   �   #         f     
   D   M   /   �              �t�bhhK ��h��R�(KK��h�C�      �         �t�bhhK ��h��R�(KK��h�Cl         	   �  �   �                                            �     =            �t�bhhK ��h��R�(KK3��h�C�      ^                  ,   �         !            	                 �   �         �         A           �   �         P   &      I      #               h           �t�bhhK ��h��R�(KK��h�C\   	      1      �  �   y     _  �        �           �                 �t�bhhK ��h��R�(KK��h�CD�              �   :     6  �     �   6   
           �t�bhhK ��h��R�(KK��h�C89       �     8     _      �   @                �t�bhhK ��h��R�(KK��h�C�  �        �        �t�bhhK ��h��R�(KK��h�CH        2   �   1     �                 5  �           �t�bhhK ��h��R�(KK	��h�C$   *  =   ^  ]   U   >        �t�bhhK ��h��R�(KK��h�C8                  {      �  �              �t�bhhK ��h��R�(KK��h�C4   5   q                    1           �t�bhhK ��h��R�(KK��h�CT   '  y                                 �         �   �   2        �t�bhhK ��h��R�(KK��h�C8        
      �   �
        �      �         �t�bhhK ��h��R�(KK��h�CH
   ;  H         <                  4      G              �t�bhhK ��h��R�(KK"��h�C��  2         G   �  [      �  h                    o   	            �  �     v   >  N     I                 �t�bhhK ��h��R�(KK��h�C0      L  #   !   
   5   �  �            �t�bhhK ��h��R�(KK��h�C@   �
     
   6      �     	   �   )      q            �t�bhhK ��h��R�(KK��h�C8      %                        {   �        �t�bhhK ��h��R�(KK��h�C      C        �t�bhhK ��h��R�(KK��h�C0   
   Z            	      �           �t�bhhK ��h��R�(KK(��h�C�      s         7     W               7     �               7      ,  �  2     �
        �     �   r     r  H         B         �t�bhhK ��h��R�(KK��h�C,e         �      f                 �t�bhhK ��h��R�(KK��h�Cl   )         
     P               I   
   �      �        R                         �t�bhhK ��h��R�(KK��h�C8      >  ,   F        �     �     1         �t�bhhK ��h��R�(KK��h�CL   :      �  m         #     w        �   �     ?          �t�bhhK ��h��R�(KK��h�C\
            w  $   �     �                  Z   
      
   ,              �t�bhhK ��h��R�(KK/��h�C�'   >   (            
         �  �     {         
      �  �  $
           .   $
     [            .      j     �  ?            4           �   C        �t�bhhK ��h��R�(KK��h�C@         �     �                @   g   G         �t�bhhK ��h��R�(KK��h�Cp!         )  �     P  �                               P   P   +      F        �        �t�bhhK ��h��R�(KK��h�C,   &           d                 �t�bhhK ��h��R�(KK��h�CH*   �        z     a   �  0            �   �     �        �t�bhhK ��h��R�(KK��h�C4      �     %   �   V         �  �        �t�bhhK ��h��R�(KK��h�Cl      �   j   4     �                 j   �              S     3   +   /   �
           �t�bhhK ��h��R�(KK��h�C          �	  �   �         �t�bhhK ��h��R�(KK��h�C             H           �t�bhhK ��h��R�(KK��h�Cd   `        =               ]  q   Q        �   O     y  	   /   �   �           �t�bhhK ��h��R�(KK%��h�C�!         W   �              Z               �     �  /     Y  f      f   l         �  �  �  �      U      �  /        �t�bhhK ��h��R�(KK��h�C4   
   �  S      �  �     b  I  @        �t�bhhK ��h��R�(KK��h�CH   	  *     r   �  g   4   �              �   �           �t�bhhK ��h��R�(KK��h�C         �         �t�bhhK ��h��R�(KK��h�CH      2      $   Y   �         %      :   n   	   �   �        �t�bhhK ��h��R�(KK��h�C,   g   �  
               0        �t�bhhK ��h��R�(KK��h�Cz           �        �t�bhhK ��h��R�(KK��h�Cl
   5     ,  `   �        2      2      2     �   &     a   P      w   �  V      A        �t�bhhK ��h��R�(KK��h�C         �        �t�bhhK ��h��R�(KK	��h�C$C   	   
         9   �        �t�bhhK ��h��R�(KK��h�C8            �     �     �                 �t�bhhK ��h��R�(KK��h�CL�  �  x                          /   5      �
  2            �t�bhhK ��h��R�(KK��h�C0   1     +     �     �     @         �t�bhhK ��h��R�(KK
��h�C(
   �   �  3   {      j
           �t�bhhK ��h��R�(KK��h�C<     W     
   �   �   �      .   �                �t�bhhK ��h��R�(KK��h�CH   e  3  _         b                    i               �t�bhhK ��h��R�(KK��h�Ch
   �      �     
   N  �      
   4      <  �     �  �  D                          �t�bhhK ��h��R�(KK��h�C   "          �t�bhhK ��h��R�(KK��h�CD      �   U   /     +   /   ?   7  �   ?   �     ,        �t�bhhK ��h��R�(KK��h�CP   G         J         \      	   z   �     �   [      0            �t�bhhK ��h��R�(KK
��h�C(         �           M        �t�bhhK ��h��R�(KK��h�CP=   ^  �      #              y      +  
   8  V      \   �        �t�bhhK ��h��R�(KK��h�C@   �     X  �         �            q   t  x        �t�bhhK ��h��R�(KK	��h�C$            �   P   �         �t�bhhK ��h��R�(KK ��h�C�                 �     	   u      �     Y      �      J  $            G         �  '                �t�bhhK ��h��R�(KK	��h�C$   q   ]  6  3      �        �t�bhhK ��h��R�(KK��h�C       &      {            �t�bhhK ��h��R�(KK��h�C|      h   a  �   S        0         
   O        
   :   �   �      5   /   B      9   L      �           �t�bhhK ��h��R�(KK��h�C     
           �        �t�bhhK ��h��R�(KK��h�C0'   >   (   g  g         �     3         �t�bhhK ��h��R�(KK��h�C@      �  U      :               {                  �t�bhhK ��h��R�(KK��h�Cu   o   s   3            �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C'     (               �t�bhhK ��h��R�(KK
��h�C(   <   �           <            �t�bhhK ��h��R�(KK��h�C40  	   ~   �  
   �   �  	   �      #         �t�bhhK ��h��R�(KK��h�C
                     �t�bhhK ��h��R�(KK��h�CL      _               �           �                      �t�bhhK ��h��R�(KK	��h�C$   )      6   5
  5  �
        �t�bhhK ��h��R�(KK��h�C0�  �           z     8   E   �	        �t�bhhK ��h��R�(KK��h�C@   B           Q         G      
   �   M            �t�bhhK ��h��R�(KK$��h�C�   �                       �  �        t	        �                       <   �   {	                             �t�bhhK ��h��R�(KK��h�C@   &   
         �	  #         �  d      
   c         �t�bhhK ��h��R�(KK��h�C4   s   �           M   1      4  3         �t�bhhK ��h��R�(KK(��h�C�            a      ,  F   +   �                       3            o   	   ?      ~     8      G  L   "      f   )      a   �         �t�bhhK ��h��R�(KK��h�C@u                  �                              �t�bhhK ��h��R�(KK��h�C<   �        *   4      �  �     r             �t�bhhK ��h��R�(KK��h�C0�  #            �        �            �t�bhhK ��h��R�(KK��h�C@      �   G            �     )                     �t�bhhK ��h��R�(KK��h�CP               "   	   �   !   �     t   �  �                    �t�bhhK ��h��R�(KK	��h�C$v           �     �        �t�bhhK ��h��R�(KK��h�C\'   >   (      &   p   *         5         $         A   	      �   7  G   �      �t�bhhK ��h��R�(KK��h�C      w            �t�bhhK ��h��R�(KK"��h�C�      n  �         �  	      p      P      8   $      ]         �         �            s     
         s        �t�bhhK ��h��R�(KK(��h�C�   7   E   ;   r      
   0     ;   	      �     	   Z      z  {           	   S     	   z   e   <   �
  v   X  �        C   -   �        �t�bhhK ��h��R�(KK4��h�C�      7   j  1  0   %   _  �        �            	         �  	   �     |         t        k     �        �  �
     -   �   �   x                             �        �t�bhhK ��h��R�(KK��h�C4      �  �         �   �     w            �t�bhhK ��h��R�(KK��h�C'   
         �   (      �t�bhhK ��h��R�(KK��h�CD   z   P      �  A         :               t            �t�bhhK ��h��R�(KK��h�C0              #   ;   
               �t�bhhK ��h��R�(KK��h�CL�  2   �  �  (  �	        U      	   �  t   v  �   &           �t�bhhK ��h��R�(KK ��h�C�   c     �  ^            �        �              "                    	   �
  ,   +   ,   �             �t�bhhK ��h��R�(KK��h�C   s      }        �t�bhhK ��h��R�(KK-��h�C�      �     	   �                 �                  �    �      t                 H           D     0            #     H  q  +            �t�bhhK ��h��R�(KK��h�Cp      A  s      /   �   `       j   �     v   {            }     )            �  I         �t�bhhK ��h��R�(KK��h�C,  �         �  �     �  �  �      �t�bhhK ��h��R�(KK
��h�C(      7      z  	   Y           �t�bhhK ��h��R�(KK��h�Ctr  m            �                  �                  B  
      �   `   $  �   '  @   !        �t�bhhK ��h��R�(KK��h�C0'   >   (   �   G         T               �t�bhhK ��h��R�(KK��h�CX   �   W  �                 �  �   S   ;     �   ,         �           �t�bhhK ��h��R�(KK��h�C4�  @   !          "   	   �              �t�bhhK ��h��R�(KK��h�Cx      C         �             C         6     )   n      �   m   �   A   .  .      I  <           �t�bhhK ��h��R�(KK��h�C
   �  3   �         �t�bhhK ��h��R�(KK��h�C<   �      
                  
   �               �t�bhhK ��h��R�(KK��h�C                     �t�bhhK ��h��R�(KK ��h�C�      )   :      q   �  �     k              �  )   �   �        t   ~   h           z   p              �t�bhhK ��h��R�(KK��h�C<        �           =   �        
            �t�bhhK ��h��R�(KK!��h�C�         :      >  W     �      j   �       <            `	        6            �   F   �                  �t�bhhK ��h��R�(KK��h�C                  �t�bhhK ��h��R�(KK%��h�C�        
             n               ]  "       3   :           �      ;        9  ?      ]  "  �   #            �t�bhhK ��h��R�(KK��h�Cp     R        R      a         �            �  h  �  K      Q        �                 �t�bhhK ��h��R�(KK��h�Ct      w         �  E   	               �	     �           �      C        U  &              �t�bhhK ��h��R�(KK	��h�C$     ,   r      ?            �t�bhhK ��h��R�(KK*��h�C�5      �   \         ~        q  �  �        +  3   +      �      $   5      I	  3   f            *	         	            g                �t�bhhK ��h��R�(KK��h�C0         3         
   �  #   i         �t�bhhK ��h��R�(KK��h�C4            s    �   +                 �t�bhhK ��h��R�(KK��h�C         9   (  [        �t�bhhK ��h��R�(KK��h�CP                C         *                     !      �        �t�bhhK ��h��R�(KK	��h�C$                  G         �t�bhhK ��h��R�(KK��h�C@   %      6        �        .   J   �  	   D        �t�bhhK ��h��R�(KK��h�C   g   �  K   �        �t�bhhK ��h��R�(KK&��h�C�   
   L            7   I     !           �     N        ~      `   �  (     v  	            
     
  	   �             �t�bhhK ��h��R�(KK%��h�C�      L                  �   p          A   
                    A     
            �               2  �  �        �t�bhhK ��h��R�(KK	��h�C$�   #   �   3  ?   �   d         �t�bhhK ��h��R�(KK��h�CTV  �     E    %  v  N   �            �         "   	   �  1         �t�bhhK ��h��R�(KK��h�C,   �     �  7        �  �
        �t�bhhK ��h��R�(KK��h�C4
   c     �      �        �  [            �t�bhhK ��h��R�(KK��h�C<         	   �   F                     �	        �t�bhhK ��h��R�(KK��h�C\�   �  
      I   	   �
                    `  �     5          �          �t�bhhK ��h��R�(KK3��h�C̋         ]   T  "   y   �  C      y      /     O      �   a                                      >     {           )      �   �   �      ?   �  	     	   �  3         �t�bhhK ��h��R�(KK��h�Ch   R   8   1      E   	                 �
       5     �  	        �              �t�bhhK ��h��R�(KK��h�CD   �     	        �     �      �   V         _         �t�bhhK ��h��R�(KK
��h�C(         �    	      �         �t�bhhK ��h��R�(KK��h�CT           �      $            a         �  -      �               �t�bhhK ��h��R�(KK
��h�C(      g      �   �  G           �t�bhhK ��h��R�(KK��h�C8!   
   �           �  
      
   �           �t�bhhK ��h��R�(KK��h�Cx            C   Y  2   �     Z     Q  F   z  +   r
           �      V         ;         �        �t�bhhK ��h��R�(KK
��h�C(                 <   �        �t�bhhK ��h��R�(KK��h�C4   b   d            L    \  �   #         �t�bhhK ��h��R�(KK��h�CD�     &      O   �   8                     �   �        �t�bhhK ��h��R�(KK5��h�C�   t   s     t   s  &   7     �  �         V
           l  �  ;      9   L   �   ;   7     �    3   �                     �     }      d     �              +               �t�bhhK ��h��R�(KK��h�CT   �  /   V         $                  m         -      �   n         �t�bhhK ��h��R�(KK(��h�C�   �
     u   |     �  F            �	           �   |                                      M  H      �   �  V                  �t�bhhK ��h��R�(KK��h�C@    
     �           W  z      �      S  �        �t�bhhK ��h��R�(KK��h�Cp   %   �   Y   	                  �            /                           <   �  �        �t�bhhK ��h��R�(KK��h�C4�  H      Q              j  2            �t�bhhK ��h��R�(KK��h�C8               O   �   �         I   o         �t�bhhK ��h��R�(KK��h�C|�              G               	   �     F   Y   
              �  �              �              �t�bhhK ��h��R�(KK��h�Ct
   �   e   �      4  �                 o  ]   
   6      [  s           p  e   #   x  �         �t�bhhK ��h��R�(KK��h�C<                  	   �      F   &               �t�bhhK ��h��R�(KK��h�CT'   >   (   �   e     �           �        
   �   #                  �t�bhhK ��h��R�(KK ��h�C�
   �   �     m     b      �   �     #   �   	   �   �   	         U     u         	            k           �t�bhhK ��h��R�(KK��h�C<!   ^  �   F   +   �  4   *         >  �  -         �t�bhhK ��h��R�(KK,��h�C�
            �     W   D  @   G               S   	   c   5  0      �  ^                    a     n            7      �     �     t   N
        �t�bhhK ��h��R�(KK(��h�C�   �   �        #  *        M         �         M      �  W         m  �         M         ;      �          �  U     }        �t�bhhK ��h��R�(KK��h�C0y  �  ]   �  y  H  �   �  @            �t�bhhK ��h��R�(KK��h�Cd     �  c      4  �                   w            `	        �      �        �t�bhhK ��h��R�(KK��h�CL      N      �  �  �  �  E                      �         �t�bhhK ��h��R�(KK��h�C 	   �  �                 �t�bhhK ��h��R�(KK��h�C<   u         �   `               2               �t�bhhK ��h��R�(KK��h�C8K      w                     �  �      9     �t�bhhK ��h��R�(KK	��h�C$%   s      �         �         �t�bhhK ��h��R�(KK	��h�C$      G   D   N  1            �t�bhhK ��h��R�(KK��h�C\   �  C  ;      �  C     k   	            �   �  	   
   �                 �t�bhhK ��h��R�(KK��h�C,�   �  
   #               �          �t�bhhK ��h��R�(KK��h�C<
   s            �        $      �   s            �t�bhhK ��h��R�(KK��h�C8t     )   9   �        	         �           �t�bhhK ��h��R�(KK��h�CD   �   �        Y      �  �     v                     �t�bhhK ��h��R�(KK��h�C,         �     �   	   T           �t�bhhK ��h��R�(KK,��h�C�   !   
   �   "   	            �          	        5   
   �      �              �              �  A   N         5      6      T   i   �        �t�bhhK ��h��R�(KK)��h�C�      O      �  `   �   &   .   z      j     2         �     	            G            �                     `   7  +   �  2   F         �t�bhhK ��h��R�(KK.��h�C�   L      �      +   �     "   	      �        	      �  �  &      �      P              6            �   A  �                  	     �              �t�bhhK ��h��R�(KK��h�C,M   :                 .  �        �t�bhhK ��h��R�(KK��h�C9   (                  �t�bhhK ��h��R�(KK��h�CT   9      �        ,   /   ;         X  7  	   M           �        �t�bhhK ��h��R�(KK1��h�C�      
   R     9        #         ?   d   	   
   �   +     S                  3      �  Y   i     3     '   >   (   g        "      �      /   �                  �t�bhhK ��h��R�(KK.��h�C�         .
        w                    	   �  z  m      %   4   �     !      :   �         F         �   ~   +   �        t   �           t            �t�bhhK ��h��R�(KK��h�C\u      �   ]   w   �	  V         �   �         u   �           �     i         �t�bhhK ��h��R�(KK��h�C,   �     �  +  A      A            �t�bhhK ��h��R�(KK��h�CT0   7   �  �      	           �  :            R   q   �     3         �t�bhhK ��h��R�(KK��h�C,     g   �        �   �  �         �t�bhhK ��h��R�(KK��h�C0
   L            9   L   "      �        �t�bhhK ��h��R�(KK	��h�C$f  g              �        �t�bhhK ��h��R�(KK
��h�C('   >   (      �     �  �        �t�bhhK ��h��R�(KK
��h�C(      �        	   z            �t�bhhK ��h��R�(KK��h�CD   A     T        b  F                  4           �t�bhhK ��h��R�(KK��h�Ct            �  �      �              ,                          �      f                  �t�bhhK ��h��R�(KK��h�C<         �   m            -         }            �t�bhhK ��h��R�(KK��h�Ct1   �  -   6   <   +  j  @   !  f   �     �  #   q   �           #            |     �  �        �t�bhhK ��h��R�(KK#��h�C�=      )  �                            
      �           5  F   G     m  �           *      =   m  �        �t�bhhK ��h��R�(KK��h�C@      	   k
  /
  	   �          �        L
        �t�bhhK ��h��R�(KK��h�C_   �      �            �t�bhhK ��h��R�(KK<��h�C�      K               
            �  +         $                +      s  �                 �                 	   �            O   U   ;      �  ;      O   U   �     �           j   �         �t�bhhK ��h��R�(KK	��h�C$
   ]   l	     
   ]   �        �t�bhhK ��h��R�(KK ��h�C�   
   Z      !      �  m        O      M            �   �  �        �   
	  	   �        4  G  �        �t�bhhK ��h��R�(KK��h�C@      H   ^   6
  y  �        E     �      \        �t�bhhK ��h��R�(KK��h�CT   	      �   !         �        b   �        C   P      :   }        �t�bhhK ��h��R�(KK��h�C0?   �  +   o           �   ,   �        �t�bhhK ��h��R�(KK��h�C0   x      S     ,  	        �        �t�bhhK ��h��R�(KK#��h�C�	   Y   	        �        �  �  	      ^            
   �         �  	      T   �  �      2   �     �  W            �t�bhhK ��h��R�(KK��h�C@
   �              @            �                 �t�bhhK ��h��R�(KK"��h�C�      B   �  	      q   �     �         2                  �         �      �            	   �      ^   �        �t�bhhK ��h��R�(KK��h�CP         �
       	         .  ;   '   >   (      +  )            �t�bhhK ��h��R�(KK��h�Cd[     X      �               �  X      ?     +   /           3   �   I   �         �t�bhhK ��h��R�(KK ��h�C�         i           5      2  ?  �      o                       M            �     �  �           �t�bhhK ��h��R�(KK��h�C`1            �     �  �   �        g      �     �  �      �                  �t�bhhK ��h��R�(KK��h�CL   7   �   &                 
     �  <  �  u      �        �t�bhhK ��h��R�(KK
��h�C(   #                           �t�bhhK ��h��R�(KK��h�C`K   �            7   I   A      N                  y                           �t�be.