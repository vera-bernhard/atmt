����      ]�(�numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i4�����R�(K�<�NNNJ����J����K t�b�C8)            '         �                    �t�bhhK ��h��R�(KK��h�C0  �                                �t�bhhK ��h��R�(KK��h�C0   �            o                    �t�bhhK ��h��R�(KK��h�C�              �t�bhhK ��h��R�(KK��h�C4     #     �     M            �        �t�bhhK ��h��R�(KK��h�CP            
              a     2        \   �      c         �t�bhhK ��h��R�(KK��h�C0'     N        �   '                 �t�bhhK ��h��R�(KK%��h�C�G   %   ]  �     �   �        �      �        �     M   g
     �   �                                                   �t�bhhK ��h��R�(KK��h�CX                                            7     b  �  �        �t�bhhK ��h��R�(KK(��h�C��         �   J   �  ]         �  �  T        V   2      �                       V         0        �  
   _                     �t�bhhK ��h��R�(KK��h�C,         �              �         �t�bhhK ��h��R�(KK
��h�C(�   ]      #  '                 �t�bhhK ��h��R�(KK��h�C8y   �     �  J   �      +  �         ]         �t�bhhK ��h��R�(KK��h�CP'       �   �        I  �                 b                  �t�bhhK ��h��R�(KK��h�Ch�      �   D  w   -      �   �     ]        %            �   �   J         �            �t�bhhK ��h��R�(KK	��h�C$#  �        ]        r      �t�bhhK ��h��R�(KK��h�C    �  �                 �t�bhhK ��h��R�(KK��h�C4               5   �           �  r      �t�bhhK ��h��R�(KK&��h�C�         4	      9   �        <              ]              ]     (                 '
     �         
      ]  �	        �t�bhhK ��h��R�(KK��h�CL�             *        %      �  	  �      b              �t�bhhK ��h��R�(KK��h�C�  9               �t�bhhK ��h��R�(KK-��h�C��         ]  g           �      �   �               �               I         �           \         �
  �       �     D	           I            �t�bhhK ��h��R�(KK��h�Cx         
      %   �  s   
          �        %               �        %                    �t�bhhK ��h��R�(KK
��h�C(   &                  r   "     �t�bhhK ��h��R�(KK��h�Cd         �  �        �	     A         a     	     D  �  #        %   5        �t�bhhK ��h��R�(KK)��h�C�   ]       
                  �      )        �         ]     �      �                                 �  C   �     [           �t�bhhK ��h��R�(KK��h�C4�   �  �         +        �   N            �t�bhhK ��h��R�(KK��h�C0         '           �               �t�bhhK ��h��R�(KK ��h�C��   ,                       %         0     
   #     �  �      %      �                    I         �t�bhhK ��h��R�(KK��h�Cd               
   �        C      0            :         �      %     �        �t�bhhK ��h��R�(KK��h�C|   �      
      �      �              �   �   v                             �                     �t�bhhK ��h��R�(KK��h�CX�   D  7  S      �     	     �      :     o  �  �         �   �         �t�bhhK ��h��R�(KK��h�CD'  5   D  �  ,        D  �          �  "      r      �t�bhhK ��h��R�(KK��h�CH�      0                                   �            �t�bhhK ��h��R�(KK��h�C`   5     %      �             �      �      S      %         �  !           �t�bhhK ��h��R�(KK��h�C�                  �t�bhhK ��h��R�(KK��h�CH   8        �               �   �   �     �      -         �t�bhhK ��h��R�(KK��h�CH            �         �     �               
  L         �t�bhhK ��h��R�(KK��h�C\            *   '     �         �      �   �            �  �               �t�bhhK ��h��R�(KK/��h�C��   W  �  
   $           "     5  �   c      �      "        �   �     �      *  #  �        I   �  ?           V         �      ]                    �t�bhhK ��h��R�(KK��h�C|               2   W     �        �   �  �                                 P  �  W              �t�bhhK ��h��R�(KK��h�CX   �                     �      .   :                  H               �t�bhhK ��h��R�(KK��h�CT  '  d  %   n  '  d        m   '           �  0  %   s            �t�bhhK ��h��R�(KK��h�CL         �   �     *   %                              r      �t�bhhK ��h��R�(KK
��h�C(�      �  ]     �  �  ]        �t�bhhK ��h��R�(KK��h�C8
   A   �           �         �  
   )        �t�bhhK ��h��R�(KK��h�Cx                             �      %   -   �                [      �  �  �         �        �t�bhhK ��h��R�(KK��h�C0           7   �                    �t�bhhK ��h��R�(KK��h�CD      �        '        '     �     '              �t�bhhK ��h��R�(KK��h�CT   '        	             �                           �  r      �t�bhhK ��h��R�(KK��h�CD         (            I	     �                        �t�bhhK ��h��R�(KK��h�C0   �        '  .  �      �            �t�bhhK ��h��R�(KK��h�C<�   �     �                                   �t�bhhK ��h��R�(KK	��h�C$      &   '     
            �t�bhhK ��h��R�(KK��h�C0                 �     �   �        �t�bhhK ��h��R�(KK#��h�C��            �         I   N      
   W           *                             C        #                    �t�bhhK ��h��R�(KK	��h�C$�              �           �t�bhhK ��h��R�(KK��h�C �   �      �               �t�bhhK ��h��R�(KK/��h�C�   �              �           �   �     e        �                          %               G   �                            *                 �t�bhhK ��h��R�(KK��h�Cd   5  '              !  �     %   .        �                                 �t�bhhK ��h��R�(KK2��h�Cȳ   �   �               �         �      
   �        '           �           �  �        �   �         o               y
        �           �  �   {
           �t�bhhK ��h��R�(KK��h�Cx      ]           A         +           �      �
          �   J   N              \  �        �t�bhhK ��h��R�(KK��h�C4#  I   �                %               �t�bhhK ��h��R�(KK��h�C      �   /              �t�bhhK ��h��R�(KK��h�C0M      .               I   �           �t�bhhK ��h��R�(KK"��h�C�      �	  �      �                    2   6                    �     �  �     t  �   �   �         �        �t�bhhK ��h��R�(KK��h�CP      7   �        	     	  �     ]     �                     �t�bhhK ��h��R�(KK��h�C`*         -  C   �            V   %   s                  >      M      �         �t�bhhK ��h��R�(KK��h�CP   �  �  �  �                        �        �              �t�bhhK ��h��R�(KK��h�C<                                             �t�bhhK ��h��R�(KK��h�CX      �  2   5        
                                            �t�bhhK ��h��R�(KK��h�C   �      9   �        �t�bhhK ��h��R�(KK��h�C4y      �     H              �   7         �t�bhhK ��h��R�(KK	��h�C$         �   #   
   :        �t�bhhK ��h��R�(KK��h�C8�      �     �  �     �   /      �           �t�bhhK ��h��R�(KK��h�C`      �     +         �           a         5        *  A   \   2   �        �t�bhhK ��h��R�(KK��h�C%      -            �t�bhhK ��h��R�(KK��h�C8�      ]        �     o                    �t�bhhK ��h��R�(KK��h�CL�   '         p        N   �                 c   �  �  r      �t�bhhK ��h��R�(KK��h�C \   H      o  �     r      �t�bhhK ��h��R�(KK��h�C                     �t�bhhK ��h��R�(KK��h�Cd             �                �      �      �     �                   �        �t�bhhK ��h��R�(KK��h�C,      V         ~      $      r      �t�bhhK ��h��R�(KK��h�C,�         �            �        �t�bhhK ��h��R�(KK��h�C,o  o            a  ]   �           �t�bhhK ��h��R�(KK��h�C�  �   �               �t�bhhK ��h��R�(KK��h�Cd�         '     �                     *   '     �           \   ]               �t�bhhK ��h��R�(KK��h�C�                     �t�bhhK ��h��R�(KK
��h�C(      �                       �t�bhhK ��h��R�(KK��h�CD�   Q            �                 
         5        �t�bhhK ��h��R�(KK��h�C,�                               �t�bhhK ��h��R�(KK��h�Cp�   /   S  �   j                  [  8     �   %      a   �     �  N   8     �     /         �t�bhhK ��h��R�(KK
��h�C(]         �     I              �t�bhhK ��h��R�(KK��h�CL            
      ]  T                 :      A   T        �t�bhhK ��h��R�(KK��h�C8'  &               #           �            �t�bhhK ��h��R�(KK��h�Ct'     (                         �      �
  %                  �         �  V               �t�bhhK ��h��R�(KK
��h�C(         H            H         �t�bhhK ��h��R�(KK��h�C`                  �                 '           �     '        *        �t�bhhK ��h��R�(KK��h�C4   '   �           �     �   ]  �	        �t�bhhK ��h��R�(KK��h�C      %               �t�bhhK ��h��R�(KK��h�CX   �      �  7         �   �  w     d  N  �                           �t�bhhK ��h��R�(KK��h�C,�         �
  �     (              �t�bhhK ��h��R�(KK
��h�C(         �     �  �  �         �t�bhhK ��h��R�(KK
��h�C(               
   A   T        �t�bhhK ��h��R�(KK1��h�CĄ	           �                       �   L         �         0         �         �  L      �     
   \   '  &         �                 �        !           �t�bhhK ��h��R�(KK��h�C<        �      �   n                          �t�bhhK ��h��R�(KK%��h�C�      \         $               \         
   $            �              ^           �   �   �      %      �   +         �t�bhhK ��h��R�(KK��h�C�   �  >            �t�bhhK ��h��R�(KK��h�C\�   �      c                  �   �      0      
      {     s   7   �        �t�bhhK ��h��R�(KK��h�C4�
     �   �     �     2                  �t�bhhK ��h��R�(KK��h�C \      T      �      r      �t�bhhK ��h��R�(KK��h�C,�   �  �            q  7   �        �t�bhhK ��h��R�(KK��h�CX   '        '  
         L   �     \      !        C         /         �t�bhhK ��h��R�(KK8��h�C�               '     H   r     R              �        �  #  '  x     R              '              �     �              �              #  '  �     #     �     �         �t�bhhK ��h��R�(KK	��h�C$        N      �           �t�bhhK ��h��R�(KK<��h�C�      
   _         ]           �  G         ]      �     \            =
     =        �        =  D                   ]      -      �                  �        d  �     �  �  %            �t�bhhK ��h��R�(KK
��h�C(�   7   g   �        �            �t�bhhK ��h��R�(KK��h�C   �      t        �t�bhhK ��h��R�(KK��h�C0�         �   �   �                     �t�bhhK ��h��R�(KK��h�C@            %   �  �      �     �      o  �        �t�bhhK ��h��R�(KK��h�C       �
     �t�bhhK ��h��R�(KK��h�C\�   �   �     �     0        o         "              �   5   <   �  "     �t�bhhK ��h��R�(KK��h�C|*   '  a  �   �         #        �   �  %   �  �                "  �      0        �      �   "        �t�bhhK ��h��R�(KK��h�Cd   *   �      �      *   �   �   �           7   v        �   �   v	     +  �        �t�bhhK ��h��R�(KK��h�Ch   L   g         W  c            
      �                 
           P  �        �t�bhhK ��h��R�(KK
��h�C(�   w           �  7            �t�bhhK ��h��R�(KK��h�Cl      W     
               �         "  �  �        V      p  j   �        \   r      �t�bhhK ��h��R�(KK��h�C@�   �       
   #           �        �   7         �t�bhhK ��h��R�(KK��h�Cx   H   A      �   �   L   
         �   \   �           0                 '                       �t�bhhK ��h��R�(KK3��h�C�   *      $  #        �                       �  `                                           *   2      
         �  '   �  ?  V   `              %            �t�bhhK ��h��R�(KK��h�C,   y     '  �           %        �t�bhhK ��h��R�(KK��h�CP                  �                    :                     �t�bhhK ��h��R�(KK��h�CP               �  
            �                 �           �t�bhhK ��h��R�(KK��h�CL         �      '     d                       �   ]         �t�bhhK ��h��R�(KK��h�C               �t�bhhK ��h��R�(KK��h�C@'  5        >        u
  �        �     �        �t�bhhK ��h��R�(KK��h�C<�                  \            �   9            �t�bhhK ��h��R�(KK��h�C`*   �   a  �      �        "  M   $                     �     Y     "        �t�bhhK ��h��R�(KK��h�C       �        d        �t�bhhK ��h��R�(KK��h�CD   '   A      n        *   %   �   �      2   5           �t�bhhK ��h��R�(KK
��h�C(�   �      ]     q  7      r      �t�bhhK ��h��R�(KK��h�C,�  J   �   �  �     �               �t�bhhK ��h��R�(KK%��h�C��     '       L         M   �            �  �      �	  W     �                           \     
   #  '  �        �t�bhhK ��h��R�(KK��h�Ch*   '  _  �  �      _  '     \   %   �        �  _  '       �  '     c           �t�bhhK ��h��R�(KK��h�C T      '  �  �            �t�bhhK ��h��R�(KK%��h�C�   �              �   %      �                  ]            �                 �  �  �         %      J   �            �t�bhhK ��h��R�(KK��h�CL�   �     �     �         �   >     �   �                     �t�bhhK ��h��R�(KK��h�CL            :                              �   +            �t�bhhK ��h��R�(KK��h�C   �               �t�bhhK ��h��R�(KK"��h�C��   �         �      �  �                     d     u        
               �      �                      �t�bhhK ��h��R�(KK��h�C<   �         q  �               �      �        �t�bhhK ��h��R�(KK��h�C@   �   �  o     ]            b                     �t�bhhK ��h��R�(KK7��h�C�   �         �   �   �      ^     %   �      0               �   �   �   b	     �   �   (        �      %   (                    (  (     �     "  �     '  5   ]     f   �  "        �t�bhhK ��h��R�(KK/��h�C��   +     '  =     ]   �   
   �     �  =     �   +     '    g
                       �
        �   w                 �   5        ]     '           �t�bhhK ��h��R�(KK	��h�C$�   '  w  c        ]        �t�bhhK ��h��R�(KK��h�Cx                                                               �                 &        �t�bhhK ��h��R�(KK��h�C4         '                 '           �t�bhhK ��h��R�(KK��h�C4   '  	     �     '                    �t�bhhK ��h��R�(KK/��h�C�        �   �            o  �  �   �          o  �        �              I   �                  o  �        �  �
  �  �            �
  �   
        �t�bhhK ��h��R�(KK��h�C<�   �     "  )           �  8                �t�bhhK ��h��R�(KK	��h�C$�   �  I         ]           �t�bhhK ��h��R�(KK��h�CH*   �  �     �     �      �      %      �  a   �  �        �t�bhhK ��h��R�(KK	��h�C$2                           �t�bhhK ��h��R�(KK��h�C8        .              �                 �t�bhhK ��h��R�(KK��h�C`      7  �  
   $               7  �  
   8                           "     �t�bhhK ��h��R�(KK��h�C   h         b        �t�bhhK ��h��R�(KK��h�C`         �        �           �
     �   �           #   �                 �t�bhhK ��h��R�(KK��h�CH                                         i   �         �t�bhhK ��h��R�(KK2��h�C�     
                     �                 *   �      V                  V                     �                             ^     �	                    �t�bhhK ��h��R�(KK��h�Cx   �  %   �                                   �                                            �t�bhhK ��h��R�(KK��h�C4   �   �      =        �   �  '            �t�bhhK ��h��R�(KK��h�CT      "        "  �  %      �   ~     :            c               �t�bhhK ��h��R�(KK!��h�C��         
      4           �     �      �      ^              �     �   !       �            �         �t�bhhK ��h��R�(KK	��h�C$   �            �           �t�bhhK ��h��R�(KK��h�C0�      �         :   �  ]      "        �t�bhhK ��h��R�(KK��h�CT         �  '             �   g
  :         �     �              �t�bhhK ��h��R�(KK��h�Cx
   �      .   �  2   �  "     "  *   2   �	     �         �   �   "     "  *   2   �	     �   ]        �t�bhhK ��h��R�(KK��h�Cp   �   I   a  �	        o                �                     2   �           0        �t�bhhK ��h��R�(KK��h�C   C                �t�bhhK ��h��R�(KK��h�CL'  �  �      �           C        �            �            �t�bhhK ��h��R�(KK��h�C0                     �     ]        �t�bhhK ��h��R�(KK'��h�C�            �      '        `        �  L                 6  c               *  C               J                        �t�bhhK ��h��R�(KK��h�C,   �                             �t�bhhK ��h��R�(KK��h�Ct�   �                                               2            �            �            �t�bhhK ��h��R�(KK��h�CP2   5                  *        �  �  �  �                   �t�bhhK ��h��R�(KK
��h�C(            Q   #  $           �t�bhhK ��h��R�(KK��h�C<      �
  S  �          +        �           �t�bhhK ��h��R�(KK��h�C@         �  7   �     �   �
        �              �t�bhhK ��h��R�(KK��h�C\�               P     �      0   �              �  6  C      0           �t�bhhK ��h��R�(KK��h�C   �            �t�bhhK ��h��R�(KK��h�C   �  �         �     �t�bhhK ��h��R�(KK��h�CP�   �        �               '     �   B      s        N         �t�bhhK ��h��R�(KK��h�C`   9         �   '     a   �                    �   
   #        i            �t�bhhK ��h��R�(KK��h�C\      �       *      �
                 *   '        0  �   '           �t�bhhK ��h��R�(KK��h�C0C        �        �   I   �   �        �t�bhhK ��h��R�(KK
��h�C(   T      #     '        r      �t�bhhK ��h��R�(KK��h�C@   �  �  +        �                              �t�bhhK ��h��R�(KK��h�C`         �   
         �   ]                 I      �     %   i   J   �        �t�bhhK ��h��R�(KK
��h�C(�   D     \                     �t�bhhK ��h��R�(KK	��h�C$               +   "        �t�bhhK ��h��R�(KK��h�C8      W  l      
      (	                    �t�bhhK ��h��R�(KK��h�Cx      '               �     
  l  �        a     %         �     
         C   �               �t�bhhK ��h��R�(KK��h�C`'    C  y  
                  '           	                    �        �t�bhhK ��h��R�(KK��h�C]      :            �t�bhhK ��h��R�(KK��h�CL'     6     �         A                 #  %      �         �t�bhhK ��h��R�(KK��h�C\         %      W  y         6  �   ]     I  �   V      
   _               �t�bhhK ��h��R�(KK��h�CD�                           �   �   V	        �        �t�bhhK ��h��R�(KK��h�CX                  !      �         %                     L   -         �t�bhhK ��h��R�(KK��h�Ch     a                        �     2               <                     r      �t�bhhK ��h��R�(KK��h�C4�   �   [     2        �        �
        �t�bhhK ��h��R�(KK��h�C|�   �         +   *            �      �  �         j     �	              �      �      �     �        �t�bhhK ��h��R�(KK$��h�C�           �              �              �         �  �  �   a                    �     o  �  a   �           �t�bhhK ��h��R�(KK��h�CT�   �     '
  d  H   �   g
     �  /            �                     �t�bhhK ��h��R�(KK��h�CL�      %                 7            
         �  �         �t�bhhK ��h��R�(KK��h�Ch   �               A        %   �   �	  :         *   %            �     9	           �t�bhhK ��h��R�(KK��h�CX   �            �      �   +              %                           �t�bhhK ��h��R�(KK��h�C\�   '                             G                        G            �t�bhhK ��h��R�(KK��h�C,%         \   2   �   �              �t�bhhK ��h��R�(KK��h�C�            �         �t�bhhK ��h��R�(KK��h�Cp                     2                        �   7         Q         2   �   n  I         �t�bhhK ��h��R�(KK	��h�C$�                           �t�bhhK ��h��R�(KK��h�C`            p      S        %   ]  P     N   
  *      �                  �t�bhhK ��h��R�(KK%��h�C��      �     �      �   �            �      ]        t  ^  +        '        M                     '        J         �t�bhhK ��h��R�(KK��h�C          �  �  �        �t�bhhK ��h��R�(KK��h�C   �   T   r      �t�bhhK ��h��R�(KK��h�C             9   �        �t�bhhK ��h��R�(KK��h�C&   '  N      r      �t�bhhK ��h��R�(KK+��h�C�   
         2   �  
  �     �  7               \   �                 \   '              c  �     \      a                 #            �t�bhhK ��h��R�(KK��h�C`                        �            �            �            �            �t�bhhK ��h��R�(KK��h�C8   �     '  5                  '  a        �t�bhhK ��h��R�(KK��h�C   %         r      �t�bhhK ��h��R�(KK��h�C<   �  o   �              �   ^     �            �t�bhhK ��h��R�(KK��h�C�      
      b        �t�bhhK ��h��R�(KK��h�C'        :   �         �t�bhhK ��h��R�(KK��h�C@%      �     %                  :      .           �t�bhhK ��h��R�(KK��h�C,\      '     =     �       r      �t�bhhK ��h��R�(KK
��h�C('     s   	           o         �t�bhhK ��h��R�(KK ��h�C�            �           �      0                          G                    I                 �t�bhhK ��h��R�(KK��h�CtH           �   �     �  �   W  b     �  '  a          $  �      �      �      �   S         �t�bhhK ��h��R�(KK��h�C4         �            �  �   �   /         �t�bhhK ��h��R�(KK��h�C@   �   �   �     &       
        �   +     �        �t�bhhK ��h��R�(KK ��h�C�   '        G   %                 �      '  0  �  �   �      �   -      f      %         G   �  K        �t�bhhK ��h��R�(KK)��h�C�   �                             W                 Y     
   <            W  [         !         <         g   C  �              �t�bhhK ��h��R�(KK��h�C\�   �   i   W                 +        �            �      M      �
        �t�bhhK ��h��R�(KK��h�CDC                        "        "  
   �         �t�bhhK ��h��R�(KK!��h�C�   �                                    �   �        �  �           �           c                    �t�bhhK ��h��R�(KK��h�C@      �   �                 2  "      
           �t�bhhK ��h��R�(KK��h�CT              '        �   �   �     �     �        B      r      �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK
��h�C(*   q  W  (     �   c   -
        �t�bhhK ��h��R�(KK.��h�C�*   ]      =  �            =  �   �   �            0              �   �   a              
      *   '     �        �   '        �  
         !         �t�bhhK ��h��R�(KK��h�Ch           �           �   H         T   (                                       �t�bhhK ��h��R�(KK��h�C �         ]               �t�bhhK ��h��R�(KK��h�CL�         :      c  �     a      S                          �t�bhhK ��h��R�(KK��h�CT         I         '  	                    �   �                  �t�bhhK ��h��R�(KK��h�C4%   �         {                          �t�bhhK ��h��R�(KK��h�Cp�      '                        �     i                 �                             �t�bhhK ��h��R�(KK��h�Ct�   �     I   '  ]           �                          '  l  �  D	  �         C  <        �t�bhhK ��h��R�(KK��h�C   `               �t�bhhK ��h��R�(KK��h�C89      �  L                                �t�bhhK ��h��R�(KK��h�C,  �      �                        �t�bhhK ��h��R�(KK&��h�C�   ]      �                  �               �            '   �   }  w         :   A                           A           �t�bhhK ��h��R�(KK��h�C4  7   �        �   �                     �t�bhhK ��h��R�(KK��h�CT   (            /                          5  c   
   ]     r      �t�bhhK ��h��R�(KK��h�C@'  a  ]   �         �  �  y   '  r                 �t�bhhK ��h��R�(KK��h�CDV      �              @           9         �         �t�bhhK ��h��R�(KK��h�C       �   #        r      �t�bhhK ��h��R�(KK��h�C@               �   �        
     �   �	           �t�bhhK ��h��R�(KK*��h�C�                  �      
      �         R              �                                         �   H         '    �           �t�bhhK ��h��R�(KK��h�C\        �         M               �      �  R        x                 �t�bhhK ��h��R�(KK��h�C       �      a           �t�bhhK ��h��R�(KK��h�CH�         �      �                    :                  �t�bhhK ��h��R�(KK��h�C�  �            �t�bhhK ��h��R�(KK ��h�C��         �
  
   B     =                 =  �      �
        I            �         \   �               �t�bhhK ��h��R�(KK
��h�C('  �                          �t�bhhK ��h��R�(KK��h�CT+                         �                       R           �t�bhhK ��h��R�(KK!��h�C�   *   �   �  "  	  �  "        �  N   �                        �           �                          �t�bhhK ��h��R�(KK$��h�C��      `
        �   c      
            �     �         
   �  �       �         �        �         �   >            �t�bhhK ��h��R�(KK��h�C@            .      l  g                           �t�bhhK ��h��R�(KK��h�C,'  >         �          �        �t�bhhK ��h��R�(KK��h�C,�   �                            �t�bhhK ��h��R�(KK��h�CL   �     ?        �                       �     
        �t�bhhK ��h��R�(KK	��h�C$'                 i         �t�bhhK ��h��R�(KK��h�CH*      -  $      �   ]     �              `      ]        �t�bhhK ��h��R�(KK&��h�C��      �   "  `     `     �   J      M            �   J   �  *        =  �  *  �
              �   J   *  I         "        �t�bhhK ��h��R�(KK��h�Cf      �        �t�bhhK ��h��R�(KK��h�Cl�                                                         
   �        +           �t�bhhK ��h��R�(KK3��h�C�      9      '              �        *                  ]  �  
      �  $         )                  �   �  $         +       "  �   �  �
        ]       "        �t�bhhK ��h��R�(KK��h�C\         ]   �      0       �                        
      ]        �t�bhhK ��h��R�(KK��h�CD  �           �          0     �  N               �t�bhhK ��h��R�(KK��h�C8�   r         �      �       7   �      r      �t�bhhK ��h��R�(KK��h�C�           �        �t�bhhK ��h��R�(KK��h�CH   �	  �     �  _     �                 �               �t�bhhK ��h��R�(KK	��h�C$      +        a   w        �t�bhhK ��h��R�(KK��h�C8m                 j      Y                 �t�bhhK ��h��R�(KK��h�C4   �  �                                �t�bhhK ��h��R�(KK��h�CT'     �                        %         �         *  B            �t�bhhK ��h��R�(KK��h�C8�      �  �                  �     �        �t�bhhK ��h��R�(KK��h�CH�      �         �               '  �                    �t�bhhK ��h��R�(KK"��h�C�                  �      �  �     
                             �        S     (                      �t�bhhK ��h��R�(KK��h�C0   ]     �
  *   �   �  i  !           �t�bhhK ��h��R�(KK��h�C@   �  z  �   N      v           �      �  �        �t�bhhK ��h��R�(KK��h�C8      2                  ]     j            �t�bhhK ��h��R�(KK��h�C   �   %        �t�bhhK ��h��R�(KK��h�C0   �                     �           �t�bhhK ��h��R�(KK(��h�C�      5               �                     Y              '      ]                      
   $   6         �   
      A         �t�bhhK ��h��R�(KK��h�C,M         .                        �t�bhhK ��h��R�(KK��h�Cl'  �               +               �   �   �               &    
                       �t�bhhK ��h��R�(KK��h�C8      w                   �  
   ]         �t�bhhK ��h��R�(KK��h�CL�   �     �  g            '  �        w  8        @        �t�bhhK ��h��R�(KK��h�C\�            �     �     �      �               �      �                  �t�bhhK ��h��R�(KK/��h�C�                  �            ]     j         �      �                \        �            \   '           �            �
           .            �t�bhhK ��h��R�(KK��h�C@   �      ;            �         �  7   �           �t�bhhK ��h��R�(KK��h�Cp*                  �  �     �         �     �           +   +   :                        �t�bhhK ��h��R�(KK��h�C,                                  �t�bhhK ��h��R�(KK��h�CH�            �     0      V            I     
            �t�bhhK ��h��R�(KK��h�C4      �     2     �         #           �t�bhhK ��h��R�(KK��h�Cl'     D	     �     �           '  �
                 '  �     �   :   I   Y           �t�bhhK ��h��R�(KK��h�C �      '     W  �  r      �t�bhhK ��h��R�(KK��h�C '        
   y           �t�bhhK ��h��R�(KK��h�Cd   �
  �      +                 �        �
  0              I   �  �	           �t�bhhK ��h��R�(KK%��h�C�*   '  �  �               '     
            �        I	       T      T   �         >        ;      a                  �t�bhhK ��h��R�(KK��h�C4�   �      o        �     �     �         �t�bhhK ��h��R�(KK��h�CH            �  �   �  �       "  :
     �     "        �t�bhhK ��h��R�(KK��h�C      ]	  �        �t�bhhK ��h��R�(KK��h�CH
               �   �         2      �  �                �t�bhhK ��h��R�(KK��h�C,�   �     �               �        �t�bhhK ��h��R�(KK��h�C         ]  �        �t�bhhK ��h��R�(KK��h�Cl�   �     t  �  
                             T     0   +            �               �t�bhhK ��h��R�(KK��h�C         ,        �t�bhhK ��h��R�(KK	��h�C$a     �         �            �t�bhhK ��h��R�(KK��h�C8   �      %                                �t�bhhK ��h��R�(KK��h�CL      �             %      �      I   �  
                 �t�bhhK ��h��R�(KK��h�C0   _     �     �      �      7         �t�bhhK ��h��R�(KK
��h�C(�   �  �   �   j                  �t�bhhK ��h��R�(KK��h�C<"           �   �          \        r   "     �t�bhhK ��h��R�(KK��h�CH      �  �        s   l         �   �      �               �t�bhhK ��h��R�(KK��h�Ch�   �  "        �   $  �     �   �                                %         "     �t�bhhK ��h��R�(KK��h�C   #  r      �t�bhhK ��h��R�(KK��h�CD         a   I   �  :   I   �      0  �                  �t�bhhK ��h��R�(KK��h�CP         '  H                  (         6  �      V            �t�bhhK ��h��R�(KK
��h�C('                    �        �t�bhhK ��h��R�(KK��h�CP+     w     �
  
            �         �      �                  �t�bhhK ��h��R�(KK��h�C@            n     �   �           �              �t�bhhK ��h��R�(KK	��h�C$              +   w         �t�bhhK ��h��R�(KK ��h�C�                    �      o          �      �                       �     �  �   l      n        �t�bhhK ��h��R�(KK	��h�C$   �        �               �t�bhhK ��h��R�(KK��h�C              j            �t�bhhK ��h��R�(KK��h�C|                       V         �            �   �  w  6  �   �  I   A      �   D     5           �t�bhhK ��h��R�(KK��h�C    �        0           �t�bhhK ��h��R�(KK��h�C0            �     '     
   �         �t�bhhK ��h��R�(KK��h�C@      �  a      �  "     "     j   "        "     �t�bhhK ��h��R�(KK��h�Co    5   �            �t�bhhK ��h��R�(KK��h�C	        �t�bhhK ��h��R�(KK��h�C                    �t�bhhK ��h��R�(KK
��h�C(�   �              �            �t�bhhK ��h��R�(KK��h�C4�     /      �           �  
   �
        �t�bhhK ��h��R�(KK��h�C�   �         Z        �t�bhhK ��h��R�(KK��h�CL      �                                                  �t�bhhK ��h��R�(KK	��h�C$%   �      N   �  ^            �t�bhhK ��h��R�(KK��h�C0            
         �              �t�bhhK ��h��R�(KK��h�C@�   �           5  ]           �   �  *           �t�bhhK ��h��R�(KK$��h�C�%                  
                  %           )            �        �   �   �              �                  �t�bhhK ��h��R�(KK��h�C@       �            �
           �     �   -         �t�bhhK ��h��R�(KK��h�C4'  5               *  ]      �
  �         �t�bhhK ��h��R�(KK(��h�C��      '     0         c   :         �               
   �      
           �            �      �  D  #  '  T   �      0   ^        �t�bhhK ��h��R�(KK��h�C@o                   ]  �                 r      �t�bhhK ��h��R�(KK��h�C<'  �   
     �   �     �  �     �      V        �t�bhhK ��h��R�(KK��h�C0   �
                    �           �t�bhhK ��h��R�(KK��h�C@]  V  �	                   �   
                 �t�bhhK ��h��R�(KK��h�CP            
   #     �  *         C    O                     �t�bhhK ��h��R�(KK	��h�C$            .  
            �t�bhhK ��h��R�(KK��h�C\         4	         �         �           �      #      "  �         �     �t�bhhK ��h��R�(KK��h�C%                  �t�bhhK ��h��R�(KK"��h�C�         Y              %         +      �      �            �        $         �   �     �                  �t�bhhK ��h��R�(KK(��h�C�   '     =  �     �   �     =                    
                    �        (   M   �      S     �         a  C            �t�bhhK ��h��R�(KK4��h�CК      '   i  ?  V   2     �      %   �  �                 �            �  �     �                    �      _     C      0  z                          �   �        �t�bhhK ��h��R�(KK��h�C4'        �        P  <                 �t�bhhK ��h��R�(KK��h�C   �         �        �t�bhhK ��h��R�(KK��h�CD%   (   +      v   #         �           
   C           �t�bhhK ��h��R�(KK��h�C0]           
   �
  =  �               �t�bhhK ��h��R�(KK��h�CL     �  �              a         �  C  {   "   T           �t�bhhK ��h��R�(KK ��h�C�            9         "        '     
                  '                 _     :      �  r   "     �t�bhhK ��h��R�(KK��h�C'  5               �t�bhhK ��h��R�(KK-��h�C�               w              9  �                       �                                        V   %         �        E  :            �t�bhhK ��h��R�(KK��h�Cp         5   '  I   �   �     �           S  j               �   �               �         �t�bhhK ��h��R�(KK��h�C,   �  %         `     `  `  �     �t�bhhK ��h��R�(KK
��h�C(      '      �                 �t�bhhK ��h��R�(KK��h�Cty  g               '    +        !                 �  �      �  �  �  n     7   �        �t�bhhK ��h��R�(KK��h�C0         �	        '  	              �t�bhhK ��h��R�(KK��h�CX'  �           �   '              o  =  :
  �                       �t�bhhK ��h��R�(KK��h�C4   7   �     '     #     �              �t�bhhK ��h��R�(KK��h�Cx   '  a  �   ]  �  �         '  a              �   �        g     #   �  \   %                  �t�bhhK ��h��R�(KK��h�C�      �           �t�bhhK ��h��R�(KK��h�C<   :     �      �            �   i        r      �t�bhhK ��h��R�(KK��h�C   ]                 �t�bhhK ��h��R�(KK ��h�C�   '  �   �     �                   %      	  �   �           C  /            %   (   7     G        �t�bhhK ��h��R�(KK��h�C<         �            +           �            �t�bhhK ��h��R�(KK!��h�C�         �     �  �     )         �  �     �      �               N            �   c   �                 �t�bhhK ��h��R�(KK��h�C   �               �t�bhhK ��h��R�(KK%��h�C��         �              �     s        #  �        �   q     
      :           "     �      #  �     �
  "        �t�bhhK ��h��R�(KK��h�Cp         '     &      0         �     �     �  �  �  �      �   
                        �t�bhhK ��h��R�(KK��h�Ct         �      1                         G             %   �                         �t�bhhK ��h��R�(KK	��h�C$         �     �            �t�bhhK ��h��R�(KK*��h�C��  '  �                        B  �           �   :      6        �  '     �   T   %      %         �        '        �  �  �  r      �t�bhhK ��h��R�(KK��h�C0         �         �     �
  �         �t�bhhK ��h��R�(KK��h�C4�                  0                    �t�bhhK ��h��R�(KK��h�C       �   �               �t�bhhK ��h��R�(KK��h�CP      +  r      a        �   �                  *   %            �t�bhhK ��h��R�(KK	��h�C$      ]                    �t�bhhK ��h��R�(KK��h�C@�   2              b
        \   H   �     �        �t�bhhK ��h��R�(KK��h�C   �     �   �	        �t�bhhK ��h��R�(KK&��h�C�   �   D           '   �      *      $           i        /   
   �           K                          �              �t�bhhK ��h��R�(KK%��h�C��   '  D     %   ]                 �      #   �            ]        #      �      %      �              �              �t�bhhK ��h��R�(KK	��h�C$  �
  6  �  �   �   �        �t�bhhK ��h��R�(KK��h�CT�           �  o     i   `     '     �        #     �  ]         �t�bhhK ��h��R�(KK��h�C,%         �	  y   %      �           �t�bhhK ��h��R�(KK��h�C4�   A	     �        
        �            �t�bhhK ��h��R�(KK��h�C<              c                     �        �t�bhhK ��h��R�(KK��h�C\     �      �                  �         �  Z                 �  r      �t�bhhK ��h��R�(KK3��h�C�)      '        #  �      a     �            >   '  �  0      
                              �   �              '  �         �       �                  �         �t�bhhK ��h��R�(KK��h�Ch'  &   �   ]   
                    '                             �
              �t�bhhK ��h��R�(KK��h�CD%      
   _         f   o   h        �         �        �t�bhhK ��h��R�(KK
��h�C(   �              '  �        �t�bhhK ��h��R�(KK��h�CT            �                  0         J  C   �   �  '           �t�bhhK ��h��R�(KK
��h�C(      �     L   �              �t�bhhK ��h��R�(KK��h�C8*   �                  �      �               �t�bhhK ��h��R�(KK��h�Cx            a              "        c      :               �     �         =                 �t�bhhK ��h��R�(KK
��h�C(   �        %      �   �        �t�bhhK ��h��R�(KK��h�C4�   s   �        ]           G   �
        �t�bhhK ��h��R�(KK��h�CD�         '  >   �  �                     Y           �t�bhhK ��h��R�(KK5��h�C�   C        C         y   %   �  �                        Q   =     �   D    =  y   %   �     �     %            &           �   �              �     D  :               �t�bhhK ��h��R�(KK��h�CT%      I   �            �      %   u
     g         C      ;   �        �t�bhhK ��h��R�(KK(��h�C��   �     o        �  c                        P           '                                �      "      �                  �t�bhhK ��h��R�(KK��h�C@               '        (      �                  �t�bhhK ��h��R�(KK��h�Cp   2   �   �         %            .      �      I              %            �      t        �t�bhhK ��h��R�(KK��h�C4   �      �               W              �t�bhhK ��h��R�(KK��h�C8   �   �         >   �  �      
   �           �t�bhhK ��h��R�(KK��h�C|R           '                          c   �   �           '  ?   ;         '     O     "        �t�bhhK ��h��R�(KK��h�Ct�   w  M   ^     d  
                 <      �   N   
   �   �           d  M   �
  �  w         �t�bhhK ��h��R�(KK��h�C<�           "              c          "        �t�bhhK ��h��R�(KK��h�CT         �      "  �                    �   �  �
     �	  "        �t�bhhK ��h��R�(KK ��h�C��   �  V     #     s   0  B   ?     �
  w      �   �           '     o  E                    �        �t�bhhK ��h��R�(KK��h�C<*      W  c   :      �  �         �     C         �t�bhhK ��h��R�(KK,��h�C��                  �   P  7            %      o     -   Y  V      �  9   
                        �           '         M        C           �t�bhhK ��h��R�(KK(��h�C�   W  Q         �  @	     '  *  
      �  '     *  
      �            �  '     *  
      =  �   �     �     �  '     �         �t�bhhK ��h��R�(KK��h�C0               �  �   7            �t�bhhK ��h��R�(KK��h�Cd        -      d  
                 �     
                  6     �        �t�bhhK ��h��R�(KK��h�CL'     i   �   �  �             �                  
        �t�bhhK ��h��R�(KK��h�C    �     '              �t�bhhK ��h��R�(KK��h�C<   o        h   �        "           "        �t�bhhK ��h��R�(KK��h�C8�                              S      \     �t�bhhK ��h��R�(KK	��h�C$2   5      6     w  
        �t�bhhK ��h��R�(KK	��h�C$   '     J      ]   �  r      �t�bhhK ��h��R�(KK��h�C\     u  =       u                    �   Q      �                     �t�bhhK ��h��R�(KK��h�C,     �   �
  �           v	  r      �t�bhhK ��h��R�(KK��h�C<�   5         ]  �  "        "  �   5            �t�bhhK ��h��R�(KK��h�C8      �   �   O     W	     %         
         �t�bhhK ��h��R�(KK��h�CD   �  �        �      �        S                    �t�bhhK ��h��R�(KK��h�C,            %   .                 �t�bhhK ��h��R�(KK,��h�C��   *   �      #                       o            �  �   �                                      #   i         �     N      	  �            �t�bhhK ��h��R�(KK)��h�C��   '  >   �  �  �  b       \   (   '                 �           �            %      ;                     �  �	  :         �  r      �t�bhhK ��h��R�(KK.��h�C�'  D     .      :   �     #              %         �            �     �              N            �      �                                      �t�bhhK ��h��R�(KK��h�C,*  �  
   %   ]                    �t�bhhK ��h��R�(KK��h�C�               r      �t�bhhK ��h��R�(KK��h�CT   �      �     $     I   =  '     �  �	     �  
      ]  �	        �t�bhhK ��h��R�(KK1��h�CĚ      �         �   �     �
        �   �     �            o     �            �         �        P                       #  %   �     I   �                 �t�bhhK ��h��R�(KK.��h�C�         �     "  �           "              �  g      2   �        *      �  W        c         �  /   :   �	        C  N           C           �t�bhhK ��h��R�(KK��h�C\o     w            �         �   w         o  �               �   �         �t�bhhK ��h��R�(KK��h�C,   	        �  #      #            �t�bhhK ��h��R�(KK��h�CTV   '   �  �        %   �     (  �           &   �  �     �         �t�bhhK ��h��R�(KK��h�C,      �  J        �  �  �        �t�bhhK ��h��R�(KK��h�C0�   D     "     �   D  #     P        �t�bhhK ��h��R�(KK	��h�C$`               �   �        �t�bhhK ��h��R�(KK
��h�C(                              �t�bhhK ��h��R�(KK
��h�C(                  (            �t�bhhK ��h��R�(KK��h�CD              �   �  c         ]        c           �t�bhhK ��h��R�(KK��h�Ct      '        L         
                              
        �     T                  �t�bhhK ��h��R�(KK��h�C<�   %      )   g      %      C         �            �t�bhhK ��h��R�(KK��h�Ct]      C   N   �      W  7   �  T            �
  �  P           �
  �        �  4              �t�bhhK ��h��R�(KK#��h�C�+  "        "        �         �         �                  �  c   �                    �   �   +              �t�bhhK ��h��R�(KK��h�C@%                        �           �            �t�bhhK ��h��R�(KK��h�C�  w     W           �t�bhhK ��h��R�(KK<��h�C�]     �               �               :                           :         �               '        '  �   �         `        '  >   a   =  '     =  '  >   a         w        
      �        �t�bhhK ��h��R�(KK	��h�C$�            �               �t�bhhK ��h��R�(KK ��h�C�   �         *        g         >      *           8   �            �  �     �        d              �t�bhhK ��h��R�(KK��h�C@      �   9   z             �  
   m              �t�bhhK ��h��R�(KK��h�CT         �  *                  s            a  +      �           �t�bhhK ��h��R�(KK��h�C0�   ?  :               #              �t�bhhK ��h��R�(KK��h�C0                                   �t�bhhK ��h��R�(KK#��h�C�   �            �        b
          9            �   �                 	  �  h         �        �            �t�bhhK ��h��R�(KK��h�C@�                  7            ]                 �t�bhhK ��h��R�(KK"��h�C�      A            �        L                             '     �      �              �     9            �t�bhhK ��h��R�(KK��h�CP"                       
   �  =              �     r   "     �t�bhhK ��h��R�(KK��h�Cd   �         �               Q               :   I   �
       �   �  �   �         �t�bhhK ��h��R�(KK ��h�C��         �      �      �  '  �     �          �                 *     '     �  
   Y              �t�bhhK ��h��R�(KK��h�C`]   �                           �   �              �      �                 �t�bhhK ��h��R�(KK��h�CL   '                        �   �   �     �  o              �t�bhhK ��h��R�(KK
��h�C(   �
     %                     �t�bhhK ��h��R�(KK��h�C`�   �           '   �   #      i                  �                           �t�be.