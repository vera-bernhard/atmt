minska (1/1)
möter (1/1)
Skatteförvaltningen (4/5) skatteförvaltningen (1)
grundskolor (4/4)
mataffärer (1/1)
inriktade (3/3)
tillbringa (1/1)
Kannus (1/1)
säga (23/23)
minskar (3/3)
Vanttauskoski (1/1)
speciellt (9/9)
utgångsläge (1/1)
ungdomen (1/1)
sina (57/57)
arbetsintyg (12/14) Arbetsintyg (2)
andelar (1/1)
varar (20/20)
företagarpensionsförsäkringenfinska (1/1)
närmare (13/13)
gammal (13/13)
affärsresa (1/1)
linkkiFörsamlingen (1/1)
energibesparingslampor (1/1)
barndom (1/1)
tas (23/23)
tilläggsdagar (1/1)
työttömyyskorvaus (2/2)
motarbeta (3/3)
människovärdet (1/1)
ting (3/3)
konst- (1/1)
översättningen (4/4)
Opintopolku.fi (3/3)
verksamheten (14/14)
elbolaget (1/1)
polisanmälan (1/1)
föräldrapenningperioden (3/3)
uppehållskort (5/5)
II (1/1)
allmän (8/9) Allmän (1)
skriver (11/11)
stadsrättigheter (1/1)
tandvården (6/6)
beskriver (5/5)
skattepengarna (1/1)
montera (1/1)
kuvataidekoulu (1/1)
vanhempainvapaa (1/1)
räntestödetfinska (1/1)
negativt (4/5) Negativt (1)
inkomstgräns (1/1)
nationalpark (2/2)
festivaler (1/1)
så (63/63)
födelsen (1/1)
berättelse (1/1)
maistraatti (16/16)
kaffesump (1/1)
kaffe (1/1)
avoin (7/7)
ålderspensionen (3/3)
bokat (4/4)
kulturstad (1/1)
akut (22/22)
webbplatser (13/13)
affärer (1/1)
registrering (20/29) Registrering (9)
fastighetsskötseln (3/3)
biljettjänstens (1/1)
sed (2/2)
egenskaper (1/1)
blanketter (1/1)
idrottsväsendet (1/1)
kuntoutuspsykoterapia (1/1)
bosättningsbaserade (1/1)
asumisoikeussopimus (1/1)
situationerna (1/1)
Migrationsverketfinska (1/1)
bokad (1/1)
felfri (1/1)
innevarande (1/1)
upphörande (2/2)
buddhism (1/1)
minipiller (1/1)
arbetsoförmåga (1/1)
föregår (1/1)
presenter (2/2)
identifieras (1/1)
heminkvartering (1/1)
oppisopimuskoulutus (1/1)
distansgymnasiet (1/1)
budskap (1/1)
återvinningsstationer (1/1)
dyra (6/6)
utgift (1/1)
pensionspremierna (1/1)
arbetarskyddschef (1/1)
planerar (10/10)
yrkesutbildningen (1/1)
ämbetsverk (1/1)
hurdan (2/2)
drogmissbruk (1/1)
handikappidrott (1/1)
personlig (8/8)
ansluta (10/10)
stulits (1/1)
tidtabellerfinska (1/1)
legaliserat (2/2)
familjeärenden (2/2)
framföra (2/2)
tillgångarna (1/1)
mobiltelefontillverkaren (1/1)
meddelanden (1/1)
planerad (1/1)
oväsen (1/1)
läckaget (1/1)
rådgivningens (1/1)
föräldramöten (2/2)
hälsovårdscentralen (7/7)
blombukett (1/1)
institut (6/6)
samtala (2/2)
hemtjänster (1/1)
livsmiljö (1/1)
ansöker (72/72)
trossamfund (5/5)
3D (1/1)
ses (1/1)
dig (368/368)
familjecentret (4/4)
bedriver (5/5)
läcker (1/1)
köping (1/1)
parkgympa (1/1)
problemet (1/1)
strävar (3/3)
osaomistusasunto (2/2)
Vanhemman (2/2)
skyddshem (15/18) Skyddshem (3)
bevara (2/2)
ungdomsgårdar (5/5)
fortsättningsvis (1/1)
honom (3/3)
toimisto.fi (1/1)
kunskapscenter (1/1)
vårens (1/1)
samtidigt (25/25)
ämnar (2/2)
tukiverkko (1/1)
underhålla (1/1)
nordiska (13/13)
senast (25/25)
flytten (7/7)
därför (5/5)
rasism (4/4)
bifogas (1/1)
hobbyklubbar (1/1)
flyttningsdagen (1/1)
Lumon (2/2)
ju (1/1)
undervisning (43/43)
HRT:s (2/2)
högskolestuderandefinska (1/1)
barnmorska (1/1)
reservationsavgifter (1/1)
moderskapspenningperiodens (1/1)
het (1/1)
uppsikt (3/3)
hamnat (2/2)
försenad (2/2)
finländsk (18/18)
verksamhetsplanen (1/1)
förhistoria (1/1)
Sovjetunionen (8/8)
företagande (12/12)
data- (1/1)
församlingarfinska (1/1)
flyttades (2/2)
tilltalar (1/1)
sammanlagda (2/2)
pensionsskyddet (2/2)
arbetsförmögen (1/1)
väst- (2/2)
helt (5/5)
problem (83/90) Problem (7)
Brottsofferjouren (4/5) brottsofferjouren (1)
pappor (1/1)
antagen (4/4)
utkommer (3/3)
middag (1/1)
administrativa (2/2)
utbildningslinjer (1/1)
Metropolia (1/1)
medling (6/6)
köpt (3/3)
bostadsansökan (3/3)
nödinkvartering (2/2)
fostret (1/1)
inleda (3/3)
CC (1/1)
familjfinska (1/1)
eventuella (7/7)
parkeringsavgiften (1/1)
intresseorganisationfinska (1/1)
tiotals (1/1)
regioner (1/1)
utvecklar (2/2)
markområden (1/1)
samlaget (1/1)
sosiaalipäivystys (1/1)
har (1057/1057)
slidmynningen (1/1)
progressivt (1/1)
hälsovårdarens (3/3)
vuxenutbildningsstöd (1/1)
fostrets (2/2)
SERI (2/2)
bosättningsort (1/1)
acceptansen (1/1)
tillverkas (2/2)
domstol (2/2)
Hanhikivi (1/1)
överenskommen (1/1)
Utbildningsstyrelsens (13/17) utbildningsstyrelsens (4)
handelskammare (2/2)
vaccineras (1/1)
kvinna (3/3)
närmaste (20/20)
förtrogen (1/1)
sjukskötarens (2/2)
resehandling (2/2)
Europaparlamentsvalet (1/1)
resekorten (1/1)
webbtjänsten (7/7)
pensioner (2/2)
mete (1/1)
förändring (1/1)
samkommunen (3/3)
elbolag (1/1)
tung (1/1)
advokatförbundfinska (1/1)
ehkäisyneuvola (1/1)
sönder (1/1)
työehtosopimukset (1/1)
tidskriften (1/1)
elbolags (1/1)
parken (1/1)
turvallisuusvirasto (1/1)
styrka (9/9)
servicepunkterna (1/1)
planer (1/1)
arbetspensionssystemet (1/1)
inbringar (2/2)
elektriska (2/2)
åtföljs (2/2)
pensionstagare (3/3)
intersexuella (1/1)
Nokia (1/1)
boendemöjligheter (1/1)
bokar (11/11)
avdragsgill (2/2)
freden (1/1)
konsulat (3/3)
litauiska (1/1)
lokaler (7/7)
köket (1/1)
kontaktspråket (1/1)
billigare (2/2)
butiken (1/1)
is (1/1)
tandvårdsjourenfinska (1/1)
idag (2/2)
underhåller (1/1)
somaliska (46/46)
slott (4/4)
tjänsteleverantörers (1/1)
utbildningen (53/53)
härkomst (4/4)
börjat (3/3)
varierande (1/1)
yta (1/1)
studiestödetfinska (1/1)
yrkeshögskolorna (2/2)
personerfinska (1/1)
tidtabellen (1/1)
nationer (1/1)
varat (5/5)
kursstart (1/1)
Pejas (2/2)
småbarnspedagogik (11/11)
Omena (4/4)
flickorfinska (2/2)
utsätta (1/1)
reseplaneraren (3/5) Reseplaneraren (2)
äktenskapsförord (4/5) Äktenskapsförord (1)
distansstudier (1/1)
Helsingforsregionen (5/5)
delägarbostadfinska (2/2)
studieplaner (1/1)
teatrar (4/4)
gardet (1/1)
Företagarna (1/1)
entrédörren (2/2)
gymnasiestudierna (2/2)
högklassiga (1/1)
deltagarna (1/1)
medelstora (1/1)
B (7/7)
inverka (1/1)
svenskspråkiga (10/10)
underhållsskyldigafinska (1/1)
bassjälvrisken (1/1)
stavelsen (1/1)
församlingen (1/1)
F (1/1)
tidsbunden (2/2)
arbetarskyddsfrågor (1/1)
nås (2/2)
resan (2/2)
verksamhetsstället (1/1)
trygghetfinska (1/1)
juni (9/9)
familjerna (1/1)
bedömning (6/6)
vintersporterna (1/1)
applikationer (1/1)
anarki (2/2)
idrottssällskap (2/2)
olika (179/179)
sjukhuskostnaderna (1/1)
skyldigheterna (2/2)
film (4/4)
närståendevårdare (1/1)
beter (2/2)
finansieringsvederlag (1/1)
dags (1/1)
flyttsakerna (1/1)
badar (4/4)
ansökanfinska (2/2)
flyttanmälan (3/3)
sittunderlag (1/1)
kortet (8/8)
medborgarnas (2/2)
akademiskt (1/1)
blankett (15/15)
mångkulturellt (2/2)
utanför (17/17)
semesterna (1/1)
Marthaförbundet (1/1)
nivå (7/7)
rättsbiträde (3/3)
karriärmentorskap (1/1)
studievägledarna (2/2)
respekteras (1/1)
registerstryrelsen (1/1)
ägodelarna (1/1)
sön (2/2)
kommunalskatt (1/1)
ungdomsgården (2/3) Ungdomsgården (1)
appen (2/2)
Näringsliv (3/3)
gymnasiumfinska (1/1)
fyllas (1/1)
prepositioner (1/1)
inflyttningen (2/2)
alkohol (6/6)
dagarna (1/1)
rehabiliteringsstöd (1/1)
medium (1/1)
chef (8/8)
pauser (2/2)
statliga (9/9)
flaggar (1/1)
pensionsanstalten (1/1)
identiska (3/3)
kreditupplysningsregistret (2/2)
självrisktid (2/2)
förtjänade (1/1)
-stiftelser (1/1)
undersida (1/1)
högst (37/37)
albanska (7/7)
norska (9/9)
varav (6/6)
seger (1/1)
universitet (43/48) Universitet (5)
övningsskola (1/1)
vandrarhem (1/1)
fisk (1/1)
examensnivån (1/1)
kesäteatterifinska (1/1)
Handikappforums (1/1)
drogs (1/1)
läroanstaltens (2/2)
kondylom (1/1)
avtog (1/1)
del (65/65)
firas (11/11)
genus (1/1)
perheneuvonta (1/1)
skattebyrå (3/3)
äktenskapshinder (6/6)
månaderna (5/5)
individualism (1/1)
hösten (9/9)
makar (2/2)
upphovsmannen (1/1)
privat (46/46)
sjukförsäkring (8/8)
nyheter (2/2)
språketfinska (6/6)
joggingbanor (1/1)
parten (3/3)
hämta (6/6)
kortvarigt (1/1)
företagarhandböcker (1/1)
bokföringen (6/6)
Mona (4/4)
redan (30/30)
simpass (1/1)
angett (1/1)
giltig (2/2)
yrken (11/11)
familjeförhållanden (4/4)
tillståndstjänstenfinska (1/1)
förekommer (2/2)
sosiaaliohjaaja (1/1)
Yle (1/1)
utställningarfinska (1/1)
elapparat (2/2)
insjuknandet (4/4)
avtalsperioden (1/1)
stödbostad (3/3)
radhuslägenheter (1/1)
barnskyddets (2/2)
utrikespolitik (1/1)
apoteket (8/8)
campingområdenfinska (1/1)
bemärkelsedagar (1/1)
kräva (10/10)
fritid (4/5) Fritid (1)
sambon (4/4)
Infopankki.fi (1/1)
Kitfinska (1/1)
bolagsmän (1/1)
tobaksprodukter (1/1)
hälsostationsläkaren (1/1)
förhandlare (1/1)
hitar (2/2)
stationen (1/1)
barndomen (1/1)
kontinuerliga (3/3)
spisen (4/4)
anmäl (2/2)
sök (1/1)
utbildningarfinska (2/2)
lyfter (1/1)
bostadslösafinska (2/2)
heltid (8/8)
AA (2/2)
föräldrapenning (3/3)
försäkringsbolag (11/11)
beskattningsbara (3/3)
hyresbeloppet (1/1)
sommaruniversitetet (2/2)
påverkar (14/14)
folks (1/1)
skyddsåldersgränsen (1/1)
slutliga (3/3)
PISA (1/1)
Infobanken (5/5)
nämn (1/1)
budget (1/1)
erbjudande (1/1)
skolgången (2/2)
läroplikt (3/3)
frånvaron (1/1)
hänt (1/1)
tron (2/2)
vårdkostnadsförsäkring (1/1)
bussbiljetter (1/1)
bl.a. (7/7)
övriga (28/28)
skrivfärdigheter (1/1)
pensionssystemen (1/1)
polisen (18/19) Polisen (1)
cykla (4/4)
förpackningsmaterial (1/1)
frivilligarbete (5/6) Frivilligarbete (1)
specialyrkesläroanstalter (1/1)
organen (1/1)
utesluta (1/1)
Asuntosäätiös (1/1)
körkortfinska (1/1)
återvänder (3/3)
pepparkakor (1/1)
ända (3/3)
polisens (8/9) Polisens (1)
lähityön (1/1)
verohallinto (1/1)
erkänns (1/1)
upplösande (1/1)
riksdagsval (2/2)
Muurola (1/1)
växelvis (1/1)
trafikförbindelser (1/1)
blåser (1/1)
pappersformulär (1/1)
asunnotfinska (1/1)
taget (3/3)
logi (1/1)
intresserade (6/6)
barnskötare (3/3)
förtagaren (1/1)
uppsägning (4/4)
gånger (13/13)
försäkrad (3/3)
kapital (2/2)
friska (1/1)
rättshjälpsbyrå (10/10)
medlemskortetfinska (1/1)
socialmyndigheters (1/1)
upphävande (1/1)
arbetslösafinska (3/3)
organiserade (1/1)
integrationsutbildning (5/5)
servicesedlar (1/1)
polisstationernafinska (1/1)
fötts (3/3)
företagarutbildningar (1/1)
arbetslösfinska (1/1)
Myrkytystietokeskus (1/1)
avbokat (1/1)
kistor (1/1)
rådgivningsbyråerna (3/3)
herpes (1/1)
beviljar (4/4)
identifierats (1/1)
förhållandet (1/1)
relativt (4/4)
uppfostrande (1/1)
köra (6/6)
placera (2/2)
alkukartoitus (2/2)
medlingen (1/1)
kinesiska (36/36)
vill (149/149)
skadan (2/2)
problemen (1/1)
växlande (1/1)
post (32/32)
regionförvaltningsverk (1/1)
anmälas (5/5)
B1 (2/2)
länderna (18/18)
brottmål (3/3)
arbetslöshetskassor (1/1)
föräldradagpenningens (1/1)
vuxenutbildning (8/8)
teckenspråkstolk (1/1)
byråerna (1/1)
lever (4/4)
arbetarskyddsinspektioner (1/1)
tillståndsansökan (4/4)
språkanvändares (2/2)
-Förbundet (1/1)
arbetstiderna (1/1)
pensionsåldern (1/1)
utfärdats (10/10)
Monikas (1/1)
bankonto (1/1)
motionsspår (1/1)
studentrabatter (1/1)
bolagsmannen (1/1)
bruksvederlag (3/3)
Karlebynejdens (2/2)
tionde (5/5)
barnrådgivningsbyrån (1/1)
undervisningstillstånd (1/1)
underlivet (1/1)
placeras (1/1)
domstolen (4/4)
vigseltillfället (1/1)
personers (3/3)
hälsomotionskalendern (1/1)
antecknar (1/1)
kyrka (5/5)
brottfinska (1/1)
Yrkenas (1/1)
välhållen (1/1)
öppettiderfinska (2/2)
filmens (1/1)
insjöarna (1/1)
Sporttikortti (1/1)
telefontjänst (11/11)
studiestödetengelska (1/1)
förälderns (3/3)
noll (1/1)
meneefinska (1/1)
bedömningsgrunder (1/1)
yrkeskunskaper (2/2)
arbetstillstånd (1/1)
tilläggsinformation (1/1)
Terveyden (1/1)
gravkvarter (1/1)
Veikko (1/1)
visas (5/5)
platsen (1/1)
hälsovårdsbranschen (1/1)
beviljandet (1/1)
tillhandahålla (2/2)
integrationsplanfinska (1/1)
barnrådgivning (1/1)
kirkko (2/2)
handelsregistret (2/2)
närskola (3/3)
ärekränkning (1/1)
läs- (1/1)
ut (113/113)
precis (2/2)
dröjsmålsränta (1/1)
förskottsuppbördsregistret (2/2)
bidrag (11/11)
myndigheter (35/35)
hushållsapparater (1/1)
att (1223/1233) Att (10)
lokaltidningar (2/2)
självfinska (2/2)
intervju (1/1)
motsätter (2/2)
ansökningsproceduren (1/1)
senioruniversitetet (2/2)
Kuntien (1/1)
fyllde (1/1)
praktiknära (2/2)
bostadsägaren (2/2)
väljs (12/12)
toimintakeskus (1/1)
mammor (1/1)
barnfinska (7/7)
genomför (1/1)
antagningen (1/1)
religionsfrihet (2/2)
mamma- (1/1)
Lichtenstein (1/1)
längs (1/1)
vandra (1/1)
påverkan (5/5)
värmesystem (1/1)
mångsidigt (1/1)
förlossningen (18/18)
förarutbildning (1/1)
allmäneuropeisk (1/1)
förpackningar (3/3)
bruksvederlaget (2/2)
elden (1/1)
inredning (1/1)
nytta (5/5)
motiverat (1/1)
ammatti- (3/3)
framhäver (1/1)
bank (4/5) Bank (1)
privatvårdsstöd (2/2)
myndiga (2/2)
vidtar (1/1)
utreds (4/4)
hindersprövningen (6/6)
beskriva (1/1)
frukter (1/1)
medborgares (7/7)
Alberga (1/1)
konfidentiellt (3/3)
nio (5/5)
veronumero (2/2)
föräldrapenningsperioden (1/1)
berätta (5/5)
tusentals (2/2)
självständiga (3/3)
överhuvudtaget (1/1)
kärnkompetens (2/2)
betalningsstörningfinska (1/1)
Gammelstadsforsen (1/1)
hyressed (1/1)
flyttningen (3/3)
avdragen (1/1)
dagvårdsstart (1/1)
friluftsmuseum (1/1)
persons (3/3)
medeltida (1/1)
gåvor (1/1)
utvecklingsstadium (1/1)
arbetslöshetsstöd (1/1)
utrikesflygen (1/1)
handlingarna (3/3)
familjeplanering (5/5)
nyttig (8/8)
Fennovoimas (1/1)
potilasasiamies (2/2)
nättjänsten (2/2)
esteiden (3/3)
karta (1/1)
samhällsvetenskaper (2/2)
hälsovårdsenhet (1/1)
skrapning (2/2)
Esbos (1/1)
sommargymnasium (1/1)
skuldfria (1/1)
Mina (4/4)
arbetslöshetsförmån (7/7)
informationen (6/6)
orolig (2/2)
hemvist (2/2)
legaliserad (2/2)
ordnas (81/81)
bedöma (3/3)
skolkuratorn (2/2)
programmet (1/1)
levnadskostnaderna (1/1)
paret (2/2)
ärlighet (3/3)
lagman (1/1)
bakgrund (5/5)
väster (2/2)
byggs (1/1)
kollektivtrafikens (5/5)
kansalaisen (1/1)
avsedd (39/39)
plast (1/1)
hätänumero (2/2)
juridiskt (2/2)
ersatts (1/1)
sammanställts (1/1)
blödningar (3/3)
yrkeshögskolestudier (1/1)
behandlingen (7/7)
CVfinska (2/2)
försörjningen (4/4)
hälsovårdsstiftelses (1/1)
lärande (4/4)
bolaget (1/1)
istiden (1/1)
deltidsarbeta (1/1)
bemött (1/1)
missnöjd (1/1)
motionsform (1/1)
åsikter (3/3)
synnerhet (1/1)
bolsjevikregeringen (1/1)
utvecklingsstörningar (1/1)
väldigt (4/4)
ingå (10/10)
gravida (8/8)
sammanträden (3/3)
förvaltas (1/1)
krisen (1/1)
näringsministeriet (8/8)
diskussioner (2/2)
avlägger (10/10)
med (667/667)
anledningarna (1/1)
telefonnummer (8/8)
giftorätten (1/1)
palvelu (1/1)
MIELI (2/2)
publicus (2/2)
brandvarnare (6/6)
samtals- (1/1)
bolagets (1/1)
sysslorna (3/3)
kallelsen (1/1)
privatläkare (4/4)
försäljningsmetoder (1/1)
1500kt (1/1)
lyckas (1/1)
må (1/1)
hotar (9/9)
studerandeengelska (1/1)
barnfamiljer (7/7)
grupperna (1/1)
häradsskrivare (1/1)
öppettider (8/8)
Jesusbarnet (1/1)
lika (15/15)
invandrarkunder (1/1)
uppgifterfinska (1/1)
Vantaan (10/10)
vädra (1/1)
Kvinnokliniken (1/1)
självständighetens (1/1)
försörjningsförutsättningen (2/2)
minderårig (2/2)
bekymrar (1/1)
tillsvidareanställning (1/1)
testamentsgåva (1/1)
inkomsten (2/2)
hälsopunkterfinska (1/1)
kyrkoherden (1/1)
krama (1/1)
pensionering (1/1)
får (399/399)
ytmaterial (1/1)
kvalifikationer (4/4)
beordra (1/1)
arbetsgivarens (4/6) Arbetsgivarens (2)
doseras (1/1)
Nettineuvola (1/1)
könsstympning (2/2)
dagpenningens (1/1)
vardagssysslor (2/2)
hälsorådgivningens (1/1)
sevärt (1/1)
prövningfinska (2/2)
fornlämningsområde (1/1)
demonstration (1/1)
enheter (2/2)
Håkansböle (6/6)
amatörteatrar (2/2)
alternativ (8/8)
städernas (1/1)
barnskyddslagenfinska (1/1)
hotat (2/2)
vila (1/1)
utgörs (3/3)
produktionsmedel (2/2)
Finlex (2/2)
tillställning (1/1)
kommun (19/19)
grupplivförsäkring (1/1)
fiskeområden (1/1)
medborgarorganisationer (1/1)
folkpensionens (1/1)
karaoke (1/1)
träning (1/1)
behovet (6/6)
bär (4/4)
ministrarna (1/1)
bildar (1/1)
utarbetas (5/5)
färdigheterna (1/1)
psykoterapi (4/4)
gifte (1/1)
spela (4/4)
allvarliga (1/1)
telefontid (1/1)
Internetberoende (1/1)
RFV (1/1)
nummer (6/6)
vårdbidrag (1/1)
farföräldrar (2/2)
tim. (1/1)
MinSkatt (3/3)
ännu (10/10)
tvisten (1/1)
läsämnena (1/1)
å (3/3)
nuortenkeskus (2/2)
flyktingstatus (16/16)
Furumo (3/3)
registreringsanmälan (1/2) Registreringsanmälan (1)
företagskulturen (2/2)
motion (26/27) Motion (1)
upprätthålls (5/5)
sluttexterna (1/1)
hemvård (6/6)
verka (2/2)
språkkurserna (1/1)
introduktion (1/1)
aktuell (4/4)
hembesök (2/2)
Museiverkets (2/2)
biblioteks (1/1)
biljettpriserna (2/2)
steril (2/2)
komplettera (2/2)
skattefriheten (1/1)
responssystemet (1/1)
faktiska (1/1)
släkting (6/6)
arbetslösa (25/25)
skivor (1/1)
skaka (1/1)
bero (1/1)
erövrats (1/1)
rättvist (3/3)
tobak (1/1)
ansökningarna (2/2)
tortyr (1/1)
exempel (355/355)
anslutning (8/8)
vårdenhet (2/2)
yrkessjukdom (1/1)
medlare (2/2)
efternamnet (2/2)
idrottsföreningar (1/1)
hotad (1/1)
lägger (2/2)
Patent- (2/3) patent- (1)
öka (2/2)
besluten (1/1)
tingsrätten (9/9)
privatsektorn (1/1)
Nordea (1/1)
nationalmuseumfinska (1/1)
kielitaito (2/2)
boendet (9/9)
Mielenterveysseura (3/3)
bindande (6/6)
diskuterar (2/2)
hyr (8/8)
punkt (1/1)
femton (1/1)
hyreshusbolaget (1/1)
inför (11/11)
amorteras (1/1)
skor (1/1)
trappan (1/1)
perustamisilmoitus (1/1)
allmänheten (2/2)
förändringsarbeten (2/2)
historiafinska (1/1)
yrkesstudier (1/1)
erhållit (2/2)
återkallar (2/2)
behärskar (2/2)
evenemangskalenderfinska (1/1)
fallen (1/1)
arbetefinska (1/1)
trygg (5/5)
webbenkäter (1/1)
integrationen (4/4)
romanifinska (1/1)
räkningar (2/2)
säätiö (1/1)
förberedande (39/41) Förberedande (2)
godkännande (1/1)
sökningen (1/1)
VAV (2/2)
rättshjälpsbyrån (4/4)
låga (4/4)
sjukledighetsdagen (1/1)
omständighet (1/1)
dyrt (1/1)
sjukdomar (8/8)
måltidsstödet (1/1)
offentligt (7/7)
naturhistoriska (1/1)
affärsverksamhetsplan (9/9)
hamnade (1/1)
genomgå (2/2)
larm (1/1)
kortare (5/5)
sommaruniversitetfinska (2/2)
företagsledning (1/1)
skada (8/8)
allmänläkare (3/3)
lånegaranti (1/1)
studielån (4/4)
tyger (1/1)
upprättandet (3/3)
språkfinska (2/2)
ll (1/1)
tåg (3/3)
instruktioner (1/1)
bensinstationer (2/2)
beräknas (10/10)
parkeringsbiljetten (1/1)
grunddagpenning (8/8)
51:a (2/2)
hemmet (36/36)
yrkesskolorna (1/1)
vidimeras (1/1)
B2 (1/1)
intervjuer (1/1)
finansierade (3/3)
följs (11/11)
barnrådgivningen (8/8)
tolkningsspråket (1/1)
osakligt (3/3)
pengarna (1/1)
Sandudd (1/1)
besöksförbudfinska (1/1)
pimpla (2/2)
personefterforskningen (1/1)
äter (4/4)
henne (4/4)
folkomröstningar (1/1)
barnen (25/25)
kyrkan (21/21)
pedagogiska (3/3)
Korso (3/3)
samhälleliga (1/1)
missbrukat (1/1)
EU- (6/6)
betald (1/1)
beräkna (3/3)
elarbeten (1/1)
biblioteksnätverket (1/1)
vardag (2/2)
någons (1/1)
dock (54/54)
vise (1/1)
terveydenhoitaja (2/2)
tävlingen (4/4)
personbeteckning (31/31)
förpackningen (1/1)
valmansförening (1/1)
begravningen (3/3)
filmfestivaler (2/2)
familjeåterföreningen (1/1)
invandrarbarn (4/4)
anser (3/3)
åligger (2/2)
kompetens (3/3)
bosniska (2/2)
näringslivet (1/1)
tämligen (1/1)
festivalerfinska (1/1)
president (4/4)
teckenspråk (3/3)
förlängning (2/2)
anstalt (2/2)
webbsidor (8/8)
individuellt (3/3)
arbetslöshetskassan (6/6)
förlorar (3/3)
upplevelser (1/1)
telefonservicefinska (1/1)
fått (44/44)
seniorineuvonta (2/2)
familjemedlemmarnas (2/2)
återförening (1/1)
upphävs (2/2)
HOAS (8/8)
pensionssystem (1/1)
nuvarande (7/7)
chattenfinska (1/1)
utmärkta (1/1)
säsongtopp (1/1)
estniska (51/51)
upprepade (1/1)
stödåtgärderfinska (1/1)
fastighetsförmedlare (1/1)
människor (37/37)
P (3/5) p (2)
partier (1/1)
mottagningscentret (1/1)
skatteförvaltningenfinska (1/1)
antecknats (3/3)
kärren (1/1)
hormonella (2/2)
skala (1/1)
erbjuds (13/13)
depressionen (1/1)
fordrar (1/1)
arbetspensionsanstalter (1/1)
förskolebarn (2/2)
maskinmästare (1/1)
erkännande (12/14) Erkännande (2)
började (6/6)
mopedkort (1/1)
döva (1/1)
material (13/13)
ledighet (4/4)
åka (5/5)
upphört (6/6)
skulden (2/2)
samboskap (1/1)
veckoslut (15/15)
tillstånd (57/57)
finansieringsalternativ (3/3)
annan (65/65)
Verla (1/1)
uppsägningsvillkor (3/3)
maximibelopp (1/1)
Schengenområdet (6/6)
kaupunki (1/1)
sammanfattning (3/3)
studiebyrå (1/1)
språkkunskapskraven (1/1)
brand (9/9)
ungdomstjänster (6/6)
moderskaps- (1/1)
arbetslivets (1/1)
telefonsamtal (1/1)
ungdomsgrupper (1/1)
utrustningen (2/2)
älv (1/1)
Väestöliitto (6/6)
fax (3/3)
eläkevakuutus (2/2)
rösten (1/1)
psykiatrisk (2/2)
arbetsavtalet (15/15)
ett (963/965) Ett (2)
tryggat (2/2)
HIVfinska (1/1)
vänta (8/8)
arbetssäkerheten (2/2)
tidsbeställning (7/7)
startade (1/1)
semesterersättning (2/2)
huvudstadsregionen (12/12)
Trapesa (2/2)
duar (3/3)
anslutningsblankett (1/1)
sjukförsäkringen (13/13)
ammattiopisto (4/4)
förväg (22/22)
revisionsbyrå (1/1)
förgiftats (1/1)
hemvården (2/2)
fördel (2/2)
övervaka (1/1)
civilståndsintyg (1/1)
hamnar (2/2)
rekrytering (1/1)
idrottsområdet (4/4)
vardagar (17/17)
käräjäoikeus (3/3)
utrikespolitiken (1/1)
sambo (17/17)
strid (1/1)
läkarpriserfinska (1/1)
töms (1/1)
tandvårdstjänster (1/1)
fotot (1/1)
förknippade (2/2)
småbarn (1/1)
YH (2/2)
yrkesläroanstalt (8/8)
sund (1/1)
hälsostationsläkare (1/1)
väsentlig (3/3)
medborgarskapsansökan (2/2)
helger (6/6)
LinkedIn (1/1)
Myrbacka (2/2)
hälsostationernas (2/2)
webbplatsfinska (4/4)
Adolf (1/1)
julsånger (1/1)
pensionens (1/1)
skattebyråns (1/1)
börjar (34/34)
tidsperioder (1/1)
folkhögskola (2/2)
vittnen (4/4)
stödformer (1/1)
fågelungar (2/2)
gemensamt (11/11)
vända (7/7)
försäkringarna (1/1)
Huvudstadens (3/3)
hyresbostäderengelska (1/1)
trafikfinska (1/1)
personal (2/2)
fackförbund (14/16) Fackförbund (2)
familjerådgivningen (18/18)
band (1/1)
bestyren (1/1)
använder (17/17)
medicinskt (1/1)
lokaltrafikens (1/1)
Chile (1/1)
gården (1/1)
FRK:s (1/1)
telegram (1/1)
regionen (3/3)
uppehållskortet (3/3)
resorna (1/1)
skötsel (2/2)
deltidsarbete (1/1)
vigselhandlingarna (1/1)
bibliotekets (3/3)
digitalbox (1/1)
självstyre (2/2)
utredningen (3/3)
Haag (1/1)
tågtidtabellerna (1/1)
färdtjänsten (1/1)
sjöar (1/1)
åringar (5/5)
förskola (2/2)
följebrev (1/1)
lämnas (13/13)
dömer (1/1)
form (11/11)
diskrimineringsombudsmannens (2/2)
inkomst (12/12)
handikapptolkar (1/1)
Nimettömät (1/1)
kalla (2/2)
skör (1/1)
förmyndarskap (2/2)
uppkommer (1/1)
alle (1/1)
grundskolanengelska (1/1)
ruokakunta (1/1)
samling (1/1)
hög (7/7)
lön (46/46)
hälsorådgivningfinska (2/2)
hela (27/27)
sociala (74/74)
teoretiskt (1/1)
borgerliga (1/1)
Korkalovaara (1/1)
köpa (32/33) Köpa (1)
kl (73/73)
vårdnadshavarens (1/1)
stödtjänsterna (2/2)
användarna (4/4)
lösas (3/3)
verksamhetsformerna (1/1)
dras (4/4)
anhörigvård (1/1)
betalningen (1/1)
varmare (1/1)
tredjelandsmedborgare (1/1)
kreditgivningfinska (1/1)
koordinatoren (1/1)
hälsostations (1/1)
ingreppet (1/1)
arbete (78/82) Arbete (4)
repetera (1/1)
hemmaarbete (1/1)
vuxengymnasier (2/2)
duger (3/3)
mor (11/11)
jämställdhetsombudsmannen (3/3)
tutkinta (1/1)
förmån (2/2)
beredning (2/2)
ringa (58/58)
hälsocentralläkarens (1/1)
Rovanapa (2/2)
konsthusen (1/1)
inledande (27/27)
upprättas (5/5)
vårdnadshavaren (1/1)
Uudenmaan (1/1)
sjukförsäkringsersättningen (1/1)
työsuojelun (1/1)
forna (1/1)
Luksia (1/1)
begravningsbyråer (2/2)
studentexamenfinska (1/1)
beteendefinska (3/3)
påtryckningar (1/1)
borta (1/1)
moderskapspenningperioden (1/1)
skolresa (1/1)
värdefull (1/1)
stadssund (1/1)
lukiopohjainen (1/1)
sidor (18/18)
elva (3/3)
exakta (3/3)
ersättningarfinska (1/1)
måltidstjänster (1/1)
befunnit (1/1)
moderskapsledighet (2/2)
motionfinska (1/1)
företagsformerfinska (1/1)
talous- (1/1)
restaurang (3/3)
inrättas (1/1)
rosoll (1/1)
handlingar (11/11)
rakt (3/3)
verkställande (1/1)
hyresbostäder (32/32)
sammanhängande (1/1)
folkhögskolanfinska (1/1)
socialskyddsförmånerna (1/1)
Wien (2/2)
sjukskrivning (1/1)
utlandsresa (1/1)
minderåriga (7/7)
patientens (2/2)
religiösa (10/10)
förslag (3/3)
utbetalat (1/1)
välkomna (3/3)
åldersspannet (1/1)
lägsta (1/1)
konstuniversitet (2/2)
stämma (3/3)
måndagar (3/3)
oktober (2/2)
befolkningen (3/3)
assistentens (1/1)
tillfrisknande (1/1)
efternamn (48/48)
idrottstjänster (5/5)
innebär (20/20)
äitiysneuvola (2/2)
boenderådgivare (1/1)
meritförteckning (5/5)
lagen (26/26)
kommunfinska (1/1)
returnera (1/1)
önskar (5/5)
hindersprövning (5/5)
A1.3 (1/1)
rutterna (1/1)
upphörde (1/1)
tulkki (1/1)
antingen (35/35)
stora (15/16) Stora (1)
flyktingens (1/1)
beskattning (6/10) Beskattning (4)
sähköinen (1/1)
alternativa (1/1)
grupp (9/9)
faderskapsledighet (3/3)
erkänts (3/3)
ledigheterna (1/1)
stressyndromfinska (1/1)
far (9/9)
biIdkonstskola (1/1)
läst (4/4)
grunder (9/9)
enhetlig (1/1)
Unescos (1/1)
tandhälsovårdenfinska (1/1)
begå (2/2)
mousserande (1/1)
miljön (3/3)
samråd (2/2)
vårdnaden (8/8)
linjen (1/1)
idrottsmöjligheter (2/2)
reseförsäkring (1/1)
ortodoxa (13/13)
läkemedlen (1/1)
tandvård (19/19)
arbetsplatsintroduktion (1/1)
bankernas (1/1)
betalningsplan (2/2)
parterapi (1/1)
söndagen (1/1)
Sparbanken (1/1)
förmånligare (9/9)
förete (1/1)
avgiften (4/4)
grundskola (1/1)
sakkunnig (2/2)
förhöjningsdelen (1/1)
rajoitetusti (1/1)
magistratfinska (1/1)
Ingående (2/3) ingående (1)
företer (1/1)
Fjällrävsstigen (1/1)
försätts (1/1)
underhålls (1/1)
japanska (6/6)
omedelbart (3/3)
receptet (1/1)
legaliserade (1/1)
oftast (22/22)
resekort (9/9)
sjukhusvård (2/2)
presidentvalfinska (1/1)
fritidsintressen (3/3)
väntat (1/1)
dateras (1/1)
vad (22/24) Vad (2)
ITE (1/1)
symboler (1/1)
arrangören (1/1)
trupper (1/1)
rätt (226/226)
handledningstjänster (1/1)
utbildats (1/1)
sitt (53/53)
ungdomslokalerna (1/1)
hanteras (2/2)
seder (5/5)
stipendiesystem (2/2)
nutidskonst (1/1)
värnpliktiga (1/1)
uppståndelse (1/1)
igen (2/2)
nattjour (3/3)
kriser (1/1)
isen (7/7)
allemansrätten (2/2)
flyttrörelsen (1/1)
husfinska (2/2)
sorg (1/1)
servicebolag (1/1)
valkretsar (1/1)
förmiddagar (1/1)
förlorat (1/1)
förmåga (2/2)
misstänks (2/2)
hantera (2/2)
representeras (1/1)
alkoholisterfinska (1/1)
Omatila (4/4)
medlas (1/1)
operation (2/2)
prov (6/6)
osuuskunta (1/1)
guiden (2/2)
motiverade (1/1)
självrisktiden (2/2)
stadgar (1/1)
skolor (18/18)
utländskt (2/2)
Grani (2/2)
hembygdsmuseerna (1/1)
känslofyllda (1/1)
hantverk (3/3)
skydd (12/12)
korrigerande (1/1)
yrkesbenämning (1/1)
A2.2 (1/1)
konsumenträttigheterfinska (1/1)
någonstans (3/3)
bostadsrättsavtalet (1/1)
liten (11/11)
kök (1/1)
hedersrelaterade (2/2)
nordliga (3/3)
matematik (1/1)
sexåringar (2/2)
Sello (1/1)
museikvarterens (1/1)
vanlig (3/3)
ungdomarna (2/2)
måltider (4/4)
uttryckligen (1/1)
Sovjetunionens (1/1)
syrjintä (1/1)
måndag (9/9)
indoeuropeiska (1/1)
vietnamesiska (7/7)
källa (1/1)
överallt (1/1)
personerlinkkiEsbo (1/1)
Hagalunds (1/1)
lukio (4/4)
kommunalt (3/3)
sjukvårdstjänsterna (4/4)
branschspecifika (1/1)
beställer (7/7)
varmaste (1/1)
gamla (8/9) Gamla (1)
mottagningen (5/5)
berättigad (2/2)
beroende (10/10)
psykologhjälp (1/1)
går (43/43)
trapphuset (2/2)
ansökningsblankett (9/9)
utbytesprogrammetengelska (1/1)
forskningen (1/1)
ledare (1/1)
tohtori (1/1)
vägg (1/1)
gångtrafiken (1/1)
socialarbetarefinska (1/1)
djuren (1/1)
ingrepp (1/1)
täckjacka (1/1)
mån.-tors. (1/1)
utsätts (1/1)
tidsgränser (1/1)
nödsamtal (1/1)
halvt (1/1)
badstränder (1/1)
ansvara (1/1)
kandidat- (1/1)
integreras (1/1)
arbetsuppgifterna (2/2)
umgänget (4/4)
använts (2/2)
inkassokostnader (1/1)
Vanda (115/115)
advokater (1/1)
anhålla (1/1)
hälsovårdaren (9/9)
centralernafinska (1/1)
avslås (1/1)
kön (22/22)
innehar (2/2)
alkoholism (1/1)
hengenvaara (1/1)
Barnskyddsförbund (4/5) barnskyddsförbund (1)
fordonsskatten (1/1)
förknippas (1/1)
släktning (1/1)
nödfall (8/8)
familjeverksamhet (1/1)
inträffat (2/2)
utnyttjande (1/1)
Takuusäätiös (1/1)
bostadsrättsavgift (1/1)
valmistava (1/1)
döda (2/2)
civilvigslar (1/1)
pensionerna (3/3)
undgås (1/1)
hälstocentralen (1/1)
uppehållsrätten (18/18)
servicerådgivningen (1/1)
sökte (1/1)
ombyggnadsarbeten (1/1)
käpp (1/1)
vitsord (5/5)
sjunga (2/2)
grundtryggheten (1/1)
kostnad (1/1)
gravområde (2/2)
överföras (1/1)
stipendium (4/4)
asylsökandefinska (2/2)
doulaverksamheten (1/1)
textade (1/1)
telefonen (2/2)
bedrivit (1/1)
fortlöpande (2/2)
kontaktar (3/3)
bo (55/55)
vårdnad (16/16)
smarttelefonen (1/1)
till (1547/1553) Till (6)
eduskunta (2/2)
Omnia (3/3)
SIMHE (4/4)
kylskåpets (1/1)
storlekar (1/1)
hette (1/1)
partiella (3/3)
Österbotten (2/2)
sjukdomstid (2/2)
utbildningsanordnare (1/1)
gått (10/10)
hälsoproblem (1/1)
sjöfästning (1/1)
ljusa (1/1)
statens (9/9)
informering (1/1)
läroanstalten (11/11)
besitter (1/1)
betalningskrav (1/1)
likabehandling (12/12)
matsäck (1/1)
tryggare (1/1)
tjänstens (2/2)
medarbetare (1/1)
upphovsmannens (1/1)
fackevenemang (1/1)
ämbetsbevis (2/2)
ArPL (1/1)
diskrimineringsfall (1/1)
hyrsvärden (1/1)
trafik (3/3)
skiljas (3/3)
seglare (1/1)
diskmaskin (1/1)
rättighet (2/2)
skogar (1/1)
intervjuerna (1/1)
biografkedjan (1/1)
mödrarådgivningar (1/1)
början (16/16)
anslutningsledning (1/1)
hyresvärd (2/2)
Lastensuojelulaki (1/1)
undervisningen (26/26)
anställningsoptioner (1/1)
förebygga (1/1)
hemkommun (104/114) Hemkommun (10)
klinikka (3/3)
behåller (2/2)
bearbetningar (1/1)
godkänd (3/3)
historiska (4/4)
förvaltningsmyndigheter (1/1)
förskott (1/1)
Helsinkis (1/1)
talar (6/6)
ganska (1/1)
Tullens (1/2) tullens (1)
Kopparbergsvägen (1/1)
festivalen (1/1)
skattar (1/1)
vattentrafiken (1/1)
byta (8/8)
ordentlig (2/2)
kran (1/1)
areal (3/3)
företagsverksamheten (9/9)
Dublinprocessen (1/1)
språkversionerna (2/2)
bostadens (9/9)
hobbyverksamhet (5/5)
konkurrera (1/1)
avlägsnande (1/1)
museer (10/10)
Hedersrelaterat (1/1)
döden (1/1)
ljudböcker (2/2)
preventivrådgivningen (1/1)
kassan (5/5)
Kyllönen (2/2)
syften (1/1)
partnern (2/2)
tidigt (6/6)
gripa (1/1)
blanketten (18/18)
julgran (1/1)
nämnden (1/1)
stadens (53/53)
livsfara (2/2)
rusmedelsberoende (1/1)
bassjälvrisk (1/1)
omsorg (2/2)
förblir (3/3)
grunddagpenningen (1/1)
perukirja (1/1)
biljettpriser (2/2)
FPA.Som (1/1)
asyl (20/20)
flyktingbakgrund (1/1)
beträda (2/2)
störa (1/1)
billigast (1/1)
yngsta (2/2)
startas (1/1)
alls (1/1)
ord (4/4)
framgår (3/3)
bostadssökande (1/1)
arbetssäkerhets- (1/1)
myndighets (1/1)
återkalla (1/1)
produktionen (1/1)
framgå (3/3)
oväntat (2/2)
enskild (4/4)
elektroniskt (11/11)
upptäcker (8/8)
Suomenlinna (1/1)
inriktningar (1/1)
kontrakt (1/1)
mataffären (1/1)
gäller (40/40)
kontaktuppgifter (6/6)
skriftliga (5/5)
skilsmässoansökan (6/6)
samfällighets (3/3)
röster (2/2)
uppfyller (5/5)
omhändertagande (1/1)
verkställer (1/1)
stilla (1/1)
nätbankkoder (1/1)
telefonabonnemang (1/1)
påföljder (1/1)
diskutera (7/7)
förtroendemannen (4/4)
ur (8/8)
turkiska (15/15)
erhöll (1/1)
tullanmälan (1/1)
anslöts (2/2)
Karlebynejden (1/1)
funktionshinder (1/1)
läggas (1/1)
roligt (1/1)
nomineras (2/2)
gymnasieutbildningen (1/1)
anvisningar (19/19)
inkomstgränsen (1/1)
fisketillståndfinska (1/1)
Residuum (2/2)
jakt (2/2)
examensdel (2/2)
prevention (5/5)
arbetslöshetsförmånfinska (1/1)
perhehoito (1/1)
vitsorden (1/1)
rekreation (1/1)
registreringen (6/6)
ovanlig (1/1)
vem (15/15)
förändrades (1/1)
beskattningenfinska (2/2)
arvolautakunta (1/1)
sjuk (20/20)
työsuojelupiiri (1/1)
stöder (8/8)
semesterresa (1/1)
ansvarsområden (1/1)
välfärds- (1/1)
telefon (38/38)
kredituppgifterna (1/1)
identitetsbevis (8/8)
skridskobanor (1/1)
työpaikat (2/2)
Jönsasvägen (1/1)
hälsorisk (1/1)
urvalsbaserade (1/1)
kremeras (1/1)
förmånligaste (1/1)
krismottagning (2/2)
bibliotekfinska (1/1)
reparationsarbeten (1/1)
integrering (1/1)
familjeförmånerna (1/1)
allmännyttiga (1/1)
EMMA (1/1)
hindi (1/1)
försvara (2/2)
arbetskraftsutbildningfinska (1/1)
dammsugaren (1/1)
utvisad (1/1)
föreningsmedlemmar (1/1)
viss (20/20)
klinikerna (1/1)
Indien (1/1)
desto (1/1)
centraliserade (3/3)
slut (4/4)
skrämma (1/1)
Määräaikainen (1/1)
krävs (32/32)
aktörerna (1/1)
tack (4/4)
tredje (6/6)
delbeslut (3/3)
avtalet (21/21)
utarbetandet (1/1)
översättning (1/1)
misstänka (1/1)
ersättningen (1/1)
Apostille (1/1)
Herman (1/1)
filmvisningarfinska (1/1)
tidigare (21/21)
Caisa (1/1)
gjort (5/5)
beslutsmakt (1/1)
restauranger (1/1)
stad (47/47)
tempel (1/1)
utkomstskyddet (4/4)
folkhögskolorfinska (1/1)
kyrkanfinska (1/1)
EK (2/3) Ek (1)
omskärelsen (2/2)
specialtillstånd (1/1)
söker (41/41)
rådgivning (54/54)
eija.kyllonen (1/1)
tillståndskort (1/1)
teknisk (1/1)
färdas (4/4)
barnlöshet (1/1)
musikverksamhet (1/1)
apoteken (1/1)
dubbade (1/1)
Uleåborgs (1/1)
Infobank (1/1)
politiskt (1/1)
passfinska (1/1)
skolgång (4/4)
alltså (25/25)
än (106/106)
vuxen (5/5)
studentexpeditionen (1/1)
tull (1/1)
jourhavande (2/2)
hemmetfinska (1/1)
regnar (1/1)
h (1/1)
asylsamtal (1/1)
packa (1/1)
några (24/24)
medborgarskapfinska (3/3)
tio (3/3)
oman (1/1)
menas (1/1)
förlorade (2/2)
start (1/1)
skolpsykologen (2/2)
upplösning (2/2)
efter (88/88)
tidsbeställningen (2/2)
torteras (1/1)
belägen (1/1)
ställe (9/9)
hjälper (63/63)
koppling (1/1)
studiemiljö (2/2)
föreningsverksamhet (2/2)
hushållets (1/1)
dricks (1/1)
hammashoitola (2/2)
arbetsför (1/1)
arbetarskyddsmyndigheter (1/1)
uppmuntras (1/1)
eKirjasto (1/1)
ställer (2/2)
erövrade (2/2)
laga (3/3)
utbetalningen (2/2)
European (1/1)
veckoslutet (2/2)
tryggt (5/5)
högskolestudier (8/8)
trafik- (1/1)
verkställa (1/1)
tillståndet (17/17)
kortfinska (1/1)
utöver (5/5)
mån. (1/1)
specialsmåbarnspedagogiken (1/1)
studiebetyg (1/1)
tag (1/1)
remixa (1/1)
äe (1/1)
bröstcancer (2/2)
arbetarinstitutet (1/1)
möjlig (2/2)
kommunerna (18/18)
matställen (1/1)
minimilöner (4/4)
grannar (1/1)
ägarbostäder (1/1)
gårdsområdet (1/1)
stat (4/4)
graviditeten (16/16)
överenskommelse (3/3)
testamentti (2/2)
därmed (2/2)
kieli (1/1)
varor (5/5)
toimeentulotuki (1/1)
inlärning (4/4)
varhaiskasvatushakemus (1/1)
telefonledes (4/4)
flerårigt (1/1)
anknutna (1/1)
socialt (1/1)
försvarsmakt (1/1)
befolkningsdatasystemet (14/14)
par (17/17)
livsåskådning (1/1)
väg (2/2)
kund (12/12)
specialiserade (1/1)
församlings (3/3)
förbudet (1/1)
Virtanen (2/2)
vin (1/1)
kvarskatten (1/1)
kurserna (16/16)
arbetslöshetsdagpenning (2/2)
besöka (35/35)
arbetssökning (1/1)
påbrå (1/1)
varainsiirtovero (1/1)
brådskande (27/27)
starkt (2/2)
tillräcklig (10/10)
marknadsföring (1/1)
utdrag (3/3)
droganvändning (1/1)
reparationer (5/5)
hälsovården (18/18)
skadligt (1/1)
källan (1/1)
bostadssidor (1/1)
befolkningsdatasystem (4/4)
hemsida (1/1)
utfärdades (1/1)
Apteekkariliitto (1/1)
anställningsavtal (1/1)
våldsam (3/3)
kartanfinska (1/1)
lugga (1/1)
synskada (1/1)
genomförandet (1/1)
Musikantitfinska (1/1)
jourtelefon (1/1)
handelstrafik (1/1)
förändras (1/1)
Yhden (2/2)
Axxell (2/2)
mylla (1/1)
matkulturenengelska (1/1)
håller (11/11)
värme (1/1)
bostadsaktiebolag (5/5)
internationella (19/21) Internationella (2)
variera (4/4)
nyttar (1/1)
ersättningsgilla (1/1)
underhållsstöd (4/4)
utgångstid (1/1)
hallen (1/1)
föder (4/4)
yrkesutbildning (35/36) Yrkesutbildning (1)
grenförbunden (1/1)
stiftas (1/1)
egenskaperna (1/1)
sektorn (10/10)
kontanter (5/5)
olycksfallsförsäkring (3/3)
meddelandekortet (1/1)
högskolexamen (1/1)
planen (1/1)
hälsomotionsgrupper (1/1)
idrottscentret (1/1)
livskompetensen (1/1)
resepti (1/1)
vrida (1/1)
terminsavgifter (1/1)
beräkning (1/1)
huvudjärnvägsstation (1/1)
flyttsak (2/2)
högklassig (1/1)
skattefritt (1/1)
försenade (2/2)
tillfoga (2/2)
betalningsdagar (1/1)
avsnitten (1/1)
Flyktingrådgivningen (3/3)
hemsjukvård (1/1)
A1.2 (1/1)
sommaren (10/10)
praktiken (5/5)
fyller (17/17)
familjedagvårdare (7/7)
ej (1/1)
hårdaste (1/1)
betänketid (2/2)
våningen (4/4)
ensamstående (3/3)
caféer (1/1)
hemvårdsstöd (13/13)
Medborgarrådgivning (1/1)
asevelvollisuus (1/1)
arvingarna (1/1)
beslutet (13/13)
lisensiaatti (1/1)
religionsutövande (1/1)
diplomingenjörsexamen (1/1)
leder (8/8)
avgiftsbelagt (4/4)
berusad (1/1)
seniorer (6/6)
fordonsföreskrifter (1/1)
dokument (4/4)
pojkens (1/1)
Folkmusik (1/1)
ägo (1/1)
förstasida (1/1)
videkvistar (1/1)
effektiva (1/1)
ändamålet (1/1)
evankelis (1/1)
EES (35/35)
ingendera (1/1)
kronologisk (2/2)
familj (22/22)
bioprogrammet (1/1)
mars (6/6)
rusmedelsbruk (1/1)
fortsättningen (1/1)
reserverad (1/1)
klarlägga (1/1)
Al (1/1)
uppstartsföretag (2/2)
sälfångst (1/1)
anmält (4/4)
Schengen (1/1)
ens (3/3)
servicestället (10/10)
rusmedels- (1/1)
bolagsvederlag (1/1)
tillgångar (4/4)
företagsläkare (1/1)
trauma (1/1)
kamratstöd (2/2)
löptid (1/1)
museet (3/3)
ordning (2/2)
socialtjänsterna (2/2)
bussar (4/4)
organisationer (15/15)
gångfinska (1/1)
gymnasiernas (1/1)
stadsmuseum (1/1)
förmedling (1/1)
indriver (1/1)
arbetskulturen (5/5)
barnpassningshjälpen (1/1)
själva (12/12)
enkla (1/1)
föräldrarnafinska (1/1)
brottsmål (1/1)
införde (2/2)
Kokkola (2/2)
tågbiljetter (1/1)
luftfartsyrken (1/1)
spelar (1/1)
gifter (4/4)
bygga (6/6)
bilda (1/1)
elinkeinotoimisto (4/4)
ljud (1/1)
yrkesbeteckning (1/1)
helheter (1/1)
sammankallas (1/1)
byggherrar (1/1)
hårdare (1/1)
Turku (1/1)
finlandssvenska (2/2)
erfarenhet (2/2)
upphöra (2/2)
ändamål (1/1)
Sveriges (2/2)
bosättning (2/2)
permanenta (2/2)
gymnasieskolans (1/1)
såväl (5/5)
Baltikum (1/1)
språkkursernas (1/1)
medlemmars (2/2)
felen (1/1)
skolans (10/10)
välartat (1/1)
kommunernafinska (2/2)
Helsingfors (169/169)
andra (185/185)
intresse (4/4)
djurskötarexamen (1/1)
överskridits (1/1)
sosiaalivirasto (1/1)
Sverige (16/16)
ägt (1/1)
avslagits (1/1)
Karlebyfinska (5/5)
inhämta (4/4)
Olofsborg (1/1)
fuktisolering (1/1)
anger (3/3)
internationellt (8/8)
museot.fi (1/1)
lämplig (14/14)
TE (73/74) te (1)
handskar (1/1)
års (16/16)
läroavtalscenterfinska (1/1)
försäkringsintyg (1/1)
fortsättningskriget (1/1)
mycket (66/66)
invandrararbete (1/1)
Konvaljvägen (1/1)
lagt (1/1)
träsliperi (1/1)
betalades (2/2)
namn (21/21)
utbildningsprogrammet (1/1)
köpebrevet (1/1)
bekräftade (1/1)
konsumenter (1/1)
linje (2/2)
stadiet (6/6)
miljö (5/5)
Avfallshantering (3/4) avfallshantering (1)
påverkat (1/1)
mallarfinska (1/1)
oikeudet (1/1)
köptjänst (1/1)
idka (4/4)
ansökningstiden (3/3)
ärendena (1/1)
missbruksvård (1/1)
stödet (12/12)
föreningens (3/3)
skaffa (26/26)
rum (4/4)
Soites (4/4)
godtagbara (1/1)
RIKU (1/1)
samboförhållandet (6/6)
arbetsgivaren (49/49)
företett (1/1)
skaffar (6/6)
näringsbyråns (9/9)
hälsoåvård (1/1)
mitt (9/9)
förlängd (1/1)
studieplatsen (1/1)
säsongsarbetsvisum (1/1)
yrkesutövning (2/2)
styrs (2/2)
beställa (14/14)
i (2699/2701) I (2)
universitetscenter (1/1)
skolläkaren (3/3)
praktiska (7/7)
mentalvårdstjänster (2/2)
skulle (9/9)
tänka (2/2)
civiltjänstgöring (1/1)
särställning (1/1)
hälsafinska (2/2)
nationernas (2/2)
husbolaget (2/2)
rådgivnings- (2/2)
tabletdator (1/1)
välja (16/16)
dagvårdsplats (8/8)
tandläkarkontroller (1/1)
handläggningsavgiften (1/1)
polikliniker (2/2)
registrerades (2/2)
hälsorelaterade (1/1)
telefonnumret (2/2)
fler (10/10)
himmelsfärdsdag (1/1)
goda (10/10)
naturcenter (1/1)
behövs (28/28)
egna (44/44)
informationstjänst (1/1)
beslutsfattarna (1/1)
socialväsen (2/2)
hjälpsystemet (1/1)
K.H.Renlunds (3/3)
kundens (2/2)
kosthållsbranschen (1/1)
kulturcentral (1/1)
debiteras (1/1)
uppgiften (3/3)
antal (4/4)
Jorv (10/10)
äktenskapsintyg (4/4)
verkar (2/2)
uppehälle (5/5)
flygplatser (1/1)
grundskolans (12/12)
folkpensionen (1/1)
nybörjare (1/1)
lättläst (1/1)
förmedlingsarvode (1/1)
barnet (160/160)
hand (60/60)
flytthjälp (1/1)
rekommenderas (2/2)
forskarefinska (1/1)
symtom (1/1)
rådgivningstjänst (5/5)
familjerådgivningfinska (1/1)
konkret (1/1)
låneräntan (1/1)
användningsdatumet (1/1)
väder (1/1)
erfarenheter (3/3)
finansierat (1/1)
barndagvård (8/8)
eläkekassa (1/1)
Europaparlamentsvalfinska (1/1)
bekänna (1/1)
frysens (1/1)
sträcker (1/1)
studieprogram (2/2)
boendekostnader (5/5)
R (1/1)
apparater (2/2)
medborgarskapsanmälan (4/4)
hoitoapupalvelu (1/1)
alltför (3/3)
elvärme (1/1)
betjänad (1/1)
lampor (2/2)
arbetarskyddsmyndigheternafinska (1/1)
ert (1/1)
alkohol- (3/3)
ordningen (1/1)
kuntoutus (2/2)
handikappadefinska (3/3)
oppilaitos (1/1)
tillgängliga (3/3)
flyttsaker (4/4)
högskolestuderande (1/1)
linjekartor (1/1)
avgifter (5/5)
långa (6/6)
filmarkiv (1/1)
möjligheten (3/3)
barnskyddfinska (1/1)
uppfattning (1/1)
arbetsinkomst (2/2)
kurator (1/1)
ökade (1/1)
sommarsolståndet (1/1)
skrivit (1/1)
begränsas (2/2)
språketengelska (1/1)
skadar (1/1)
avsnitt (5/5)
specialdiet (1/1)
rekommendationer (1/1)
praktik (4/4)
motionsevenemang (1/1)
tempus (1/1)
stödpersonen (1/1)
hyresgästerna (1/1)
skolämnen (1/1)
utbildningsväsendetfinska (1/1)
studentkort (1/1)
betjänar (29/29)
äta (1/1)
nödvändiga (5/5)
vägra (7/7)
bestämd (4/4)
avgörande (3/3)
läsa (16/16)
helhetsbetonat (1/1)
Opiskelija (4/4)
orsaker (8/8)
klasser (5/5)
helgdagar (4/4)
dagpenning (13/13)
språk- (3/3)
stadissa.fi (2/2)
fallet (2/2)
ledigheten (1/1)
ansökningstider (2/2)
utses (3/3)
patienter (1/1)
tjänsterfinska (9/9)
gymnasiet (21/21)
G (1/1)
klarläggs (1/1)
arbetsoförmögenhet (2/2)
utvisning (1/1)
temadagar (1/1)
pensionsanstalt (3/3)
Ohjaamo (1/1)
erbjuda (3/3)
bebott (3/3)
förfaringssätten (1/1)
gången (2/2)
sorani (3/3)
disk- (1/1)
servicecentret (1/1)
höger (1/1)
utsidan (1/1)
löner (2/2)
poliklinik (1/1)
hen (28/28)
tolkningstjänsten (1/1)
anmälan (25/25)
vardagkvällar (1/1)
km2 (5/5)
psykisk (3/5) Psykisk (2)
lähetetty (1/1)
bereda (1/1)
genetiska (1/1)
överenskommelsen (3/3)
lantdagsmannen (1/1)
kartläggningar (1/1)
invaliditetspension (6/6)
lastenneuvola (5/5)
förtroendeuppdrag (1/1)
begravningsplatsfinska (1/1)
människorna (3/3)
små (15/15)
vinnare (2/2)
vandring (2/2)
konstnären (1/1)
psykologi (1/1)
hälsostationerna (10/10)
invandringsfrågor (1/1)
pedagoger (2/2)
lågstadiet (2/2)
webben (2/2)
underhållsskyldiga (1/1)
företagsrådgivning (2/4) Företagsrådgivning (2)
kostnadsfri (12/12)
månad (24/24)
kopia (4/4)
föreslog (1/1)
medverkar (2/2)
åker (5/5)
sjukdomsfall (1/1)
upptäcka (1/1)
utbildningstiden (2/2)
InfoFinland (21/21)
svårare (4/4)
Kaustby (2/2)
fortbildning (5/5)
bekymmer (1/1)
stöd- (2/3) Stöd- (1)
krismottagningen (1/1)
lovat (2/2)
lähestymiskielto (1/1)
Norge (7/7)
yhtiö (1/1)
scenkonst (1/1)
februari (5/5)
minimivillkor (1/1)
specialbibliotek (1/1)
webbsidorna (1/1)
knappsatsen (1/1)
uppfylla (3/3)
käsiraha (1/1)
minnestest (1/1)
byggplats (1/1)
kallade (3/3)
diabetesfinska (1/1)
inletts (1/1)
arbetskollektivavtal (1/1)
ingriper (1/1)
inredningsarkitekt (1/1)
lånat (1/1)
Begravningbyråers (1/1)
tvingades (1/1)
postadress (1/1)
sexuell (5/5)
här (32/32)
ungdomsväsendet (1/1)
Perho (1/1)
vederbörligt (1/1)
sambor (5/5)
många (143/143)
felaktiga (3/3)
bostadsköpet (1/1)
biljetter (2/2)
uppgift (8/8)
barnskyddsmyndigheten (2/2)
Spafinska (2/2)
ansökningsförfarandena (1/1)
lokaltrafiken (1/1)
barnrådgivningens (1/1)
renkött (1/1)
befrämjande (1/1)
trafikknutpunkt (1/1)
vårdande (1/1)
kommunalval (9/9)
olyckor (2/2)
intresserad (8/8)
bostadsaktiebolagets (2/2)
WC:n (1/1)
hörselskadade (5/5)
hyresetta (1/1)
reparation (1/1)
separat (23/23)
personalen (5/5)
syfte (2/2)
mandatperioder (1/1)
befinner (5/5)
väntar (6/6)
Vionojas (1/1)
köparens (1/1)
ordningsreglerna (7/7)
originalexemplaren (5/5)
tolk (40/40)
anställningsavtalets (1/1)
aikuiskoulutustuki (1/1)
förmedlare (1/1)
måltiden (1/1)
parter (1/1)
underhållsbehov (3/3)
förtjänat (1/1)
intjänade (3/3)
Vionoja (1/1)
anknyter (4/4)
kommissionen (1/1)
årskurs (5/5)
köparen (2/2)
organisationens (2/2)
vuxenutbildningen (1/1)
allmäneuropeiskt (1/1)
hissa (1/1)
underhyresgäst (3/3)
löpt (2/2)
stapelrättigheter (1/1)
behovsprövad (3/3)
startandet (1/1)
SOA (1/1)
samlas (3/3)
cyklister (1/1)
tillåtelse (1/1)
kypsyysnäyte (1/1)
verifiera (1/1)
framgångsrikt (1/1)
åldrarna (2/2)
kunskap (2/2)
barnlöshetsklinik (1/1)
omfattar (24/24)
hemort (17/17)
fre (22/22)
kortkurser (1/1)
skiftesvård (1/1)
antas (3/3)
Päihdelinkki (2/2)
fulla (1/1)
just (4/4)
makens (4/5) Makens (1)
lunchsedlar (1/1)
diskriminerad (1/1)
Alkoholistit (1/1)
garanti (2/2)
läder- (1/1)
yrkeshögskolorfinska (4/4)
åldringar (4/4)
Lapplands (21/21)
yrkeshögskolan (9/10) Yrkeshögskolan (1)
utbildnings (1/1)
ungdomsgårdarna (4/4)
släckningsfilt (2/2)
inkräktar (1/1)
ekonomin (1/1)
skatteprocenten (2/2)
Sanomat (1/1)
invandrarungdomar (1/1)
VAU (1/1)
samboförhållande (14/16) Samboförhållande (2)
rekryteringsevenemang (1/1)
överskrids (1/1)
auttamisjärjestelmä (1/1)
identiteten (2/2)
EVK (1/1)
elpriserfinska (1/1)
kansli (7/7)
följa (19/19)
avsnittet (1/1)
pensionsförsäkring (3/3)
slogs (1/1)
vistelsen (4/4)
el (3/3)
högtidlig (1/1)
genomgått (1/1)
vigselförrättningen (1/1)
sairaalan (1/1)
psykiatriskötare (1/1)
paddling (1/1)
hyötyliikunta (1/1)
serviceboendet (2/2)
börja (16/16)
verk (1/1)
Korset (6/6)
Rovaniemen (2/2)
rehabiliteringfinska (5/5)
länken (3/3)
frivillig (5/5)
fortsätta (8/8)
tidpunkten (5/5)
nu (1/1)
riket (1/1)
typer (4/4)
kaikille (1/1)
universitetsexamen (2/2)
avgiftsbelagda (9/9)
orsakat (4/4)
metspö (3/3)
extra (4/4)
läroplikten (2/2)
Pyhäjoki (1/1)
begära (14/14)
mångsidiga (3/3)
fadernfinska (1/1)
arbetspensionsanstalt (1/1)
integrationfinska (1/1)
ansökan (145/147) Ansökan (2)
gäster (1/1)
jobbannonsen (3/3)
barnbidrag (8/9) Barnbidrag (1)
flexibla (1/1)
hälsosam (1/1)
särbehandlas (2/2)
vårdas (8/8)
Förenta (1/1)
grundandet (1/1)
integritetsskydd (1/1)
rörelsenedsättning (2/2)
tukiasuminen (1/1)
arbetskraftsmyndigheten (1/1)
affärsverksamhet (3/3)
hälsorådgivningen (2/2)
mervärdesskatt (3/3)
gymnasieskolor (2/2)
ge (23/23)
socialskyddsavtal (2/2)
Rovalan (7/7)
sanning (1/1)
uthyrning (1/1)
självständighetsdagen (1/1)
avslutar (1/1)
kontakta (116/116)
betalningspåminnelse (1/1)
kartläggningfinska (1/1)
matkakortti (2/2)
leksaker (2/2)
självständigheten (1/1)
reparera (1/1)
färdmedel (1/1)
vinterskor (1/1)
receptfinska (1/1)
räkna (2/2)
Giftinformationscentralen (1/1)
områden (17/17)
familjeträningen (1/1)
speciella (1/1)
gör (30/30)
osakliga (1/1)
skatteavdrag (1/1)
storfurstendömets (1/1)
öppnas (1/1)
bolagsman (2/2)
Rovaniemiområdet (1/1)
at (3/3)
affärspartner (1/1)
väderleksrapporterna (1/1)
mening (1/1)
sosiaali- (4/6) Sosiaali- (2)
babyskydd (1/1)
avlider (4/4)
värden (1/1)
turvakoti (4/6) Turvakoti (2)
täcka (5/5)
flyktingen (1/1)
vägledning (5/5)
förnamn (1/1)
rekommendera (2/2)
investerare (1/1)
skoldagarna (1/1)
pojkar (4/4)
företagsrådgivningscentra (1/1)
sekajäte (1/1)
avvägs (1/1)
vaccinationsprogrammet (1/1)
demokrati (1/1)
familjen (49/49)
yrkesinstitut (8/8)
humanistiska (4/6) Humanistiska (2)
Soldatskär (1/1)
språket (50/50)
ärende (3/3)
anordnar (1/1)
regeringen (2/2)
begravning (4/4)
företagstjänsterna (1/1)
sjöfartsbranschen (1/1)
fackets (1/1)
vet (6/6)
våning (4/4)
utlänningar (19/19)
förbindelse (2/2)
egendom (28/28)
jobbet (3/3)
universitetet (19/19)
affärsidén (2/2)
Äkta (1/2) äkta (1)
dubbelrum (1/1)
parförhållandet (14/14)
råd (89/89)
frånvarande (2/2)
nedan (1/1)
värdesätts (4/4)
var (48/56) Var (8)
tolv (6/6)
registrerade (6/6)
vårdsystemet (1/1)
toiminimi (2/2)
verksamhetfinska (3/3)
återbetalas (1/1)
feber (1/1)
anordnad (2/2)
Kotoutumiskeskus (1/1)
daghem (34/34)
anställningen (9/9)
rör (40/40)
yliopisto (4/4)
spel (4/4)
hälsovårdstjänsterna (21/21)
genom (47/47)
serviceställena (1/1)
resurscenter (1/1)
drogproblemfinska (1/1)
julen (2/2)
studieområde (1/1)
verokortti (3/3)
godkänner (4/4)
ägarbostad (17/20) Ägarbostad (3)
depression (2/2)
verksamma (5/5)
ifrågavarande (4/4)
parförhållandets (1/1)
asunto (2/2)
psykoterapeut (1/1)
inga (9/9)
näringsbyrån (40/40)
slutat (1/1)
koulu- (1/1)
biologi (1/1)
annonserar (1/1)
Ristrand (1/1)
respektive (2/2)
buss (1/1)
utförandet (5/5)
Erasmus (2/2)
nya (40/40)
Hyvin (1/1)
rädsla (1/1)
lapsettomuusklinikka (1/1)
busslinjer (2/2)
arbetstagarefinska (1/1)
daghemmet (7/7)
prepaid (2/2)
bekanta (6/6)
30l (1/1)
föräldrarfinska (1/1)
bostadsbidrag (20/25) Bostadsbidrag (5)
kunnanvaltuusto (1/1)
körkort (11/11)
simhallen (1/1)
skötare (5/5)
API (1/1)
ålder (13/13)
individuella (1/1)
invandrarmänfinska (1/1)
avgörs (1/1)
mångkulturell (3/3)
förbereder (3/3)
sommar- (1/1)
lokalerna (1/1)
utrustning (3/3)
barnlöshetspolikliniken (1/1)
utbildningfinska (2/2)
bedömningen (1/1)
veckovisa (1/1)
servicepunkten (3/3)
högskoleutbildning (5/5)
asunnot (6/12) Asunnot (6)
understöd (10/10)
ungdomarnas (2/2)
informationfinska (1/1)
dödsfallet (1/1)
vårdfinska (1/1)
judiska (1/1)
caféerna (1/1)
rummet (1/1)
beaktar (2/2)
brandlarm (1/1)
skattepliktiga (1/1)
idkas (2/2)
jobbsökningenfinska (1/1)
vikens (1/1)
kränkande (1/1)
beakta (7/7)
ägare (6/6)
tillhörande (1/1)
resesättet (1/1)
strykjärnet (1/1)
allvarligt (4/4)
slås (1/1)
uppgår (1/1)
statsborgen (1/1)
bok (1/1)
läkare (35/35)
livet (11/12) Livet (1)
mångfaldigades (1/1)
webbtjänstfinska (1/1)
specialvårdpenning (2/2)
branscher (10/10)
människogrupp (1/1)
Raumo (1/1)
bokföring (1/1)
biograferna (1/1)
Barnkliniken (3/3)
Karl (1/1)
identitetskort (7/7)
studieresor (1/1)
kommuntillägg (4/4)
brottsmisstänkta (3/3)
svensk (1/1)
förhållanden (2/2)
Mannerheims (2/2)
oartigt (3/3)
integrationsspråk (1/1)
lägenhetshotell (2/2)
meningar (1/1)
nödsituation (11/11)
jobbsajterfinska (1/1)
längden (1/1)
ni (42/42)
åtalsprövning (1/1)
farligt (4/4)
försöka (1/1)
populärare (1/1)
lärt (3/3)
anskaffningspris (1/1)
industristad (1/1)
nytt (26/26)
boendeservice (2/2)
smittsamma (2/2)
cykelvägar (2/2)
styr (1/1)
notaries (1/1)
integrationsåtgärderna (1/1)
apteekki (1/1)
kontrollera (19/19)
roll (2/2)
vänskap (1/1)
parkerna (1/1)
kurser (36/36)
sysselsättnings- (1/1)
byråfinska (1/1)
fågelbon (2/2)
utbildnings- (1/1)
otrogenhet (1/1)
fyllning (1/1)
kollektivtrafiken (4/4)
operera (1/1)
ditt (254/254)
Nyföretagarcentral (1/1)
Juristförbunds (2/2)
PUK (1/1)
säker (5/5)
stödundervisningen (1/1)
kristendomen (1/1)
symtomen (1/1)
straffpåföljd (1/1)
männen (1/1)
Räckhals (1/1)
avsikt (2/2)
miljöer (1/1)
frispråkighet (1/1)
gymnasieböckerna (3/3)
uppehållstillstånden (1/1)
poliklinikka (3/3)
engelska (783/783)
säljer (9/9)
köpeanbudet (2/2)
områdeskoordinatorn (1/1)
ägda (1/1)
intill (3/3)
skattedeklarationen (6/6)
maahanmuuttajapalvelut (1/1)
farföräldrarna (1/1)
flyttar (86/86)
besvarar (2/2)
etnisk (2/2)
jordbruks- (1/1)
skäl (14/14)
flytta (16/21) Flytta (5)
färdtjänst (7/7)
servicestyrcentral (1/1)
giltighetstid (1/1)
aikuisopisto (6/7) Aikuisopisto (1)
hit (1/1)
kö (1/1)
äldrefinska (1/1)
talet (15/15)
brandsläckare (1/1)
huvudsyssla (3/3)
integrationsstöd (1/1)
musiikkiopisto (1/1)
cykeln (1/1)
sådan (9/9)
ängre (1/1)
förflutit (1/1)
arvodet (1/1)
offentliga (56/56)
sopkärlen (1/1)
riksdagsledamot (1/1)
tolkförbund (2/2)
Hyresboende (1/1)
växter (1/1)
Konsumentförbund (1/1)
sommaruniversitetetfinska (1/1)
vähennykset (1/1)
turistersvenska (1/1)
nationell (1/1)
ökar (1/1)
yrittäjien (1/1)
ingåtts (5/5)
työtulo (1/1)
Genève- (2/2)
Familjeledighet (2/4) familjeledighet (2)
Salutorget (1/1)
familjedagvård (2/2)
tjänstemannafinska (1/1)
röstningsställe (1/1)
hemvårdsstödets (1/1)
ansökt (4/4)
batteri (2/2)
obligatoriska (4/4)
arbetslöshetskassafinska (1/1)
äktenskap (52/54) Äktenskap (2)
familjemedlemmarna (2/2)
åldrar (5/5)
delar (11/11)
förverkligandet (1/1)
center (5/5)
ifyllda (3/3)
bekräftas (1/1)
kilometer (2/2)
definieras (4/4)
månaders (5/5)
förvärvat (2/2)
läsas (2/2)
knöt (1/1)
månader (71/71)
juristens (1/1)
överförda (1/1)
tidsbestämt (8/8)
datumet (2/2)
utreda (5/5)
fest (3/3)
populär (1/1)
insamlingsställen (1/1)
daghemmen (3/3)
mellanrum (4/4)
storfurstendöme (1/1)
engelskspråkig (6/6)
anställningar (4/4)
annars (5/5)
besöket (3/3)
överföringen (1/1)
egendomen (16/16)
specialiserat (2/2)
anledningar (1/1)
agerar (1/1)
friluftsliv (4/4)
vidaredistribuera (1/1)
sättet (4/4)
gav (2/2)
barnatillsyningsmännen (1/1)
dagvårdens (2/2)
förrätta (1/1)
industri (2/2)
utrikeshandel (1/1)
påvisas (1/1)
parrådgivning (1/1)
yrkesprov (1/1)
TTS (1/1)
företagets (8/8)
dyrast (1/1)
bland (38/38)
neuvola (4/4)
lovade (1/1)
arkitektur (2/2)
preventivmetoder (1/1)
begränsningarna (4/4)
trappuppgången (1/1)
bedöms (7/7)
runtom (3/3)
hygienpass (1/1)
psykoterapeutti (1/1)
förlossningsdatumet (3/3)
skollov (1/1)
tolkar (2/2)
studerandena (1/1)
parterna (7/7)
läsesal (1/1)
samboende (1/1)
medlemskommunernas (1/1)
pappersblanketter (1/1)
klass (5/5)
orsak (7/7)
pappaledig (1/1)
Business (5/5)
perheneuvola (6/6)
syn (2/2)
funktionalitet (1/1)
äventyra (1/1)
torsdag (2/2)
närundervisning (1/1)
över (82/82)
ammatillinen (3/3)
sällskapar (1/1)
ordböckerfinska (2/2)
arbetsintyget (2/2)
dödsorsaken (2/2)
sistnämnda (1/1)
samborna (3/3)
jobbsökning (4/4)
levereras (1/1)
sopsortering (1/1)
hälsovårdssamkommun (7/7)
islamska (1/1)
färdtjänster (1/1)
uppleva (1/1)
förmåner (28/28)
rumänska (12/12)
församlingfinska (1/1)
lönespecifikationen (2/2)
man (251/251)
behandling (9/9)
statsgaranti (2/2)
kansalaisuusilmoitus (2/2)
utbilda (5/5)
specialyrkesexamen (3/3)
jobbsökande (2/2)
kejsarsnitt (3/3)
riskabelt (1/1)
färdigheter (22/22)
fallit (3/3)
ladda (7/7)
känner (12/12)
Suomessa (2/2)
närvarande (3/3)
skapandet (1/1)
överklaga (7/7)
arbetslivetfinska (1/1)
alternativen (1/1)
bilteknik (1/1)
överens (43/43)
tukipiste (2/2)
förorter (1/1)
peruskoulupohjainen (1/1)
urval (1/1)
pendlar (1/1)
intressant (2/2)
linkkiMiljöministeriet (1/1)
familjeförhållandena (1/1)
grundlagen (2/2)
in (81/85) In (4)
matkulturer (1/1)
församlingssammansutning (1/1)
val (13/16) Val (3)
korkein (1/1)
fem (24/24)
studera (89/89)
aborten (1/1)
utbildningsprogrammen (2/2)
VSB (1/1)
redogörelse (5/5)
hudfärg (3/3)
människovärde (1/1)
mån.-fre. (4/4)
vuxenutbildningsinstitut (4/4)
beskattningsbeslut (1/1)
ränta (1/1)
försäkringar (9/9)
statsstöd (1/1)
insjöar (1/1)
lättare (6/6)
traumatiska (1/1)
Kyrkbacken (1/1)
något (71/71)
vården (11/11)
himmelsfärd (1/1)
studenthem (1/1)
problemfinska (2/2)
anslagstavlor (1/1)
komma (53/53)
fackliga (1/1)
föräldradagpenning (5/5)
smärtlindring (1/1)
stängd (1/1)
slutarbete (2/2)
työkyvyttömyyseläke (1/1)
innehållits (1/1)
århundradet (1/1)
arbetskontrakt (1/1)
specialundervisning (5/5)
skal (1/1)
kollektivavtalet (14/14)
Gustav (3/3)
förnya (4/4)
rörelser (1/1)
rådgivningsbyråer (6/6)
originalhandlingen (1/1)
delägare (1/1)
sköter (23/23)
utgöra (4/4)
välbefinnandeområden (1/1)
magisterstudierna (1/1)
lokalförvaltningfinska (1/1)
innefattar (1/1)
kulturella (1/1)
övernatta (5/5)
fullgjort (1/1)
återvinning (6/6)
måltid (2/2)
smälter (1/1)
industrialiseringen (2/2)
rättvisa (1/1)
storindustrin (1/1)
C2 (1/1)
ingen (22/22)
huruvida (7/7)
personligen (11/11)
delat (1/1)
taitavan (1/1)
byråerfinska (1/1)
styrgrupp (1/1)
obegränsad (2/2)
krigsskadeståndet (1/1)
lite (11/11)
velkaneuvonta (1/1)
dagtid (3/3)
seniorrådgivningen (4/5) Seniorrådgivningen (1)
MB (10/10)
MERCURIA (1/1)
rådgivningstelefon (1/1)
ångest (1/1)
länderfinska (1/1)
konfessionslösa (2/2)
mödrahemsverksamheten (1/1)
nätbankskoderna (1/1)
skolhälsovårdarna (1/1)
medborgarorganisation (1/1)
bra (54/54)
brottsanmälanfinska (1/1)
medicinska (2/2)
idrott (3/3)
förtrogna (1/1)
bokbussar (1/1)
försvunnit (1/1)
tidningar (9/9)
vetenskaplig (1/1)
biblioteketfinska (2/2)
Tyskland (1/1)
sjukförsäkrad (2/2)
arbetskamraterna (1/1)
centrum (9/9)
hoidon (1/1)
kommunernas (4/4)
familjepension (5/5)
huvudstadsregionens (3/3)
Steinerskola (2/2)
garanterar (1/1)
penningunderstöd (2/2)
ansökningar (4/4)
arbetsavtalslagen (2/2)
hoitoraha (2/2)
espoo.fi (1/1)
Saarnio (2/3) saarnio (1)
översättningarna (1/1)
jämställda (3/3)
flickor (5/5)
språkkurser (3/3)
guldåldern (1/1)
tjänsteprocesserna (1/1)
åtalas (1/1)
skolväsendet (1/1)
militärunderstöd (1/1)
handelsläroanstalten (1/1)
bioprogram (1/1)
insjuknade (1/1)
teoretiska (1/1)
kollegor (3/3)
kouluterveydenhoitaja (1/1)
viga (1/1)
äts (1/1)
sysslor (1/1)
grupper (11/11)
upphängningsbygel (1/1)
resekostnaderna (2/2)
binder (2/2)
delges (1/1)
bilplatser (1/1)
sydkusten (1/1)
fritidsverksamhet (1/1)
anlitar (1/1)
arbetsplatsens (4/4)
mössa (1/1)
anlita (14/14)
könssjukdom (3/3)
studentbostad (2/2)
centralförbund (1/2) Centralförbund (1)
arbetsmarknadsstödet (1/1)
hot (12/12)
lösa (2/2)
lekparker (3/3)
ehkäisyneuvonta (1/1)
Brottsofferjourens (2/2)
församling (7/7)
biträdande (1/1)
Iso (5/5)
statsförvaltningens (5/5)
Schengenländer (1/1)
förmånen (1/1)
integrationsplaner (1/1)
arbetspensionsutdrag (1/1)
tulkkaus (1/1)
utföras (3/3)
representera (1/1)
framstegsvänligt (1/1)
kommunvalfinska (1/1)
verksamhetssätt (1/1)
sålt (1/1)
läkemedel (25/29) Läkemedel (4)
förlänga (3/3)
kemiska (1/1)
kontakter (2/2)
innehåll (5/5)
långfredagen (1/1)
fungera (2/2)
invalidpension (4/4)
skapa (7/7)
noga (13/13)
teckenspråket (1/1)
opetuksen (1/1)
Stensvik (1/1)
testamente (5/5)
fråga (68/68)
beskickningarna (1/1)
Kelviå (5/5)
seurakunnan (1/1)
föbund (1/1)
grund (122/122)
statligt (1/1)
firma (1/1)
företagshälsovårdenfinska (1/1)
besvärsanvisning (1/1)
tillnyktrings- (1/1)
Itä (1/1)
julafton (2/2)
handeln (4/4)
peruskoulutukseen (1/1)
elevernas (3/3)
byggnader (2/2)
inomhus (1/1)
påbyggnadsnivå (1/1)
Versofinska (1/1)
mental (8/9) Mental (1)
följaktligen (1/1)
representerade (4/4)
medverka (1/1)
tillfrågad (1/1)
överlåter (2/2)
åldern (11/11)
territorium (2/2)
åtgärdande (1/1)
tusen (2/2)
utbudet (3/3)
stadsdirektörer (1/1)
nätverk (9/9)
sägs (1/1)
skolorna (5/5)
arvsskattfinska (1/1)
Kafnetin (1/1)
barnkapning (1/1)
webbtjänster (2/2)
avbrott (9/9)
varandras (1/1)
västländerna (1/1)
vårdpenning (10/10)
gränssnittet (1/1)
förbundets (2/2)
arrangerar (1/1)
chatten (2/2)
fruktan (1/1)
kt (5/5)
taxin (1/1)
skolbarnfinska (3/3)
samarbete (4/4)
juridiska (6/6)
avgift (2/2)
ägaren (1/1)
Health (1/1)
användaren (2/2)
bevisa (6/6)
kroatiska (4/4)
sätter (2/2)
utan (101/101)
köpta (1/1)
datoranvändningen (1/1)
faderskapet (12/12)
bevisar (2/2)
föräldrapenningperiodens (1/1)
skattepengar (1/1)
flit (1/1)
måltidsstöd (1/1)
Inkomstregistrets (1/1)
provar (1/1)
handikapporganisationer (1/1)
RAOS (1/1)
familjeplaneringsrådgivningen (1/1)
kunnat (2/2)
världskriget (2/2)
fullständigt (1/1)
hemsidor (2/2)
hemförsäkringen (4/4)
förmånliga (3/3)
regel (7/7)
skicka (27/27)
utredning (15/15)
anställningstiden (1/1)
USA (4/4)
skickar (12/12)
visering (1/1)
skyddskårerna (1/1)
tjänste- (1/1)
underhållsbidrag (8/8)
skol- (1/1)
sagts (1/1)
driver (3/3)
smarta (1/1)
kompletteringsutbildning (1/1)
avtala (1/1)
respons (6/6)
grundas (3/3)
verksamheter (1/1)
natt (1/1)
sparas (2/2)
researrangemangen (1/1)
grädde (1/1)
adoption (3/3)
återflyttningfinska (1/1)
jag (54/54)
studiemöjligheter (5/5)
skiftarbetstillägg (1/1)
händelsen (1/1)
webbplatsens (1/1)
jobbsajt (1/1)
påsken (1/1)
Lahtis (1/1)
ungdomspolitiken (1/1)
mental- (2/2)
hotfull (1/1)
responslänk (1/1)
franska (60/60)
arvo (1/1)
insinööri (1/1)
vinster (1/1)
yrkesexamenfinska (1/1)
perheasioiden (2/2)
utevistelser (2/2)
skild (1/1)
centralsjukhus (3/3)
handpenningen (1/1)
värde (1/1)
skedda (1/1)
välsignas (1/1)
uppdragsgivare (1/1)
Maahanmuuttajanuorten (1/1)
fastlagen (1/1)
nätverket (1/1)
könssjukdomarfinska (1/1)
utför (4/4)
läkarstation (14/14)
myhelsinki.fi (1/1)
centraliserat (1/1)
religioner (3/4) Religioner (1)
missbruk (2/2)
reseersättning (1/1)
nätetfinska (1/1)
mångfald (2/2)
utsatta (2/2)
föreningen (12/14) Föreningen (2)
familjemedlem (28/30) Familjemedlem (2)
affärsidé (1/1)
kullfallna (1/1)
rimligt (2/2)
övningar (1/1)
pensionsinkomster (1/1)
hör (26/26)
eventuellt (11/11)
maksuhäiriömerkintä (1/1)
arbetskraftsutbildningen (2/2)
förbrukning (3/3)
förskolanfinska (1/1)
brottet (1/1)
vanligen (46/46)
skuldrådgivarefinska (1/1)
perustoimeentulotuki (1/1)
OYS (1/1)
änkling (2/2)
föräldradagpenningar (3/3)
tandborstar (2/2)
skyddshemmet (5/5)
insikt (1/1)
text (1/1)
anmärkning (2/2)
fängelsestraff (3/3)
enlighet (7/7)
jäte (1/1)
fackförbundet (5/5)
upplöses (1/1)
intyg (26/26)
demokratin (1/1)
delaktig (1/1)
vilka (37/37)
växelverkan (2/2)
AKAVA (1/2) Akava (1)
Rovaniemifinska (2/2)
vigselceremonin (1/1)
förvaltningsrätten (1/1)
aktiviteter (10/10)
rutter (5/5)
beredd (1/1)
orten (4/4)
hälsostation (37/37)
funktionsnedsättning (7/7)
Pääkaupungin (2/2)
uppsägningen (1/1)
hälsofrämjande (1/1)
Kampen (2/2)
familjecenter (1/1)
tillväxtföretagare (2/2)
kulturföreningar (2/2)
-lokaler (1/1)
avsätta (1/1)
motionstjänsternafinska (1/1)
utlåtande (9/9)
husbolagets (2/2)
språkexamen (10/10)
tiden (25/25)
undersöker (3/3)
myndigheterna (16/16)
hälsovårdstjänsterfinska (1/1)
förskottsskatt (1/1)
begravas (3/3)
skyldighet (7/7)
under (232/232)
subventionerade (1/1)
missbruksproblem (6/7) Missbruksproblem (1)
gruppfamiljedaghem (4/4)
Elfvik (1/1)
viktigt (30/30)
tillträde (2/2)
Nylandfinska (1/1)
helsingforsare (1/1)
registreringsblanketten (1/1)
idrottsanläggningarna (1/1)
lönesystemet (1/1)
webbläsarinställningar (1/1)
invånare (45/45)
studentbostadsstiftelser (1/1)
sent (4/4)
motsvarighet (2/2)
lastensuojelu (1/1)
presidenten (3/3)
finansrådgivningen (1/1)
läsårsavgiften (2/2)
förvaltningen (2/2)
kejsare (1/1)
etc (1/1)
enfas (2/2)
arbetstider (5/5)
arbetstagarens (5/5)
förskottsuppbördsregister (1/1)
applikationsbutiken (1/1)
minimibelopp (1/1)
dagen (15/15)
familjeträning (1/1)
visumfritt (2/2)
inlärnings- (1/1)
arbetsförsök (1/1)
förbjudet (2/2)
skilt (3/3)
skåp (1/1)
Noux (1/1)
tillstånden (1/1)
vardagsum (1/1)
takt (2/2)
inkassobyrån (1/1)
författningar (1/1)
grundlagenfinska (1/1)
turvakaukalo (1/1)
välgrundad (3/3)
arbetsavtal (8/8)
menyn (1/2) Menyn (1)
handelsregisterutdraget (1/1)
brottsligt (1/1)
SOS (1/1)
krav (4/4)
akuta (5/5)
kierrätys.info (1/1)
Mariegatan (1/1)
akutvården (1/1)
Nuorisoasuntoliitto (1/1)
handarbete (4/4)
oikeus (1/1)
ositus (1/1)
nedsättande (2/2)
invandrararbetefinska (1/1)
finskt (30/34) Finskt (4)
hända (2/2)
ställas (3/3)
Akademi (1/1)
regionkontor (1/1)
hälsotillstånd (7/7)
underskrift (2/2)
Villa (1/1)
snittbetyg (1/1)
handikapptjänster (2/2)
ägodelar (2/2)
makans (1/1)
verksamhet (40/40)
Västerkulla (1/1)
urologiska (1/1)
vårdinrättning (2/2)
posta (3/3)
webbplatserna (1/1)
moderskapsunderstöd (6/6)
flaskor (1/1)
serviceproducent (1/1)
bibliotekarienfinska (1/1)
innehåller (14/14)
latauspiste (1/1)
skrift (1/1)
ställena (1/1)
närliggande (2/2)
sjukvård (8/8)
asumisoikeusmaksu (1/1)
tills (16/16)
förstår (1/1)
infödda (1/1)
förstå (2/2)
tillsvidare (6/6)
holländska (10/10)
bromsas (1/1)
hallitus (1/1)
avlönat (1/1)
poliisi (1/1)
högutbildade (1/1)
infektion (1/1)
bristfälliga (1/1)
akademiska (1/1)
avlyssnas (1/1)
bilplats (1/1)
naturhuset (1/1)
sömnskola (1/1)
justitieministeriets (2/2)
Ylikylä (1/1)
rullstol (1/1)
familjer (25/28) Familjer (3)
tillhandahåller (19/19)
orättvist (1/1)
natur (1/1)
svenskan (2/2)
pensionärsrabatten (1/1)
guld (1/1)
avtalad (2/2)
stadslotsen (1/1)
C1 (1/1)
dåligt (1/1)
keskus (1/1)
sex (22/22)
MoniNets (4/4)
motionsslingorna (1/1)
metall (1/1)
avausleikkaus (2/2)
fortbildar (1/1)
MoniNet (4/4)
förråd (1/1)
grundskolorna (1/1)
barnlöst (1/1)
bastuugn (2/2)
måla (1/1)
semester (4/4)
säkerhets- (1/1)
landet (32/32)
begravningfinska (1/1)
regeringenfinska (1/1)
trafiken (2/3) Trafiken (1)
likaså (2/2)
undernivåer (1/1)
invånarantal (1/1)
familjepensionen (1/1)
arbetat (10/10)
drogfritt (1/1)
utträda (1/1)
enkelt (2/2)
Uusi (1/1)
expertråd (1/1)
skattmyndigheten (1/1)
skyldigheter (23/23)
gravkontor (1/1)
ELY (1/1)
bidraget (2/2)
lyhytkurssi (1/1)
öppet (38/39) Öppet (1)
inträdesprov (2/2)
nämna (1/1)
övertygelse (5/5)
investerat (1/1)
fattar (15/15)
grundats (2/2)
riksdagenfinska (1/1)
invandrafamiljer (1/1)
godtar (1/1)
Koivuhaan (1/1)
räntan (2/3) Räntan (1)
populäraste (1/1)
Romppu (1/1)
myndighetens (2/2)
tvingande (2/2)
basis (11/11)
underhållsförmåga (2/2)
bostadsbidraget (3/3)
internetionellt (1/1)
tydliga (1/1)
skräpa (1/1)
ena (16/16)
bytas (1/1)
järnvägsstation (1/1)
kortvariga (2/2)
grundat (2/2)
drabbats (1/1)
aluekoordinaattori (2/2)
lånet (7/7)
jämlikt (4/4)
slutar (9/9)
receptbelagda (1/1)
förbjuden (2/2)
dagstidningar (2/2)
invandrareleverna (1/1)
diskriminerings- (2/2)
Seremoniat (1/1)
ikäihmisten (1/1)
allmänhet (10/10)
tillkalla (1/1)
borgen (6/6)
undrar (1/1)
webbaserade (1/1)
också (308/308)
rundvandringar (2/2)
sak (5/5)
tjänstetid (2/2)
daghemsföreståndarna (2/2)
invandrarföreningar (3/3)
lääkinnällinen (1/1)
sydkust (1/1)
skolbarns (4/4)
kraftig (1/1)
Studenternas (1/1)
landsvägsförbindelsermed (1/1)
tingsrätt (3/3)
työ- (3/4) Työ- (1)
riskfaktorer (1/1)
företagsformen (3/3)
dörrklocka (1/1)
hänsyn (5/5)
situationer (32/32)
bostadslösas (1/1)
kommunikationen (1/1)
kalkyleras (1/1)
lagstadgad (2/2)
kontrollen (1/1)
borgensmän (1/1)
överklagan (1/1)
samorganisation (1/1)
lågstadiets (1/1)
nödnumretfinska (1/1)
tillfällig (9/9)
samlats (1/1)
katolska (2/2)
finansiering (12/12)
närserviceprincipen (2/2)
yrkesutbildningfinska (4/4)
upprättade (1/1)
ändå (25/25)
utkomst (6/6)
mellannivån (1/1)
kuntoutuspäätös (1/1)
jouren (6/6)
inbrottstjuvar (1/1)
yrkesinstitutet (1/1)
familjerådgivningsbyråerna (1/1)
öster (2/2)
föråldrade (1/1)
gymnasie- (1/1)
isännöitsijä (1/1)
lära (21/21)
oikeusaputoimisto (4/4)
yrkesvägledning (1/1)
vigselintyg (1/1)
exempelvis (15/15)
medgivande (3/3)
Schengenvisumfinska (1/1)
rekisteröintitodistus (2/2)
juridik (2/2)
Apostilleintyg (1/1)
läkarmottagningen (3/3)
nordiskt (7/7)
Tavastehus (1/1)
anmälningsblankett (1/1)
lönar (17/17)
gjorde (1/1)
antagning (1/1)
ryskspråkiga (1/1)
tillsammans (56/56)
kortfattad (1/1)
servicebostäder (1/1)
dygn (3/3)
vakuus (1/1)
funderar (5/5)
väestötietojärjestelmä (1/1)
työntekijä (1/1)
tvärvetenskapliga (1/1)
handelsplats (1/1)
reservera (4/4)
konfidentiell (1/1)
museerna (4/4)
nättjänst (1/1)
värderingar (1/1)
stadshuset (2/2)
särskild (6/6)
besiktigas (1/1)
invandrarkvinnor (10/10)
perhe (1/1)
stads (61/61)
detta (95/95)
jobbsajter (2/2)
socialtjänst (1/1)
Anon (1/1)
individer (1/1)
arbetsvillkoret (2/2)
kansalaisopisto (2/2)
lottar (1/1)
obekvämt (1/1)
slutexamen (1/1)
vittna (1/1)
Garantistiftelsen (1/1)
tandvårdstjänsterna (1/1)
tutkiminen (2/2)
oikeusturvavakuutus (1/1)
sökanden (3/3)
Barnsjukhuset (2/3) barnsjukhuset (1)
energiavfall (2/2)
kastrullock (1/1)
flyttning (1/1)
religion (31/31)
inleds (8/8)
socialhandledarna (1/1)
överenskommit (1/1)
hjälp (183/183)
beslutat (2/2)
utsända (1/1)
lekparksträffar (1/1)
möblerade (1/1)
Suomipassi (1/1)
gonorré (1/1)
snabel (1/1)
trivsamt (1/1)
funktionellt (1/1)
pris (6/6)
terapeuten (1/1)
pågår (16/16)
skiljer (5/5)
stadsdirektören (1/1)
torgsidan (1/1)
andelslagets (3/3)
samfällighet (3/3)
av (1120/1120)
familjedagvården (2/2)
kring (9/9)
ibland (11/11)
yläkoulu (1/1)
baserade (1/1)
ung (7/7)
likadant (1/1)
koncentrationssvårigheter (1/1)
inkomstbeskattningfinska (1/1)
finlandssvenskarna (1/1)
ändring (1/1)
hav (1/1)
röstning (2/2)
Silkesportens (1/1)
visumansökan (1/1)
koder (1/1)
obetalda (2/2)
vänskapsförening (1/1)
kalendermånad (2/2)
apotek (4/4)
kostnadsersättningfinska (1/1)
cykel (1/1)
medlemsavgift (2/2)
belägna (3/3)
försämrar (1/1)
teaterstad (1/1)
webbtjänst (9/9)
september (3/3)
programmeringsgränssnitt (1/1)
giftorätt (1/1)
vuxengymnasiums (1/1)
älvar (1/1)
lågkonjunkturen (1/1)
uppföljning (1/1)
näringsbyråeran (1/1)
morbror (1/1)
offret (1/1)
bilskatten (1/1)
migration (1/1)
industriprodukter (1/1)
medborgarinstitutet (1/1)
responsen (1/1)
linkkiBybiblioteken (1/1)
idrottshallar (2/2)
slutade (1/1)
inkorporerade (1/1)
kommunikationsteknik (1/1)
frihet (1/1)
Ullava (3/3)
tjära (3/3)
boendetfinska (1/1)
vi (11/15) Vi (4)
kollektivbostäder (1/1)
Trafi (1/1)
medlem (20/20)
sjukledigheten (3/3)
ansökningens (1/1)
gemensamma (37/37)
harkinnanvarainen (1/1)
bosättningsland (1/1)
kroppsaga (2/2)
innehavarkort (1/1)
återvändande (1/1)
Veroprosentti (1/1)
brutit (2/2)
emot (13/13)
helhet (3/3)
månatligen (2/2)
ungdomsevenemang (1/1)
Estland (1/1)
Välkommen (1/1)
fiska (2/2)
utbildning (87/92) Utbildning (5)
slutbetyget (1/1)
plastföremål (1/1)
gravt (1/1)
rättigheterfinska (1/1)
viktigaste (9/9)
sig (184/184)
öppning (1/1)
konsumentens (3/3)
enklast (1/1)
Kylämaja (1/1)
politik (1/1)
räknar (1/1)
familjevåldfinska (2/2)
universitetets (2/2)
arbetslandet (1/1)
mentalvårdsenheten (1/1)
flykting (8/9) Flykting (1)
helhetsbetonade (1/1)
underteckna (4/4)
växer (2/2)
nackdel (1/1)
telefonrådgivning (3/3)
Wilma (6/6)
arbetsverksamhet (2/2)
femte (2/2)
finsk (51/51)
meta (1/1)
avstängda (1/1)
privatskolor (1/1)
vuxna (33/33)
spisfläkten (1/1)
Sveaborgs (1/1)
allaktivitetscentret (1/1)
skadegörelse (1/1)
grunderna (2/2)
åtta (3/3)
beaktande (2/2)
hyresgäster (3/3)
utgående (8/8)
fredagar (2/2)
vattenskada (5/5)
vuxenstuderande (4/4)
problematiskt (1/1)
intressebevakningsorganisation (3/3)
veronpalautus (2/2)
turistbyrå (1/1)
flera (61/61)
utfärda (6/6)
avdrag (5/5)
ekonomisk (1/1)
riksdagens (1/1)
skiljasfinska (1/1)
fyllt (29/29)
ersätta (8/8)
legalisering (2/2)
Nyland (8/8)
A1.1 (1/1)
uppförandet (1/1)
övertid (2/2)
arbetserfarenheten (1/1)
personbeskattning (1/1)
svårt (17/17)
grannmedlingscentret (1/1)
handlägger (1/1)
dagpenningen (4/4)
Torggatan (1/1)
socialservice (1/1)
elev (2/2)
åsikt (8/8)
kielenä (1/1)
Espoon (7/7)
högsommarens (1/1)
reda (22/22)
studerandefinska (5/5)
ersättas (1/1)
anställningens (3/3)
kommunikationsfärdigheter (1/1)
utomlandsfinska (2/2)
yrke (16/16)
surfplatta (1/1)
tandvårdens (2/2)
livssituationen (1/1)
premier (1/1)
musikundervisning (1/1)
förtida (3/3)
stödperson (4/4)
To (4/4)
Ab (2/2)
utfärdas (1/1)
bulgariska (6/6)
resedokument (3/3)
vederbörliga (2/2)
bild (2/2)
utrymme (1/1)
bygg (1/1)
hälsovårdsministeriets (3/3)
bereds (1/1)
uträtta (3/3)
läggning (6/6)
avancemang (2/2)
ämnet (6/6)
medlemsfamiljerna (1/1)
jourmottagning (1/1)
polikliniken (8/8)
anspråkslöshet (1/1)
saknas (2/2)
registrerat (12/12)
visumansökningsblankett (1/1)
asukastila (1/1)
tidpunkt (2/2)
papparollen (1/1)
bostadsrådgivning (1/1)
undersökas (1/1)
lunchpaus (1/1)
särskilt (15/15)
Esbo (100/100)
uppehålla (1/1)
tidsbokningssystem (1/1)
lyftanordningar (1/1)
halvsyskon (1/1)
cirka (31/31)
månadsskift (1/1)
aktiebolag (4/4)
ASE (7/7)
rutten (1/1)
överlåtits (1/1)
renoveringen (1/1)
redaktör (1/1)
finskakurs (1/1)
moder (1/1)
då (82/82)
terapi (2/2)
betraktats (1/1)
förföljelse (2/2)
låter (1/1)
högersinnade (1/1)
födelseattest (6/6)
handelsflotta (1/1)
kollektivavtal (4/4)
näringsbyråerfinska (1/1)
resa (7/7)
hyreskontrakt (2/2)
dina (112/113) Dina (1)
yrkesskola (1/1)
när (196/202) När (6)
inlärningen (1/1)
settlementföreningen (1/1)
uppvärmningen (1/1)
pyssel (1/1)
kulturcenter (1/1)
kl. (1/1)
tjänstestyrningen (1/1)
wc (1/1)
farförälder (2/2)
grannkommuner (1/1)
tidsbokning (11/11)
museums (1/1)
grundade (2/2)
önskemål (6/6)
allt (17/17)
nivån (5/5)
upptäckt (1/1)
religiöst (9/9)
beslutar (13/13)
yhdistys (1/1)
ingås (5/5)
kansainvälinen (1/1)
repertoar (1/1)
riktad (1/1)
föräldrarnas (10/10)
dagars (1/1)
uppgå (2/2)
leta (7/7)
gårdsområden (1/1)
Kunta (5/5)
ansökningsblanketter (2/2)
Grankulla (40/40)
framförd (1/1)
papper (5/5)
girering (1/1)
invandrarbyrå (2/2)
inledningsvis (1/1)
upplevt (1/1)
församlingssammanslutnings (2/2)
bostadslånet (3/3)
Religionerna (1/1)
därifrån (1/1)
officiell (4/4)
kära (1/1)
valomgången (3/3)
redaktioner (1/1)
fredag (8/8)
knapp (1/1)
postadressen (1/1)
mobilabonnemang (1/1)
vore (2/2)
utländska (17/20) Utländska (3)
torka (1/1)
hyresbostad (33/35) Hyresbostad (2)
entreprenörskap (5/5)
avioliiton (2/2)
ramen (1/1)
arbetsplatserfinska (1/1)
barnfostran (1/1)
framställningen (2/2)
instanser (2/2)
paluun (1/1)
tar (52/52)
Strandväg (1/1)
länsbaserade (1/1)
jobbfinska (1/1)
borgare (1/1)
läkarintyg (5/5)
hemkommunen (3/3)
erfarenhetstillägg (1/1)
läkemedelsförpackningen (1/1)
ställt (2/2)
hyresgästenfinska (1/1)
stickkontakt (1/1)
hjälpt (1/1)
förskoleundervisningen (13/13)
dessafinska (1/1)
kommunen (34/34)
inspiration (1/1)
principerna (1/1)
kulturcentret (1/1)
fortsatta (9/9)
Befolkningsregistercentralen (1/1)
Marthaförbundetfinska (1/1)
konstruktioner (2/2)
begravningsplatser (4/4)
försäljningsställen (1/1)
först (50/50)
hyresvärden (18/18)
förutsättningar (3/3)
Metropolias (1/1)
bostadsrättsavgifter (1/1)
familjeförhållande (1/1)
familjebostäder (1/1)
betyg (4/4)
typ (4/4)
sjukvårdstjänster (5/5)
hemresan (2/2)
strategier (1/1)
enhet (7/7)
sö (1/1)
tävlingsdeltagaren (1/1)
sysselsättning (5/5)
dagligen (1/1)
440kt (1/1)
päiväkoti (2/2)
egendomsfördelning (1/1)
granskas (1/1)
granska (1/1)
yliopistollinen (1/1)
delgivits (1/1)
kväv (1/1)
mentorprogram (1/1)
råder (2/2)
verkliga (2/2)
rederiverksamheten (1/1)
sysselsättningsplan (4/4)
undervisar (4/4)
gardinerna (1/1)
skidor (2/2)
redogörs (1/1)
ser (8/8)
ingenjör (1/1)
språkkunniga (1/1)
stadgarna (1/1)
elevens (8/8)
förmynderskap (2/2)
bruttoinkomster (1/1)
valdagen (8/8)
varsel (1/1)
pensionerad (1/1)
Bio (1/1)
välmående (3/3)
fungerande (1/1)
födelsedagar (1/1)
produkter (5/5)
etablerades (2/2)
samtalsklubbar (1/1)
liv (15/15)
kliniken (7/8) Kliniken (1)
boendeform (1/1)
koncentrerad (1/1)
forststyrelsens (1/1)
bristen (2/2)
faderskap (4/4)
baserat (4/4)
kontaktperson (1/1)
kommunala (18/18)
publicerats (3/3)
finansieringsandelar (1/1)
beskickningen (14/14)
beslut (47/47)
ordkonst (1/1)
vigseln (9/9)
klinikstiftelsens (2/2)
biografer (3/3)
husets (8/8)
funktionsförmåga (1/1)
vapaaehtoisen (1/1)
servicebostadsgrupp (1/1)
sträckte (1/1)
värdesätter (3/3)
respektera (1/1)
sättas (1/1)
faktum (1/1)
ärendehantering (2/2)
patientavgift (1/1)
bortföranden (1/1)
V (2/2)
kvotflyktingens (1/1)
Myyrinkis (1/1)
löfte (1/1)
upprättat (3/3)
intressebevakningsorganisationer (1/1)
veckor (12/12)
servicepunkt (1/1)
avses (16/16)
arabiska (59/59)
kommunicerar (1/1)
familjebandfinska (2/2)
operationen (5/5)
engångskaraktär (1/1)
snön (1/1)
idrottsplaner (2/2)
auktoriserad (1/1)
lönetillägg (1/1)
anställda (45/45)
full (4/4)
dator (5/5)
arvonlisävero (1/1)
identitetsnummer (1/1)
tvätt (1/1)
skönhetsvård (1/1)
myndighetstjänst (1/1)
kulturförening (1/1)
drivas (1/1)
hoppat (1/1)
ungdomsbostäder (5/5)
bastulaven (1/1)
växte (1/1)
tillämpas (6/6)
kuntoutuslaitos (1/1)
finnas (10/10)
baseras (1/1)
äldre- (1/1)
verkets (1/1)
gymnasiekurser (1/1)
abortti (1/1)
arrangerades (1/1)
utgifter (5/5)
helgerna (2/2)
Väestöliittos (2/2)
nämnda (3/3)
er (8/8)
farliga (2/2)
vardagen (7/7)
sosiaalineuvonta (1/1)
följ (1/1)
partiellt (2/2)
vederlagets (1/1)
visum (20/20)
nödvändigt (4/4)
slutsyn (1/1)
avgifterna (1/1)
magistratens (7/7)
brottsmålsvittnen (1/1)
skatten (2/2)
uppsägningstiden (7/7)
socialbyrå (2/2)
forskning (5/5)
hautaustoimisto (2/2)
föreslå (2/2)
vardagliga (4/4)
Silkinportin (1/1)
hem (34/34)
portugisiska (18/18)
sairauspäiväraha (2/2)
kansliet (1/1)
sökfält (1/1)
tandvårdsjouren (1/1)
kvotflyktingar (8/8)
missbrukstjänster (1/1)
tal (1/1)
Danmark (1/1)
uppge (5/5)
Andelsbanken (1/1)
integrationsrelaterade (4/4)
förbättra (12/12)
mognadsprov (2/2)
föräldraskapet (4/4)
medborgarefinska (11/11)
kunnig (1/1)
hälsovårdstjänster (23/26) Hälsovårdstjänster (3)
upplevs (1/1)
utbetalas (9/9)
vattenkonsumtionen (1/1)
företagaren (5/5)
snabba (1/1)
medborgarinstituten (1/1)
betänketiden (5/5)
statsministern (2/2)
grunderfinska (1/1)
boendefrågor (1/1)
Runeberg (1/1)
kulturevenemang (1/1)
Dövas (3/3)
nuorisoasema (1/1)
äitiysraha (2/2)
tolka (1/1)
busstation (1/1)
januari (12/12)
svårigheter (3/3)
integrationsplanen (9/9)
uppdrag (3/3)
agera (1/1)
hyresavtal (16/18) Hyresavtal (2)
volontärarbete (1/1)
erityisäitiysraha (1/1)
arbetsmiljö (1/1)
konkurrerar (2/2)
tillvalsämnen (1/1)
öva (2/2)
fördröjas (1/1)
krissituationer (8/8)
www.kopiosto.fi (1/1)
kunna (38/38)
opetustoimi (1/1)
Sammallahdenmäki (1/1)
ofta (44/44)
fristående (9/9)
Kaustarviken (1/1)
klicka (1/1)
identifiering (2/2)
esiopetus (3/3)
isländska (1/1)
grannarna (1/1)
grannen (1/1)
kedja (1/1)
huvudhälsostation (1/1)
tjänsteställen (1/1)
gällande (6/6)
beredningen (1/1)
joustava (1/1)
förteckning (5/5)
misstänkt (1/1)
kandiderar (1/1)
kväll (1/1)
förmodligen (1/1)
denna (22/23) Denna (1)
fanns (3/3)
papprullar (1/1)
parentes (1/1)
polska (13/13)
betalning (1/1)
arbetssökande (25/25)
papperslösa (6/6)
resekostnader (1/1)
uppgöra (1/1)
två (97/97)
hälft (1/1)
narkomaner (2/2)
psykoterapitjänst (1/1)
dokumentmallar (1/1)
treårigt (2/2)
utlandetfinska (1/1)
användarpanel (2/2)
grammatikövningar (1/1)
Rinteenkulmafinska (1/1)
tillsyn (1/1)
utnyttja (13/13)
bostadsrättsbostaden (1/1)
Infobankens (3/3)
bostadslånfinska (1/1)
utveckla (12/12)
toimisto (4/4)
könsidentitet (3/3)
beskickningar (10/10)
alltid (66/66)
fiskeavfall (1/1)
konsumtionsskatt (1/1)
lagarfinska (1/1)
fre. (1/1)
orterna (1/1)
peruspäiväraha (1/1)
skolpsykologerna (1/1)
närmotion (1/1)
undantagsfall (4/4)
våldet (1/1)
diskrimineringen (1/1)
familjefrågorfinska (2/2)
Nuorten (3/3)
hjälpbehovet (2/2)
beskattningsbeslutet (4/4)
byar (1/1)
når (1/1)
stödpersoner (1/1)
patientjournalen (1/1)
årfinska (2/2)
kvarter (1/1)
möbler (4/4)
arbetskraft (2/2)
Konsumentförbunds (1/1)
hälscentralsavgifter (1/1)
slovakiska (1/1)
tillfälliga (3/3)
badrum (1/1)
gatan (1/1)
valet (3/3)
pengar (10/10)
Global (7/7)
aktörer (1/1)
hon (47/47)
haft (7/7)
region (2/2)
stadinasunnot.fi (1/1)
filosofi (1/1)
bodelningsman (2/2)
finskakurser (3/3)
delägarbostäder (4/4)
territoriet (3/3)
Mt (2/2)
grundlag (2/2)
grundare (2/2)
tiderna (1/1)
vattenmätare (1/1)
asylansökan (15/15)
lång (17/17)
Smith (2/2)
heltidsstuderande (1/1)
återvinningsstation (1/1)
efternamnen (1/1)
servicecenter (1/1)
ansikte (2/2)
driftställe (1/1)
Lumo (1/1)
ärver (2/2)
informationsservice (1/1)
brett (1/1)
larmar (1/1)
redovisning (2/2)
brotten (1/1)
tidningarna (1/1)
finländarna (19/19)
bokbussarna (1/1)
makthavaren (1/1)
häxor (1/1)
invånarnas (1/1)
köpas (6/6)
Kiinteistöyhtiö (1/1)
tilläggsundervisning (2/2)
ansiotulovähennys (1/1)
motionsalternativfinska (1/1)
ämnena (1/1)
behöva (6/6)
siktar (1/1)
licentiatexamen (1/1)
Inre (4/4)
politiska (6/6)
köksskåpen (1/1)
högskolors (1/1)
nyligen (5/5)
tvillingar (1/1)
kalendern (1/1)
utkomststödfinska (1/1)
symptom (2/2)
normal (2/2)
cykelkarta (1/1)
kursen (4/4)
ovannämnda (1/1)
minuter (1/1)
märkts (1/1)
frågar (2/2)
ogift (3/3)
läge (1/1)
läkartid (4/4)
bekostas (1/1)
muntligt (2/2)
busstidtabellerna (1/1)
förhand (19/19)
hemspråksundervisning (5/5)
stärker (1/1)
östra (2/3) Östra (1)
beskattningsbeslutfinska (1/1)
byggdes (1/1)
långtidssjuka (2/2)
kvadratmeter (2/2)
persiska (25/25)
hobbymöjligheter (2/2)
pappersrecept (1/1)
sägas (2/2)
sysselsättningen (1/1)
universitets- (1/1)
kontorenfinska (1/1)
överklagar (1/1)
textfält (1/1)
bekosta (3/3)
munsjukdomar (1/1)
ungdom (1/1)
människohandelfinska (1/1)
sopbehållare (1/1)
upptäckande (1/1)
uttrycka (2/2)
sådant (16/16)
skapar (1/1)
lö (1/1)
ryskaryska (1/1)
funderingar (1/1)
kriisipalvelu (1/1)
tuki (5/5)
yhdenvertaisuus- (1/1)
diskriminerande (2/2)
vårdnadshavare (23/23)
ensam (15/15)
kollaps (1/1)
ungdomstjänsterfinska (1/1)
dagvårdenfinska (1/1)
viseringspliktigt (1/1)
anställningsvillkoren (2/2)
övernattar (1/1)
hörsel (2/2)
näringsidkare (5/5)
lekparkerna (1/1)
städa (1/1)
läsåret (2/2)
jympa (1/1)
förlossningsavdelningen (1/1)
diskmaskinen (2/2)
pålitligt (3/3)
opetus (2/2)
teckna (9/9)
startsida (1/1)
livsåskådningskunskap (2/2)
avvisa (2/2)
tecknar (2/2)
äidinkielen (1/1)
redskapet (1/1)
fås (14/14)
begränsat (1/1)
grundutbildning (2/2)
erityisammattioppilaitos (1/1)
tidsbeställningfinska (1/1)
psykiatrian (1/1)
medborgare (138/139) Medborgare (1)
arbetsmarknadsstöd (4/4)
format (4/4)
minoriteter (3/3)
om (1845/1851) Om (6)
klart (1/1)
Resultatenheten (1/1)
män (25/25)
handikappservice (2/2)
Advokatförbunds (1/1)
rätta (4/4)
självständighet (2/2)
bilaga (1/1)
separeras (1/1)
finskspråkiga (14/14)
Unionin (1/1)
näyttötutkinto (4/4)
tonåringar (1/1)
mig (3/3)
stödtjänster (6/6)
nätbankskoder (4/4)
kierratys.info (2/2)
hemhjälpfinska (1/1)
utbildningens (1/1)
ängarna (1/1)
registrerad (3/3)
förlossningssjukhuset (2/2)
enspråkiga (2/2)
Informationscentralen (2/2)
närståendevård (6/6)
evenemang (9/9)
vårdare (1/1)
bosatta (16/16)
lagringsavgifter (1/1)
modersmålsundervisning (1/1)
kommandiittiyhtiö (1/1)
arbetsplatsen (25/25)
föreningsmöten (1/1)
vårdanstalter (1/1)
kb (4/5) kB (1)
namnskylt (1/1)
möjliggör (1/1)
köpingen (1/1)
affärsmodell (1/1)
innehållen (1/1)
köpeanbud (1/1)
centralmuseetfinska (1/1)
centralen (2/2)
trots (6/6)
kommunfullmäktige (5/5)
högskola (7/7)
Osviitta (1/1)
vägar (1/1)
specifikationsdel (2/2)
Havukoski (1/1)
besökarna (1/1)
makten (4/4)
besöken (1/1)
giftermål (1/1)
skolresestödetfinska (1/1)
on (2/2)
översätta (1/1)
högskolornas (3/3)
småbarnspedagogisk (1/1)
för (1620/1622) För (2)
arbetarskydd (2/3) Arbetarskydd (1)
identitet (14/14)
byggnaderna (1/1)
sommarkollon (1/1)
serviceboende (12/12)
avoimet (2/2)
medlemskap (2/2)
förvärvsinkomstavdrag (1/1)
målarfärg (1/1)
övervakar (10/10)
E101 (2/2)
stödfunktioner (1/1)
rad (1/1)
magisterexamen (3/3)
efterskott (4/4)
modern (20/20)
proffs (2/2)
yhdenvertaisuusvaltuutettu (1/1)
jourmottagningen (17/17)
laddat (1/1)
AUS (1/1)
Begravningsbyråers (1/1)
hinner (3/3)
ungdomar (27/27)
mer (418/418)
belönas (1/1)
samhällsvetenskapliga (3/3)
söderifrån (1/1)
Yhdenvertaisuuslaki (1/2) yhdenvertaisuuslaki (1)
preventionen (1/1)
stor (10/10)
berättigar (2/2)
koulumatkatuki (1/1)
daghemfinska (1/1)
jokamiehen (1/1)
nummerserie (1/1)
föräldralediga (1/1)
Laureas (1/1)
babyn (3/3)
skilsmässan (5/5)
prick (1/1)
skapade (1/1)
elektroniska (5/5)
direkt (55/55)
ersättning (16/16)
långvarig (3/3)
väl (8/8)
avslutade (2/2)
universitetssjukhus (2/2)
vindruta (1/1)
jämlika (1/1)
använd (2/2)
inträde (3/3)
vartannat (3/3)
förödmjukande (1/1)
förklarade (1/1)
någonting (2/2)
juristhjälp (1/1)
mat (18/18)
beskattningsrätt (1/1)
judarna (1/1)
kärnkraftverket (3/3)
urspråken (1/1)
arbetslöshetskassa (9/10) Arbetslöshetskassa (1)
varken (1/1)
Vasagatan (1/1)
Vionojafinska (1/1)
kollektivavtalen (3/3)
möjlighet (23/23)
vårdartiklar (1/1)
arbetstagaren (16/16)
ordningsnummer (1/1)
armé (1/1)
tillståndsenhet (1/1)
lokal (1/1)
fullsatta (1/1)
mall (1/1)
avancerade (1/1)
Rovalas (1/1)
Ruokavirasto (1/1)
sjukhusjouren (1/1)
mångfacetterad (1/1)
kranvatten (1/1)
skrivas (3/3)
underleveransarbete (1/1)
Inkomstregistret (1/1)
recept (15/15)
öppnad (1/1)
studiepenning (2/2)
företagshälsovården (7/8) Företagshälsovården (1)
yttre (1/1)
minimilönerna (1/1)
A2.1 (1/1)
övervåningen (1/1)
läkarintyget (1/1)
siviilisäätytodistus (1/1)
Varia (3/3)
tors (5/5)
allmänna (18/18)
stödjer (5/5)
betalar (71/71)
kunnandet (2/2)
barnlösheten (1/1)
ring (10/12) Ring (2)
försäljningen (4/4)
yngre (5/5)
rådgivningen (23/23)
besvären (4/4)
betraktar (1/1)
tandläkarkontroll (2/2)
län (3/3)
invid (1/1)
betala (88/88)
läroavtalsutbildning (5/5)
finansieringen (4/4)
löntagare (1/1)
livsmedel (2/2)
dubbelexamen (1/1)
företagsform (2/2)
omständigheterna (1/1)
dennes (4/4)
ras (2/2)
penningbelopp (1/1)
ungafinska (8/8)
ogiltigt (1/1)
grundundervisningenfinska (1/1)
fadern (10/10)
bilen (6/6)
bort (4/4)
arbetsgivarförbunden (1/1)
ritualer (1/1)
kännas (1/1)
årligen (1/1)
praktiskt (1/1)
förening (9/9)
graviditet (10/10)
publiceras (1/1)
kesäyliopisto (1/1)
födelsedatum (3/3)
avsätts (1/1)
minns (4/4)
språkexaminafinska (4/4)
webbsidan (1/1)
mark (3/3)
biljettkontoren (1/1)
grannmedling (1/1)
kommunalvalet (2/2)
familjemedlems (1/1)
rådgivningstjänster (4/4)
Kervo (2/2)
kommunerer (1/1)
Päivystysapu (1/1)
krig (4/4)
FPA (94/108) Fpa (14)
bostadslån (7/7)
flytväst (1/1)
kan (1874/1875) Kan (1)
luthersk (1/1)
central (2/2)
vuxengymnasiet (5/5)
musikhus (1/1)
anhöriga (10/10)
idrottsplatser (5/5)
löneintyg (4/4)
vattenkran (1/1)
privatpersoner (8/8)
veroilmoitus (1/1)
aktiva (5/5)
sång (1/1)
Centria (1/1)
återflyttarefinska (1/1)
preventivmedelsrådgivningens (1/1)
utbildningsstöd (1/1)
ugnen (1/1)
underhållsskyldighet (2/2)
lån (23/23)
skyddshusfinska (2/2)
mielenterveysseuran (1/1)
tre (83/83)
tillståndsärenden (4/4)
representerar (6/6)
hälsostationen (38/38)
Danske (1/1)
hurudan (2/2)
sjukvårdskostnader (2/2)
fort (8/8)
teknik (2/2)
hyresavtalet (16/16)
uppehållstillståndskortet (1/1)
språken (5/5)
Hilma (1/1)
begåtts (2/2)
sevärdheter (1/1)
anrika (1/1)
specialdiakoner (1/1)
administration (1/1)
länder (36/36)
föräldraledigheten (7/7)
asuntosäätiö (2/2)
hinder (15/15)
ungdomsledarna (1/1)
misslyckades (1/1)
allmänbildande (3/3)
anmäler (14/14)
pojkes (1/1)
viktiga (7/9) Viktiga (2)
hyresgarantin (2/2)
skyldiga (4/4)
distansundervisning (1/1)
regent (1/1)
sjukdomsattack (1/1)
alla (120/120)
meddelar (4/4)
barnskyddslagen (1/1)
vapaarahoitteinen (1/1)
Startup (1/1)
kielitutkinto (3/3)
folkmängd (1/1)
biljettpriset (1/1)
öst (2/2)
lettiska (1/1)
socialverk (2/2)
glaset (1/1)
byråer (3/3)
förvärvsinkomst (2/2)
verksamhetsställen (9/9)
centralsjukhuset (1/1)
arbetarinstitutets (1/1)
avlidit (1/1)
klasserna (1/1)
varmt (2/2)
textinnehåll (1/1)
närvara (1/1)
ABC (2/2)
personbeteckningar (1/1)
förra (1/1)
HelsingforsRegionen.fi (1/2) Helsingforsregionen.fi (1)
hälsocentraler (1/1)
Apotekareförbundets (1/1)
fira (1/1)
spelproblemfinska (1/1)
arkivet (1/1)
framtidens (1/1)
studerande (52/54) Studerande (2)
intressanta (1/1)
flerfaldigt (5/5)
indelat (4/4)
lämnats (3/3)
betyder (24/24)
rimliga (1/1)
sjukvården (11/11)
tvåspråkigt (2/2)
följeslagare (1/1)
befolkning (2/2)
invånarlokalen (1/1)
belastad (1/1)
gynekologiska (2/2)
meddelandet (2/2)
sluta (6/6)
hörde (2/2)
folk (2/2)
vissa (88/88)
områdets (2/2)
stödboende (3/3)
80:e (1/1)
servicen (1/1)
utbytesstudent (2/2)
familjeledigheten (2/2)
smidig (1/1)
arbetsplatssajtfinska (1/1)
tacka (2/2)
simma (1/1)
personförsäkring (1/1)
instrument (2/2)
internet (40/61) Internet (21)
lånesumman (1/1)
inhemska (3/3)
skriftligt (27/27)
fritiden (1/1)
området (18/18)
motionsmöjligheter (2/2)
fatta (5/5)
bastuugnen (3/3)
diskriminering (37/39) Diskriminering (2)
asylansökningsblankett (1/1)
partnerskap (2/2)
godta (1/1)
insjuknat (1/1)
hälsovård (3/3)
Karlebys (2/2)
utvecklingsstörda (3/3)
kliniker (2/2)
examensinriktad (1/1)
karneval (1/1)
samarbetsområdet (1/1)
bör (18/18)
hjälpsystem (1/1)
kollektiv (1/1)
terapeut (1/1)
kopiera (2/2)
Kehitysvammahuollon (1/1)
arbetslagstiftningen (2/2)
säljas (1/1)
underskrifterna (1/1)
pensionärerfinska (1/1)
lediga (12/12)
missbrukarproblem (2/2)
stegen (1/1)
grader (3/3)
brottsoffer (1/1)
utmattade (1/1)
Dickursby (4/4)
kvarskatt (3/3)
tandläkare (8/8)
be (44/44)
fackföreningsverksamhet (1/1)
mån (16/16)
ämnesområden (1/1)
Karleby (56/56)
reliefbilder (1/1)
tips (3/3)
färdigt (2/2)
lagarna (5/5)
fött (3/3)
vårdtillägg (1/1)
livmodern (1/1)
viseringsfria (1/1)
insamlingskärl (2/2)
behandlas (28/28)
förmögen (1/1)
gränsen (1/1)
hans (10/10)
summa (4/4)
MTV3 (1/1)
Vandakanalen (1/1)
högljutt (3/3)
tolksbehovet (1/1)
flyttservice (1/1)
fackförbundsverksamhetfinska (2/2)
bostäderfinska (2/2)
frånskild (1/1)
danskonst (1/1)
cykelleder (1/1)
stödspråkfinska (1/1)
yrkesinriktad (31/31)
Vuxeninstitut (1/1)
kymppiluokka (2/2)
bilskatt (1/1)
snöa (1/1)
personaltjänsteföretag (1/1)
rehabiliteringstjänster (1/1)
undersökningar (4/4)
inkorporerades (1/1)
vågar (2/2)
äktenskapet (29/29)
Esbobor (1/1)
sopsäck (1/1)
fuktproblem (1/1)
tätskikt (1/1)
församlingens (1/1)
motioner (1/1)
databank (1/1)
Ryssland (9/9)
ungdomsbostadsföreningen (1/1)
datorn (1/1)
graviditetsmånaden (5/5)
Finnishcourses.fi (2/4) finnishcourses.fi (2)
sommartid (1/1)
släktens (1/1)
pauserna (1/1)
metron (2/2)
Chydeniusfinska (1/1)
pensionsärenden (1/1)
Centralförbundet (1/1)
läraren (3/3)
arbetslöshetsförmåner (1/1)
förälder (36/36)
högteknologiska (1/1)
missbruksfrågor (1/1)
umgängesrätt (6/6)
landfinska (1/1)
bestraffas (1/1)
kotivakuutus (1/1)
löften (1/1)
Insurance (1/1)
regionutvecklingen (1/1)
almanacksbyrå (2/2)
lapsikaappaus (1/1)
valuta (4/4)
ljus (2/2)
flest (2/2)
mannen (5/5)
Medelhavet (1/1)
säsongsarbete (2/2)
sjukdagpenningfinska (2/2)
lider (2/2)
mottagning (4/4)
behärska (1/1)
saker (27/27)
kommuner (20/20)
släkten (1/1)
kansanopisto (2/2)
tvingar (1/1)
avgångsbetyget (1/1)
serviceställe (5/5)
tvinga (8/8)
mödra- (8/8)
visa (12/12)
yrkeshögskolafinska (3/3)
CD- (1/1)
tillgängligheten (1/1)
uppsägningstid (2/2)
bostadsförmedlaren (4/4)
katastrofer (1/1)
måsta (1/1)
överenskommits (3/3)
ändras (4/4)
naken (1/1)
stödcentretfinska (1/1)
bidragen (1/1)
specialvårdspenning (1/1)
inskolning (3/3)
Mielenterveys (1/1)
Finavia (1/1)
domstolsbeslut (4/4)
havsvik (1/1)
ansvariga (5/5)
religionen (2/2)
lägre (9/9)
examina (8/8)
lönekvittona (1/1)
behörig (1/1)
äitiysavustus (2/2)
kyrkliga (5/5)
ståt (1/1)
biografens (1/1)
kristelefon (3/3)
lov (1/1)
RAMK (2/2)
säkert (3/3)
föräldrars (2/2)
befogade (1/1)
trafikeras (1/1)
byråns (13/13)
omhändertas (1/1)
slottfinska (1/1)
rubriken (8/8)
par- (1/1)
möjligt (41/41)
resekortet (2/2)
hushållfinska (1/1)
förskoleundervisningfinska (3/3)
flyktingar (14/14)
rättshjälp (5/5)
motionslokaler (1/1)
påbyggnadsutbildning (4/4)
linkkiRovaniemi (3/3)
skötseln (6/6)
Finlands (67/67)
alkuomavastuu (1/1)
tillhandahållas (1/1)
stället (2/2)
avfallet (5/5)
avlagt (38/38)
Finland (1008/1008)
diskrimineringfinska (1/1)
Livräddningsförbund (1/1)
riksdagen (2/2)
psykiskt (1/1)
förorsakat (1/1)
kort (21/22) Kort (1)
gruppmöten (1/1)
utrikesministeriets (4/4)
Ateneum (1/1)
sälja (6/6)
förutsättning (1/1)
djur (1/1)
anges (11/11)
frågorna (1/1)
festföremålet (1/1)
kunde (2/2)
ry. (1/1)
HIV (2/2)
sökandena (1/1)
nödnumret (32/32)
enheten (4/4)
utvisas (2/2)
skede (5/5)
skadats (4/4)
mångsidig (2/2)
återflyttning (1/1)
skyldigheterfinska (1/1)
källskattekort (1/1)
morgonen (7/7)
höja (4/4)
lagrar (1/1)
tingsrättfinska (2/2)
aktier (2/2)
producerar (1/1)
kontakttolkcentral (1/1)
KOSEKs (1/1)
fisket (1/1)
tisdagar (3/3)
muovi (1/1)
skyddar (1/1)
banker (3/3)
skydda (3/3)
frivilliga (4/4)
tillrådligt (1/1)
graviditetsintyg (1/1)
delen (10/10)
könssjukdomar (8/8)
pass (23/23)
samband (10/10)
språkcaféerna (2/2)
särskilda (5/5)
Vantaa (1/1)
språkkunskaper (27/28) Språkkunskaper (1)
papperspåse (1/1)
från (235/235)
andelslaget (1/1)
minst (61/61)
bibehålls (1/1)
påse (1/1)
vigseltiden (1/1)
gymnasiestudier (6/6)
rehabiliteringsbeslut (1/1)
läkarrecept (3/3)
tillståndsärende (1/1)
hade (7/7)
uppstartsföretagare (11/11)
rätten (11/11)
Klockarmalmens (1/1)
förhandla (2/2)
telefonabonnemangfinska (1/1)
lätta (1/1)
synskadadefinska (1/1)
förplikta (1/1)
EMMAfinska (1/1)
webbankkoder (4/4)
ambassad (1/1)
hurdana (6/6)
App (1/1)
Vvo (1/2) VVO (1)
hjälptelefonen (2/2)
höghusfinska (1/1)
ylioppilaskokeet (1/1)
atmosfär (1/1)
hitta (28/28)
smärtor (3/3)
ger (82/83) GER (1)
Utbildningsstyrelsen (3/3)
modersmålsprovet (2/2)
mödrahemmet (2/2)
samtal (4/4)
lääkärintodistus (1/1)
födelsedatumet (1/1)
kallelse (1/1)
ändra (6/6)
inloggning (1/1)
lättföretagande (1/1)
högt (4/4)
försörja (3/3)
skola (18/18)
ungdomscentralen (1/1)
Nödcentralsverkets (1/1)
Psykologiförbund (1/1)
konditionen (2/2)
regionkontorfinska (1/1)
livmoderhalscancer (2/2)
moderskapsförpackning (1/1)
livssituation (7/7)
säkerhetsanvisningar (1/1)
utsökningfinska (1/1)
tingsdomare (1/1)
byrån (54/54)
arabisktalande (1/1)
svars (1/1)
myndigheterfinska (1/1)
gemensam (8/8)
rusmedelsberoendefinska (2/2)
ansökningen (7/7)
välfungerande (1/1)
gårdsbyggnader (1/1)
oavbrutet (1/1)
Nuppi (3/3)
uppehållstillstånd (269/274) Uppehållstillstånd (5)
vårdkostnader (1/1)
jaktfinska (1/1)
inverkar (6/6)
väst (2/2)
undersöka (1/1)
medicineringen (1/1)
gymnasieskolorna (2/2)
oumbärliga (1/1)
avbryts (3/3)
stadgas (3/3)
uppföljningen (1/1)
Sporttia (1/1)
verklig (2/2)
toisena (1/1)
skolors (1/1)
användarråd (1/1)
somliga (1/1)
anpassningsbara (1/1)
lääkäri (2/2)
boendetid (1/1)
trästadshelheter (1/1)
teckenspråketfinska (1/1)
bilhandlare (1/1)
svarar (6/6)
löper (4/4)
säkerhet (11/11)
studielivet (1/1)
sjukvårdfinska (1/1)
språkinlärning (1/1)
aikuislukio (4/4)
patientförening (1/1)
HelsingforsHels (1/1)
förlängas (3/3)
Haartmanska (4/4)
registerstyrelsens (1/1)
klient (1/1)
flygstationen (1/1)
återvändandefinska (1/1)
utflykter (6/6)
rädda (1/1)
skolelever (1/1)
inleddes (2/2)
familjerfinska (3/3)
initiala (2/2)
småstad (1/1)
föras (2/2)
förvärvsarbete (2/2)
tatarerna (1/1)
balansera (1/1)
eftermiddagsverksamhet (3/3)
autonomt (1/1)
täcker (3/3)
krissituation (5/5)
exakt (2/2)
listan (2/2)
rehabiliteringar (1/1)
universitetfinska (6/6)
sjukdagpenning (11/11)
yrkesutbildningar (1/1)
sista (6/6)
motsvarar (11/11)
begränsar (2/2)
fastställts (5/5)
tisdag (1/1)
institution (1/1)
sexuellt (7/7)
standardblanketter (1/1)
innehas (2/2)
planeras (1/1)
myndigheten (18/18)
gick (2/2)
godkännas (1/1)
suomi (1/2) Suomi (1)
lägg (2/2)
postfack (1/1)
Project (1/1)
sin (75/75)
laitos (2/2)
lämpar (2/2)
tasa (2/3) Tasa (1)
kända (1/1)
prövas (2/2)
bostadssökandet (1/1)
graviditetstest (2/2)
planera (2/2)
motions- (1/1)
jobbsökningscoachning (1/1)
festmat (1/1)
ons. (1/1)
varandra (16/16)
-eller (1/1)
Nordplus (1/1)
dröjsmål (1/1)
hemförlossning (1/1)
koululaisten (1/1)
jurister (4/4)
fastighetsägare (1/1)
framställning (1/1)
oktoberrevolutionen (1/1)
samtalar (3/3)
samarbetar (1/1)
öppningsoperation (3/3)
tulosyksikkö (1/1)
fattas (10/10)
godtas (1/1)
kontonummerfinska (1/1)
arbetarskyddet (2/2)
eleverna (5/5)
handikappet (1/1)
skolornas (2/2)
Clinic (7/7)
köa (1/1)
bostadslösa (5/5)
obligatoriskt (3/3)
Halloween (1/1)
studielinjer (1/1)
webbplatsen (19/19)
sökandens (2/2)
skilja (3/3)
uppväxtmiljö (1/1)
kielikahvila (1/1)
brott (48/50) Brott (2)
penningspelproblemfinska (1/1)
Tammerfors (2/2)
skryter (1/1)
rödbetssallad (1/1)
märkningen (1/1)
ungdomsstationen (3/3)
kommunallagen (1/1)
kursutbudet (1/1)
metodstudier (2/2)
midsommareldar (1/1)
Tullrådgivningen (1/1)
småbarnspedagogiken (12/12)
bokhandlar (1/1)
Karlebystödet (1/1)
varifrån (1/1)
bedömningar (1/1)
främjande (2/2)
jämställdheten (1/1)
finansiera (1/1)
arvsskatt (1/1)
handikappservicen (2/2)
villasamhället (1/1)
vita (4/4)
närbibliotek (1/1)
intyget (11/11)
handikapptjänsternafinska (1/1)
Tullen (1/1)
polisstation (1/1)
anställdas (5/5)
nationella (2/2)
beviljas (36/36)
fördelning (2/2)
Domus (1/1)
rekommendabelt (1/1)
kulturhistoria (2/2)
sköterskan (1/1)
betydande (1/1)
vardags- (1/1)
förändringar (2/2)
utbildningskoncern (1/1)
visumcentral (1/1)
islam (1/1)
babyns (1/1)
hanke (1/1)
nia (2/2)
staten (8/8)
umgängesarrangemanget (1/1)
Schengenvisum (1/1)
hindrar (1/1)
intagning (1/1)
hotell (1/1)
specialfinansieringsbolag (1/1)
neutral (1/1)
missbruks- (1/1)
arbetarinstitutens (1/1)
närståendevårdfinska (6/6)
barnrådgivningsbyråns (1/1)
blev (17/17)
företagsekonomi (1/1)
grundinformation (1/1)
tandkirurgi (1/1)
bevilja (1/1)
gränssnittetfinska (1/1)
mäklararvode (1/1)
offentlig (8/8)
nyföretagarcentralerna (1/1)
resor (2/2)
ledd (5/5)
Punaisen (2/2)
färdighetsnivå (2/2)
privata (45/45)
placerar (2/2)
överlåtelse (1/1)
invandrarenheten (2/2)
äger (11/11)
startar (5/5)
handläggningsavgift (1/1)
född (1/1)
informationsmöten (3/3)
bådas (2/2)
tullmyndigheterna (1/1)
starta (17/17)
resväg (1/1)
examen (68/68)
medel (17/17)
Varias (1/1)
bostadsform (1/1)
jämnt (5/5)
fordonfinska (1/1)
faktorer (2/2)
pompa (1/1)
vanligt (9/9)
efterhand (5/5)
kommer (62/62)
livshotande (2/2)
seudun (3/3)
punktlighet (3/3)
FPA:s (55/57) Fpa:s (2)
presidentens (1/1)
årervinns (1/1)
näringsbyråerna (4/4)
utfärder (2/2)
ägande (1/1)
centraler (1/1)
oavsett (7/7)
giltiga (2/2)
register (1/1)
ersätter (12/12)
denne (3/3)
Clubs (1/1)
Aalto (2/2)
gjorda (1/1)
våldsamt (3/3)
päivystys (3/3)
rörande (3/3)
översatt (2/2)
upplagan (1/1)
luopumisilmoitus (1/1)
olycksfall (5/5)
sköta (21/21)
april (4/4)
landskommunen (1/1)
regelbundna (3/3)
Folkdans (1/1)
klassificerats (1/1)
sökmotorns (2/2)
studentkårens (1/1)
modersmålsundervisningen (1/1)
bostadsaktiebolaget (6/6)
Hörselförbundetfinska (1/1)
skattas (1/1)
tillgodoräknas (2/2)
bibehålla (2/2)
km (1/1)
Firmaxifinska (1/1)
förberedelserna (2/2)
sorgfinska (1/1)
onsdagar (4/4)
krävande (5/5)
musikgrupper (1/1)
kvällarna (1/1)
dagstidning (1/1)
Konsumentrådgivningen (1/2) konsumentrådgivningen (1)
kvällen (4/4)
stadsdelfinska (3/3)
känna (6/6)
seurakuntien (1/1)
godkänt (4/4)
Rosatom (1/1)
bilens (1/1)
International (2/2)
avgångsbetyg (5/5)
arbetspraktik (3/3)
Ambassader (2/2)
hyrt (1/1)
beskrivningar (1/1)
godkänts (3/3)
Kiasmafinska (1/1)
hälften (1/1)
riksdag (1/1)
bredvid (1/1)
syssla (2/2)
vilket (44/44)
människohandel (12/12)
nätterna (3/3)
mobilcertifikat (3/3)
staden (32/32)
rådgivare (1/1)
sjukvårdsdistrikt (3/3)
kör (1/1)
ny (12/12)
uppdatera (2/2)
kallt (3/3)
emellertid (9/9)
läkemedelfinska (1/1)
faktureringstjänst (1/1)
ökat (3/3)
Ammatilliseen (1/1)
skuldrådgivningen (1/1)
matka.fi (1/1)
utser (3/3)
ledamöter (5/5)
kommersiella (2/2)
dela (5/5)
arbetsintygfinska (1/1)
Petäjävesi (1/1)
specialfall (1/1)
gett (2/2)
diplomi (1/1)
socialarbetaren (2/2)
glasförpackningar (1/1)
onyktert (1/1)
kranen (1/1)
fasta (3/3)
tis. (1/1)
glasögon (1/1)
specialgymnasier (1/1)
uppdragsavtal (2/2)
föreningarfinska (1/1)
stadsfullmäktige (7/7)
omfattande (6/6)
växande (1/1)
bortgång (1/1)
arbetsförhållanden (3/3)
kulturell (1/1)
styrelse (2/2)
du (2752/2757) Du (5)
tema (1/1)
beskattningsärenden (1/1)
fortsatte (1/1)
miljötjänster (1/1)
rehabiliteringsbehovet (1/1)
heltidsarbete (2/2)
lager (1/1)
företagarutbildning (4/4)
litet (6/6)
förtroende (1/1)
skald (1/1)
korttidsvård (1/1)
invandrat (2/2)
elektronisk (5/5)
hobbymöjligheterna (1/1)
rf (11/11)
underuthyrning (1/1)
oklarheter (3/3)
lisä (1/1)
födelseattester (3/3)
arbetsplatserna (7/7)
makarfinska (1/1)
och (2619/2619)
serbokroatiska (1/1)
bolagsordningen (1/1)
självrisk (1/1)
motivera (1/1)
högtid (1/1)
delaktighet (1/1)
säkerheter (1/1)
besegrat (1/1)
Översättningar (1/1)
söka (138/138)
päivystysajanvaraus (1/1)
återhämtningen (3/3)
förmedlingsarvodet (3/3)
tjänst (11/11)
arbetsintervju (1/1)
förvaltning (1/1)
församlingarna (4/4)
mest (3/3)
musikskolor (1/1)
ansöks (4/4)
bebiskläder (1/1)
missbrukarefinska (2/2)
yrkenfinska (1/1)
förvärvsarbeta (3/3)
tidsbegränsat (2/2)
krigsskadestånd (1/1)
former (4/4)
diskriminera (3/3)
socialarbete (6/6)
huvudstad (3/3)
högskolor (12/13) Högskolor (1)
tidsbundet (7/7)
svenskafinska (2/2)
miljoner (1/1)
broschyren (1/1)
betydelse (1/1)
skulder (10/10)
miljöministeriet (1/1)
bytet (1/1)
ofrånkomliga (1/1)
skyddsbehov (1/1)
jobbansökan (5/5)
tagit (2/2)
arbetslöshetspenning (1/1)
tidtabeller (2/2)
tyst (3/3)
skatt (21/21)
skolbarn (2/2)
ordningsnummerfinska (1/1)
stiftelser (3/3)
invånarna (10/10)
enas (2/2)
inbyggd (1/1)
lånas (1/1)
klagar (1/1)
vintrarna (1/1)
naturvetenskapliga (2/2)
bostad (102/102)
påverkas (7/7)
verkligen (3/3)
namnändring (3/3)
hundra (1/1)
lyssna (2/2)
Rovaniemi (42/42)
inhämtat (1/1)
marknadsundersökning (1/1)
arbetets (2/2)
utbud (1/1)
musikinstitut (3/3)
hemsidorfinska (1/1)
boendefinska (1/1)
medicinsk (13/13)
hälsotjänster (3/3)
tidskrifter (3/3)
hobbygrupper (1/1)
barnförhöjningen (1/1)
onsdag (1/1)
botas (1/1)
akutmottagningen (1/1)
hälsovårdsstationen (1/1)
skrivs (4/4)
paddlare (1/1)
tillståndsansökningarfinska (1/1)
läkarstationfinska (1/1)
juridisk (7/7)
tvätten (1/1)
handpenning (1/1)
noggrant (2/2)
förskolan (4/4)
arrangeras (4/4)
åtgärder (4/4)
räknare (1/1)
firandet (1/1)
insjuknar (10/10)
arbetet (49/49)
utveckling (15/18) Utveckling (3)
påverka (25/25)
rörelsehindradefinska (1/1)
helst (23/23)
konkurrenter (1/1)
flertal (1/1)
framtid (2/2)
republiken (1/1)
övrigt (2/2)
mentalvårdstjänsterna (1/1)
resmålen (1/1)
bilskola (1/1)
avloppet (1/1)
mor- (4/4)
tidsfrist (2/2)
jobbsökningen (11/11)
strejk (1/1)
bostadsområde (4/4)
mitten (3/3)
hälso- (20/20)
kristen (1/1)
flyktinghjälp (3/3)
opiskeluterveydenhoitajat (1/1)
skäliga (4/4)
Konstskolanfinska (1/1)
studentteaters (1/1)
stiftar (1/1)
myndig (5/5)
via (103/103)
bestämmanderätt (1/1)
Kristinestad (1/1)
motionshobbyer (1/1)
avträdelseanmälan (1/1)
tuberkulosfinska (2/2)
sparat (1/1)
snabbköp (1/1)
volontärarbetefinska (1/1)
Tölö (2/2)
halsduk (1/1)
skattskyldiga (1/1)
yttra (1/1)
omänsklig (1/1)
grannländer (2/2)
kvotflyktingarfinska (1/1)
leda (1/1)
sjuksköterska (2/2)
somrarna (1/1)
bostadsförmedlingar (1/1)
musikinstitutet (1/1)
hyra (21/21)
barnpassningsservicen (1/1)
värmeaggregat (1/1)
4:e (2/2)
förbereda (2/2)
damm (1/1)
familjerådgivning (5/5)
läkar- (1/1)
familjeförening (2/2)
ungdomsväsende (1/1)
hävas (2/2)
ekonomi- (3/3)
vattendrag (3/3)
nyttiga (2/2)
Poikien (1/1)
Ceremonier (1/1)
Maahanmuuttovirasto (9/9)
skärgård (1/1)
länkar (5/5)
publicerades (1/1)
slå (3/3)
ambulans (1/1)
närstående (20/20)
voimavarakeskus (1/1)
samfundet (1/1)
uppskatta (4/4)
anor (1/1)
Simundervisnings- (1/1)
landskapsmuseumfinska (1/1)
Yritys (2/2)
sannolikt (2/2)
transvestiter (1/1)
problemsituationer (1/1)
förmånlig (2/2)
asiointipiste (1/1)
Utvecklingsstörning (1/2) utvecklingsstörning (1)
Schengenländerna (1/1)
installera (1/1)
oroliga (1/1)
arbetsgivarförbundet (1/1)
invandrartjänster (1/1)
museets (1/1)
översättas (3/3)
arbetstid (10/10)
uttryck (2/2)
värdegrunden (1/1)
initiativ (1/1)
kommanditbolaget (1/1)
äldsta (2/2)
ansökningsprocessen (1/1)
doktorsexamen (4/4)
toalettstolen (1/1)
reseplanerare (1/1)
avsedda (27/27)
familjerådgivningscentral (3/4) Familjerådgivningscentral (1)
elatustuki (1/1)
helsinki.fi (1/1)
butiker (2/2)
osittainen (1/1)
studentmössor (1/1)
blind (1/1)
föda (3/3)
transport (1/1)
utbetalad (2/2)
meddelats (1/1)
kostar (12/12)
gravid (7/7)
tågen (1/1)
lista (7/9) Lista (2)
kvinnans (2/2)
försörjer (1/1)
rådgivningsbyråns (1/1)
kuljetuspalvelu (1/1)
upphovsrättsavgifter (1/1)
år (260/260)
tjänstekollektivavtal (1/1)
kommuntilläggfinska (1/1)
sjukdagpenningen (3/3)
högskoleexamen (18/18)
före (52/52)
abikurssi (1/1)
ungdomsledare (1/1)
Böle (4/4)
rahoitusvastike (1/1)
ettdera (1/1)
körning (1/1)
Asokoditfinska (2/2)
Studieinfo.fi (9/9)
socialservicecenter (1/1)
träd (3/3)
pensionskassor (2/2)
remiss (12/12)
personligt (6/6)
studentbostadsstiftelse (6/6)
jourtidsbeställning (1/1)
pojken (2/2)
arktiska (3/3)
miljö- (1/1)
arbetspensionsanstalten (3/3)
sjukdom (20/20)
styrelsemedlem (1/1)
tjänstekollektivavtalet (1/1)
namnen (3/3)
bruksföremål (1/1)
äktenskapfinska (2/2)
språkkunskapskrav (1/1)
registrerar (7/7)
åtagit (1/1)
kvinnan (5/5)
hyresgaranti (1/1)
IHH (1/1)
uppstartsföretagarefinska (1/1)
min (5/7) Min (2)
flicka (1/1)
bostadsrättsbostadfinska (1/1)
slutföra (1/1)
lönen (16/16)
samlingar (3/3)
tolkförbunds (1/1)
affären (1/1)
tfn (16/17) Tfn (1)
sätta (1/1)
norra (2/2)
festlokal (1/1)
definierar (1/1)
integritet (3/3)
ytan (1/1)
utlandsprefix (1/1)
studiepenningen (1/1)
Kanada (1/1)
IT (1/1)
pilkning (1/1)
besök (8/8)
driva (5/5)
studiepenningens (1/1)
studieort (1/1)
hyresstöd (2/2)
sjukpenning (1/1)
rekreationsområde (1/1)
skriven (1/1)
datum (2/2)
spelberoende (3/3)
igenom (5/5)
haltijakohtainen (1/1)
sjukvårdskortetfinska (2/2)
tvungen (8/8)
daggymnasiet (1/1)
samtalspriset (1/1)
fastställs (15/15)
loss (1/1)
berättar (9/9)
stugan (1/1)
en (1442/1442)
biograf (2/2)
utgår (3/3)
förmånligast (1/1)
samt (81/81)
kvinnorfinska (1/1)
spelande (3/3)
görs (37/37)
observera (3/3)
sjukhusen (1/1)
personbeteckningen (7/7)
yrkesval (1/1)
skolan (43/43)
heller (14/14)
betjäning (3/3)
fortsätter (2/2)
preparaten (1/1)
assistans (1/1)
bestäms (6/6)
tillhandahålls (9/9)
villkor (18/18)
rf:s (3/3)
samjouren (1/1)
internetsidor (1/1)
produkt (1/1)
vuxenläroanstalter (2/2)
bistår (2/2)
finländskt (5/5)
turneringar (1/1)
betalningstiden (3/3)
bank- (1/1)
Vinge (2/2)
statsrådet (2/2)
dolda (1/1)
skyddshuset (1/1)
insatt (2/2)
brottsoffret (1/1)
kvälls- (2/2)
amatörer (1/1)
yrkesläroanstalterfinska (1/1)
värnplikt (1/1)
kunden (6/6)
grundskolebaserad (4/4)
tillräckligt (25/25)
fenomen (1/1)
barnets (93/94) Barnets (1)
preventivrådgivning (1/1)
ovanligt (1/1)
trafikreglerna (2/2)
reaali (1/1)
linkkiFörbundet (1/1)
utöka (2/2)
dagliga (12/12)
publicera (1/1)
kulturgrupper (1/1)
thai (10/10)
kundrådgivningen (1/1)
parkeringsbiljett (1/1)
halt (2/2)
uppges (3/3)
själv (93/93)
räkningen (5/5)
skaffas (1/1)
vars (20/20)
förmögnare (1/1)
transporttjänst (1/1)
sökt (3/3)
förvärvsinkomster (1/1)
tillverkningen (1/1)
turist (2/2)
föreningar (13/14) Föreningar (1)
vårdåtgärder (1/1)
samfund (17/17)
bevittnat (1/1)
det (475/476) Det (1)
handredskapsavgiften (1/1)
instans (3/3)
skeden (2/2)
EHIC (1/1)
skötandet (2/2)
olycksfallsstation (2/2)
vokabulär- (1/1)
familjens (21/21)
huvudsakliga (1/1)
detsamma (1/1)
universitetetfinska (1/1)
plan (1/1)
sortering (1/1)
utrikes (1/1)
prövotiden (2/2)
chefer (1/1)
paus (1/1)
Avara (2/2)
fönstren (2/2)
sjukhuset (17/17)
arbetslöshetsförsäkringen (2/2)
beredskap (1/1)
Twitter (1/1)
förbereds (1/1)
utmätning (3/3)
grundexamen (7/7)
kunskapscentret (1/1)
Nöteborgsfreden (1/1)
genomsnitt (4/4)
anställning (21/21)
deltid (5/5)
sjukdomen (1/1)
undertrycka (1/1)
trottoaren (1/1)
internationell (2/3) Internationell (1)
befolkningsregistret (5/5)
minimikraven (1/1)
undervisningsspråket (7/7)
anmälningsblanketten (2/2)
handledning (21/21)
prata (12/12)
filmer (8/8)
inhemsk (1/1)
NA (1/1)
skolgångsbiträde (1/1)
språkstudier (1/1)
äänioikeusrekisteri (1/1)
fingeravtryck (1/1)
jourmottagningfinska (1/1)
någondera (3/3)
bemanningsbolag (1/1)
boenderegistret (2/2)
fri (1/1)
frysen (1/1)
plastförpackningar (1/1)
synskadade (4/4)
dialekterfinska (1/1)
nivåer (7/7)
näringstjänsten (1/1)
serveras (3/3)
skaffat (1/1)
toimintaohjelma (1/1)
TyEL (1/1)
lönesättning (1/1)
handikappservicefinska (4/4)
betalda (1/1)
måste (206/206)
tälta (1/1)
köp (5/5)
social- (26/26)
PB (1/1)
psykoterapifinska (1/1)
barnförhöjning (1/1)
hel (1/1)
rundvandringarna (1/1)
vårdledigheten (2/2)
urologisk (1/1)
höga (1/1)
näst (1/1)
handelsstad (2/2)
Martinus (1/1)
finskakunskaper (1/1)
rättsväsendet (1/1)
företagsekonomiska (1/1)
platser (5/5)
västerut (1/1)
batterierna (1/1)
läser (8/8)
anonymt (2/2)
opintotuki (2/2)
studietiden (1/1)
plastleksaker (1/1)
centrala (8/8)
Helsingforstilläggetfinska (1/1)
anhörig (9/9)
systemet (1/1)
Tysklands (1/1)
kontrolleras (3/3)
gränsövergång (2/2)
medlemskommuner (1/1)
kartläggning (17/17)
jordbruk (1/1)
automatik (1/1)
innerstad (1/1)
Trafiksäkerhetsverkets (1/1)
europeiskt (2/2)
förbinder (1/1)
underskridas (1/1)
följeslagartjänstfinska (2/2)
kortvarig (4/4)
tolken (13/13)
dagvårdplats (1/1)
menar (1/1)
annorlunda (2/2)
nej (1/1)
oroar (1/1)
konstämnen (3/3)
rättshjälpfinska (1/1)
arbetsolycksfall (1/1)
Väestörekisterikeskus (1/1)
tillståndsenheter (1/1)
eld (2/2)
flyktingarfinska (3/3)
romerna (1/1)
pågå (1/1)
tingsrättenfinska (1/1)
försäkringen (4/4)
uppvisa (1/1)
fiskeredskap (1/1)
huset (4/4)
hemvårdsavgiften (1/1)
startpeng (5/5)
grekiska (2/2)
estetiska (1/1)
fientlig (1/1)
Pulkamontiefinska (1/1)
toleransen (1/1)
motionsslingor (3/3)
trivas (1/1)
kurdiska (24/24)
förutom (2/2)
notarius (1/1)
brottsanmälan (7/7)
promenader (1/1)
skyldig (10/10)
upprättar (3/3)
gång (14/14)
belysta (1/1)
talas (8/8)
räkning (3/3)
känslor (1/1)
öppnar (11/11)
rusmedelsmottagning (1/1)
flyttgodsfinska (1/1)
juristen (1/1)
underlättar (6/6)
makarnas (6/6)
sjunde (1/1)
flaggan (2/2)
både (24/24)
samfunden (1/1)
lekverksamhet (1/1)
preventivmedels- (1/1)
mottagningscenter (1/1)
jobba (2/2)
livmoderns (1/1)
kommunsidorna (1/1)
flyktingkvoten (1/1)
genomgår (1/1)
samarbetsmöjligheter (1/1)
makarna (18/18)
livligare (1/1)
hyresdeposition (2/2)
rådfråga (2/2)
bekräfta (1/1)
frånvaro (1/1)
organisera (1/1)
tandhälsan (1/1)
familjemedlemmen (1/1)
arbetslivsguide (1/1)
disponenten (3/3)
uppringd (2/2)
lekar (1/1)
invandrares (2/2)
vårdar (16/16)
fördela (2/2)
Eira (1/1)
kyrklig (2/2)
umgänge (2/2)
efterlevande (2/2)
lokaltidningen (3/3)
medicinerna (1/1)
innanför (1/1)
färger (1/1)
speciell (2/2)
funktionsförmågan (2/2)
kopior (2/2)
tryggaste (2/2)
samtycke (4/4)
koulukuraattorit (1/1)
samtalsstöd (1/1)
räntorna (1/1)
svarat (1/1)
årstiderna (2/2)
avgjorts (1/1)
hallinto (1/1)
isär (3/3)
närmast (5/5)
fördelas (1/1)
bidra (2/2)
rättegång (1/1)
tidsbokningstjänst (1/1)
mödrarådgivning (1/1)
institutioner (2/2)
kulturkontor (1/1)
låg (1/1)
formulerad (1/1)
oss (1/1)
sjukskötare (6/6)
biografen (1/1)
fysiskt (1/1)
nödläge (1/1)
kvinnorna (3/3)
familjehus (1/1)
stred (2/2)
föräldrar (37/37)
klubbar (6/6)
adresserna (1/1)
företedde (1/1)
utlänningars (1/1)
förlora (7/7)
äventyras (1/1)
socialstationen (1/1)
lampa (1/1)
fackman (1/1)
ingick (1/1)
sjukhus (31/31)
ungdomsstation (1/1)
bevåg (1/1)
föräldraskap (2/2)
nycklarna (1/1)
förläggning (1/1)
villkoren (15/15)
styrkorna (1/1)
dagverksamhet (4/4)
situation (31/31)
samjour (1/1)
intressebevakning (1/1)
födelse (10/10)
ärvs (1/1)
näringsidkande (1/1)
freelancer (1/1)
Gloet (2/2)
erkände (1/1)
arbetstagare (32/33) Arbetstagare (1)
Flerspråkiga (2/2)
vokabulär (2/2)
handikappbidrag (5/5)
närskolan (2/2)
aldrig (2/2)
parternas (1/1)
garantipensionens (1/1)
såvida (1/1)
händer (2/2)
gren (1/1)
lönearbete (3/3)
korrigerar (1/1)
Abfinska (1/1)
syns (4/4)
texttelefon (1/1)
familjelivet (1/1)
karttjänstfinska (1/1)
detalj (1/1)
social (12/12)
läkarremiss (2/2)
handarbeten (3/3)
Suomenkielisen (1/1)
utreder (10/10)
förts (1/1)
regelbundet (5/5)
Kipinä (2/2)
läroämnen (4/4)
dagar (35/35)
bostadsrättsavtal (1/1)
lektioner (2/2)
organisation (4/4)
Banvägen (1/1)
vårdledig (3/3)
specialist (6/6)
grenarna (1/1)
pedagogiskt (1/1)
Finnvera (3/3)
nyfödda (1/1)
blir (59/59)
förrättas (14/14)
invandrarmän (3/3)
fakturera (2/2)
språk (85/85)
Rösa (1/1)
österut (1/1)
upplever (7/7)
Vandafinska (1/1)
bostadsort (2/2)
sysselsättningstjänster (1/1)
hemlig (1/1)
invandrarbakgrund (5/5)
ekonomi (4/4)
tätorterna (1/1)
håll (10/10)
kombineras (1/1)
ämne (3/3)
plötsligt (4/4)
ekonomiska (22/24) Ekonomiska (2)
grannkommunen (1/1)
sidan (36/36)
Vasa (6/6)
stödja (2/2)
stridig (1/1)
2:a (1/1)
serviceplanen (1/1)
stunderna (1/1)
mamman (1/1)
stipendier (4/4)
kaksoistutkinto (1/1)
tolktjänsterna (4/4)
valts (1/1)
hjärtat (1/1)
Isyyden (1/1)
dagvård (10/11) Dagvård (1)
ambassaden (1/1)
Konttisen (1/1)
skolhälsovårdenfinska (1/1)
inkomstrelaterat (1/1)
ungdomars (1/1)
Handelsbanken (1/1)
avslag (2/2)
månatliga (1/1)
stödengelska (1/1)
www.infopankki.fi (1/1)
motionera (1/1)
hemifrån (2/2)
buffert (1/1)
letar (5/5)
kunder (5/5)
psykoterapeutens (1/1)
bostäder (38/38)
lands (5/5)
redogörelsen (1/1)
jourmottagningarna (1/1)
längd (3/3)
likvärdigt (4/4)
tjänstebehörighet (2/2)
intagna (1/1)
garantin (1/1)
kierrätyspiste (1/1)
socialbyrån (15/15)
ställs (5/5)
död (2/2)
Spa (1/1)
taasengelska (1/1)
redaktion (2/2)
Schengenland (1/1)
postfinska (1/1)
bostadsvisning (2/2)
lekpark (2/2)
skolanfinska (2/2)
flygresor (1/1)
belagt (1/1)
fots (2/2)
avboka (2/2)
skyddfinska (4/4)
flexibel (7/7)
ersättningsgill (1/1)
avbokar (1/1)
byarna (1/1)
studierfinska (2/2)
förlossningsavdelning (1/1)
uppehållstillståndet (14/14)
förhandsmeddelande (1/1)
Röda (10/15) röda (5)
arbetarskyddsfullmäktige (2/2)
företagare (51/54) Företagare (3)
Monde (1/1)
sammanslutning (1/1)
Kilo (2/2)
skyddshus (10/10)
socialskyddet (3/3)
yrkeskvalifikationer (1/1)
tunnustaminen (1/1)
näromgivning (2/2)
ansvarar (12/12)
förenings (1/1)
trafikerar (1/1)
arbetsuppgifter (8/8)
ryska (146/146)
rådgivningsbyrå (2/2)
svår (5/5)
café (1/1)
bibliotekarien (2/2)
återflyttare (2/2)
problemavfall (1/1)
varvid (1/1)
pappa (1/1)
utom (4/4)
existensminimum (2/2)
&quot; (14/14)
markägarna (1/1)
ansvarig (4/4)
presenteras (3/3)
metalli (1/1)
Företagsfinlands (2/3) FöretagsFinlands (1)
områdena (1/1)
strängare (1/1)
yrkeskunskap (1/1)
närtågen (1/1)
hittar (202/202)
Villenpirtti (1/1)
fyll (4/4)
väcker (3/3)
förbjuder (5/5)
riksväg (1/1)
Miehen (6/6)
storlek (16/16)
yrket (1/1)
toimipiste (1/1)
Företagsfinland (1/1)
sökfunktionen (1/1)
byggd (1/1)
säger (12/12)
Fpas (1/1)
utvidgar (1/1)
tjänsteman (1/1)
korrigera (1/1)
annonser (4/4)
perintövero (1/1)
aptit (1/1)
per (60/60)
-motion (1/1)
vare (5/5)
stadsbibliotek (7/7)
skidspår (2/2)
nattetid (1/1)
kontakt (51/51)
visumcentralen (1/1)
makan (8/8)
varningsmärke (1/1)
ägarskapet (1/1)
anhörigafinska (1/1)
vice (1/1)
samma (72/72)
ansökningspraxis (1/1)
teaterföreställningar (2/2)
ungdomsverksamheten (1/1)
intressen (7/7)
förpliktelser (1/1)
Sport (5/7) sport (2)
avkoppling (1/1)
kunnallisvaalit (1/1)
minderårigt (4/4)
familjsvenska (1/1)
inriktning (1/1)
Nupoli (4/4)
våldssituationer (1/1)
uttalas (1/1)
understöds (1/1)
kemikaler (1/1)
serbiska (1/1)
andel (6/6)
lutherska (19/19)
alternativt (2/2)
studiekraven (1/1)
koncernen (1/1)
Chydenius (2/2)
DVD (1/1)
adress (27/27)
Kivenkolo (5/5)
NewCo (5/5)
metallindustrin (1/1)
arbetslivsfärdigheter (2/2)
penningunderstödfinska (1/1)
synagoga (1/1)
självständig (2/2)
huvuddukar (1/1)
broschyrer (2/2)
se (16/16)
svara (1/1)
förmögenhet (3/3)
läkemedlet (3/3)
andraspråk (3/3)
födseln (4/4)
umgängesrättfinska (2/2)
slutet (14/14)
bifoga (7/7)
notering (1/1)
jämställdhet (12/14) Jämställdhet (2)
officiella (5/5)
mängd (5/5)
fara (6/6)
Norden (1/1)
semesterpenning (1/1)
västliga (1/1)
avbryta (2/2)
giltigt (12/12)
gift (12/12)
vaarallinen (1/1)
utvecklades (2/2)
vattenkranarna (1/1)
vilken (39/39)
pappersblankett (5/5)
antibiotika (1/1)
vanliga (12/12)
hyresgäst (1/1)
polisstationen (6/6)
ntresserad (1/1)
kopplas (2/2)
yttrandefrihet (1/1)
stiftelsen (2/2)
batteriinsamlingslådor (1/1)
suppleanter (1/1)
posttraumatiskt (2/2)
Mårtensdal (1/1)
munhälsovårdfinska (1/1)
detaljerna (1/1)
böcker (16/16)
varuhus (1/1)
teatrarnas (2/2)
bostadsbehov (4/4)
avlidna (4/4)
chefredaktör (2/2)
ursprung (12/12)
frivilligarbeta (1/1)
specialkompetens (1/1)
rättelserna (2/2)
Familjeledigheter (1/1)
skilsmässafinska (2/2)
stärka (1/1)
undertecknade (1/1)
egentliga (4/4)
könsminoriteterfinska (1/1)
säljs (6/6)
lokalförvaltning (3/3)
studentkår (1/1)
ansvar (8/8)
skriftligen (2/2)
Finnish (2/2)
förgiftningfinska (1/1)
era (2/2)
stämning (1/1)
rekreationsdagar (1/1)
omgivningen (1/1)
mellan (40/40)
uppenbart (1/1)
ta (117/117)
konst (11/12) Konst (1)
säkerheten (3/3)
familjeåterförening (6/6)
serviceboendefinska (1/1)
uppgjort (1/1)
översättningstjänsterfinska (1/1)
bestämmelser (2/2)
ansökte (2/2)
webbapotek (1/1)
motsvarande (5/5)
trähus (1/1)
föreningarna (1/1)
metrostationer (1/1)
telefonnumren (1/1)
hos (167/167)
Ounasälv (1/1)
rasistiska (2/2)
igång (2/2)
kaavinta (1/1)
Petikkos (1/1)
Ihmiskaupan (1/1)
servicehus (5/5)
studieresultat (1/1)
Institutet (2/3) institutet (1)
ändrade (1/1)
drogbruk (1/1)
hälsan (13/13)
läsning (2/2)
nätbankskoderfinska (1/1)
läroavtal (3/3)
förs (3/3)
uppfattas (1/1)
Internetfinska (8/10) internetfinska (2)
varannan (1/1)
bärbar (1/1)
täydennyskoulutus (1/1)
nybörjareengelska (1/1)
beroendeproblem (1/1)
uppmärksammar (1/1)
cycling (1/1)
Tankkari (1/1)
stadigvarande (45/45)
slags (17/17)
kortti (2/2)
ungas (26/26)
antagits (2/2)
posten (2/2)
vintern (7/7)
följd (5/5)
hushållspapper (2/2)
samkönade (2/2)
träffarna (1/1)
Pensionsskyddscentralen (6/6)
kultur (13/13)
servicerådgivning (1/1)
semesterdagar (1/1)
förtroendeman (4/4)
köpare (2/2)
tandklinikerna (1/1)
Rysslands (2/2)
grammatikengelska (1/1)
vårdutgifterna (1/1)
spara (2/2)
tull- (1/1)
numret (9/9)
utförs (4/4)
ungdomarfinska (2/2)
arbetarskyddfinska (2/2)
skärgårdenfinska (1/1)
storleken (4/4)
sända (1/1)
kvotflyktingarna (1/1)
övrig (2/2)
arbets- (58/59) Arbets- (1)
bostadsrättsbostad (10/11) Bostadsrättsbostad (1)
specialtjänster (1/1)
familjeförmåner (2/2)
tåg- (1/1)
förvärvats (1/1)
friare (1/1)
risker (2/2)
konserter (1/1)
uppstod (1/1)
löneutbetalningen (4/4)
utgång (1/1)
studieområden (4/4)
densamma (1/1)
stödtjänsterfinska (1/1)
lärandet (1/1)
kyrkor (1/1)
ris (1/1)
den (588/602) Den (14)
ramper (1/1)
hyresvärdar (5/5)
traditionsarbetefinska (1/1)
turistbyrån (1/1)
kotikunta (6/6)
skattenumret (3/3)
lag (37/37)
arbetsgivares (1/1)
han (44/44)
surfplattan (1/1)
vilkas (1/1)
återförenas (1/1)
Myyringin (1/1)
studierna (26/26)
beräknade (6/6)
Olkkari (1/1)
tystnadsplikt (2/2)
bilagor (6/6)
partiregistret (1/1)
trafikverkets (1/1)
make (27/27)
myndighetsärenden (1/1)
verkstäder (1/1)
lekens (1/1)
arbetsplats (27/27)
förslossningsdatumet (1/1)
gardena (1/1)
ockuperade (1/1)
studentkårer (2/2)
perioden (2/2)
sjuk- (1/1)
yrkeshögskola (18/18)
församlingars (1/1)
klarspråk (1/1)
kosthålls- (2/2)
myndighetshandlingen (1/1)
työttömyysturvan (1/1)
brottmålet (1/1)
giltighetstiden (2/2)
mödrahem (2/2)
vistats (6/6)
direktör (1/1)
hobbyer (4/4)
idrottsklubbar (6/6)
rehabiliteringspenning (2/2)
fullt (1/1)
fortfarande (9/9)
työeläkelaitokset (1/1)
bara (13/13)
undervisnings- (1/1)
bidragens (1/1)
bemötande (3/3)
servicetorget (1/1)
noggrann (2/2)
mottagit (1/1)
kulturhistorisk (1/1)
yrkesläroanstalter (6/6)
kundtjänsten (7/7)
narkotika (1/1)
kopplat (1/1)
företaget (18/18)
gränserna (2/2)
juli (7/7)
arbetssätt (1/1)
populära (4/4)
transformera (1/1)
flyg (3/3)
skilts (1/1)
upprepa (1/1)
höstens (1/1)
rötterna (1/1)
centralerna (1/1)
volym (1/1)
tjänat (1/1)
torra (2/2)
bodelning (1/1)
yrkesutbildningenfinska (1/1)
besökare (1/1)
työvoimakoulutus (1/1)
asylsökande (22/22)
abort (8/9) Abort (1)
Köpcentret (1/1)
förflyttningstillstånd (1/1)
säsongsarbetefinska (1/1)
vakuutus (2/2)
drar (1/1)
föreningsmötet (1/1)
intelligenta (1/1)
föremål (2/2)
dagvården (13/13)
fysioterapeut (1/1)
arbetslöshetskassorfinska (1/1)
kista (1/1)
förhållande (1/1)
delegation (1/1)
återresa (2/2)
orsaken (6/6)
klassen (4/4)
läsår (4/4)
anvisning (1/1)
höst (1/1)
bättre (5/5)
besökt (3/3)
servicesställen (1/1)
överväger (7/7)
samhörighet (1/1)
sköts (4/4)
fullgjorts (2/2)
fiskebyn (1/1)
sjukvårdsersättningar (1/1)
skattemedel (1/1)
garantipension (2/2)
lönerna (3/3)
arbetskraftsutbildning (18/19) Arbetskraftsutbildning (1)
kustregionerna (1/1)
Kokkolan (1/1)
ytterligare (9/9)
kvällstid (4/4)
karens (1/1)
långt (4/4)
hörselnfinska (1/1)
TV:n (1/1)
hyresförhållandet (2/2)
könen (2/2)
starka (2/2)
språkexamina (5/5)
Sportkort (1/1)
part (5/5)
startpaket (1/1)
grannmedlingfinska (1/1)
tillfälle (1/1)
leva (6/6)
nationalitet (9/9)
arbetsförmåga (1/1)
Sininauha (1/1)
försöker (6/6)
högsta (8/8)
tidigast (2/2)
lekparkernas (1/1)
pakolainen (1/1)
hurdant (4/4)
offer (24/24)
nationalparker (1/1)
uppskattar (4/4)
uppvisande (1/1)
vederlag (2/2)
livlig (1/1)
minnas (2/2)
hyreslägenheten (1/1)
storstäderna (1/1)
företags (1/1)
samarbetsavtal (2/2)
återkallande (1/1)
underhållsbidraget (4/4)
bildats (2/2)
försäljning (1/1)
positiva (1/1)
företag (101/101)
Östersjön (1/1)
yöpäivystys (2/2)
invånarantalet (1/1)
överklagas (1/1)
Spektr (1/1)
anhörigas (1/1)
händelser (5/5)
främja (9/9)
spis (1/1)
tillslutas (1/1)
Lapset (1/1)
känns (1/1)
unionenfinska (1/1)
strax (1/1)
ledamöterna (1/1)
hoppas (1/1)
rehabiliteringen (5/5)
främjar (5/5)
västeuropéer (1/1)
kultur- (2/2)
sinsemellan (1/1)
skuldrådgivare (1/1)
hårt (1/1)
gynekolog (4/4)
tycker (1/1)
salu (3/3)
näringsbyrå (14/14)
yrkena (1/1)
vikt (1/1)
varan (1/1)
ned (6/6)
nekande (1/1)
interna (1/1)
Sodankylä (1/1)
klockslaget (1/1)
inträdesprovet (2/2)
mödrarådgivningen (8/8)
omfattning (5/5)
högtidligt (1/1)
bruk (3/3)
möten (6/6)
uskonnonvapaus (1/1)
fryser (1/1)
besiktningsstationer (2/2)
kaffepaus (2/2)
socialskyddsförmåner (1/1)
tvunget (1/1)
terminen (1/1)
allmänt (6/6)
mobbad (1/1)
filmerfinska (1/1)
hemhjälp (1/1)
återvinns (1/1)
tidningsannonser (2/2)
arbetslöshetsförmånen (2/2)
cookies (1/1)
danska (2/2)
realiseringen (1/1)
skattekort (20/20)
asiointi (1/1)
tandkliniken (3/3)
arbetsuppgiften (4/4)
enligt (53/53)
musiker (1/1)
planering (2/2)
breddgraderna (1/1)
gammalt (6/6)
hyresdepositionen (3/3)
Schweiz (31/31)
chefen (1/1)
förebyggande (6/6)
sairaala (2/2)
ske (2/2)
dagvårdsavgifter (2/2)
jämlikhet (4/6) Jämlikhet (2)
föreskrivas (1/1)
herraväldet (1/1)
vistelse (9/9)
vakuutusyhtiö (1/1)
genomtänkta (1/1)
anmäla (40/40)
kompletterar (2/2)
undervisningstjänster (2/2)
arbetslagstiftningenfinska (1/1)
Setlementti (7/7)
startande (1/1)
högskolorna (7/7)
hjälptelefon (3/3)
ställningen (1/1)
familjepensionsskydd (1/1)
Monika (3/3)
jämkning (1/1)
transportera (1/1)
rösträttsregistret (6/6)
bistånd (1/1)
problematiska (5/6) Problematiska (1)
vinterlov (1/1)
sosiaalitoimisto (3/3)
möjliga (1/1)
anses (10/10)
där (110/110)
kommunikationssvårigheter (1/1)
billigaste (1/1)
regiontrafiken (1/1)
Helsingforsregionens (10/10)
informations- (2/2)
okomplicerat (1/1)
projektet (1/1)
kommunens (18/18)
namnlag (1/1)
flyktingarna (2/2)
roliga (1/1)
välityspalkkio (1/1)
disponibla (3/3)
Bredvikens (1/1)
kontorstjänster (1/1)
tigga (1/1)
ryssarna (1/1)
regeringarna (1/1)
nettolönen (1/1)
åren (6/6)
person (64/64)
magistraternafinska (1/1)
lastenvalvoja (3/3)
markägarens (1/1)
Mellersta (11/13) mellersta (2)
möjligheter (11/11)
nätverka (1/1)
adopterar (1/1)
plastförpackningarna (1/1)
koulukuraattori (1/1)
endera (4/4)
enskilde (1/1)
utlandet (13/13)
reglerna (4/4)
sjukförsäkringskort (1/1)
god (11/12) God (1)
konstarter (3/3)
språkkaféerna (1/1)
vattenånga (1/1)
midsommartraditionerna (1/1)
aning (1/1)
Sinettä (1/1)
högskolekoncern (1/1)
perioder (5/5)
midsommar (1/1)
förskrivningsrätt (1/1)
bakgaller (1/1)
fall (62/62)
muslimska (1/1)
läkemedelsbutikerna (1/1)
slussar (1/1)
sekretessplikt (2/2)
rehabiliterande (2/2)
slussa (1/1)
fysiska (4/4)
bett (2/2)
åtminstone (13/13)
Tallinn (2/2)
bostadslös (3/3)
hemförsäkring (5/5)
obegränsat (1/1)
arbetsplatser (13/13)
textning (1/1)
godkänns (3/3)
hälsa (63/69) Hälsa (6)
sommaruniversitet (2/2)
fastställer (2/2)
parkera (1/1)
mathjälp (1/1)
brännskador (1/1)
drivs (5/5)
bemötts (1/1)
yrityksen (1/1)
regiontaxi (1/1)
helgdag (1/1)
intrång (1/1)
Renlund (1/1)
antecknas (4/4)
behörighet (4/4)
omedelbar (5/5)
mot (36/36)
konstundervisningfinska (1/1)
universitetsutbildningfinska (1/1)
verksamhetsställe (6/6)
republik (2/2)
tulkkikeskus (1/1)
läget (1/1)
Luetaan (1/1)
dagvårdstjänster (2/2)
vägguttaget (1/1)
plågor (1/1)
anställdafinska (1/1)
päivälukio (1/1)
mångformigt (1/1)
tvåspråkighet (1/1)
registreras (20/20)
anställningsförhållande (1/1)
Israel (1/1)
samman (2/2)
annat (135/135)
legalisera (1/1)
gruppera (1/1)
assistent (1/1)
intygen (1/1)
Renlunds (1/1)
klinikens (5/5)
organisationen (1/1)
beloppet (5/5)
studeranden (7/7)
grundlagfinska (1/1)
insamlingsställe (1/1)
politisk (2/2)
tryggar (8/8)
Kieppi (2/2)
lör (1/1)
förlängs (3/3)
bokas (1/1)
samtliga (11/11)
trygga (8/8)
missgynnas (1/1)
ovanför (2/2)
inslag.Om (1/1)
hävs (1/1)
förbundet (2/3) Förbundet (1)
klädregler (1/1)
förbjuda (1/1)
avled (1/1)
arbetsgivarförbund (1/1)
handikapp (18/18)
kosta (1/1)
vårdplats (3/3)
utbildningssystemet (1/1)
sammanhang (2/2)
restaurangbranschen (1/1)
lyder (1/1)
befann (1/1)
stadgade (1/1)
automatiskt (7/7)
understiger (1/1)
finns (411/411)
inslag (1/1)
affärsmannen (1/1)
verben (1/1)
måltidservice (1/1)
hälsotjänsterna (3/4) Hälsotjänsterna (1)
U2 (1/1)
euro (23/23)
förfallodagen (2/2)
rehabiliteringscenter (1/1)
omständigheter (4/4)
norrsken (3/3)
naturskyddsområde (2/2)
fick (12/12)
kommuns (3/3)
visumets (1/1)
anställd (15/15)
familjepensionfinska (1/1)
upphör (18/18)
järnvägsstationer (1/1)
dess (18/18)
tillhörighet (3/3)
fåglar (1/1)
talets (1/1)
besvärlig (1/1)
bistå (2/2)
parkeringsautomat (1/1)
spanska (37/37)
största (16/16)
tietopankki (1/1)
verkosto (1/1)
mentor (2/2)
tandläkaren (3/3)
IB (1/1)
familjemedlemmar (21/21)
vårdledighet (4/4)
handledd (2/2)
webblanketten (1/1)
arbetsgivarna (4/4)
vinterkriget (1/1)
Björkby (2/2)
intressebevakningsorganisationfinska (1/1)
civiltjänstgörare (2/2)
huvudsakligen (2/2)
sitter (3/3)
partner (12/12)
Flyktingrådgivningens (1/1)
tjänstestället (11/11)
skatteräknare (1/1)
Sveaborg (2/2)
verovelvollisen (1/1)
kris (2/2)
fastställa (1/1)
ammattitutkinto (1/1)
minnesbilderna (1/1)
dyrare (11/11)
varierar (18/18)
skolarbete (1/1)
bussbolag (1/1)
försäljningsmetoderna (1/1)
plastkasse (2/2)
offentliggöra (1/1)
lämningar (1/1)
maj (1/1)
höghus (10/10)
stadsbiblioteken (1/1)
läger (3/3)
resmålet (1/1)
kontakttolkar (1/1)
landsbygden (3/3)
mödrarådgivningstjänsterna (1/1)
publikationer (1/1)
arbeten (1/1)
integrations- (2/2)
riksomfattande (4/4)
arbetarna (2/2)
finansieringsbolag (1/1)
rättigheterna (2/2)
progressiv (4/4)
Förbund (5/5)
dagvårdsplatserfinska (1/1)
utbildningskoncernfinska (1/1)
magistraten (87/88) Magistraten (1)
köpte (1/1)
anvisar (2/2)
egnahemshus (5/5)
anvisa (1/1)
tidiga (3/3)
näringsbyråer (2/2)
hyvinvoinnin (1/1)
kotoutumissuunnitelma (1/1)
filmfestival (1/1)
motionärer (1/1)
biojäte (1/1)
r.f. (4/4)
städer (22/26) Städer (4)
utformas (1/1)
rådgivningsbyrån (21/21)
mamma (1/1)
solen (3/3)
ålderspensionsålder (1/1)
konstaktiviteter (1/1)
företagarens (3/4) Företagarens (1)
stort (8/8)
projekt (3/3)
socialjouren (2/2)
turvapaikkapuhuttelu (1/1)
tänkande (1/1)
hälsocentralsjouren (1/1)
utlänningarengelska (1/1)
banken (11/11)
pedagogik (5/5)
andelslag (6/6)
grunden (5/5)
välbefinnande (1/1)
invandrarkvinnorfinska (1/1)
lösgjorde (1/1)
kränker (1/1)
säkring (1/1)
brann (1/1)
åt (22/22)
åldersgränser (1/1)
kontaktinformation (1/1)
-kuntayhtymä (1/1)
givet (1/1)
inlärningssvårigheter (1/1)
yrkes- (2/2)
göras (29/29)
utexaminerats (1/1)
bransch (9/9)
förlossningssjukhus (1/1)
ortodoksinen (1/1)
tjänsterna (31/31)
tävlingsarrangören (1/1)
heltidsarbetande (1/1)
flyttfirmorna (1/1)
enda (1/1)
kartläggningen (14/14)
Rinteenkulma (1/1)
vetenskaps- (3/3)
preparat (1/1)
Skatteförvaltningens (9/12) skatteförvaltningens (3)
internationalisering (1/1)
misstag (1/1)
insulin (1/1)
sidorna (9/9)
Sanduddsgatan (1/1)
familjebidrag (1/1)
synnerligen (1/1)
läkemedelskostnaderna (1/1)
levt (1/1)
kartor (1/1)
springa (1/1)
fyra (26/26)
kvalitet (2/2)
stämman (1/1)
världsarven (1/1)
Bottniska (2/2)
sjukfall (3/3)
rådgivningstjänsten (1/1)
matlagning (3/3)
handläggarna (1/1)
priserna (5/5)
konkurs (3/3)
snöar (1/1)
fyrverkerierna (1/1)
ca (4/4)
valmentava (1/1)
skuldrådgivning (3/3)
löntagar- (1/1)
kommunaval (1/1)
papperspåsar (1/1)
servicehandledaren (1/1)
värkjouren (1/1)
läkarundersökning (4/4)
familjefrågor (4/4)
utländsk (15/16) Utländsk (1)
medför (1/1)
kung (4/4)
bostadfinska (3/3)
baltiska (1/1)
genomsnittliga (1/1)
tidsbokningen (5/5)
Akatemia (3/3)
pyntas (1/1)
invånarverksamheten (1/1)
kyrkans (3/4) Kyrkans (1)
medeltalet (1/1)
annonsen (2/2)
gård (1/1)
upphovsrätts- (1/1)
burmesiska (1/1)
barnens (7/7)
hoitotakuu (1/1)
medelhög (1/1)
boende (44/48) Boende (4)
utexamineras (1/1)
dansa (3/3)
arbetslöshetstförmån (1/1)
avgör (3/3)
Loktorget (2/2)
Helsingforsfinska (9/9)
varorna (1/1)
ungerska (8/8)
evenemangskalendrarna (3/3)
formen (1/1)
Kärlek (1/1)
hus (7/7)
viken (3/3)
fortsatt (13/15) Fortsatt (2)
ungdomspsykiatriska (1/1)
fiske (3/3)
utvecklas (2/2)
resedokumentfinska (1/1)
yrkeskunnighet (7/7)
bostadsförmedlingen (1/1)
servicehandledning (1/1)
hemkommunens (1/1)
hälsoundersökning (1/1)
pratar (4/4)
lånekort (1/1)
bikulturellt (1/1)
illegalt (1/1)
nuorisoasunnot (2/2)
medborgaren (1/1)
skedet (1/1)
arbetssökandefinska (2/2)
ögonkontakt (2/2)
förmedlar (2/2)
hyresvärdens (2/2)
lastensairaala (1/1)
rabatt (5/5)
företagarefinska (6/6)
grannskapet (1/1)
löpning (1/1)
semestrar (3/3)
behöver (266/270) Behöver (4)
lönebesked (1/1)
elavtal (4/4)
demensfinska (1/1)
minnesproblemen (1/1)
lånetiden (1/1)
salar (1/1)
utbytesstudier (1/1)
användningen (6/6)
kommunikation (4/4)
ansvarsområde (1/1)
klockan (10/10)
kraftiga (1/1)
inkomstrelaterade (5/5)
verksamhetscenter (2/2)
hemlands (4/4)
garantipensionen (2/2)
bästa (11/11)
tingsrätts (2/2)
mötesplatsen (1/1)
säkerhetstjänster (1/1)
tillverkning (1/1)
nedtecknas (2/2)
avfallshanteringen (1/1)
invånarinitiativ (1/1)
dagpenningenfinska (1/1)
svag (1/1)
samerna (1/1)
hittat (3/3)
förövaren (1/1)
prövotid (1/1)
omfatta (5/5)
fram (13/13)
visar (2/2)
rådgivningsbyråernas (2/2)
massörexamen (1/1)
ugriska (1/1)
återfå (1/1)
omfattas (43/43)
bröllopsdagen (1/1)
rättsskyddsförsäkring (1/1)
uppdateringen (1/1)
förseningsavgift (1/1)
ombeds (1/1)
röst (3/3)
starttiraha (1/1)
smärtjouren (1/1)
klär (1/1)
hjälpen (8/8)
högstadiet (4/4)
närståendevåld (1/1)
hemland (20/20)
ställen (3/3)
kommunal (6/6)
tillfällen (1/1)
lagenliga (1/1)
läroboken (1/1)
utomlands (61/61)
nedsatt (1/1)
biblioteken (6/6)
köpet (4/4)
rehabilitering (42/43) Rehabilitering (1)
kämpades (1/1)
cirkuskonst (2/2)
virkatodistus (1/1)
batterier (1/1)
personbolag (1/1)
fastställande (2/2)
åring (1/1)
kämpade (1/1)
ändrat (1/1)
miljöcentralerna (1/1)
medlemsland (1/1)
ungdomsarbetet (3/3)
undervisas (3/3)
förhindra (1/1)
uppbära (1/1)
rehabiliteringsplan (2/2)
samarbeta (1/1)
inresa (1/1)
Jesu (3/3)
efteråt (1/1)
ansökningstiderna (2/2)
Kylämajafinska (1/1)
kommanditbolag (4/4)
Fulbright (2/2)
sju (8/8)
förväntar (5/5)
stadenfinska (3/3)
flyktingfinska (1/1)
obetald (1/1)
dagvårdsproducenten (1/1)
skjuta (1/1)
löneperioden (1/1)
beskattas (2/2)
ljudet (1/1)
övertidstillägg (1/1)
hemlandet (2/2)
mobiltelefonens (1/1)
köper (13/13)
branschen (2/2)
sommaruniversitetets (1/1)
individuell (1/1)
livförsäkring (1/1)
ändringsarbeten (2/2)
finskspråkigt (2/2)
står (11/11)
mediciner (2/2)
bedrevs (1/1)
beskickning (16/16)
vårda (1/1)
personuppgifter (5/5)
organisationers (2/2)
vanligaste (8/8)
undertecknas (1/1)
verotoimisto (3/3)
döma (1/1)
pensionfinska (1/1)
hälsovårdenfinska (1/1)
utarbetats (1/1)
program (8/8)
ljust (1/1)
kyrkoherdeämbetet (1/1)
ofött (1/1)
arbetarskyddsdistriktet (1/1)
jobbar (1/1)
munhälsans (1/1)
avgöras (1/1)
underlättas (1/1)
missbruksproblemfinska (2/2)
utbildningsväsendet (2/2)
augusti (6/6)
traditioner (1/1)
könummer (4/4)
förvärvar (1/1)
preventivmedel (12/12)
timmarna (1/1)
skilsmässa (50/54) Skilsmässa (4)
D (1/1)
statsöverhuvud (1/1)
betjänas (1/1)
mindre (24/24)
fönstret (1/1)
betjäna (1/1)
ammattiliitto (1/1)
CV:t (2/2)
konventioner (1/1)
stöd (81/92) Stöd (11)
utvecklingsidéer (1/1)
Nuorisosäätiö (2/2)
socialväsendet (1/1)
skattekortet (6/6)
boendekostnaderna (6/6)
examenfinska (1/1)
Myyrinki (1/1)
öppna (55/55)
Quebec (1/1)
STTK (1/1)
fordon (1/1)
stambyte (1/1)
utlänningsbyrån (3/3)
producera (3/3)
namnet (2/2)
kulturarvet (1/1)
Oma (1/1)
räknas (10/10)
löneanspråk (1/1)
företagsservicecentralerna (1/1)
inskärper (1/1)
stängt (6/6)
konsertsalar (1/1)
Liechtenstein (12/12)
naturen (11/11)
arbetslöshetsförmånerfinska (1/1)
förhandlar (1/1)
Esbotillägget (1/1)
fett (1/1)
äktenskapslagenfinska (1/1)
marknaden (1/1)
yrkesutbildade (1/1)
flygplatsen (1/1)
nyttigt (2/2)
Perheiden (2/2)
förutsatt (1/1)
suomi.fi (2/3) Suomi.fi (1)
dragits (1/1)
registrerats (3/3)
servicevägledning (1/1)
tryggad (3/3)
tilläggsutbildning (3/3)
bibliotekstjänstfinska (1/1)
skador (3/3)
gentemot (2/2)
stater (2/2)
narkomaanit (1/1)
farfinska (1/1)
ålders- (1/1)
Grankullafinska (1/1)
ville (2/2)
bankärendenfinska (1/1)
företagstjänster (1/1)
svenskspråkig (8/8)
ber (1/1)
mörkare (1/1)
administrerar (1/1)
Rex (2/2)
Regionförvaltningsverket (2/2)
sorteras (1/1)
arbetarskyddsmyndigheterna (3/3)
terapibesök (1/1)
integritetsskyddet (1/1)
parförhållanden (3/3)
upplysningar (2/2)
t.ex. (18/18)
finansiärer (2/2)
äitiyspakkaus (1/1)
undersökningarna (5/5)
vårdkostnaderna (1/1)
peruskoulu (3/3)
fel (12/12)
året (19/19)
uppehållstillståndfinska (6/6)
itsehoitolääke (1/1)
ute (3/3)
följande (48/48)
materialet (4/4)
makas (4/4)
föräldrarna (51/51)
nioårig (1/1)
eftersom (19/19)
kontinuerlig (1/1)
sortera (1/1)
hyresbostaden (2/2)
barn (315/319) Barn (4)
firar (1/1)
skatterna (1/1)
tapaturmavakuutus (1/1)
julens (1/1)
beviljande (1/1)
fart (1/1)
experter (3/3)
saknar (6/6)
läs (2/2)
arbetslivet (20/20)
utlämnad (1/1)
frågorfinska (1/1)
Nylands (10/10)
utarbeta (3/3)
personen (9/9)
informellt (1/1)
vanligtvis (47/47)
centret (5/5)
högskolenivå (1/1)
huvudsak (3/3)
blommor (2/2)
bli (27/29) Bli (2)
stödåtgärder (1/1)
vattenavgift (1/1)
Livsmedelsverket (1/1)
bekantar (1/1)
Pakolaisneuvonta (2/2)
examensnivåerna (1/1)
ammattikorkeakoulu (4/4)
försvarandet (1/1)
låta (7/7)
blödande (1/1)
reser (5/5)
Åbo (7/7)
idkandet (1/1)
föds (18/18)
ombord (1/1)
kontaktuppgifterfinska (7/7)
delta (35/35)
tror (2/2)
torsdagar (2/2)
innebära (1/1)
teaterfinska (1/1)
diakoniarbetaren (1/1)
S2 (4/4)
arbetsdagen (2/2)
tillgänglig (2/2)
seniorrådgivning (1/1)
trädgårdsskötsel (1/1)
läroinrättning (2/2)
begränsad (4/4)
världen (2/2)
första (40/40)
vammaistuki (2/2)
bildkonstskolor (1/1)
banklån (4/4)
självrisken (2/2)
avstånd (1/1)
städerna (7/7)
Kela (11/11)
primärhälsovård (2/2)
motionsrutter (1/1)
handling (4/4)
bestraffning (2/2)
stjälande (1/1)
barnskyddsmyndigheterna (2/2)
företagshälsovårdens (1/1)
kapitalinkomst (1/1)
appar (2/2)
Tavataan (1/1)
nättjänsterna (2/2)
arbetafinska (2/2)
grundläggande (43/45) Grundläggande (2)
ortodox (4/4)
beträffande (2/2)
bostadsförsäljningsannonser (2/2)
räddningsverk (1/1)
behandlar (4/4)
Sveaborgsfärjorna (2/2)
upphovsrätt (6/6)
skattebyrån (13/13)
reglerar (1/1)
bibliotekskort (7/7)
åkrarna (1/1)
anknytning (2/2)
Novgorod (2/2)
industrialisering (1/1)
behålla (1/1)
sökandes (1/1)
besöksförbud (3/3)
täckande (1/1)
centralt (1/1)
sätt (44/44)
sår (1/1)
underhåll (5/5)
ry (16/16)
därom (1/1)
viitekehys (1/1)
norr (1/1)
återhämtar (3/3)
avtalade (2/2)
ihop (1/1)
existerande (1/1)
anpassa (1/1)
tomt (1/1)
museum (3/3)
huvudbiblioteket (1/1)
handikappat (8/8)
lämnar (12/12)
sökande (6/6)
maken (10/10)
Hakunilan (1/1)
uppehållstiden (1/1)
studiemiljön (1/1)
informera (1/1)
huvudpolisstation (1/1)
utlänning (2/2)
huvudstaden (2/2)
städning (1/1)
växa (2/2)
FIRMAXI (1/1)
hyrs (9/9)
besvaras (2/2)
talo (2/2)
användande (1/1)
personliga (3/3)
förkortat (1/1)
biblioteket (17/17)
utskrivna (1/1)
anställer (1/1)
kostnadsfria (11/11)
samarbetet (2/2)
varhaiskasvatuspäällikkö (1/1)
Karlebystöd (1/1)
harmoniska (1/1)
ägs (9/9)
patienten (4/4)
anställningsskyddet (1/1)
ålderfinska (1/1)
boka (57/57)
kulturer (6/6)
tjänstemän (1/1)
därefter (12/12)
faderskapserkännande (1/1)
representant (2/2)
asuntoa (2/2)
artigt (2/2)
försäkring (7/7)
följas (1/1)
besvara (1/1)
skolåldern (21/21)
medlemsländer (1/1)
könumret (1/1)
invånarparker (1/2) Invånarparker (1)
för- (1/1)
tittar (1/1)
handleder (8/8)
UNHCR:s (3/3)
Europaparlamentsval (4/4)
åriga (10/10)
landsomfattande (1/1)
rådgivningsställe (1/1)
hemlika (1/1)
tungt (1/1)
relationsrådgivning (2/2)
hushållsmaskin (1/1)
hyresboendefinska (1/1)
biometriska (1/1)
lönespecifikation (1/1)
finska (348/355) Finska (7)
familjehem (2/2)
simhallar (4/4)
bedömer (16/16)
leverans- (1/1)
byggen (1/1)
lärokurs (5/5)
påskdagen (1/1)
olaglig (1/1)
yrkeshögskolanfinska (2/2)
gravplats (1/1)
kiinteistövero (1/1)
servicepunkter (1/1)
riktnummer (1/1)
rutt (4/4)
på (1686/1687) På (1)
webbplats (174/174)
kartlägga (2/2)
hobbyverksamheter (2/2)
Nuortennettifinska (1/1)
valkrets (1/1)
texter (1/1)
avgår (2/2)
eventuell (2/2)
bekant (2/2)
motionsdosen (1/1)
veta (4/4)
tvättstuga (2/2)
dåliga (1/1)
tillåter (3/3)
kommunsidor (1/1)
vara (146/146)
landskapsplanerare (1/1)
kontot (1/1)
folkhögskolafinska (1/1)
behandlingsmetoder (1/1)
kontinuerligt (8/8)
krishjälp (1/1)
baserad (2/2)
tillsätter (1/1)
Nationalgalleriet (1/1)
Vantaalla.info (1/1)
stiftelsens (2/2)
möte (5/5)
inskrivet (1/1)
krisjour (3/3)
avsluta (1/1)
efterfrågan (1/1)
yrkeshögskolor (9/12) Yrkeshögskolor (3)
garantipensionerna (1/1)
avslutas (1/1)
tiotusentals (2/2)
avlopp (2/2)
vigselfinska (2/2)
Creative (1/1)
röra (20/20)
genomförs (2/2)
uppehållsrätt (28/28)
borde (2/2)
finländska (60/64) Finländska (4)
biljetten (1/1)
informationsförmedlare (1/1)
gruppen (5/5)
linkkiLaNuti (1/1)
änka (2/2)
bostadsaktie (2/2)
finskspråkig (3/3)
uppförs (1/1)
Valviras (1/1)
invånaren (1/1)
hundratals (1/1)
fyllda (1/1)
hemvårdsstödet (3/3)
anordnas (5/5)
ha (119/119)
svenska (890/890)
regler (5/5)
stadsbor (1/1)
Easyfinnishfinska (1/1)
de (328/335) De (7)
Reittiopas (2/2)
rekryteringen (1/1)
Ajovarmas (2/2)
dör (6/6)
tatarer (1/1)
betalningsanmärkningar (2/2)
finsk- (1/1)
kulturtjänster (2/2)
barnomsorgen (1/1)
ulkomaalaisten (1/1)
barnatillsyningsmannen (10/10)
föddes (1/1)
erforderliga (1/1)
nöjd (1/1)
Valvira (3/3)
försök (1/1)
Jourhjälpen (1/1)
EU:s (2/2)
studiematerial (1/1)
förvalta (2/2)
familjehusen (1/1)
servicenivån (1/1)
elektrisk (2/2)
frukta (1/1)
digital (1/1)
krisområden (1/1)
arbetarskyddsföreskrifterna (2/2)
inreseförbud (2/2)
läroverket (1/1)
jobbsökningfinska (1/1)
fruktar (2/2)
nordlig (1/1)
handelsmän (1/1)
lämnade (4/4)
hänvisa (1/1)
vuxensocialarbetetfinska (1/1)
enkel- (1/1)
hemma (39/39)
integrera (2/2)
etniska (3/3)
mossa (1/1)
telefonjouren (1/1)
arbetar- (1/1)
klädskåp (1/1)
institutets (7/7)
utlåtandet (3/3)
hänvisas (1/1)
resenärerfinska (1/1)
slidan (1/1)
fritt (14/14)
eleven (2/2)
avfallsåtervinningfinska (1/1)
klarar (11/11)
bestämmer (4/4)
handläggningen (2/2)
handel (1/1)
pdf (25/26) PDF (1)
göra (73/73)
påverkafinska (3/3)
hemkommuns (3/3)
förman (1/1)
nödcentralen (2/2)
försörjning (12/12)
hammashoidon (3/3)
maistraatti.fi (2/2)
korrekta (3/3)
skattedeklaration (1/1)
folkpensionerna (1/1)
baserar (1/1)
konstmuseum (2/2)
annons (1/1)
hushåll (7/7)
magisterprogram (4/4)
byggas (1/1)
behov (38/38)
bildas (4/4)
patients (1/1)
dött (2/2)
idrottshobbyer (1/1)
Kors (9/11) kors (2)
verket (9/9)
träna (1/1)
prövning (11/13) Prövning (2)
Finlandfinska (28/28)
Liikenteen (1/1)
försiktig (1/1)
fukt (2/2)
kvällar (6/6)
turism- (2/2)
studerar (21/21)
barnfamiljerfinska (2/2)
tillräckliga (25/25)
stödundervisning (3/3)
handikapprådgivningen (2/2)
viktigare (1/1)
l (3/3)
andras (3/3)
ner (4/4)
flaggdagarna (1/1)
familjerådgivningscentralen (1/1)
råkar (7/7)
mellanskillnaden (1/1)
återgå (3/3)
information (337/342) Information (5)
utövar (7/7)
studiekamrater (1/1)
bedrivs (1/1)
avlidnes (2/2)
semestern (2/2)
avlidne (4/4)
universitetskurser (1/1)
påbörjas (2/2)
kejsaren (1/1)
studieprogrammet (1/1)
närarbetets (1/1)
enskilda (6/6)
semesterresor (1/1)
kylskåpet (2/2)
fortsättare (1/1)
Liitto (4/4)
staterna (1/1)
Bostadslöshet (1/1)
förlikning (2/2)
älvarna (1/1)
Fernissan (1/1)
finansierar (1/1)
finländare (11/11)
vidare (10/10)
dekorerat (1/1)
organisationsverksamhet (1/1)
kompletteras (2/2)
timmar (14/14)
sen (1/1)
anledning (5/5)
vädret (2/2)
Pro (3/3)
låneräknare (1/1)
yrkeshögskoleexamina (1/1)
etableringsanmälan (2/2)
ordnade (1/1)
brinna (3/3)
upprätthåll (1/1)
Soite (5/5)
Europaskolan (1/1)
såsom (23/23)
betraktas (5/5)
diskuteras (1/1)
även (347/347)
nettopalkka (1/1)
kvotflykting (4/4)
möjligtvis (1/1)
skidåkning (2/2)
myndighet (11/11)
överklagande (1/1)
bekostat (1/1)
jobb (55/55)
kielioppi (1/1)
samhällsmedlem (1/1)
ordnades (1/1)
tvåspråkig (1/1)
väljas (4/4)
hälsovårdsverket (1/1)
återkallas (6/6)
privatsfär (1/1)
video (2/2)
europeiska (11/18) Europeiska (7)
lagstiftningen (6/6)
avgiftsfria (8/8)
eftermiddagen (2/2)
lyckades (2/2)
fakturor (1/1)
anspråkslös (1/1)
arbetsmarknaden (1/1)
Oulun (1/1)
förfaller (2/2)
kännedom (1/1)
status (1/1)
ihåg (25/25)
större (13/13)
webbläsare (1/1)
vaccinationerna (2/2)
Lochteå (1/1)
bolagsavtal (1/1)
föreskriver (1/1)
meddelande (4/4)
begravningsbidrag (1/1)
ämnen (10/10)
tingsrättens (5/5)
södra (5/5)
rådgivningspunkt (1/1)
sida (270/270)
affärsverksamhetsplanen (5/5)
historia (6/6)
förlossning (8/8)
böter (4/4)
omkring (1/1)
punktskriftsböcker (1/1)
privatskola (2/2)
karriären (1/1)
könsminoriteters (1/1)
franskan (1/1)
formella (1/1)
varderas (1/1)
utbildningsplats (2/2)
storprojekt (1/1)
barnuppfostran (1/1)
inkomsterna (6/6)
Komihåglista (2/4) komihåglista (2)
nybörjarkurser (1/1)
läkarutlåtande (2/2)
yrkesbevis (1/1)
tvätta (2/2)
konventionsstaterna (1/1)
Alexandersgatan (1/1)
dömas (5/5)
säsongsarbetstillstånd (1/1)
daghemsdagen (1/1)
kräver (21/21)
förföljd (2/2)
kaupunginvaltuusto (1/1)
työväenopisto (4/4)
garantier (1/1)
skolhälsovården (2/2)
tretton (1/1)
vidimera (1/1)
ärva (2/2)
smärtan (1/1)
skogsmuseumfinska (1/1)
tekniska (1/1)
påverkanfinska (1/1)
förvaltningsdomstolen (5/5)
slutfört (1/1)
luggas (1/1)
Migrationsverkets (27/27)
båtlivfinska (1/1)
England (1/1)
vetenskapsbibliotek (1/1)
integration (13/18) Integration (5)
vardera (2/2)
lagligt (5/5)
upp (67/67)
korttidsrehabilitering (1/1)
hälsovårdscentraler (1/1)
årstider (2/2)
kunskaper (27/27)
lyfta (3/3)
rättsliga (1/1)
flyktingläger (2/2)
förhandsröstningstiden (1/1)
bastu (6/6)
Esbofinska (3/3)
undervisningssektorn (1/1)
audiovisuella (1/1)
huvudansvaret (1/1)
stöds (1/1)
kommande (1/1)
betalningsanmärkning (2/2)
YTHS (1/1)
stängda (2/2)
röstar (2/2)
lunch (3/3)
lånekostnaderna (1/1)
upprätthållande (1/1)
Kuluttajansuojalaki (1/1)
sukupuolitauti (1/1)
bondgård (1/1)
sammanlagt (2/2)
stödmottagarens (1/1)
Navigatorn (5/5)
arbetspensionsutdragen (1/1)
egenfinansieringsandel (1/1)
byggbranschen (1/1)
hälsovårdare (19/19)
kartläggs (1/1)
porten (1/1)
anställningsvillkor (1/1)
Facebook (1/1)
swahili (2/2)
husdjur (1/1)
magistratet (1/1)
föräldraledig (3/3)
anställningsrådgivningen (1/1)
snabb (1/1)
Backas (1/1)
Kompetenscentret (1/1)
gymnasier (6/6)
erityishoitoraha (1/1)
råkat (4/4)
ovanliga (1/1)
jobbförmedlingssidor (2/2)
Ungdomspolikliniken (1/1)
bolag (6/6)
som (1265/1266) Som (1)
pääkaupunkiseudun (1/1)
vecka (7/7)
tvätt- (1/1)
affärsverksamheten (2/2)
Kasabergsområdet (1/1)
flygeln (1/1)
barnpassning (1/1)
åldringspension (1/1)
näringfinska (1/1)
innan (75/75)
utlänningarfinska (3/3)
Sato (2/2)
ulosotto (1/1)
nuorisopsykiatrian (1/1)
yrkesinriktade (6/6)
lagakraftvunnet (1/1)
likvidation (1/1)
lindras (1/1)
olja (1/1)
kursavgiften (2/2)
turism (4/4)
prat (2/2)
uppgifter (37/39) Uppgifter (2)
studiefärdigheter (1/1)
skogsbruksingenjör (1/1)
oppisopimustoimisto (1/1)
äldre (14/19) Äldre (5)
maka (31/31)
punktligt (1/1)
årskurser (1/1)
Eija (2/2)
egenföretagare (1/1)
verifierats (1/1)
teaterfestivaler (1/1)
gårdar (1/1)
Hautaustoimistojen (1/1)
måltidstjänst (1/1)
adresser (3/3)
svartsjuka (1/1)
vetenskap (1/1)
religionssamfunds (2/2)
priser (5/5)
-trivsel (1/1)
ansökning (5/5)
system (3/3)
studiestöd (8/8)
barns (19/23) Barns (4)
skogsindustrin (1/1)
gynekologisk (1/1)
medverkat (4/4)
uppsökande (3/3)
överbefälhavare (1/1)
elapparater (1/1)
uppskattning (2/2)
försvar (1/1)
ordnar (66/66)
vistas (35/35)
skattenummer (5/5)
alkoholdrycker (2/2)
utbildar (2/2)
kondition (1/1)
österifrån (1/1)
vattenkannor (1/1)
oåterkalleligt (1/1)
Avia (1/1)
responsiv (1/1)
gymnasieelever (1/1)
ennakonpidätys (2/2)
vuxengymnasium (12/13) Vuxengymnasium (1)
markägaren (1/1)
bouppteckningen (3/3)
cirkus (1/1)
bifaller (1/1)
tvingats (1/1)
läkaren (20/20)
sjukhusavgifter (1/1)
förhöjd (1/1)
lägga (5/5)
valt (1/1)
ska (417/417)
intagen (1/1)
kombinerat (5/5)
jourtid (1/1)
utövat (2/2)
privatvårdsstödet (1/1)
discipliner (1/1)
avvisas (1/1)
grundande (3/3)
saken (9/9)
liikenne (1/1)
läkarens (2/2)
sommarlov (1/1)
Svartskär (1/1)
styrker (2/2)
rökfria (1/1)
hålls (8/8)
berör (5/5)
empirestil (1/1)
webbankkoderna (1/1)
utbildningar (7/7)
slutit (1/1)
Kehitysvammaliittos (1/1)
länge (27/27)
tjänstemännen (2/2)
parktanterna (1/1)
vilja (1/1)
arbetspensionsutdraget (1/1)
dubbelnamn (1/1)
hemfriden (1/1)
lokala (8/8)
programmeringsgränssnittfinska (1/1)
rådgivningstjänsterna (3/3)
registerstyrelsen (5/5)
begravningsplats (8/8)
kommunicera (1/1)
spårvagnarna (1/1)
uppförande (1/1)
flyttade (6/6)
arbetslösheten (4/4)
rättegången (2/2)
frivilligt (8/8)
skattefria (1/1)
gjorts (1/1)
sairausvakuutus (4/4)
skidåkningfinska (1/1)
fördelningen (3/3)
disponent (2/2)
lyftandet (1/1)
krigen (2/2)
erbjuder (79/79)
tand- (1/1)
Europafinska (1/1)
lägenheter (1/1)
cykling (4/4)
säljaren (7/7)
land (140/140)
källskatt (1/1)
kallare (1/1)
info (8/8)
marken (1/1)
gäst (2/2)
handikappad (4/4)
registreringsintyg (2/2)
undervisningenfinska (2/2)
ungdomsgård (2/2)
insamlat (2/2)
museiområden (1/1)
kommersiellt (1/1)
förskoleenheter (1/1)
mentala (12/12)
inresereglerna (1/1)
är (1322/1322)
kielenkäyttäjän (2/2)
legaliseras (4/4)
upprätthåller (4/4)
miljöområdet (2/2)
registrera (36/36)
ländernafinska (1/1)
jaga (1/1)
situationen (14/14)
hyresvärdarnas (1/1)
rabatter (1/1)
böckerna (1/1)
hygienföreskrifter (1/1)
profil (2/2)
förutsätta (1/1)
anhörigfinska (1/1)
konstindustri (2/2)
övertidsarbete (1/1)
anlänt (2/2)
Naiset (1/1)
delägarbostad (2/3) Delägarbostad (1)
löneinkomster (2/2)
R3 (2/2)
ympärileikkaus (3/3)
känt (1/1)
lokaltidningarna (1/1)
tillbaka (6/6)
packas (2/2)
universiteten (3/3)
kiosker (4/4)
jakttillstånd (1/1)
Celia (1/1)
emigranter (2/2)
Kalkkers (1/1)
rädd (3/3)
samhället (14/14)
överlåtelseskatt (3/3)
höjs (1/1)
skadad (1/1)
utrikesministeriet (2/2)
församlingenfinska (1/1)
inleder (6/6)
anställa (3/3)
äktenskapslagen (1/1)
blivit (30/30)
tillgång (5/5)
färdig (1/1)
Linja (7/10) linja (3)
hektar (1/1)
omsorgsfullt (2/2)
höra (5/5)
socialnämnden (1/1)
rörlighet (3/3)
fysik (1/1)
vårdenheter (1/1)
HSL (2/2)
utredningar (5/5)
inlärningsresultaten (1/1)
työttömyyskassa (1/1)
bekänner (2/2)
nätet (13/13)
hobbyutbud (1/1)
kulturhus (1/1)
gymnasium (13/14) Gymnasium (1)
förvärvsarbetar (2/2)
släktband (1/1)
lokal- (1/1)
beror (42/42)
Rooska (1/1)
kallad (2/2)
barntillsynsmannen (1/1)
används (7/7)
allvarlig (1/1)
trygghet (13/13)
tilläggsstudier (1/1)
sysselsättningsstöd (2/2)
expert (1/1)
område (28/28)
startpenning (5/5)
vänner (6/7) Vänner (1)
Seniorinfo (1/1)
Laurea (2/2)
adressen (10/10)
invaliditet (1/1)
behandlats (1/1)
hjälpmedel (18/18)
studiestödfinska (1/1)
musikskolorna (1/1)
E303 (1/1)
lätt (5/5)
vägnar (1/1)
konstskola (1/1)
Australien (1/1)
backe (1/1)
Helsingforsbor (1/1)
tyska (38/38)
dagvårdsplatsen (1/1)
reklammedel (1/1)
Rovala (2/2)
gymnasieutbildningfinska (1/1)
kandidater (1/1)
heder (1/1)
medborgarna (2/2)
smidigt (1/1)
nordligaste (2/2)
koulupsykologit (1/1)
medlemmar (15/15)
språktest (1/1)
grundval (1/1)
vuxenutbildningscentra (1/1)
Foreigners (2/2)
Verso (1/1)
tvärtom (1/1)
Centralorganisation (1/1)
ekonomibranschen (2/2)
skuldrådgivningfinska (1/1)
ansöka (206/206)
moderns (7/7)
förvänta (1/1)
avfall (10/10)
utvecklingsstördafinska (1/1)
fungerar (5/5)
visumärenden (1/1)
uppehållstillståndetfinska (1/1)
kostnader (9/9)
stadigt (1/1)
utsatt (23/23)
dygnet (25/25)
begäran (6/6)
ändringar (6/6)
hemstad (2/2)
utförande (1/1)
advokat (1/1)
arbetstagarnas (5/5)
ons (3/3)
förebyggandet (1/1)
universitets (3/3)
syskon (4/4)
rullator (1/1)
ateriatuki (1/1)
fastställas (3/3)
perustuslaki (1/1)
närheten (4/4)
terveysasema (13/13)
yksityisen (1/1)
kunderna (10/10)
boendetjänster (2/2)
asylprocessens (1/1)
ingår (23/23)
faderns (4/4)
vän (7/7)
eller (1301/1301)
kurs (4/4)
förutsätter (5/5)
förverkligas (3/3)
priset (2/2)
översättar- (3/3)
klubbarfinska (1/1)
psykolog (3/3)
Vandatillägget (1/1)
lös (1/1)
gratis (22/22)
hota (1/1)
hälsocentral (1/1)
samtalet (5/5)
studietid (1/1)
sälj (1/1)
kontaktuppgifterna (15/15)
korta (4/4)
treårig (1/1)
kamratförening (1/1)
invånarhusen (1/1)
religionstillhörigheten (1/1)
Anonyymit (1/1)
liknande (2/2)
asuminen.fifinska (2/2)
välfärd (6/6)
läroanstalterna (2/2)
kerho (1/1)
yrkeshögskoleexamen (10/10)
startpengen (1/1)
tideräkningen (1/1)
kapitalinkomsten (1/1)
arbetslös (34/34)
Mejlansvägen (1/1)
tillväxt (4/4)
skriva (16/16)
tidtabellerna (1/1)
Clinic:s (1/1)
fastighet (4/4)
anslutet (2/2)
fisketillstånd (3/3)
slag (2/2)
barnskyddet (4/4)
nog (1/1)
arbetsinkomster (2/2)
identitetshandling (6/6)
uppriktighet (1/1)
letade (1/1)
utvecklingen (5/5)
bekräftande (1/1)
ärenden (58/58)
mobbning (1/1)
studenthälsovårdarna (1/1)
ingripa (3/3)
studieregisterutdrag (1/1)
längre (23/23)
työterveyshuolto (1/1)
arbetsmarknadsstödets (1/1)
betalas (44/44)
-årigt (1/1)
lämpliga (2/2)
få (338/338)
Startpunkter (1/1)
läkarcentral (1/1)
erhålla (3/3)
ansökningstid (1/1)
Vailla (1/1)
passa (1/1)
högteknologisk (1/1)
läroanstalternas (2/2)
humanitärt (1/1)
Kemi (1/2) kemi (1)
situationerfinska (1/1)
avliden (1/1)
rektorn (1/1)
bestämma (10/10)
royaltyn (1/1)
kriisipäivystys (3/3)
utbetald (1/1)
bokfinska (1/1)
inbördeskrig (1/1)
länders (5/5)
säkerställa (5/5)
psykiska (6/6)
beviljades (3/3)
räknats (1/1)
samverkan (1/1)
bostadsbyrå (1/1)
hobby (7/7)
inkludera (1/1)
men (71/71)
skorna (1/1)
språkcaféer (2/2)
kulturproducenter (1/1)
ledig (1/1)
procent (26/26)
försäkringspremier (1/1)
överenskomna (2/2)
vån (14/14)
tysta (4/4)
dagvårdsplatser (1/1)
ventilationssystem (1/1)
UNHCR (4/4)
läroavtalsbyrån (1/1)
opintolinja (1/1)
unga (72/72)
arbetsmotivation (1/1)
fiskelov (1/1)
yrkesexamen (11/11)
kartong (1/1)
kulturen (10/10)
rättshjälpen (1/1)
veckan (4/4)
fester (3/3)
samtalshjälp (4/4)
affärsförhandlingar (1/1)
bakgrundsmusik (2/2)
vaccinerar (1/1)
gott (7/7)
infödd (4/4)
aurora (1/1)
graviditetsprevention (2/2)
återvända (5/5)
upptäcks (2/2)
befriats (2/2)
fundera (8/8)
ylioppilastutkinto (1/1)
modersmål (35/35)
stöttar (1/1)
prövningsbaserat (1/1)
nationellt (1/1)
gruppfamiljedagvården (1/1)
betalat (10/10)
tolkning (3/3)
studentskrivningarna (1/1)
undantag (4/5) Undantag (1)
bollplaner (1/1)
förlovningen (1/1)
skyddshemfinska (3/3)
beslutsorganet (1/1)
majoriteten (1/1)
äktenskapengelska (1/1)
makes (5/5)
sopsorterar (1/1)
stödhandtag (1/1)
vardagsmotion (1/1)
ventilation (1/1)
undertecknar (4/4)
utgången (4/4)
utkomstskydd (9/11) Utkomstskydd (2)
tillåtna (2/2)
avläggs (1/1)
består (8/8)
yhteispäivystys (1/1)
högerextrema (1/1)
adoptera (1/1)
begått (4/4)
relationsrådgivningstjänsterfinska (1/1)
uppfylls (4/4)
betalats (3/3)
temperaturen (2/2)
medelst (2/2)
sagotimmar (1/1)
samkommunens (1/1)
överstiga (2/2)
hemfrid (1/1)
bindestreck (1/1)
övergår (1/1)
återkallats (2/2)
lär (16/16)
ibruktagande (1/1)
fast (10/10)
flesta (29/29)
verksamhetsspråk (1/1)
picknick (1/1)
hammashoito (1/1)
navigator (1/1)
House (2/2)
licentiat- (1/1)
gottgörelse (1/1)
studielinjerna (1/1)
människohandelns (2/2)
konkreta (1/1)
nästan (12/12)
period (5/5)
avstå (1/1)
slottets (1/1)
separation (1/1)
oljevärme (1/1)
ensikoti (1/1)
industrin (1/1)
tydlig (1/1)
praktikant (1/1)
Europaparlamentet (4/4)
självständighetsdagens (1/1)
ry:s (2/2)
eläke (1/1)
företagsformer (2/3) Företagsformer (1)
besiktningskontor (1/1)
steg (5/5)
företagarkurser (1/1)
camping (1/1)
skolkuratorerna (2/2)
palveluohjaaja (1/1)
Duo (1/1)
bestämda (1/1)
nöjaktiga (3/3)
utfärdat (1/1)
arbetsinkomsten (1/1)
sorteringen (1/1)
personer (96/96)
förhandsröstningsställe (1/1)
Vandas (2/2)
servicenummer (1/1)
avslå (1/1)
föregående (1/1)
bastun (4/4)
lämnat (3/3)
utbyten (1/1)
vuokrasopimus (1/1)
annanstans (10/10)
dit (6/6)
arbetsavtalfinska (1/1)
skötaren (2/2)
företagarnas (6/6)
sukupuolitautien (1/1)
lönenivån (1/1)
biogas (1/1)
rötter (1/1)
utbildningenfinska (1/1)
kontor (4/4)
bärande (1/1)
införd (1/1)
spänning (2/2)
skolresor (1/1)
bedömningsskalan (1/1)
musik (18/18)
karensen (1/1)
månaden (6/6)
angelägenheter (5/5)
videon (1/1)
parts (1/1)
undervisningsväsendet (1/1)
-svenska (1/1)
arbetarinstituten (2/2)
hur (93/94) Hur (1)
växel (1/1)
taxa (1/1)
arbetsgivare (63/63)
Internetuppkoppling (1/1)
karttjänsten (2/2)
dag (27/27)
socken (1/1)
aktiv (2/2)
brandsläckaren (1/1)
styrkor (1/1)
ja (19/19)
bankgiroblankett (1/1)
sommarteatern (1/1)
YEL (1/1)
kvar (10/10)
beslutsfattande (3/3)
gymnasiebaserad (2/2)
turvatalo (3/3)
lekparksverksamhetfinska (1/1)
fritidsaktiviteterna (1/1)
alakoulu (1/1)
mekanisk (1/1)
finskundervisning (2/2)
responssystemfinska (1/1)
pääomatulo (1/1)
skatteprocent (6/6)
kvinnor (34/34)
tid (148/148)
tvättmaskinen (1/1)
undersökning (8/8)
tillfrågas (1/1)
palveluasuminen (1/1)
utsänd (1/1)
praxis (1/1)
Optia (1/1)
undervisningsgrupper (1/1)
klubben (2/2)
avser (6/6)
underlätta (2/2)
socialarbetare (10/10)
autonoma (1/1)
Commons (1/1)
kandidat (4/4)
bisyssla (2/2)
försvårar (1/1)
delvis (10/10)
satsat (1/1)
kotihoito (1/1)
samtalskostnad (1/1)
oljud (3/3)
fostras (2/2)
tecknat (1/1)
avfallshanteringfinska (1/1)
tvingas (5/5)
ort (5/5)
kompetensbaserat (2/2)
idrotts- (1/1)
identifiera (2/2)
matburkar (1/1)
borgerlig (2/2)
sorts (2/2)
handikappråd (1/1)
nödcentraloperatörens (1/1)
inhyste (1/1)
www.infofinland.fi (1/1)
separata (4/4)
Kvarkens (1/1)
lek (2/2)
ledande (2/2)
nationalspråk (2/2)
ID (5/5)
telefoner (1/1)
konflikter (5/5)
EU (117/117)
hobbystudier (2/2)
vaginalt (2/2)
slidmynning (1/1)
sexuella (6/6)
grupps (1/1)
traditionell (2/2)
apotekets (3/3)
radhus (3/3)
arbetstiden (4/4)
fotografi (1/1)
demokratiska (1/1)
läroavtalscenter (3/3)
tis (2/2)
hautausavustus (1/1)
tillväga (1/1)
lånord (1/1)
brev (5/5)
yhdenvertaisuus (1/1)
kuntoutustuki (1/1)
konstaterar (1/1)
märker (1/1)
fastän (5/5)
förekomma (2/2)
bönder (1/1)
temperaturerna (1/1)
institutfinska (1/1)
intressebevakare (1/1)
lådor (1/1)
samfundfinska (2/2)
undervisningfinska (2/2)
självständigt (14/14)
terminsavgift (1/1)
uhrien (1/1)
församlingar (10/10)
sidoapotek (1/1)
normalt (4/4)
riskerna (1/1)
platsansökan (1/1)
foto (1/1)
sämre (3/3)
delarna (2/2)
mål (3/3)
resten (3/3)
relationer (1/1)
kravet (3/3)
oavlönat (1/1)
söks (4/4)
examenstillfällen (1/1)
verifieras (1/1)
Studentkårers (1/1)
ledda (2/2)
mödravården (2/2)
vart (10/10)
utställningar (7/7)
vigslar (2/2)
skarvsladd (1/1)
mannens (1/1)
oavlönad (3/3)
krisarbetare (1/1)
verksamhetsprogram (1/1)
bekräftats (2/2)
genast (9/9)
förutsättningarna (3/3)
förskottsinnehållning (2/2)
yrkeshögskoleexamenfinska (1/1)
fortbildningfinska (1/1)
slotten (2/2)
existerar (3/3)
högljudd (1/1)
flyktingorganisation (2/2)
engelskspråkiga (3/3)
kom (18/18)
väderförhållanden (1/1)
inom (99/99)
kontoutdrag (1/1)
Pojkarnas (1/1)
fullmäktiges (2/2)
Arbetseffektivitetsföreningen (2/2)
familjeplaneringsrådgivningarna (1/1)
utvecklingsplan (2/2)
kommunikationskanal (1/1)
resmål (1/1)
rollen (1/1)
ljusaste (1/1)
fortare (1/1)
itsenäisen (1/1)
abonnemang (4/4)
utvisningfinska (1/1)
ungefär (16/16)
neuvontapalvelu (1/1)
förstörs (2/2)
Yrittäjät (1/1)
vidimerad (1/1)
fördjupa (1/1)
Enter (26/26)
Dödsfall (1/1)
spårvagnar (1/1)
illegala (1/1)
erillinen (1/1)
häva (2/2)
mellanmål (1/1)
Korsets (1/1)
Oodi (2/2)
Arctica (3/3)
deltar (6/6)
plötsliga (1/1)
användning (2/2)
exemplar (1/1)
telefontjänster (1/1)
talen (2/2)
jämkas (1/1)
kristna (3/3)
FPA.I (1/1)
kemikalier (2/2)
visning (1/1)
begäras (2/2)
framför (1/1)
faktor (1/1)
medier (3/4) Medier (1)
Olkkarifinska (1/1)
telefonservice (2/2)
VALMA (13/13)
samhällelig (1/1)
midnattssolens (1/1)
trafikförsäkring (1/1)
Isyysraha (1/1)
avsett (10/10)
närarbetefinska (1/1)
varit (22/22)
ålderdom (1/1)
kollektivtrafikförbindelser (4/4)
sakkunniga (1/1)
oberoende (5/5)
motionsplatserna (1/1)
autovero (1/1)
fattats (4/4)
dessa (56/56)
Västra (8/11) västra (3)
säkerställer (1/1)
slutligen (1/1)
födas (1/1)
titta (5/5)
panelen (2/2)
framsteg (1/1)
hyrestiden (3/3)
ylempi (1/1)
förskoleundervisningenfinska (3/3)
vuxengymnasierna (1/1)
Kluuvi (1/1)
asylansökanfinska (1/1)
framhävs (2/2)
träffpunkten (1/1)
aktiveringsmodellen (1/1)
pimpelfiske (1/1)
samhällsgrupp (2/2)
grammatikfinska (1/1)
koulunkäyntiavustaja (1/1)
ansökningsblanketten (3/3)
klinikkaan (1/1)
drag (1/1)
Clinicin (1/1)
paperi (1/1)
färdighetsnivåerna (1/1)
A (25/26) a (1)
stunder (1/1)
ekonomiplaneringen (1/1)
flytt (8/8)
ekonominfinska (1/1)
licensen (2/2)
immateriella (1/1)
kassakvittot (1/1)
bostadsrättsavgiften (4/4)
ställning (9/9)
rokotus (1/1)
stå (1/1)
Nelonen (1/1)
lämna (39/39)
skoldagen (3/3)
upptagna (1/1)
journumret (2/2)
College (1/1)
resurser (2/2)
FRK (1/1)
universitetsutbildningar (1/1)
läkarhjälp (1/1)
pappersformat (1/1)
familjeskäl (4/4)
sjöstad (1/1)
handikappade (35/36) Handikappade (1)
ålderspension (5/5)
mikrovågsugnen (1/1)
högskolan (4/4)
tullanmäla (1/1)
utkomststöd (18/18)
handlingen (2/2)
kallas (12/12)
rättshjälpsbyråer (1/1)
dagvårdsplatsfinska (2/2)
brottsoffrets (1/1)
Barnskydd (1/1)
psykiater (1/1)
samlar (1/1)
huvudhälsostationen (1/1)
facket (1/1)
service (2/3) Service (1)
integrationsplan (14/14)
sexualitetfinska (1/1)
bekantskaper (1/1)
trakasserier (2/2)
for (2/2)
familjeband (25/25)
examensnivå (1/1)
befogad (1/1)
tillverka (1/1)
Ludvig (1/1)
beaktas (14/14)
idrottsgrenar (3/3)
värd (1/1)
aktivt (4/4)
begär (2/2)
engelskspråkigt (1/1)
italienska (15/15)
meriterna (1/1)
högskolexamenfinska (1/1)
mentalvårdstjänsternafinska (1/1)
hörseln (1/1)
psykiatriska (1/1)
långvarigt (1/1)
konstruktionen (1/1)
inkluderar (1/1)
Arbisfinska (1/1)
skadas (1/1)
utfärdad (1/1)
betonat (1/1)
viktigast (1/1)
bygg- (1/1)
Anders (1/1)
skatteåterbäring (4/4)
din (511/511)
utfärdar (2/2)
fastställt (1/1)
bott (22/22)
medborgarinstitut (8/8)
Card (1/1)
lasi (1/1)
mörkt (1/1)
våld (57/61) Våld (4)
skrivna (1/1)
hennes (9/9)
unionens (2/2)
civil (2/2)
Suomen (12/13) suomen (1)
r.f (1/1)
kost (2/2)
nära (13/13)
klä (4/4)
tolkcentral (3/3)
yrkeshögskolekurser (1/1)
Jakobstad (2/2)
företagfinska (2/2)
raskauden (1/1)
miljon (1/1)
yleinen (3/3)
gå (36/36)
studerandehälsovården (2/2)
avvika (3/3)
straffbart (2/2)
medborgarskapet (1/1)
någon (71/71)
kursernas (1/1)
bostadsrättsbostäder (4/4)
konfidentiella (2/2)
påfrestande (2/2)
koulu (2/2)
unionen (6/6)
automat (1/1)
moderskapsledigheten (5/5)
skolelevers (1/1)
åtal (1/1)
områdeskoordinatorerna (1/1)
varje (35/35)
kraft (13/13)
Ristin (2/2)
FöretagsEsbo (1/1)
uteblir (1/1)
uträttar (3/3)
lärokursen (2/2)
palvelutalo (1/1)
tjänster (128/133) Tjänster (5)
människa (2/2)
sörja (4/4)
doula (1/1)
klara (16/16)
Europa (3/3)
länk (3/3)
omskärelse (6/6)
ansiotulo (1/1)
besöker (10/10)
kommunstyrelsen (1/1)
beviljats (11/11)
begår (4/4)
prioriteten (1/1)
Kaapatut (1/1)
lapsilisä (1/1)
oljemängden (1/1)
musicera (1/1)
Nordisk (3/4) nordisk (1)
kommunsida (1/1)
kauniainen.fi (1/1)
behovsprövat (2/2)
friluftsleder (1/1)
länkarna (2/2)
skattemyndigheten (3/3)
kommit (12/12)
faderskapsledigheten (3/3)
oleskeluoikeuden (1/1)
ordningsnumret (1/1)
insjukna (1/1)
flyttas (1/1)
postpositioner (1/1)
SHVS (1/1)
finansiärerna (1/1)
valkretsen (1/1)
komposteras (1/1)
erityisammattitutkinto (1/1)
marker (1/1)
invandrarefinska (20/20)
borealis (1/1)
lähikoulu (1/1)
bouppteckningfinska (1/1)
bodelningen (4/4)
beslutas (5/5)
Schengenstat (1/1)
Myrbackahuset (1/1)
belopp (23/23)
vandringfinska (1/1)
krisjouren (11/11)
InfoFinlands (289/289)
olycka (10/10)
ges (42/42)
bikulturella (1/1)
oavslutad (1/1)
webbsida (2/2)
arbetsoförmögen (2/2)
lokaltrafik (1/1)
elev- (1/1)
söder (1/1)
inget (21/21)
sjukvårdskort (1/1)
vuxnafinska (3/3)
uppstå (1/1)
smittats (1/1)
hembygdsmuseer (1/1)
regelbunden (2/2)
vakinaista (2/2)
uppstår (5/5)
utbildningsprogram (8/8)
hamnverksamheten (1/1)
annans (2/2)
skolkuratorer (1/1)
kostnadsfritt (5/5)
diabetes (2/2)
ringer (13/13)
kvinnlig (2/2)
databas (1/1)
besluta (10/10)
faderlöst (2/2)
registret (1/1)
narkos (1/1)
LUVA (3/3)
bedriva (1/1)
sakerna (1/1)
kontaktade (1/1)
förmiddagen (1/1)
arbetspensionsförsäkringarna (1/1)
Peijaksen (2/2)
webbundervisning (1/1)
händerna (1/1)
gymnasieutbildning (6/6)
hygienen (1/1)
flyttat (9/9)
omskurits (2/2)
lähdevero (1/1)
museidagen (1/1)
Helsingin (5/5)
etniskt (7/7)
Mundus (1/1)
plats (26/26)
finansieras (1/1)
Nivavaara (1/1)
hyresbostadfinska (1/1)
medborgarinstitutets (4/4)
vårt (2/2)
ovan (4/4)
kundtjänstfinska (1/1)
språkkaféer (1/1)
tog (3/3)
rester (1/1)
byrå (17/17)
matfinska (1/1)
utöva (8/8)
grenar (3/3)
utifrån (10/10)
efterlevandes (1/1)
varför (4/4)
språkversioner (1/1)
Stenängens (1/1)
dagvårdfinska (3/3)
avvecklas (1/1)
gränser (2/2)
påsen (2/2)
YouTube (2/2)
farlig (1/1)
luterilainen (1/1)
hyresgästen (4/4)
sakkunskap (1/1)
hemvårdsstödfinska (2/2)
hemsjukvården (1/1)
bryter (4/4)
fostran (18/21) Fostran (3)
stranden (1/1)
ehkäisy (1/1)
Tyttöjen (1/1)
sorggrupper (1/1)
dagsgymnasierna (1/1)
möjligheterna (3/3)
utgör (2/2)
ansluter (4/4)
badrumsrenovering (1/1)
helgons (3/3)
ingått (6/6)
förvärvsarbetande (1/1)
studieförmåga (1/1)
Migrationsverket (28/31) migrationsverket (3)
kortfattade (1/1)
socialskydd (1/1)
tvingade (1/1)
webbutik (1/1)
taket (1/1)
Kronoby (1/1)
invandrarens (1/1)
boendeträffpunkter (1/1)
universitetsstudier (3/3)
servicerådgivare (1/1)
anstaltsvårdenfinska (1/1)
babyresa (1/1)
lagar (13/13)
religionssamfund (4/4)
lönsamheten (1/1)
antalet (5/5)
serviceställen (2/2)
straffa (1/1)
skriftlig (7/7)
handlar (2/2)
nödsituationer (8/8)
germanska (1/1)
fyrverkerier (1/1)
FPAfinska (1/1)
ingång (3/3)
december (6/6)
bilagorna (4/4)
tjeckiska (1/1)
studier (80/81) Studier (1)
bygget (1/1)
vattenledningar (2/2)
avgiftsfritt (3/3)
handläggning (1/1)
vård (57/57)
A1 (5/5)
FIRST (1/1)
straffas (1/1)
HelMet (3/4) Helmet (1)
initiativtagande (1/1)
framskrider (3/3)
maximitiden (1/1)
bioavfall (2/2)
bortfaller (1/1)
kläder (6/6)
friluftsmuseumfinska (1/1)
tryckta (1/1)
betalt (2/2)
videoklippet (12/12)
kärnkraftverksprojekt (1/1)
absolut (1/1)
barnklubbar (3/3)
naturkunskap (1/1)
gränsöverskridande (1/1)
arvolaki (1/1)
påvisa (3/3)
Lappland (6/6)
samhällslivet (1/1)
rösträtt (13/13)
organ (1/1)
stöda (4/4)
rörelsehandikappad (1/1)
vatten (4/4)
patientombudsmannen (2/2)
åldringshem (1/1)
tillfälligt (21/22) Tillfälligt (1)
Tulli (1/1)
läroanstalter (17/17)
Oy:s (6/6)
Celsiusgrader (3/3)
härsken (1/1)
träffa (8/8)
grundskolan (33/33)
kunnande (16/16)
bankkonto (14/14)
bor (84/84)
internettjänsten (1/1)
isdubbar (1/1)
lärare (4/4)
träffar (1/1)
uppträder (2/2)
senaste (9/9)
droger (5/5)
terveysministeriö (2/2)
civilstånd (1/1)
jourtelefonen (2/2)
statlig (1/1)
befolkningsdataregistret (1/1)
ungdomsarbetare (1/1)
besvärstillstånd (2/2)
bäst (9/9)
hyresvärder (1/1)
grundundervisning (2/2)
påminnelse- (1/1)
förvärvsrelaterad (1/1)
faderskapspenningdagar (4/4)
läskunnighet (1/1)
bostadsrätten (2/2)
nationalmuseum (1/1)
d.v.s. (14/14)
gälla (2/2)
friluftsområden (1/1)
rättigheter (40/41) Rättigheter (1)
piller (2/2)
vuotiaan (1/1)
mobil (1/1)
elledningar (2/2)
ständigt (1/1)
NTM (3/3)
begränsa (1/1)
legitimerad (1/1)
bereder (2/2)
barnatillsyningsmännenfinska (2/2)
anmälningsdagen (2/2)
samiska (8/8)
folkpension (6/6)
jurist (14/14)
tala (14/14)
sådana (14/14)
betalningar (3/3)
utvecklingsstörd (3/3)
tillhör (11/11)
stiger (4/4)
Yrittäjän (1/1)
förnyas (1/1)
sedan (11/11)
kompetensområden (1/1)
pålitlig (3/3)
rösta (16/16)
hälsovårdens (1/1)
ärendet (11/11)
litar (1/1)
pappret (1/1)
Åboregionen (1/1)
vattenavgiften (3/3)
polisanmäla (1/1)
studieplats (29/29)
redaktionen (1/1)
vräka (1/1)
sederengelska (1/1)
hyrorna (1/1)
hörselundersökning (1/1)
telefontjänsten (6/6)
vak (1/1)
CV (13/13)
pojkvän (1/1)
modersmålet (6/6)
gärna (3/3)
utevistelse (1/1)
monteringsarbetsplats (1/1)
lördagar (1/1)
vårdens (1/1)
exceptionellt (2/2)
snitt (1/1)
Flickornas (2/2)
inkomster (34/34)
Matkahuoltos (4/4)
uppehållstillståndsärenden (1/1)
Island (7/7)
inlärningsgrupp (1/1)
grad (1/1)
framskrida (1/1)
akutpreventivmedel (1/1)
konflikterna (2/2)
typen (1/1)
föreslår (3/3)
uppfyllas (1/1)
pappersansökan (1/1)
ordna (23/23)
trakasserar (1/1)
pysyvä (1/1)
internetanslutning (1/2) Internetanslutning (1)
anställningsintervju (1/1)
varma (4/4)
hotfullt (1/1)
skogsbruksområden (1/1)
vite (1/1)
kulturministeriet (4/4)
rusmedel (2/2)
företagsverksamhet (15/15)
sjukt (6/6)
Nuorisoasiainkeskus (1/1)
döms (1/1)
dörrar (1/1)
lantdag (1/1)
seniorerfinska (1/1)
parförhållande (24/24)
föräldern (23/23)
icke (5/6) Icke (1)
försvunna (1/1)
experterna (1/1)
lagstadgade (1/1)
hens (1/1)
parets (1/1)
arbetserfarenhet (10/10)
årskurserna (12/12)
VR (1/1)
värmeelement (1/1)
nivåerna (2/2)
dans (6/6)
klienter (8/8)
visst (6/6)
uppgifterna (12/12)
avsevärt (3/3)
koulutus (3/3)
gymnasiestudierfinska (1/1)
examensstuderande (2/2)
www.gramex.fi (1/1)
medeltiden (1/1)
föreskrivs (2/2)
bostadsaktier (1/1)
originalspråk (1/1)
järnaffärer (1/1)
viseringsskyldiga (1/1)
fakulteten (1/1)
e (29/30) E (1)
relationerna (3/3)
minoritetsspråk (1/1)
orsakar (4/4)
stannar (5/5)
arbetarinstitut (11/11)
accepterade (1/1)
tidsbokningfinska (1/1)
levnadskostnader (2/2)
utbytesstudenter (1/1)
brinnande (1/1)
stanna (10/10)
gymnasierna (2/2)
orsaka (5/5)
van (1/1)
konventionerna (2/2)
vaccination (1/1)
referensramen (1/1)
religionsundervisningen (2/2)
idrottsanläggningar (1/1)
bostäderna (4/4)
utföra (9/9)
hel.fi (2/2)
intervjuar (1/1)
plastprodukter (2/2)
universitetens (1/1)
ange (8/8)
beslutsfattandet (6/6)
syskonrabatt (1/1)
normala (1/1)
skilda (1/1)
punkten (1/1)
påtryckning (1/1)
rubrik (1/1)
sker (14/14)
högre (26/26)
idkar (1/1)
jämföra (4/4)
ekonomiskt (4/5) Ekonomiskt (1)
undersökningen (3/3)
guidade (3/3)
riksdagsledamöter (1/1)
pensionärer (4/4)
present (1/1)
industrialiserades (1/1)
Kejsardömet (1/1)
elever (9/9)
tjänsteleverantör (1/1)
ansökningsbilagorna (6/6)
specialdagvård (1/1)
brottsofferfinska (2/2)
republikens (1/1)
avtal (30/30)
förskoleplats (4/4)
förlossningsdatum (1/1)
www.teosto.fi (1/1)
ligger (22/22)
Hollihaan (1/1)
Arbetslöshetsförsäkring (5/9) arbetslöshetsförsäkring (4)
portfölj (1/1)
snabbare (3/3)
preliminär (1/1)
tillgången (2/2)
avancerad (1/1)
skatterelaterade (1/1)
24h (3/3)
tätorter (2/2)
värms (1/1)
november (4/4)
organisationerna (1/1)
Asianajajaliitto (1/1)
invandrarbyrån (4/4)
exporterade (2/2)
intyga (1/1)
ohälsa (1/1)
avgiftningsvård (1/1)
socialtjänster (4/4)
Apostilleavtaletengelska (1/1)
emellan (1/1)
sällskapande (3/3)
specialundervisningen (1/1)
skett (1/1)
originalspråket (1/1)
bildkonst (8/8)
Opetushallitus (5/7) opetushallitus (2)
utvecklat (1/1)
väljer (10/10)
Työväen (2/2)
likvärdiga (2/2)
professionella (1/1)
morgon (2/2)
halvvägs (1/1)
frilansarefinska (1/1)
försäkringspremierna (4/4)
landskapsbibliotek (3/3)
sjunger (1/1)
kraven (2/2)
mottagningar (2/2)
linkkiLapplands (1/1)
tänker (2/2)
HNS (3/3)
påsk (1/1)
julstjärnor (1/1)
vigsel (11/11)
bevisas (4/4)
uppmuntrar (2/2)
ylletröja (1/1)
boningsort (1/1)
utomstående (3/3)
brister (3/3)
eget (62/62)
relaterade (1/1)
förhållandena (1/1)
natten (2/2)
avger (1/1)
osasairauspäiväraha (1/1)
mera (5/5)
Naapuruussovittelun (1/1)
tolktjänster (5/5)
skickas (8/8)
bosatt (19/19)
installeras (1/1)
medeltemperaturen (1/1)
InfoFinland.fi (2/2)
ombud (1/1)
flygplats (7/7)
specialboende (1/1)
renoveringskostnaden (1/1)
svenskspråkigt (4/4)
nödvändigtvis (10/10)
Oy (9/9)
småbarnsfostran (4/4)
svar (1/1)
Oikarainen (1/1)
deras (36/36)
räcker (11/11)
stödcentret (3/3)
ansvaret (9/9)
gifta (23/23)
yttranderätt (1/1)
arbetsprov (2/2)
sökmotorer (1/1)
bilder (3/3)
Tukiliittos (1/1)
bygger (1/1)
revisionsbyråer (1/1)
kontaktspråk (1/1)
rådgivningarna (2/2)
tv (5/6) TV (1)
öppen (13/13)
hemkommunfinska (1/1)
beskrivs (2/2)
original (6/6)
fastlagsbullar (1/1)
kristelefonfinska (1/1)
kundtjänst (1/1)
läroanstalt (12/12)
abonnemanget (1/1)
finskafinska (2/2)
Estnäs (1/1)
avlagda (1/1)
undervisningstimmar (1/1)
skenäktenskap (1/1)
svalt (2/2)
Kafnettis (1/1)
Finnkinos (1/1)
loven (1/1)
moderna (1/1)
hälsomyndighet (1/1)
bibliotekskunderna (1/1)
fritidsaktiviteter (3/3)
studentexamen (7/7)
Kehitysvammaisten (1/1)
parkeringsautomater (1/1)
kuntoutussuunnitelma (1/1)
betalningssvårigheter (1/1)
psykologen (2/2)
utbetalning (4/4)
integrationsutbildningen (2/2)
dra (3/3)
klienten (2/2)
skoltiden (1/1)
järnvägsstationerna (1/1)
asylprocessen (1/1)
svagheterna (1/1)
ägarbostäderfinska (2/2)
fakulteterna (1/1)
graviditetenfinska (1/1)
isolering (1/1)
arbetsliv (1/1)
kostnaderna (15/15)
Struves (1/1)
upphovsrättsliga (1/1)
bekostar (1/1)
diskriminerat (2/2)
aktuella (6/6)
samtycker (2/2)
systerdotter (1/1)
medlemmarna (3/3)
Österbottens (17/17)
partiell (9/9)
hyresbostäderfinska (5/5)
pension (16/17) Pension (1)
varieteter (1/1)
folkhögskolan (3/3)
dvs. (3/3)
grundar (6/6)
officiellt (11/15) Officiellt (4)
svåra (2/2)
guidar (1/1)
grunda (31/31)
matkakortin (1/1)
kreditgivning (1/1)
positivt (4/4)
olydiga (1/1)
avtalas (1/1)
musikhobby (1/1)
dari (2/2)
varumärkesrätt (1/1)
använda (79/79)
innehållet (4/7) Innehållet (3)
fylla (19/19)
kondomer (1/1)
tillförlitligt (2/2)
tillväxten (1/1)
oleskelulupa (1/1)
upprätta (6/6)
öppenvården (1/1)
försäkringsbolaget (1/1)
främmande (9/9)
käyttövastike (1/1)
arbetspension (6/6)
Kansa (1/1)
bekräftar (5/5)
användas (6/6)
Uunofinska (1/1)
nattcaféet (1/1)
färre (1/1)
kotihoidon (2/2)
hemspråksundervisningfinska (1/1)
permanent (17/17)
anslutna (1/1)
föra (12/12)
åstadkomma (1/1)
Seure (1/1)
taxitjänster (1/1)
makars (1/1)
föreläsningsserier (1/1)
Internetanslutningar (1/1)
Eiran (1/1)
studiemetoder (1/1)
byggherren (1/1)
näringslivstjänsterna (1/1)
tryggheten (61/61)
arbeta (80/82) Arbeta (2)
passar (7/7)
reglerade (4/4)
omavastuuaika (2/2)
tandklinik (4/4)
arbetar (40/40)
hålla (4/4)
VR:s (2/2)
olägenhet (1/1)
studerat (3/3)
snabbt (11/11)
släktingar (9/9)
hämtas (1/1)
angående (3/3)
snart (1/1)
föräldraledighet (2/2)
spelproblem (4/4)
bankerna (1/1)
liksom (2/2)
digital- (1/1)
terapin (2/2)
underhållet (1/1)
misstanken (1/1)
läggs (1/1)
uppväxt (4/4)
allra (2/2)
faderskapsärendet (1/1)
privatpersoners (1/1)
jämte (1/1)
rasistiskt (5/5)
arbetstagarna (3/3)
inkvartering (2/2)
studietakt (1/1)
fars (1/1)
evangelisk (17/17)
målsättningar (1/1)
teater (8/8)
etälukio (1/1)
källorna (1/1)
öarna (2/2)
skick (7/7)
krävas (1/1)
frågor (51/51)
regionförvaltningsverken (1/1)
Klimatet (1/2) klimatet (1)
ombes (1/1)
hälsostationens (1/1)
papperslöshetfinska (1/1)
linkkiFinnkino (1/1)
ungdomsarbete (3/3)
godtagbar (3/3)
tagalog (1/1)
tidsbegränsade (1/1)
kreditkort (3/3)
barnatillsynsmannen (1/1)
löneutbetalningfinska (1/1)
grund- (1/1)
motorfordon (3/3)
smal (1/1)
bevis (4/4)
bibliotek (16/17) Bibliotek (1)
vaccinationer (4/4)
förskoleundervisning (14/15) Förskoleundervisning (1)
civilvigsel (1/1)
bönestund (1/1)
vitas (1/1)
funktionell (1/1)
passfoto (2/2)
avläggas (5/5)
tider (10/10)
bestå (6/6)
misstänker (11/11)
nödvändig (3/3)
stödnät (1/1)
psykoterapin (1/1)
Uskonnot (2/2)
utmärkt (1/1)
videoklipp (3/3)
mödrar (1/1)
läroplanen (1/1)
kompletterande (2/2)
bröstsmärtor (1/1)
landets (6/6)
skolhälsovårdaren (4/4)
avgiftsbelagd (12/12)
handelscentra (1/1)
lämplighet (1/1)
efternamnfinska (1/1)
filmvisningar (1/1)
sjöss (3/3)
priserfinska (1/1)
Närpes (1/1)
följer (12/12)
diskrimineringsombudsmannen (2/3) Diskrimineringsombudsmannen (1)
läkarstationer (4/4)
lilla (1/1)
blivande (3/3)
främst (5/5)
bildkonstskola (1/1)
skogen (2/2)
näringstjänsterfinska (2/2)
cykel- (1/1)
avlägga (56/56)
aikuiskoulutuskeskus (1/1)
förarexamen (1/1)
naturstigar (1/1)
tjänsteställe (11/11)
näring (1/1)
ställa (6/6)
sökordet (1/1)
landsbygd (1/1)
begagnade (1/1)
brandvarnaren (2/2)
viktig (15/15)
tyngdpunkt (1/1)
hjälpa (26/26)
magistrat (4/4)
dessutom (25/25)
umgås (1/1)
Vandainfo (1/1)
tel (2/2)
startpenningen (1/1)
synskadades (1/1)
införskaffat (1/1)
rekisterihallitus (1/1)
stadshus (2/2)
vägande (5/5)
Lapin (1/1)
sjukvårdskortet (6/6)
uppsöka (1/1)
Tukinainen (1/1)
hälsovårdsministeriet (3/3)
HRT (3/3)
arbetssökanden (1/1)
stämmor (1/1)
stressyndrom (1/1)
beskattningen (24/24)
socialhandledningfinska (1/1)
företagshälsovård (8/9) Företagshälsovård (1)
hälsostationer (10/10)
dem (64/64)
äktenskapsförordet (2/2)
anställningsintervjun (1/1)
granne (6/6)
jour (1/1)
hobbyredskap (1/1)
tandkliniker (4/4)
översättare (4/4)
frånluftsventilerna (1/1)
ersättningar (1/1)
hörselskada (3/3)
undgår (1/1)
kanaler (5/5)
runt (29/29)
elevverksamhet (1/1)
sovittelu (2/2)
böjs (2/2)
hyran (14/14)
sökmotor (6/6)
jämställdhetsnämnden (4/4)
dagvårdsenhet (1/1)
julskinka (1/1)
familjeplaneringfinska (2/2)
demonstrationer (1/1)
båda (20/20)
Vardagslivet (1/1)
www.tuotos.fi (1/1)
människors (5/5)
samlat (1/1)
siffror (1/1)
välbefinnandet (1/1)
avslår (2/2)
erövrades (1/1)
sistone (1/1)
folkhögskolor (3/3)
syn- (1/1)
umgängetfinska (1/1)
Takuusäätiö (3/3)
tillåtet (6/6)
Tammerforsregionen (1/1)
Finlandengelska (6/6)
världsarv (2/2)
fullföljer (1/1)
snö (1/1)
båtliv (1/1)
snöskottande (1/1)
specialutbildning (1/1)
enbart (3/3)
kust (1/1)
Patentti- (1/1)
gåva (1/1)
avtalats (2/2)
mottagningscentral (4/4)
tolkningen (8/8)
stadiluotsi (1/1)
Pensionsskyddscentralens (1/1)
vid (450/450)
tävlingens (3/3)
avtalat (4/4)
Kriscentret (1/2) kriscentret (1)
utbildade (4/4)
arbetslöshetsersättning (10/10)
senare (11/11)
orter (20/20)
medborgarskap (70/70)
peruskielitaito (1/1)
vuxensocialarbetet (1/1)
leker (1/1)
diskrimineras (6/6)
yhdessä (1/1)
apotekens (1/1)
lämplighetsprov (1/1)
satt (2/2)
hälsocentralen (2/2)
arbetsamhet (1/1)
skatter (9/9)
fjärde (13/13)
Galoppbrinken (1/1)
reglerat (4/4)
krisjourenfinska (2/2)
vändagen (2/2)
heltidsstudier (4/4)
mångkulturella (6/6)
bokföringsskyldighet (1/1)
arbetslöshet (2/2)
dispens (2/2)
drog- (1/1)
linor (1/1)
arbetspensionsutdragfinska (1/1)
Helsinki (11/11)
ansökningssättet (1/1)
kölapp (1/1)
överinspektören (1/1)
osäker (2/2)
tvåspråkiga (4/4)
kropps (1/1)
delas (15/15)
hemvårdens (5/5)
skuld (1/1)
lönsam (3/3)
FöPL (1/1)
nätter (1/1)
bil (12/12)
avgiftsfri (10/10)
flerfaldiga (1/1)
invandrarförening (1/1)
moderskapsledig (3/3)
Advokatförbund (1/2) advokatförbund (1)
sökas (4/4)
ifrån (5/5)
egnahemshuset (1/1)
målet (4/4)
flyga (1/1)
arv (2/2)
oppisopimus (1/1)
grundskoleinstitutionen (1/1)
tjänsten (64/64)
ungdomsfullmäktige (1/1)
jourens (1/1)
regnbågsfamiljerfinska (1/1)
meddela (18/18)
utrymmen (1/1)
obligatorisk (2/2)
näringar (1/1)
självständighetsdag (1/1)
tolkcentraler (2/2)
inte (661/661)
uppgett (1/1)
glömde (1/1)
Ilmonet.fi (1/1)
meddelas (8/8)
granskningar (1/1)
konto (13/13)
skattepliktig (2/2)
-flickor (1/1)
borgarna (1/1)
sigfinska (1/1)
egen (83/83)
rehabiliteringsinrättning (1/1)
pensionstagarefinska (1/1)
BY (2/2)
moderskapspenning (9/9)
A2 (2/2)
Förbundfinska (1/1)
midsommaren (1/1)
företagarguider (1/1)
invandrare (86/86)
underhållsbehovet (1/1)
familjeterapi (1/1)
likaberättigandefinska (1/1)
målsättningen (1/1)
vårdnadshavares (1/1)
ammattikorkeakoulututkinto (1/1)
hemskickad (1/1)
inkomstrelaterad (9/9)
invandrarfamiljer (1/1)
närvarar (1/1)
vårdnadshavarna (2/2)
skräp (1/1)
informerar (5/5)
Stadin (4/4)
bostadsrättskontraktet (1/1)
livscykel (1/1)
aktiivimalli (1/1)
rasismi (1/1)
låna (10/10)
rikt (1/1)
skuldlinjen (1/1)
religiös (5/5)
spalt (1/1)
bekantat (1/1)
medan (5/5)
faderskapspenning (3/3)
ordföranden (3/3)
pitkä (1/1)
tolktjänst (2/2)
underrättelse (2/2)
återhämta (2/2)
egenvårdsläkemedel (1/1)
osakeyhtiö (1/1)
företagsrådgivningen (4/4)
Vuokra (1/1)
helgjour (1/1)
all (1/1)
Advisor (1/1)
presidentval (4/4)
terrängen (1/1)
medlemsländerna (1/1)
studiepoäng (2/2)
infopankki (1/1)
haku (1/1)
skillnad (1/1)
endast (44/44)
våren (14/14)
Alkoholister (2/3) alkoholister (1)
ordningsregler (2/2)
integrationsprocessen (1/1)
kriget (4/4)
bostaden (62/62)
milda (1/1)
gym (3/3)
prioriteras (2/2)
pappfabrik (1/1)
pensionen (2/2)
servicenumret (1/1)
kontrollerar (1/1)
hjälpmedlen (2/2)
valtion (1/1)
