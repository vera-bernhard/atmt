Grundläggande information
Historia
Trafik
Religion
Beslutsfattande och påverkan
Grundläggande information
Karleby finns i Mellersta Österbotten invid Bottniska viken.
Karleby stad är grundad 1620 och hette då Gamlakarleby.
Senare blev Kokkola stadens finska namn.
Vid Karleby centrum finns en av landets mest omfattande historiska trästadshelheter.
Stadsplanen är från 1650-talet.
Den omfattar 12 kvarter med hundratals trähus och gårdsbyggnader.
De äldsta av dessa är från 1600-talet.
Karleby är en kulturstad med mycket att se och uppleva.
Karleby hamn ligger i stadsdelen Yxpila och är en av Finlands mest trafikerade godshamnar.
Grunden för näringslivet i Karleby är den internationella storindustrin.
I Karleby är den kemiska industrin och industri i anslutning till denna särskilt viktig.
Karleby är även en betydande handelsstad.
Information om Karlebyfinska _ svenska _ engelska
Historia
Redan under medeltiden fanns det hamn, båtbygge och handelsplats i Karleby.
Landhöjningen har varit en central faktor i Karlebys historia.
Den har format omgivningen i hög grad och bland annat påverkat utvecklingen av hamnverksamheten och handeln.
Handel bedrevs längs med Bottniska vikens kust och jordbruk, jakt, fiske och sälfångst var även viktiga näringar.
Exporten av tjära, som blev mycket viktig för Karlebys historia, inleddes redan på 1500-talet.
Den sjunde september 1620 undertecknade Sveriges kung Gustav II Adolf en handling som gav den lilla jordbruks- och fiskebyn vid Ristrand status som stad.
Dagens stadssund var då en smal havsvik som sträckte sig ända till Kyrkbacken.
Sakta men säkert blev Karleby en viktig stad för sjöfart och skeppsbygge.
Skeppsvarv fanns bland annat i Kaustarviken, Svartskär och Soldatskär.
Inledningsvis seglade man endast till Åbo och Stockholm, eftersom Karleby som s.k. uppstad inte fick bedriva utrikeshandel.
År 1765 erhöll staden stapelrättigheter, dvs. rätt till fri utrikeshandel, främst tack vare den aktiva kyrkoherden och lantdagsmannen Anders Chydenius.
Karleby blev snabbt en förmögen stad i början av 1800-talet tack vare just handeln med tjära och rederiverksamheten.
Stadens borgare köpte tjära av bönder och exporterade den, ofta till hamnar vid Medelhavet och i England.
Karleby handelsflotta var under perioder Finlands största.
Den snabba ekonomiska utvecklingen avtog i mitten av 1800-talet, men tog ny fart i slutet av århundradet tack vare industrialiseringen.
Karleby blev en viktig industristad främst tack vare läder- och metallindustrin.
Karlebys historiafinska _ svenska _ engelska
Trafik
Karleby har goda trafikförbindelser.
Via Karleby löper riksväg 8 och 13.
Järnvägsstationen finns i stadens centrum.
Restiden med tåg till Helsingfors är cirka fyra timmar.
Flygplatsen finns i Kronoby på endast 22 kilometers avstånd från Karleby centrum.
Stadsborna erbjuds även ett tryggt, omfattande, fungerande och trivsamt nätverk för den lätta trafiken.
Karleby har satsat på att förbättra förhållandena för cyklister.
Lokalbussarna trafikerar de olika delarna av staden på vardagar.
Läs mer: Trafik.
Gator och trafikfinska _ svenska
Kollektivtrafikfinska _ svenska
linkkiVR:
Tågtidtabellerfinska _ svenska _ engelska _ ryska
Busstidtabellerfinska _ svenska _ engelska
Flyg från Karleby-Jakobstad flygplatsfinska _ svenska _ engelska
Religion
I Karleby finns flera olika religiösa samfund.
I tjänsten Uskonnot Suomessa (Religioner i Finland) finns information om religiösa samfund enligt ort.
Den evangelisk-lutherska kyrkan har fyra finskspråkiga församlingar och en svenskspråkig församling i Karleby.
Läs mer på Karleby kyrkliga samfällighets webbplats.
I Karleby finns en ortodox kyrka.
Mer information om den ortodoxa församlingens verksamhet i Karleby finns på Vasa ortodoxa församlings webbplats.
Läs mer: Kulturer och religioner i Finland.
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiVasa ortodoxa församling:
Vasa ortodoxa församlingfinska _ engelska _ ryska
Beslutsfattande och påverkan
Den högsta beslutsfattande makten i Karleby stad innehas av stadsfullmäktige.
Fullmäktigeledamöterna och deras suppleanter väljs vid kommunalval vart fjärde år.
På stadens webbplats finns information om stadsfullmäktige och dess beslut.
Invånarna kan påverka stadens beslutsfattande redan då beslut bereds.
Information om olika sätt att delta och påverka finns på stadens webbplats.
Kommunens invånare har enligt kommunallagen rätt att lämna in motioner till kommunen i ärenden som gäller dess verksamhet.
I Karleby finns ungdomsfullmäktige, äldre- och handikappråd samt ett råd för kulturell mångfald.
Läs mer: Finlands förvaltning, Val och röstning i Finland
Beslutsfattandefinska _ svenska _ engelska
Grundläggande information
Historia
Trafik
Religion
Beslutsfattande och påverkan
Grundläggande information
Karleby finns i Mellersta Österbotten invid Bottniska viken.
Karleby stad är grundad 1620 och hette då Gamlakarleby.
Senare blev Kokkola stadens finska namn.
Vid Karleby centrum finns en av landets mest omfattande historiska trästadshelheter.
Stadsplanen är från 1650-talet.
Den omfattar 12 kvarter med hundratals trähus och gårdsbyggnader.
De äldsta av dessa är från 1600-talet.
Karleby är en kulturstad med mycket att se och uppleva.
Karleby hamn ligger i stadsdelen Yxpila och är en av Finlands mest trafikerade godshamnar.
Grunden för näringslivet i Karleby är den internationella storindustrin.
I Karleby är den kemiska industrin och industri i anslutning till denna särskilt viktig.
Karleby är även en betydande handelsstad.
Information om Karlebyfinska _ svenska _ engelska
Historia
Redan under medeltiden fanns det hamn, båtbygge och handelsplats i Karleby.
Landhöjningen har varit en central faktor i Karlebys historia.
Den har format omgivningen i hög grad och bland annat påverkat utvecklingen av hamnverksamheten och handeln.
Handel bedrevs längs med Bottniska vikens kust och jordbruk, jakt, fiske och sälfångst var även viktiga näringar.
Exporten av tjära, som blev mycket viktig för Karlebys historia, inleddes redan på 1500-talet.
Den sjunde september 1620 undertecknade Sveriges kung Gustav II Adolf en handling som gav den lilla jordbruks- och fiskebyn vid Ristrand status som stad.
Dagens stadssund var då en smal havsvik som sträckte sig ända till Kyrkbacken.
Sakta men säkert blev Karleby en viktig stad för sjöfart och skeppsbygge.
Skeppsvarv fanns bland annat i Kaustarviken, Svartskär och Soldatskär.
Inledningsvis seglade man endast till Åbo och Stockholm, eftersom Karleby som s.k. uppstad inte fick bedriva utrikeshandel.
År 1765 erhöll staden stapelrättigheter, dvs. rätt till fri utrikeshandel, främst tack vare den aktiva kyrkoherden och lantdagsmannen Anders Chydenius.
Karleby blev snabbt en förmögen stad i början av 1800-talet tack vare just handeln med tjära och rederiverksamheten.
Stadens borgare köpte tjära av bönder och exporterade den, ofta till hamnar vid Medelhavet och i England.
Karleby handelsflotta var under perioder Finlands största.
Den snabba ekonomiska utvecklingen avtog i mitten av 1800-talet, men tog ny fart i slutet av århundradet tack vare industrialiseringen.
Karleby blev en viktig industristad främst tack vare läder- och metallindustrin.
Karlebys historiafinska _ svenska _ engelska
Trafik
Karleby har goda trafikförbindelser.
Via Karleby löper riksväg 8 och 13.
Järnvägsstationen finns i stadens centrum.
Restiden med tåg till Helsingfors är cirka fyra timmar.
Flygplatsen finns i Kronoby på endast 22 kilometers avstånd från Karleby centrum.
Stadsborna erbjuds även ett tryggt, omfattande, fungerande och trivsamt nätverk för den lätta trafiken.
Karleby har satsat på att förbättra förhållandena för cyklister.
Lokalbussarna trafikerar de olika delarna av staden på vardagar.
Läs mer: Trafik.
Gator och trafikfinska _ svenska
Kollektivtrafikfinska _ svenska
linkkiVR:
Tågtidtabellerfinska _ svenska _ engelska _ ryska
Busstidtabellerfinska _ svenska _ engelska
Flyg från Karleby-Jakobstad flygplatsfinska _ svenska _ engelska
Religion
I Karleby finns flera olika religiösa samfund.
I tjänsten Uskonnot Suomessa (Religioner i Finland) finns information om religiösa samfund enligt ort.
Den evangelisk-lutherska kyrkan har fyra finskspråkiga församlingar och en svenskspråkig församling i Karleby.
Läs mer på Karleby kyrkliga samfällighets webbplats.
I Karleby finns en ortodox kyrka.
Mer information om den ortodoxa församlingens verksamhet i Karleby finns på Vasa ortodoxa församlings webbplats.
Läs mer: Kulturer och religioner i Finland.
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiVasa ortodoxa församling:
Vasa ortodoxa församlingfinska _ engelska _ ryska
Beslutsfattande och påverkan
Den högsta beslutsfattande makten i Karleby stad innehas av stadsfullmäktige.
Fullmäktigeledamöterna och deras suppleanter väljs vid kommunalval vart fjärde år.
På stadens webbplats finns information om stadsfullmäktige och dess beslut.
Invånarna kan påverka stadens beslutsfattande redan då beslut bereds.
Information om olika sätt att delta och påverka finns på stadens webbplats.
Kommunens invånare har enligt kommunallagen rätt att lämna in motioner till kommunen i ärenden som gäller dess verksamhet.
I Karleby finns ungdomsfullmäktige, äldre- och handikappråd samt ett råd för kulturell mångfald.
Läs mer: Finlands förvaltning, Val och röstning i Finland
Beslutsfattandefinska _ svenska _ engelska
Grundläggande information
Historia
Trafik
Religion
Beslutsfattande och påverkan
Grundläggande information
Karleby finns i Mellersta Österbotten invid Bottniska viken.
Karleby stad är grundad 1620 och hette då Gamlakarleby.
Senare blev Kokkola stadens finska namn.
Vid Karleby centrum finns en av landets mest omfattande historiska trästadshelheter.
Stadsplanen är från 1650-talet.
Den omfattar 12 kvarter med hundratals trähus och gårdsbyggnader.
De äldsta av dessa är från 1600-talet.
Karleby är en kulturstad med mycket att se och uppleva.
Karleby hamn ligger i stadsdelen Yxpila och är en av Finlands mest trafikerade godshamnar.
Grunden för näringslivet i Karleby är den internationella storindustrin.
I Karleby är den kemiska industrin och industri i anslutning till denna särskilt viktig.
Karleby är även en betydande handelsstad.
Information om Karlebyfinska _ svenska _ engelska
Historia
Redan under medeltiden fanns det hamn, båtbygge och handelsplats i Karleby.
Landhöjningen har varit en central faktor i Karlebys historia.
Den har format omgivningen i hög grad och bland annat påverkat utvecklingen av hamnverksamheten och handeln.
Handel bedrevs längs med Bottniska vikens kust och jordbruk, jakt, fiske och sälfångst var även viktiga näringar.
Exporten av tjära, som blev mycket viktig för Karlebys historia, inleddes redan på 1500-talet.
Den sjunde september 1620 undertecknade Sveriges kung Gustav II Adolf en handling som gav den lilla jordbruks- och fiskebyn vid Ristrand status som stad.
Dagens stadssund var då en smal havsvik som sträckte sig ända till Kyrkbacken.
Sakta men säkert blev Karleby en viktig stad för sjöfart och skeppsbygge.
Skeppsvarv fanns bland annat i Kaustarviken, Svartskär och Soldatskär.
Inledningsvis seglade man endast till Åbo och Stockholm, eftersom Karleby som s.k. uppstad inte fick bedriva utrikeshandel.
År 1765 erhöll staden stapelrättigheter, dvs. rätt till fri utrikeshandel, främst tack vare den aktiva kyrkoherden och lantdagsmannen Anders Chydenius.
Karleby blev snabbt en förmögen stad i början av 1800-talet tack vare just handeln med tjära och rederiverksamheten.
Stadens borgare köpte tjära av bönder och exporterade den, ofta till hamnar vid Medelhavet och i England.
Karleby handelsflotta var under perioder Finlands största.
Den snabba ekonomiska utvecklingen avtog i mitten av 1800-talet, men tog ny fart i slutet av århundradet tack vare industrialiseringen.
Karleby blev en viktig industristad främst tack vare läder- och metallindustrin.
Karlebys historiafinska _ svenska _ engelska
Trafik
Karleby har goda trafikförbindelser.
Via Karleby löper riksväg 8 och 13.
Järnvägsstationen finns i stadens centrum.
Restiden med tåg till Helsingfors är cirka fyra timmar.
Flygplatsen finns i Kronoby på endast 22 kilometers avstånd från Karleby centrum.
Stadsborna erbjuds även ett tryggt, omfattande, fungerande och trivsamt nätverk för den lätta trafiken.
Karleby har satsat på att förbättra förhållandena för cyklister.
Lokalbussarna trafikerar de olika delarna av staden på vardagar.
Läs mer: Trafik.
Gator och trafikfinska _ svenska
Kollektivtrafikfinska _ svenska
linkkiVR:
Tågtidtabellerfinska _ svenska _ engelska _ ryska
Busstidtabellerfinska _ svenska _ engelska
Flyg från Karleby-Jakobstad flygplatsfinska _ svenska _ engelska
Religion
I Karleby finns flera olika religiösa samfund.
I tjänsten Uskonnot Suomessa (Religioner i Finland) finns information om religiösa samfund enligt ort.
Den evangelisk-lutherska kyrkan har fyra finskspråkiga församlingar och en svenskspråkig församling i Karleby.
Läs mer på Karleby kyrkliga samfällighets webbplats.
I Karleby finns en ortodox kyrka.
Mer information om den ortodoxa församlingens verksamhet i Karleby finns på Vasa ortodoxa församlings webbplats.
Läs mer: Kulturer och religioner i Finland.
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiVasa ortodoxa församling:
Vasa ortodoxa församlingfinska _ engelska _ ryska
Beslutsfattande och påverkan
Den högsta beslutsfattande makten i Karleby stad innehas av stadsfullmäktige.
Fullmäktigeledamöterna och deras suppleanter väljs vid kommunalval vart fjärde år.
På stadens webbplats finns information om stadsfullmäktige och dess beslut.
Invånarna kan påverka stadens beslutsfattande redan då beslut bereds.
Information om olika sätt att delta och påverka finns på stadens webbplats.
Kommunens invånare har enligt kommunallagen rätt att lämna in motioner till kommunen i ärenden som gäller dess verksamhet.
I Karleby finns ungdomsfullmäktige, äldre- och handikappråd samt ett råd för kulturell mångfald.
Läs mer: Finlands förvaltning, Val och röstning i Finland
Beslutsfattandefinska _ svenska _ engelska
Detta innehåll finns inte på det språk som du har valt.
Välj något annat språk.
Finska
Detta innehåll finns inte på det språk som du har valt.
Välj något annat språk.
Finska
Detta innehåll finns inte på det språk som du har valt.
Välj något annat språk.
Finska
Bibliotek
Motion
Att röra sig i naturen
Teater och film
Museer
Hobbyer för barn och unga
Föreningar
Karleby är en gammal sjöstad som erbjuder mångsidiga möjligheter för utfärder och friluftsliv.
Personer ntresserad av friluftsliv bör läsa mer om allemansrätten under rubriken ”Att röra sig i naturen” i denna tjänst.
Flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet.
Föreningar och organisationer samt hobbygrupper och kommunala institut erbjuder kurser i idrott och kultur samt bl.a. språk och hantverk.
I Snellman-salen och i stadens övriga kulturlokaler erbjuds kulturevenemang av varierande slag.
Årliga evenemang i Karleby är bland annat Veneziansk afton i slutet av sommaren, Kokkola Cup för fotbollsjuniorer, Stadsfestivalen Karleby sommarveckor, Lochteå kyrkomusikfest samt Vinterdans i Karleby och festivalen Karleby Vinterharmonika.
Mer information om fritidstjänsterna i Karleby finns på Karleby stads webbplats.
På stadens webbplats finns även en länk till Evenemangskalendern med daglig information om stadens kultur- och motionsevenemang.
Läs mer: Fritid.
Evenemangskalenderfinska
Kulturtjänsterfinska _ svenska _ engelska
Idrottstjänsterfinska _ svenska _ engelska
Bibliotek
Karleby stadsbibliotek finns i stadens centrum.
Närbiblioteken finns i Björkhagen, Kelviå, Lochteå samt Ullava kyrkby och Rahkonen.
Information om bibliotekets öppettider och tjänster finns på dess webbplats.
Biblioteket finns även på nätet.
Där kan kunderna bläddra i bibliotekets samlingar, reservera material, förnya sina lån, beställa fjärrlån och låna e-böcker under alla tider på dygnet.
Tack vare det effektiva biblioteksnätverket i Finland är nästan alla finländska biblioteks samlingar tillgängliga för bibliotekskunderna i Karleby.
Karleby stadsbibliotek/huvudbiblioteket
Storgatan 3, 67100 Karleby
Telefon: 040 806 5124, 040 806 5133
Läs mer: Bibliotek.
Bibliotekstjänsterfinska _ svenska _ engelska
Motion
I Karleby finns mångsidiga motionsmöjligheter året runt.
Staden anordnar ledda aktiviteter i Simcentret VesiVeijari och motionshallarna.
Dessutom finns det gym av flera olika slag.
Gym anpassade för äldre finns i Furuåsens aktivitetscenter och Kuusikumpu servicehus.
Staden underhåller cykelvägar, motionsrutter, joggingbanor, skidspår, badstränder, bollplaner och skridskobanor samt platser för närmotion.
I Karlebynejdens instituts nättjänst finns information om institutets mångsidiga motionsutbud.
I Karleby finns nära på hundra idrottsföreningar för olika grenar samt föreningar som arrangerar övrig motion.
Mer information om motionsmöjligheter i Karleby finns på Karleby stads webbplats.
Läs mer:
Motion.
Idrottstjänsterfinska _ svenska _ engelska
Motionsplatserfinska _ svenska
Gym för äldrefinska
Karlebynejdens institutfinska _ svenska
Att röra sig i naturen
Att röra sig i naturen är en traditionell och populär form av avkoppling för finländarna under alla årstider.
I Finland kan man med stöd av allemansrätten plocka bär och svamp i skogen och röra sig till fots, med cykel eller skidor vintertid.
Det är inte tillåtet att beträda folks gårdar utan lov.
För fiske krävs fiskelov, med undantag för mete och pilkning.
Även jakt fordrar jakttillstånd.
Allemansrätten ger inte rätt att skräpa ner i naturen, skada träd eller växter, störa eller skada fågelbon eller fågelungar, köra motorfordon utan markägarens tillstånd eller bygga ens tillfälliga byggen.
Mer information om motionsrutterna, rastplatser, möjligheter till fiske och båtliv samt exempelvis fågeltorn i Karleby finns på stadens webbplats.
Rutterna för camping, paddling, vandring, cykling och övriga rutter i Karleby finns i karttjänsten på nätet.
I karttjänsten visas även var största delen av motionsplatserna finns.
Du kan köpa friluftskartor över Karleby hos Karleby Turism: Salutorget 5, 67100 Karleby.
Läs mer: Att röra sig i naturen.
linkkiMiljöförvaltningen:
Allemansrättenfinska _ svenska _ engelska _ ryska
Motionskarta över Karlebyfinska _ svenska
Motionsrutter i Karlebyfinska _ svenska
Teater och film
Karleby är en teaterstad med långa anor, som erbjuder scenkonst på hög nivå framförd av både proffs och amatörer.
Karleby stadsteater finns i det stämningsfulla Vartiolinna (Torggatan 48).
Du kan läsa mer om amatörteatrarnas verksamhet på deras webbplats och i evenemangskalendern.
I Karleby finns biografen Bio Rex, vars två salar använder digital- och 3D-teknik.
Bio Rex program finns under länken här intill.
Läs mer: Teater och film.
Stadsteaternfinska
Biograffinska
Teater och danskonst i Karlebyfinska _ svenska _ engelska
Evenemangskalenderfinska
Museer
I hjärtat av staden, i det anrika Rooska gården, finns K.H.Renlunds museum.
Karleby stad grundade museet 1909 utgående från en testamentsgåva av affärsmannen Karl Herman Renlund (1850–1908) .
På museet finns Renlunds samling av finländsk konst från guldåldern och tillfälliga utställningar i en kulturhistorisk miljö.
Även i museikvarterens övriga byggnader finns utställningar om stadens kulturhistoria och utställningar med ITE-konst.
På K.H.Renlunds museums webbplats finns mer information om museets tjänster, utställningar samt aktuell verksamhet.
Utöver K.H.Renlunds museum lönar det sig att besöka det naturhistoriska museet Kieppi (Kieppi är stängt tills vidare på grund av brand) samt de många hembygdsmuseerna och övriga de historiska resmålen i regionen.
Exempelvis i Konst-Vionoja-centret presenteras konstnären Veikko Vionojas verk.
I Kelviå, ca 10 km norrut från Karleby, finns Toivonen djurpark och drängmuseum.
Mer information om dessa museer finns under länkarna här intill.
Läs mer: Museer.
Museer och traditionsarbetefinska _ svenska _ engelska
K.H. Renlunds museum - Mellersta Österbottens landskapsmuseumfinska _ svenska _ engelska
Kieppi, Karleby naturvetenskapliga museumfinska _ svenska _ engelska
linkkiToivonens djurpark och drängmuseum :
Toivonens djurpark och drängmuseum finska _ svenska _ engelska
Konst Vionojafinska
Hobbyer för barn och unga
Flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet.
Flera olika föreningar samt kommunala institut ger unga möjlighet att studera idrott och kultur samt bl.a. språk och hantverk.
Barn och unga kan delta i grundläggande undervisning i musik, dans, bildkonst och hantverk.
Dessutom erbjuder stadens ungdomstjänster en rockskola.
Stadens ungdomstjänster driver sju ungdomsgårdar runt om i Karleby.
De rusmedels- och rökfria ungdomslokalerna erbjuder handledd verksamhet för barn i årskurserna 3–6 och unga i åldern 13–17 år i olika delar av Karleby.
Information om hobbyverksamheter för barn och unga finns på stadens webbplats.
Rådgivningen vid Ungdomsgården Vinge ger aktuell information om bl.a. internationalisering, studier, arbetsliv, hälsa, hobbyverksamhet och boende.
Karlebynejdens institut erbjuder barn och unga olika former av hobbyverksamhet, exempelvis i konstämnen och musik.
Kontrollera vilka kurser som är aktuella i institutets webbtjänst.
Karleby evangelisk-lutherska församlingar erbjuder även hobbyverksamhet för barn och unga, såsom lekparksträffar, klubbar, musikverksamhet och läger.
Mer information om verksamheten finns på Karleby församlingssammanslutnings webbplats.
Ungdomsgården Vinge
67100 Karleby
Läs mer: Hobbyer för barn och unga.
Övrig undervisning i Karlebyfinska _ svenska
Ungdomstjänsterfinska _ svenska _ engelska
Karlebynejdens institutfinska _ svenska
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
Föreningar
Karleby har ett aktivt och mångsidigt föreningsliv för invånare i alla åldrar.
Läs mer: Föreningar.
Bibliotek
Motion
Att röra sig i naturen
Teater och film
Museer
Hobbyer för barn och unga
Föreningar
Karleby är en gammal sjöstad som erbjuder mångsidiga möjligheter för utfärder och friluftsliv.
Personer ntresserad av friluftsliv bör läsa mer om allemansrätten under rubriken ”Att röra sig i naturen” i denna tjänst.
Flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet.
Föreningar och organisationer samt hobbygrupper och kommunala institut erbjuder kurser i idrott och kultur samt bl.a. språk och hantverk.
I Snellman-salen och i stadens övriga kulturlokaler erbjuds kulturevenemang av varierande slag.
Årliga evenemang i Karleby är bland annat Veneziansk afton i slutet av sommaren, Kokkola Cup för fotbollsjuniorer, Stadsfestivalen Karleby sommarveckor, Lochteå kyrkomusikfest samt Vinterdans i Karleby och festivalen Karleby Vinterharmonika.
Mer information om fritidstjänsterna i Karleby finns på Karleby stads webbplats.
På stadens webbplats finns även en länk till Evenemangskalendern med daglig information om stadens kultur- och motionsevenemang.
Läs mer: Fritid.
Evenemangskalenderfinska
Kulturtjänsterfinska _ svenska _ engelska
Idrottstjänsterfinska _ svenska _ engelska
Bibliotek
Karleby stadsbibliotek finns i stadens centrum.
Närbiblioteken finns i Björkhagen, Kelviå, Lochteå samt Ullava kyrkby och Rahkonen.
Information om bibliotekets öppettider och tjänster finns på dess webbplats.
Biblioteket finns även på nätet.
Där kan kunderna bläddra i bibliotekets samlingar, reservera material, förnya sina lån, beställa fjärrlån och låna e-böcker under alla tider på dygnet.
Tack vare det effektiva biblioteksnätverket i Finland är nästan alla finländska biblioteks samlingar tillgängliga för bibliotekskunderna i Karleby.
Karleby stadsbibliotek/huvudbiblioteket
Storgatan 3, 67100 Karleby
Telefon: 040 806 5124, 040 806 5133
Läs mer: Bibliotek.
Bibliotekstjänsterfinska _ svenska _ engelska
Motion
I Karleby finns mångsidiga motionsmöjligheter året runt.
Staden anordnar ledda aktiviteter i Simcentret VesiVeijari och motionshallarna.
Dessutom finns det gym av flera olika slag.
Gym anpassade för äldre finns i Furuåsens aktivitetscenter och Kuusikumpu servicehus.
Staden underhåller cykelvägar, motionsrutter, joggingbanor, skidspår, badstränder, bollplaner och skridskobanor samt platser för närmotion.
I Karlebynejdens instituts nättjänst finns information om institutets mångsidiga motionsutbud.
I Karleby finns nära på hundra idrottsföreningar för olika grenar samt föreningar som arrangerar övrig motion.
Mer information om motionsmöjligheter i Karleby finns på Karleby stads webbplats.
Läs mer:
Motion.
Idrottstjänsterfinska _ svenska _ engelska
Motionsplatserfinska _ svenska
Gym för äldrefinska
Karlebynejdens institutfinska _ svenska
Att röra sig i naturen
Att röra sig i naturen är en traditionell och populär form av avkoppling för finländarna under alla årstider.
I Finland kan man med stöd av allemansrätten plocka bär och svamp i skogen och röra sig till fots, med cykel eller skidor vintertid.
Det är inte tillåtet att beträda folks gårdar utan lov.
För fiske krävs fiskelov, med undantag för mete och pilkning.
Även jakt fordrar jakttillstånd.
Allemansrätten ger inte rätt att skräpa ner i naturen, skada träd eller växter, störa eller skada fågelbon eller fågelungar, köra motorfordon utan markägarens tillstånd eller bygga ens tillfälliga byggen.
Mer information om motionsrutterna, rastplatser, möjligheter till fiske och båtliv samt exempelvis fågeltorn i Karleby finns på stadens webbplats.
Rutterna för camping, paddling, vandring, cykling och övriga rutter i Karleby finns i karttjänsten på nätet.
I karttjänsten visas även var största delen av motionsplatserna finns.
Du kan köpa friluftskartor över Karleby hos Karleby Turism: Salutorget 5, 67100 Karleby.
Läs mer: Att röra sig i naturen.
linkkiMiljöförvaltningen:
Allemansrättenfinska _ svenska _ engelska _ ryska
Motionskarta över Karlebyfinska _ svenska
Motionsrutter i Karlebyfinska _ svenska
Teater och film
Karleby är en teaterstad med långa anor, som erbjuder scenkonst på hög nivå framförd av både proffs och amatörer.
Karleby stadsteater finns i det stämningsfulla Vartiolinna (Torggatan 48).
Du kan läsa mer om amatörteatrarnas verksamhet på deras webbplats och i evenemangskalendern.
I Karleby finns biografen Bio Rex, vars två salar använder digital- och 3D-teknik.
Bio Rex program finns under länken här intill.
Läs mer: Teater och film.
Stadsteaternfinska
Biograffinska
Teater och danskonst i Karlebyfinska _ svenska _ engelska
Evenemangskalenderfinska
Museer
I hjärtat av staden, i det anrika Rooska gården, finns K.H.Renlunds museum.
Karleby stad grundade museet 1909 utgående från en testamentsgåva av affärsmannen Karl Herman Renlund (1850–1908) .
På museet finns Renlunds samling av finländsk konst från guldåldern och tillfälliga utställningar i en kulturhistorisk miljö.
Även i museikvarterens övriga byggnader finns utställningar om stadens kulturhistoria och utställningar med ITE-konst.
På K.H.Renlunds museums webbplats finns mer information om museets tjänster, utställningar samt aktuell verksamhet.
Utöver K.H.Renlunds museum lönar det sig att besöka det naturhistoriska museet Kieppi (Kieppi är stängt tills vidare på grund av brand) samt de många hembygdsmuseerna och övriga de historiska resmålen i regionen.
Exempelvis i Konst-Vionoja-centret presenteras konstnären Veikko Vionojas verk.
I Kelviå, ca 10 km norrut från Karleby, finns Toivonen djurpark och drängmuseum.
Mer information om dessa museer finns under länkarna här intill.
Läs mer: Museer.
Museer och traditionsarbetefinska _ svenska _ engelska
K.H. Renlunds museum - Mellersta Österbottens landskapsmuseumfinska _ svenska _ engelska
Kieppi, Karleby naturvetenskapliga museumfinska _ svenska _ engelska
linkkiToivonens djurpark och drängmuseum :
Toivonens djurpark och drängmuseum finska _ svenska _ engelska
Konst Vionojafinska
Hobbyer för barn och unga
Flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet.
Flera olika föreningar samt kommunala institut ger unga möjlighet att studera idrott och kultur samt bl.a. språk och hantverk.
Barn och unga kan delta i grundläggande undervisning i musik, dans, bildkonst och hantverk.
Dessutom erbjuder stadens ungdomstjänster en rockskola.
Stadens ungdomstjänster driver sju ungdomsgårdar runt om i Karleby.
De rusmedels- och rökfria ungdomslokalerna erbjuder handledd verksamhet för barn i årskurserna 3–6 och unga i åldern 13–17 år i olika delar av Karleby.
Information om hobbyverksamheter för barn och unga finns på stadens webbplats.
Rådgivningen vid Ungdomsgården Vinge ger aktuell information om bl.a. internationalisering, studier, arbetsliv, hälsa, hobbyverksamhet och boende.
Karlebynejdens institut erbjuder barn och unga olika former av hobbyverksamhet, exempelvis i konstämnen och musik.
Kontrollera vilka kurser som är aktuella i institutets webbtjänst.
Karleby evangelisk-lutherska församlingar erbjuder även hobbyverksamhet för barn och unga, såsom lekparksträffar, klubbar, musikverksamhet och läger.
Mer information om verksamheten finns på Karleby församlingssammanslutnings webbplats.
Ungdomsgården Vinge
67100 Karleby
Läs mer: Hobbyer för barn och unga.
Övrig undervisning i Karlebyfinska _ svenska
Ungdomstjänsterfinska _ svenska _ engelska
Karlebynejdens institutfinska _ svenska
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
Föreningar
Karleby har ett aktivt och mångsidigt föreningsliv för invånare i alla åldrar.
Läs mer: Föreningar.
Bibliotek
Motion
Att röra sig i naturen
Teater och film
Museer
Hobbyer för barn och unga
Föreningar
Karleby är en gammal sjöstad som erbjuder mångsidiga möjligheter för utfärder och friluftsliv.
Personer ntresserad av friluftsliv bör läsa mer om allemansrätten under rubriken ”Att röra sig i naturen” i denna tjänst.
Flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet.
Föreningar och organisationer samt hobbygrupper och kommunala institut erbjuder kurser i idrott och kultur samt bl.a. språk och hantverk.
I Snellman-salen och i stadens övriga kulturlokaler erbjuds kulturevenemang av varierande slag.
Årliga evenemang i Karleby är bland annat Veneziansk afton i slutet av sommaren, Kokkola Cup för fotbollsjuniorer, Stadsfestivalen Karleby sommarveckor, Lochteå kyrkomusikfest samt Vinterdans i Karleby och festivalen Karleby Vinterharmonika.
Mer information om fritidstjänsterna i Karleby finns på Karleby stads webbplats.
På stadens webbplats finns även en länk till Evenemangskalendern med daglig information om stadens kultur- och motionsevenemang.
Läs mer: Fritid.
Evenemangskalenderfinska
Kulturtjänsterfinska _ svenska _ engelska
Idrottstjänsterfinska _ svenska _ engelska
Bibliotek
Karleby stadsbibliotek finns i stadens centrum.
Närbiblioteken finns i Björkhagen, Kelviå, Lochteå samt Ullava kyrkby och Rahkonen.
Information om bibliotekets öppettider och tjänster finns på dess webbplats.
Biblioteket finns även på nätet.
Där kan kunderna bläddra i bibliotekets samlingar, reservera material, förnya sina lån, beställa fjärrlån och låna e-böcker under alla tider på dygnet.
Tack vare det effektiva biblioteksnätverket i Finland är nästan alla finländska biblioteks samlingar tillgängliga för bibliotekskunderna i Karleby.
Karleby stadsbibliotek/huvudbiblioteket
Storgatan 3, 67100 Karleby
Telefon: 040 806 5124, 040 806 5133
Läs mer: Bibliotek.
Bibliotekstjänsterfinska _ svenska _ engelska
Motion
I Karleby finns mångsidiga motionsmöjligheter året runt.
Staden anordnar ledda aktiviteter i Simcentret VesiVeijari och motionshallarna.
Dessutom finns det gym av flera olika slag.
Gym anpassade för äldre finns i Furuåsens aktivitetscenter och Kuusikumpu servicehus.
Staden underhåller cykelvägar, motionsrutter, joggingbanor, skidspår, badstränder, bollplaner och skridskobanor samt platser för närmotion.
I Karlebynejdens instituts nättjänst finns information om institutets mångsidiga motionsutbud.
I Karleby finns nära på hundra idrottsföreningar för olika grenar samt föreningar som arrangerar övrig motion.
Mer information om motionsmöjligheter i Karleby finns på Karleby stads webbplats.
Läs mer:
Motion.
Idrottstjänsterfinska _ svenska _ engelska
Motionsplatserfinska _ svenska
Gym för äldrefinska
Karlebynejdens institutfinska _ svenska
Att röra sig i naturen
Att röra sig i naturen är en traditionell och populär form av avkoppling för finländarna under alla årstider.
I Finland kan man med stöd av allemansrätten plocka bär och svamp i skogen och röra sig till fots, med cykel eller skidor vintertid.
Det är inte tillåtet att beträda folks gårdar utan lov.
För fiske krävs fiskelov, med undantag för mete och pilkning.
Även jakt fordrar jakttillstånd.
Allemansrätten ger inte rätt att skräpa ner i naturen, skada träd eller växter, störa eller skada fågelbon eller fågelungar, köra motorfordon utan markägarens tillstånd eller bygga ens tillfälliga byggen.
Mer information om motionsrutterna, rastplatser, möjligheter till fiske och båtliv samt exempelvis fågeltorn i Karleby finns på stadens webbplats.
Rutterna för camping, paddling, vandring, cykling och övriga rutter i Karleby finns i karttjänsten på nätet.
I karttjänsten visas även var största delen av motionsplatserna finns.
Du kan köpa friluftskartor över Karleby hos Karleby Turism: Salutorget 5, 67100 Karleby.
Läs mer: Att röra sig i naturen.
linkkiMiljöförvaltningen:
Allemansrättenfinska _ svenska _ engelska _ ryska
Motionskarta över Karlebyfinska _ svenska
Motionsrutter i Karlebyfinska _ svenska
Teater och film
Karleby är en teaterstad med långa anor, som erbjuder scenkonst på hög nivå framförd av både proffs och amatörer.
Karleby stadsteater finns i det stämningsfulla Vartiolinna (Torggatan 48).
Du kan läsa mer om amatörteatrarnas verksamhet på deras webbplats och i evenemangskalendern.
I Karleby finns biografen Bio Rex, vars två salar använder digital- och 3D-teknik.
Bio Rex program finns under länken här intill.
Läs mer: Teater och film.
Stadsteaternfinska
Biograffinska
Teater och danskonst i Karlebyfinska _ svenska _ engelska
Evenemangskalenderfinska
Museer
I hjärtat av staden, i det anrika Rooska gården, finns K.H.Renlunds museum.
Karleby stad grundade museet 1909 utgående från en testamentsgåva av affärsmannen Karl Herman Renlund (1850–1908) .
På museet finns Renlunds samling av finländsk konst från guldåldern och tillfälliga utställningar i en kulturhistorisk miljö.
Även i museikvarterens övriga byggnader finns utställningar om stadens kulturhistoria och utställningar med ITE-konst.
På K.H.Renlunds museums webbplats finns mer information om museets tjänster, utställningar samt aktuell verksamhet.
Utöver K.H.Renlunds museum lönar det sig att besöka det naturhistoriska museet Kieppi (Kieppi är stängt tills vidare på grund av brand) samt de många hembygdsmuseerna och övriga de historiska resmålen i regionen.
Exempelvis i Konst-Vionoja-centret presenteras konstnären Veikko Vionojas verk.
I Kelviå, ca 10 km norrut från Karleby, finns Toivonen djurpark och drängmuseum.
Mer information om dessa museer finns under länkarna här intill.
Läs mer: Museer.
Museer och traditionsarbetefinska _ svenska _ engelska
K.H. Renlunds museum - Mellersta Österbottens landskapsmuseumfinska _ svenska _ engelska
Kieppi, Karleby naturvetenskapliga museumfinska _ svenska _ engelska
linkkiToivonens djurpark och drängmuseum :
Toivonens djurpark och drängmuseum finska _ svenska _ engelska
Konst Vionojafinska
Hobbyer för barn och unga
Flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet.
Flera olika föreningar samt kommunala institut ger unga möjlighet att studera idrott och kultur samt bl.a. språk och hantverk.
Barn och unga kan delta i grundläggande undervisning i musik, dans, bildkonst och hantverk.
Dessutom erbjuder stadens ungdomstjänster en rockskola.
Stadens ungdomstjänster driver sju ungdomsgårdar runt om i Karleby.
De rusmedels- och rökfria ungdomslokalerna erbjuder handledd verksamhet för barn i årskurserna 3–6 och unga i åldern 13–17 år i olika delar av Karleby.
Information om hobbyverksamheter för barn och unga finns på stadens webbplats.
Rådgivningen vid Ungdomsgården Vinge ger aktuell information om bl.a. internationalisering, studier, arbetsliv, hälsa, hobbyverksamhet och boende.
Karlebynejdens institut erbjuder barn och unga olika former av hobbyverksamhet, exempelvis i konstämnen och musik.
Kontrollera vilka kurser som är aktuella i institutets webbtjänst.
Karleby evangelisk-lutherska församlingar erbjuder även hobbyverksamhet för barn och unga, såsom lekparksträffar, klubbar, musikverksamhet och läger.
Mer information om verksamheten finns på Karleby församlingssammanslutnings webbplats.
Ungdomsgården Vinge
67100 Karleby
Läs mer: Hobbyer för barn och unga.
Övrig undervisning i Karlebyfinska _ svenska
Ungdomstjänsterfinska _ svenska _ engelska
Karlebynejdens institutfinska _ svenska
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
Föreningar
Karleby har ett aktivt och mångsidigt föreningsliv för invånare i alla åldrar.
Läs mer: Föreningar.
Problem med uppehållstillstånd
Brott
Våld
Diskriminering och rasism
Behöver du en jurist?
Död
Problem i äktenskap eller parförhållande
Skilsmässa
Problem med den mentala hälsan
Missbruksproblem
I en krissituation kan du ringa nödcentralen på numret 112.
De slussar vid behov dig vidare till socialjouren.
Du ska endast ringa nödcentralen i brådskande nödsituationer, där liv, egendom eller miljön är i fara.
Problem med uppehållstillstånd
Om du har problem eller oklarheter med ditt uppehållstillstånd kan du kontakta Migrationsverket.
Migrationsverket
Korsholmsesplanaden 45
Vasa
Läs mer: Problem med uppehållstillstånd.
Brott
Om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112.
Ring inte nödnumret om det inte är fråga om en nödsituation.
Du kan göra en polisanmälan på nätet.
Mer information finns på Polisens webbplats.
Du kan även skriva ut anmälningsblanketten på nätet och lämna in den till polisstationen.
Karleby polisstation
Karlebygatan 74
67100 Karleby
Läs mer: Brott.
Tidsbokningfinska _ svenska _ engelska
Polisamälanfinska _ svenska _ engelska
Våld
Om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112.
Läs mer: Våld.
Diskriminering och rasism
Om du misstänker att du blivit utsatt för diskriminering då du sökt arbete eller på arbetsplatsen ska du först ta upp detta på din arbetsplats.
Om saken inte kan lösas på arbetsplatsen ska du kontakta arbetarskyddet vid Regionförvaltningsverket i Västra och Inre Finland.
Besöksadress:
Regionförvaltningsverket i Västra och Inre Finland
Wollfskavägen 35
65101 Vasa
Telefon: 0295 018 450
Om du utsätts för diskriminering kan du be om hjälp av Diskrimineringsombudsmannen.
Om du fallit offer för ett rasistiskt motiverat brott kan du göra en polisanmälan på nätet eller polisstationen.
Läs mer: Diskriminering och rasism.
linkkiRegionförvaltningsverket i Västra och Inre Finland:
Regionförvaltningsverket i Västra och Inre Finlandfinska _ svenska _ engelska
Hjälp och information för personer som drabbats av etnisk diskrimineringfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Behöver du en jurist?
Juridiska tjänster är avgiftsbelagda men om du har små eller medelstora inkomster, kan du få helt eller delvis avgiftsfri rättshjälp från statens rättshjälpsbyrå.
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
Besöksadress: Ämbetshuset, Torggatan 40, 67100 Karleby
Telefon: 029 566 1270
Information om enskilda jurister finns bland annat på Finlands Advokatförbunds webbplats.
Läs mer:
Behöver du en jurist?
linkkiFinlands advokatförbund:
Finlands advokatförbundfinska _ svenska _ engelska
Död
Den evangelisk-lutherska kyrkans församlingars begravningsplatser fungerar som allmänna begravningsplatser.
Där kan även avlidna som inte är medlemmar i kyrkan begravas.
De är alltså avsedda för alla invånare i staden.
Mer information finns på Karleby kyrkliga samfällighets webbplats.
Om en närstående plötsligt dör kan du söka krishjälp vid din egen hälsostation, eller utanför tjänstetid vid samjouren för Mellersta Österbottens centralsjukhus.
De evangelisk-lutherska församlingarna i Karlebynejden erbjuder även sorggrupper.
Även församlingarnas diakonimottagningar erbjuder samtalshjälp för sorgearbetet.
Läs mer: Död.
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Problem i äktenskap eller parförhållande
Vid problem i äktenskap eller parförhållande får du hjälp av Mellersta Österbottens familjerådgivningscentral som underhålls av Karleby kyrkliga samfällighets och Mellersta Österbottens social- och hälsovårdssamkommun Soites familjerådgivning.
Familjerågivningscentralen
Telefon: 050 3147 464.
Karleby familjerådgivning
67100 Karleby
tel. 044 730 7640
Läs mer: Problem i äktenskap eller parförhållande.
linkkiMellersta Österbottens Familjerådgivningscentral:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
Skilsmässa
Skilsmässa kan sökas av kvinnan, av mannen eller av båda makarna tillsammans.
Man ansöker om skilsmässa i tingsrätten.
Till att börja med görs en skriftlig skilsmässoansökan.
Österbottens tingsrätt Karleby kansli
Besöksadress: Karlebygatan 27, 67100 Karleby
Telefon: 029 56 49294
Läs mer: Skilsmässa.
Hälsovårdaren på barnrådgivningsbyrån ger råd i frågor som gäller små barns hälsa, tillväxt och utveckling.
Barnrådgivningsbyrån ger information om platser som erbjuder hjälp vid behov.
Vid problem hos unga i skolåldern hjälper exempelvis skolans hälsovårdare eller skolkuratorn.
Läs mer: Barns och ungas problem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Skolhälsovårdfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barnrådgivningarfinska _ svenska
Du kan ta upp problem med hälsovårdaren på skolan eller studieplatsen eller vuxna på ungdomsgården.
Mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats.
Föräldrar eller unga själva kan kontakta familjerådgivningen.
Där kan man tala om problem och få hjälp och stöd.
Mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats.
Familjerådgivningens telefonnummer: 044 730 7640.
Läs mer: Barns och ungas problem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Studerandehälsovårdfinska _ svenska
Ungdomsgårdar och -lokaler finska _ svenska
Problem med den mentala hälsan
Om du behöver hjälp och stöd för din mentala hälsa kan du boka en läkartid vid hälsostationen.
Läkaren bedömer situationen.
Vid behov skriver läkaren en remiss till psykiatrisk specialsjukvård.
Läs mer: Mental hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Mentalvårdstjänsterfinska _ svenska
Om du har ekonomiska problem kan du be om råd hos Mellersta Österbottens social- och hälsovårdssamkommun Soites enheter för socialarbete eller utkomststöd, tfn 040 806 5095 eller tjänstestyrningen, tfn 040 806 5093.
Om du har problem med skulder, kontakta rättshjälpsbyrån.
Du kan anlita vilken som helst rättshjälpsbyrå oberoende av din hemkommun.
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
Telefon: 029 566 1270
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Servicehandledningfinska _ svenska
Missbruksproblem
Om du har problem med alkohol, droger, läkemedel eller hasardspel kan du få vård och rehabilitering vid Porten, Mellersta Österbottens social- och hälsovårdssamkommun Soites center för missbruksproblem.
Du kan ta upp problemet med proffs inom hälsovården eller företagshälsovården, som kan slussa dig vidare i vårdsystemet, eller direkt kontakta Soites missbrukstjänster, tfn 040 8068 101.
För tillnyktrings- och avgiftningsvård debiteras en patientavgift liksom även för korttidsrehabilitering, öppen rehabilitering är gratis.
Även Karleby evangelisk-lutherska församlingssammanslutnings specialdiakoner erbjuder samtalshjälp vid missbruksproblem.
Kontaktuppgifter
Hälsovägen 4
67200 Karleby
Telefon: 040 806 8101
Läs mer: Missbruksproblem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Service för missbrukarefinska _ svenska
linkkiKarleby evangelisk-lutherska församlingssammansutning:
Karleby evangelisk-lutherska församlings arbete bland missbrukarefinska _ svenska
Problem med uppehållstillstånd
Brott
Våld
Diskriminering och rasism
Behöver du en jurist?
Död
Problem i äktenskap eller parförhållande
Skilsmässa
Problem med den mentala hälsan
Missbruksproblem
I en krissituation kan du ringa nödcentralen på numret 112.
De slussar vid behov dig vidare till socialjouren.
Du ska endast ringa nödcentralen i brådskande nödsituationer, där liv, egendom eller miljön är i fara.
Problem med uppehållstillstånd
Om du har problem eller oklarheter med ditt uppehållstillstånd kan du kontakta Migrationsverket.
Migrationsverket
Korsholmsesplanaden 45
Vasa
Läs mer: Problem med uppehållstillstånd.
Brott
Om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112.
Ring inte nödnumret om det inte är fråga om en nödsituation.
Du kan göra en polisanmälan på nätet.
Mer information finns på Polisens webbplats.
Du kan även skriva ut anmälningsblanketten på nätet och lämna in den till polisstationen.
Karleby polisstation
Karlebygatan 74
67100 Karleby
Läs mer: Brott.
Tidsbokningfinska _ svenska _ engelska
Polisamälanfinska _ svenska _ engelska
Våld
Om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112.
Läs mer: Våld.
Diskriminering och rasism
Om du misstänker att du blivit utsatt för diskriminering då du sökt arbete eller på arbetsplatsen ska du först ta upp detta på din arbetsplats.
Om saken inte kan lösas på arbetsplatsen ska du kontakta arbetarskyddet vid Regionförvaltningsverket i Västra och Inre Finland.
Besöksadress:
Regionförvaltningsverket i Västra och Inre Finland
Wollfskavägen 35
65101 Vasa
Telefon: 0295 018 450
Om du utsätts för diskriminering kan du be om hjälp av Diskrimineringsombudsmannen.
Om du fallit offer för ett rasistiskt motiverat brott kan du göra en polisanmälan på nätet eller polisstationen.
Läs mer: Diskriminering och rasism.
linkkiRegionförvaltningsverket i Västra och Inre Finland:
Regionförvaltningsverket i Västra och Inre Finlandfinska _ svenska _ engelska
Hjälp och information för personer som drabbats av etnisk diskrimineringfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Behöver du en jurist?
Juridiska tjänster är avgiftsbelagda men om du har små eller medelstora inkomster, kan du få helt eller delvis avgiftsfri rättshjälp från statens rättshjälpsbyrå.
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
Besöksadress: Ämbetshuset, Torggatan 40, 67100 Karleby
Telefon: 029 566 1270
Information om enskilda jurister finns bland annat på Finlands Advokatförbunds webbplats.
Läs mer:
Behöver du en jurist?
linkkiFinlands advokatförbund:
Finlands advokatförbundfinska _ svenska _ engelska
Död
Den evangelisk-lutherska kyrkans församlingars begravningsplatser fungerar som allmänna begravningsplatser.
Där kan även avlidna som inte är medlemmar i kyrkan begravas.
De är alltså avsedda för alla invånare i staden.
Mer information finns på Karleby kyrkliga samfällighets webbplats.
Om en närstående plötsligt dör kan du söka krishjälp vid din egen hälsostation, eller utanför tjänstetid vid samjouren för Mellersta Österbottens centralsjukhus.
De evangelisk-lutherska församlingarna i Karlebynejden erbjuder även sorggrupper.
Även församlingarnas diakonimottagningar erbjuder samtalshjälp för sorgearbetet.
Läs mer: Död.
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Problem i äktenskap eller parförhållande
Vid problem i äktenskap eller parförhållande får du hjälp av Mellersta Österbottens familjerådgivningscentral som underhålls av Karleby kyrkliga samfällighets och Mellersta Österbottens social- och hälsovårdssamkommun Soites familjerådgivning.
Familjerågivningscentralen
Telefon: 050 3147 464.
Karleby familjerådgivning
67100 Karleby
tel. 044 730 7640
Läs mer: Problem i äktenskap eller parförhållande.
linkkiMellersta Österbottens Familjerådgivningscentral:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
Skilsmässa
Skilsmässa kan sökas av kvinnan, av mannen eller av båda makarna tillsammans.
Man ansöker om skilsmässa i tingsrätten.
Till att börja med görs en skriftlig skilsmässoansökan.
Österbottens tingsrätt Karleby kansli
Besöksadress: Karlebygatan 27, 67100 Karleby
Telefon: 029 56 49294
Läs mer: Skilsmässa.
Hälsovårdaren på barnrådgivningsbyrån ger råd i frågor som gäller små barns hälsa, tillväxt och utveckling.
Barnrådgivningsbyrån ger information om platser som erbjuder hjälp vid behov.
Vid problem hos unga i skolåldern hjälper exempelvis skolans hälsovårdare eller skolkuratorn.
Läs mer: Barns och ungas problem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Skolhälsovårdfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barnrådgivningarfinska _ svenska
Du kan ta upp problem med hälsovårdaren på skolan eller studieplatsen eller vuxna på ungdomsgården.
Mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats.
Föräldrar eller unga själva kan kontakta familjerådgivningen.
Där kan man tala om problem och få hjälp och stöd.
Mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats.
Familjerådgivningens telefonnummer: 044 730 7640.
Läs mer: Barns och ungas problem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Studerandehälsovårdfinska _ svenska
Ungdomsgårdar och -lokaler finska _ svenska
Problem med den mentala hälsan
Om du behöver hjälp och stöd för din mentala hälsa kan du boka en läkartid vid hälsostationen.
Läkaren bedömer situationen.
Vid behov skriver läkaren en remiss till psykiatrisk specialsjukvård.
Läs mer: Mental hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Mentalvårdstjänsterfinska _ svenska
Om du har ekonomiska problem kan du be om råd hos Mellersta Österbottens social- och hälsovårdssamkommun Soites enheter för socialarbete eller utkomststöd, tfn 040 806 5095 eller tjänstestyrningen, tfn 040 806 5093.
Om du har problem med skulder, kontakta rättshjälpsbyrån.
Du kan anlita vilken som helst rättshjälpsbyrå oberoende av din hemkommun.
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
Telefon: 029 566 1270
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Servicehandledningfinska _ svenska
Missbruksproblem
Om du har problem med alkohol, droger, läkemedel eller hasardspel kan du få vård och rehabilitering vid Porten, Mellersta Österbottens social- och hälsovårdssamkommun Soites center för missbruksproblem.
Du kan ta upp problemet med proffs inom hälsovården eller företagshälsovården, som kan slussa dig vidare i vårdsystemet, eller direkt kontakta Soites missbrukstjänster, tfn 040 8068 101.
För tillnyktrings- och avgiftningsvård debiteras en patientavgift liksom även för korttidsrehabilitering, öppen rehabilitering är gratis.
Även Karleby evangelisk-lutherska församlingssammanslutnings specialdiakoner erbjuder samtalshjälp vid missbruksproblem.
Kontaktuppgifter
Hälsovägen 4
67200 Karleby
Telefon: 040 806 8101
Läs mer: Missbruksproblem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Service för missbrukarefinska _ svenska
linkkiKarleby evangelisk-lutherska församlingssammansutning:
Karleby evangelisk-lutherska församlings arbete bland missbrukarefinska _ svenska
Problem med uppehållstillstånd
Brott
Våld
Diskriminering och rasism
Behöver du en jurist?
Död
Problem i äktenskap eller parförhållande
Skilsmässa
Problem med den mentala hälsan
Missbruksproblem
I en krissituation kan du ringa nödcentralen på numret 112.
De slussar vid behov dig vidare till socialjouren.
Du ska endast ringa nödcentralen i brådskande nödsituationer, där liv, egendom eller miljön är i fara.
Problem med uppehållstillstånd
Om du har problem eller oklarheter med ditt uppehållstillstånd kan du kontakta Migrationsverket.
Migrationsverket
Korsholmsesplanaden 45
Vasa
Läs mer: Problem med uppehållstillstånd.
Brott
Om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112.
Ring inte nödnumret om det inte är fråga om en nödsituation.
Du kan göra en polisanmälan på nätet.
Mer information finns på Polisens webbplats.
Du kan även skriva ut anmälningsblanketten på nätet och lämna in den till polisstationen.
Karleby polisstation
Karlebygatan 74
67100 Karleby
Läs mer: Brott.
Tidsbokningfinska _ svenska _ engelska
Polisamälanfinska _ svenska _ engelska
Våld
Om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112.
Läs mer: Våld.
Diskriminering och rasism
Om du misstänker att du blivit utsatt för diskriminering då du sökt arbete eller på arbetsplatsen ska du först ta upp detta på din arbetsplats.
Om saken inte kan lösas på arbetsplatsen ska du kontakta arbetarskyddet vid Regionförvaltningsverket i Västra och Inre Finland.
Besöksadress:
Regionförvaltningsverket i Västra och Inre Finland
Wollfskavägen 35
65101 Vasa
Telefon: 0295 018 450
Om du utsätts för diskriminering kan du be om hjälp av Diskrimineringsombudsmannen.
Om du fallit offer för ett rasistiskt motiverat brott kan du göra en polisanmälan på nätet eller polisstationen.
Läs mer: Diskriminering och rasism.
linkkiRegionförvaltningsverket i Västra och Inre Finland:
Regionförvaltningsverket i Västra och Inre Finlandfinska _ svenska _ engelska
Hjälp och information för personer som drabbats av etnisk diskrimineringfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Behöver du en jurist?
Juridiska tjänster är avgiftsbelagda men om du har små eller medelstora inkomster, kan du få helt eller delvis avgiftsfri rättshjälp från statens rättshjälpsbyrå.
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
Besöksadress: Ämbetshuset, Torggatan 40, 67100 Karleby
Telefon: 029 566 1270
Information om enskilda jurister finns bland annat på Finlands Advokatförbunds webbplats.
Läs mer:
Behöver du en jurist?
linkkiFinlands advokatförbund:
Finlands advokatförbundfinska _ svenska _ engelska
Död
Den evangelisk-lutherska kyrkans församlingars begravningsplatser fungerar som allmänna begravningsplatser.
Där kan även avlidna som inte är medlemmar i kyrkan begravas.
De är alltså avsedda för alla invånare i staden.
Mer information finns på Karleby kyrkliga samfällighets webbplats.
Om en närstående plötsligt dör kan du söka krishjälp vid din egen hälsostation, eller utanför tjänstetid vid samjouren för Mellersta Österbottens centralsjukhus.
De evangelisk-lutherska församlingarna i Karlebynejden erbjuder även sorggrupper.
Även församlingarnas diakonimottagningar erbjuder samtalshjälp för sorgearbetet.
Läs mer: Död.
linkkiKarleby kyrkliga samfällighet:
Karleby kyrkliga samfällighetfinska _ svenska _ engelska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Hälsostationernafinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Problem i äktenskap eller parförhållande
Vid problem i äktenskap eller parförhållande får du hjälp av Mellersta Österbottens familjerådgivningscentral som underhålls av Karleby kyrkliga samfällighets och Mellersta Österbottens social- och hälsovårdssamkommun Soites familjerådgivning.
Familjerågivningscentralen
Telefon: 050 3147 464.
Karleby familjerådgivning
67100 Karleby
tel. 044 730 7640
Läs mer: Problem i äktenskap eller parförhållande.
linkkiMellersta Österbottens Familjerådgivningscentral:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
Skilsmässa
Skilsmässa kan sökas av kvinnan, av mannen eller av båda makarna tillsammans.
Man ansöker om skilsmässa i tingsrätten.
Till att börja med görs en skriftlig skilsmässoansökan.
Österbottens tingsrätt Karleby kansli
Besöksadress: Karlebygatan 27, 67100 Karleby
Telefon: 029 56 49294
Läs mer: Skilsmässa.
Hälsovårdaren på barnrådgivningsbyrån ger råd i frågor som gäller små barns hälsa, tillväxt och utveckling.
Barnrådgivningsbyrån ger information om platser som erbjuder hjälp vid behov.
Vid problem hos unga i skolåldern hjälper exempelvis skolans hälsovårdare eller skolkuratorn.
Läs mer: Barns och ungas problem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Skolhälsovårdfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Barnrådgivningarfinska _ svenska
Du kan ta upp problem med hälsovårdaren på skolan eller studieplatsen eller vuxna på ungdomsgården.
Mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats.
Föräldrar eller unga själva kan kontakta familjerådgivningen.
Där kan man tala om problem och få hjälp och stöd.
Mer information finns på Mellersta Österbottens social- och hälsovårdssamkommun Soites webbplats.
Familjerådgivningens telefonnummer: 044 730 7640.
Läs mer: Barns och ungas problem.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Familjerådgivningfinska _ svenska
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Studerandehälsovårdfinska _ svenska
Ungdomsgårdar och -lokaler finska _ svenska
Problem med den mentala hälsan
Om du behöver hjälp och stöd för din mentala hälsa kan du boka en läkartid vid hälsostationen.
Läkaren bedömer situationen.
Vid behov skriver läkaren en remiss till psykiatrisk specialsjukvård.
Läs mer: Mental hälsa.
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Mentalvårdstjänsterfinska _ svenska
Om du har ekonomiska problem kan du be om råd hos Mellersta Österbottens social- och hälsovårdssamkommun Soites enheter för socialarbete eller utkomststöd, tfn 040 806 5095 eller tjänstestyrningen, tfn 040 806 5093.
Om du har problem med skulder, kontakta rättshjälpsbyrån.
Du kan anlita vilken som helst rättshjälpsbyrå oberoende av din hemkommun.
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Karleby verksamhetsställe
Telefon: 029 566 1270
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
Servicehandledningfinska _ svenska
Missbruksproblem
Om du har problem med alkohol, droger, läkemedel eller hasardspel kan du få vård och rehabilitering vid Porten, Mellersta Österbottens social- och hälsovårdssamkommun Soites center för missbruksproblem.
Du kan ta upp problemet med proffs inom hälsovården eller företagshälsovården, som kan slussa dig vidare i vårdsystemet, eller direkt kontakta Soites missbrukstjänster, tfn 040 8068 101.
För tillnyktrings- och avgiftningsvård debiteras en patientavgift liksom även för korttidsrehabilitering, öppen rehabilitering är gratis.
Även Karleby evangelisk-lutherska församlingssammanslutnings specialdiakoner erbjuder samtalshjälp vid missbruksproblem.
Kontaktuppgifter
