offentlig tandvård
du kan använda de kommunala tandläkartjänsterna om du har hemkommun i Esbo .
i nödfall kan du använda kommunala tjänster även om Esbo inte är din hemkommun .
du kan boka tid hos en tandläkare på Esbo tandklinikers gemensamma nummer .
Tandklinikernas tidsbeställning
tfn ( 09 ) 816.30300
du kan ringa numret på vardagar .
om du behöver besöka tandläkaren snabbt , ta kontakt med social- och hälsostationen i Kilo .
social- och hälsostationen i Kilo
Trillagatan 5
tfn ( 09 ) 816.35900
tidsbeställning på vardagar .
om du behöver akut tandläkarvård kvällstid eller under veckoslut , kan du kontakta Haartmanska sjukhuset i Helsingfors .
jourmottagningen vid Haartmanska sjukhuset har öppet vardagar kl . 14 @-@ 21 och lö @-@ sö kl . 8 @-@ 21 .
tfn ( 09 ) 310.49999 .
linkkiEsbo stad :
Mun- och tandhälsovårdenfinska _ svenska _ engelska
privat tandvård
i Esbo finns också privata tandläkare .
du kan gå till en privat tandläkare även om du inte har rätt att använda den offentliga hälsovårdens tjänster .
privat tandvård är dyrare än offentlig tandvård .
Läs mer : tandvård .
Sök tandläkarefinska
mental hälsa
om du behöver hjälp eller stöd i mental- och / eller missbruksfrågor , boka tid till en psykiatriskötare .
du kan boka tid vardagar kl . 8 @-@ 16 på numret 09.816.31300 .
linkkiEsbo stad :
information om mentalvårdstjänsternafinska _ svenska _ engelska
Psykiatriskötarna har mottagning på hälsostationerna .
mottagning för unga finns vid Nupoli .
du kan även besöka mottagningen vid kliniken för mental- och missbruksvård på servicetorget i Iso Omena utan tidsbokning måndag till fredag kl . 8.30 @-@ 10.30 och dessutom måndag till torsdag kl . 13 @-@ 14.30 .
adress : Finnviksvägen 1 , Köpcentret Iso Omena .
om du behöver krishjälp snabbt , ta kontakt med Esbo social- och krisjour ( Espoon sosiaali- ja kriisipäivystys ) .
social- och krisjouren
Åbovägen 150
tfn ( 09 ) 816.42439
öppet alla dagar dygnet runt .
linkkiEsbo stad :
social- och krisjourenfinska _ svenska _ engelska
Läs mer : mental hälsa .
linkkiFöreningen för mental hälsa i Finland :
krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
information om mentalvårdstjänsternafinska _ svenska _ engelska
sexuell hälsa
vid hälsostationernas preventivrådgivning ( ehkäisyneuvola ) får du hjälp med graviditetsprevention och familjeplanering .
ungdomar kan diskutera frågor kring sexuell hälsa med hälsovårdaren vid sin egen skola .
linkkiEsbo stad :
Preventivrådgivningsbyråerfinska _ svenska _ engelska
om du behöver en gynekologisk undersökning , ta kontakt med hälsostationen .
du kan också boka tid vid hälsostationen om du behöver ett recept för preventivmedel eller om du överväger abort .
hälsostationernas kontaktuppgifter finns på Esbo stads webbplats .
linkkiEsbo stad :
Hälsostationernafinska _ svenska _ engelska
könssjukdomar behandlas i huvudstadsregionen på polikliniken för könssjukdomar i Helsingfors .
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS :
polikliniken för könssjukdomarfinska _ svenska _ engelska
när du väntar barn
kontakta rådgivningen ( neuvola ) när du upptäcker att du är gravid .
vid rådgivningen följs moderns , fostrets och hela familjens hälsotillstånd under graviditeten .
i Esbo finns flera rådgivningsbyråer på olika håll i staden .
du kan boka tid vid alla rådgivningsbyråer på samma nummer .
rådgivning och tidsbeställning vid rådgivningsbyrån
tfn ( 09 ) 816.22800
Läs mer : när du väntar barn .
linkkiEsbo stad :
rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
förlossning
i Esbo finns Jorv sjukhus där man kan föda barn .
om du vill kan du även föda barnet på något annat sjukhus inom samkommunen Helsingfors och Nylands sjukvårdsdistrikt ( HNS ) .
mer information hittar du på HNS webbplats .
Läs mer : förlossning .
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS :
Förlossningfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt :
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
handikappade personer
Esbo stad ordnar olika tjänster för handikappade , till exempel dagverksamhet och färdtjänster .
personer som har sin hemkommun i Esbo har rätt till dessa tjänster .
du kan ansöka om tjänster och stödfunktioner hos stadens socialarbetare .
mer information om tjänsterna för handikappade hittar du på Esbo stads handikappservice .
Esbo handikappservice
Kamrersvägen 2 A , vån . 4
tfn ( 09 ) 816.45285
Läs mer : handikappade personer
linkkiEsbo stad :
kontaktuppgifter till socialarbetarefinska _ svenska _ engelska
linkkiEsbo stad :
stödtjänster för handikappadefinska _ svenska _ engelska
ett handikappat barn
om du har ett handikappat barn kan du kontakta socialarbetaren vid handikappservicen för ditt eget område vammaispalvelut ( at ) espoo.fi .
frågor som rör skolgången för ett handikappat barn kan du ställa till skolväsendet ( opetustoimi ) samt till servicehandledaren för skolelever ( koululaisten palveluohjaaja ) .
Läs mer : ett handikappat barn
linkkiEsbo stad :
kontaktuppgifter till utbildningsväsendetfinska _ engelska
hälsovårdstjänsterna i Esbo
tandvården
mental hälsa
sexuell hälsa
när du väntar barn
handikappade personer
ring nödnumret 112 om det är fråga om en brådskande nödsituation .
ring nödnumret till exempel vid en allvarlig olycka eller när någon drabbas av en sjukdomsattack .
ring inte nödnumret om det inte är en nödsituation .
om du har din hemkommun i Esbo kan du utnyttja de offentliga hälsovårdstjänsterna .
offentliga hälsovårdstjänster tillhandahålls vid hälsostationer , tandkliniker , rådgivningsbyråer och sjukhus .
om du inte har rätt till de offentliga hälsovårdstjänsterna , kan du söka hjälp på en privat läkarstation .
på en privat läkarstation måste du betala samtliga kostnader själv .
Läs mer : hälsa .
hälsovårdstjänsterna i Esbo
offentliga hälsovårdstjänster tillhandahålls av hälsostationerna ( terveysasema ) .
hälsostationerna har öppet vardagar klockan 8 @-@ 16 .
på hälsostationerna finns vanligtvis läkarens , sjukskötarens och hälsovårdarens mottagningar .
du kan boka tid på hälsostationen per telefon .
på Esbo stads webbplats finns kontaktuppgifterna och telefonnumren till hälsostationerna .
när du ringer hälsostationen , besvaras ditt samtal inte nödvändigtvis omedelbart .
ditt nummer sparas dock i en automat och du blir uppringd .
kom i tid till mottagningen .
om du inte kan komma till mottagningen , kom ihåg att avboka din tid senast föregående vardag före klockan 14 .
om du behöver första hjälpen snabbt , kan du komma till hälsostationen utan tidsbeställning .
linkkiEsbo stad :
Hälsostationernafinska _ svenska _ engelska
linkkiEsbo stad :
Hälsovårdscentralsavgifterfinska _ svenska
privata hälsovårdstjänster
Vem som helst kan gå till en privat hälsostation .
också de personer som inte har rätt till den offentliga hälsovården i Finland kan besöka privata hälsostationer .
på en privat hälsostation måste kunden själv betala samtliga kostnader .
i Esbo finns flera privata läkarstationer .
kontaktuppgifter till privata läkare hittar du till exempel på Internet .
linkkietsilaakari.fi :
privata hälsovårdstjänsterfinska
privat läkarstationfinska _ svenska _ engelska
privat läkarstationfinska _ svenska _ engelska
läkemedel
information om köp av läkemedel hittar du på InfoFinlands sida Läkemedel .
hälsovård för papperslösa
i Helsingfors finns Global Clinic , där personer som vistas i Finland utan tillstånd kan få primärhälsovård .
tjänsterna vid Global Clinic är avgiftsfria för kunderna .
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter .
för att skydda kunderna uppges inte klinikens adress eller öppettider offentligt .
telefonnumret till Global Clinic i Helsingfors är 044.977.4547 .
Samtalet besvaras av en sjukskötare eller en läkare .
hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Läs mer : hälsovårdstjänster i Finland
kvällstid och under veckoslut har hälsostationen stängt .
då vårdas akuta sjukfall och olycksfall på jourmottagningen ( päivystys ) .
den närmaste jourmottagningen för vuxna finns vid Jorv sjukhus .
ring den kostnadsfria Jourhjälpen på tfn 116.117 innan du kommer till jourmottagningen .
jourmottagningen vid Jorv sjukhus
Åbovägen 150
tfn ( 09 ) 4711
Jourmottagningar för barn under 16 år finns i Jorv och på Barnkliniken i Helsingfors .
du behöver inte boka tid på jourmottagningen .
linkkiEsbo stad :
Jourmottagningarfinska _ svenska _ engelska
Läs mer : hälsovårdstjänster i Finland
barns hälsa
i hälsovården av 1 @-@ 6 @-@ åriga barn får man hjälp av rådgivningsbyråns ( neuvola ) hälsovårdare och läkare .
dem kan du fråga om råd och få hjälp med fostran av barn .
på rådgivningsbyrån följs att barnet är friskt och växer som det ska .
i Esbo finns flera rådgivningsbyråer på olika håll i staden .
rådgivningsbyråernas kontaktuppgifter finns på Esbo stads webbplats .
du kan boka tid vid alla rådgivningsbyråer på samma nummer .
om ett barn blir sjukt och behöver snabbt vård , ta kontakt med hälsostationen ( terveysasema ) .
Skolhälsovårdaren har hand om skolbarns hälsa .
under kvällar och veckoslut finns jourmottagningen för barn under 16 år vid Jorv sjukhus och på Barnkliniken i Helsingfors .
du kan också ta ditt barn till en privat läkarstation .
Läs mer : barns hälsa .
linkkiEsbo stad :
Barnrådgivningsbyråernas tjänsterfinska _ svenska _ engelska
linkkiEsbo stad :
rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
linkkiEsbo stad :
Hälsostationernafinska _ svenska _ engelska
linkkiEsbo stad :
information om hälsovården för skolbarnfinska _ svenska _ engelska
linkkiEsbo stad :
Jourmottagningarfinska _ svenska _ engelska
tandvården
offentlig tandvård
du kan använda de kommunala tandläkartjänsterna om du har hemkommun i Esbo .
i nödfall kan du använda kommunala tjänster även om Esbo inte är din hemkommun .
du kan boka tid hos en tandläkare på Esbo tandklinikers gemensamma nummer .
Tandklinikernas tidsbeställning
tfn ( 09 ) 816.30300
du kan ringa numret på vardagar .
om du behöver besöka tandläkaren snabbt , ta kontakt med social- och hälsostationen i Kilo .
social- och hälsostationen i Kilo
Trillagatan 5
tfn ( 09 ) 816.35900
tidsbeställning på vardagar .
om du behöver akut tandläkarvård kvällstid eller under veckoslut , kan du kontakta Haartmanska sjukhuset i Helsingfors .
jourmottagningen vid Haartmanska sjukhuset har öppet vardagar kl . 14 @-@ 21 och lö @-@ sö kl . 8 @-@ 21 .
tfn ( 09 ) 310.49999 .
linkkiEsbo stad :
Mun- och tandhälsovårdenfinska _ svenska _ engelska
privat tandvård
i Esbo finns också privata tandläkare .
du kan gå till en privat tandläkare även om du inte har rätt att använda den offentliga hälsovårdens tjänster .
privat tandvård är dyrare än offentlig tandvård .
Läs mer : tandvård .
Sök tandläkarefinska
mental hälsa
om du behöver hjälp eller stöd i mental- och / eller missbruksfrågor , boka tid till en psykiatriskötare .
du kan boka tid vardagar kl . 8 @-@ 16 på numret 09.816.31300 .
linkkiEsbo stad :
information om mentalvårdstjänsternafinska _ svenska _ engelska
Psykiatriskötarna har mottagning på hälsostationerna .
mottagning för unga finns vid Nupoli .
du kan även besöka mottagningen vid kliniken för mental- och missbruksvård på servicetorget i Iso Omena utan tidsbokning måndag till fredag kl . 8.30 @-@ 10.30 och dessutom måndag till torsdag kl . 13 @-@ 14.30 .
adress : Finnviksvägen 1 , Köpcentret Iso Omena .
om du behöver krishjälp snabbt , ta kontakt med Esbo social- och krisjour ( Espoon sosiaali- ja kriisipäivystys ) .
social- och krisjouren
Åbovägen 150
tfn ( 09 ) 816.42439
öppet alla dagar dygnet runt .
linkkiEsbo stad :
social- och krisjourenfinska _ svenska _ engelska
Läs mer : mental hälsa .
linkkiFöreningen för mental hälsa i Finland :
krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
information om mentalvårdstjänsternafinska _ svenska _ engelska
sexuell hälsa
vid hälsostationernas preventivrådgivning ( ehkäisyneuvola ) får du hjälp med graviditetsprevention och familjeplanering .
ungdomar kan diskutera frågor kring sexuell hälsa med hälsovårdaren vid sin egen skola .
linkkiEsbo stad :
Preventivrådgivningsbyråerfinska _ svenska _ engelska
om du behöver en gynekologisk undersökning , ta kontakt med hälsostationen .
du kan också boka tid vid hälsostationen om du behöver ett recept för preventivmedel eller om du överväger abort .
hälsostationernas kontaktuppgifter finns på Esbo stads webbplats .
linkkiEsbo stad :
Hälsostationernafinska _ svenska _ engelska
könssjukdomar behandlas i huvudstadsregionen på polikliniken för könssjukdomar i Helsingfors .
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS :
polikliniken för könssjukdomarfinska _ svenska _ engelska
när du väntar barn
kontakta rådgivningen ( neuvola ) när du upptäcker att du är gravid .
vid rådgivningen följs moderns , fostrets och hela familjens hälsotillstånd under graviditeten .
i Esbo finns flera rådgivningsbyråer på olika håll i staden .
du kan boka tid vid alla rådgivningsbyråer på samma nummer .
rådgivning och tidsbeställning vid rådgivningsbyrån
tfn ( 09 ) 816.22800
Läs mer : när du väntar barn .
linkkiEsbo stad :
rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
förlossning
i Esbo finns Jorv sjukhus där man kan föda barn .
om du vill kan du även föda barnet på något annat sjukhus inom samkommunen Helsingfors och Nylands sjukvårdsdistrikt ( HNS ) .
mer information hittar du på HNS webbplats .
Läs mer : förlossning .
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS :
Förlossningfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt :
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
handikappade personer
Esbo stad ordnar olika tjänster för handikappade , till exempel dagverksamhet och färdtjänster .
personer som har sin hemkommun i Esbo har rätt till dessa tjänster .
du kan ansöka om tjänster och stödfunktioner hos stadens socialarbetare .
mer information om tjänsterna för handikappade hittar du på Esbo stads handikappservice .
Esbo handikappservice
Kamrersvägen 2 A , vån . 4
tfn ( 09 ) 816.45285
handikappade personerlinkkiEsbo stad :
linkkiEsbo stad :
stödtjänster för handikappadefinska _ svenska _ engelska
ett handikappat barn
om du har ett handikappat barn kan du kontakta socialarbetaren vid handikappservicen för ditt eget område vammaispalvelut ( at ) espoo.fi .
frågor som rör skolgången för ett handikappat barn kan du ställa till skolväsendet ( opetustoimi ) samt till servicehandledaren för skolelever ( koululaisten palveluohjaaja ) .
Läs mer : ett handikappat barn
linkkiEsbo stad :
kontaktuppgifter till utbildningsväsendetfinska _ engelska
hälsovårdstjänsterna i Esbo
tandvården
mental hälsa
sexuell hälsa
när du väntar barn
handikappade personer
ring nödnumret 112 om det är fråga om en brådskande nödsituation .
ring nödnumret till exempel vid en allvarlig olycka eller när någon drabbas av en sjukdomsattack .
ring inte nödnumret om det inte är en nödsituation .
om du har din hemkommun i Esbo kan du utnyttja de offentliga hälsovårdstjänsterna .
offentliga hälsovårdstjänster tillhandahålls vid hälsostationer , tandkliniker , rådgivningsbyråer och sjukhus .
om du inte har rätt till de offentliga hälsovårdstjänsterna , kan du söka hjälp på en privat läkarstation .
på en privat läkarstation måste du betala samtliga kostnader själv .
Läs mer : hälsa .
hälsovårdstjänsterna i Esbo
offentliga hälsovårdstjänster tillhandahålls av hälsostationerna ( terveysasema ) .
hälsostationerna har öppet vardagar klockan 8 @-@ 16 .
på hälsostationerna finns vanligtvis läkarens , sjukskötarens och hälsovårdarens mottagningar .
du kan boka tid på hälsostationen per telefon .
på Esbo stads webbplats finns kontaktuppgifterna och telefonnumren till hälsostationerna .
när du ringer hälsostationen , besvaras ditt samtal inte nödvändigtvis omedelbart .
ditt nummer sparas dock i en automat och du blir uppringd .
kom i tid till mottagningen .
om du inte kan komma till mottagningen , kom ihåg att avboka din tid senast föregående vardag före klockan 14 .
om du behöver första hjälpen snabbt , kan du komma till hälsostationen utan tidsbeställning .
linkkiEsbo stad :
Hälsostationernafinska _ svenska _ engelska
linkkiEsbo stad :
Hälsovårdscentralsavgifterfinska _ svenska
privata hälsovårdstjänster
Vem som helst kan gå till en privat hälsostation .
också de personer som inte har rätt till den offentliga hälsovården i Finland kan besöka privata hälsostationer .
på en privat hälsostation måste kunden själv betala samtliga kostnader .
i Esbo finns flera privata läkarstationer .
kontaktuppgifter till privata läkare hittar du till exempel på Internet .
linkkietsilaakari.fi :
privata hälsovårdstjänsterfinska
privat läkarstationfinska _ svenska _ engelska
privat läkarstationfinska _ svenska _ engelska
läkemedel
information om köp av läkemedel hittar du på InfoFinlands sida Läkemedel .
hälsovård för papperslösa
i Helsingfors finns Global Clinic , där personer som vistas i Finland utan tillstånd kan få primärhälsovård .
tjänsterna vid Global Clinic är avgiftsfria för kunderna .
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter .
för att skydda kunderna uppges inte klinikens adress eller öppettider offentligt .
telefonnumret till Global Clinic i Helsingfors är 044.977.4547 .
Samtalet besvaras av en sjukskötare eller en läkare .
hälsotjänster för papperslösafinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Läs mer : hälsovårdstjänster i Finland
kvällstid och under veckoslut har hälsostationen stängt .
då vårdas akuta sjukfall och olycksfall på jourmottagningen ( päivystys ) .
den närmaste jourmottagningen för vuxna finns vid Jorv sjukhus .
ring den kostnadsfria Jourhjälpen på tfn 116.117 innan du kommer till jourmottagningen .
jourmottagningen vid Jorv sjukhus
Åbovägen 150
tfn ( 09 ) 4711
Jourmottagningar för barn under 16 år finns i Jorv och på Barnkliniken i Helsingfors .
du behöver inte boka tid på jourmottagningen .
linkkiEsbo stad :
Jourmottagningarfinska _ svenska _ engelska
Läs mer : hälsovårdstjänster i Finland
barns hälsa
i hälsovården av 1 @-@ 6 @-@ åriga barn får man hjälp av rådgivningsbyråns ( neuvola ) hälsovårdare och läkare .
dem kan du fråga om råd och få hjälp med fostran av barn .
på rådgivningsbyrån följs att barnet är friskt och växer som det ska .
i Esbo finns flera rådgivningsbyråer på olika håll i staden .
rådgivningsbyråernas kontaktuppgifter finns på Esbo stads webbplats .
du kan boka tid vid alla rådgivningsbyråer på samma nummer .
om ett barn blir sjukt och behöver snabbt vård , ta kontakt med hälsostationen ( terveysasema ) .
Skolhälsovårdaren har hand om skolbarns hälsa .
under kvällar och veckoslut finns jourmottagningen för barn under 16 år vid Jorv sjukhus och på Barnkliniken i Helsingfors .
du kan också ta ditt barn till en privat läkarstation .
Läs mer : barns hälsa .
linkkiEsbo stad :
Barnrådgivningsbyråernas tjänsterfinska _ svenska _ engelska
linkkiEsbo stad :
rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
linkkiEsbo stad :
Hälsostationernafinska _ svenska _ engelska
linkkiEsbo stad :
information om hälsovården för skolbarnfinska _ svenska _ engelska
linkkiEsbo stad :
Jourmottagningarfinska _ svenska _ engelska
tandvården
offentlig tandvård
du kan använda de kommunala tandläkartjänsterna om du har hemkommun i Esbo .
i nödfall kan du använda kommunala tjänster även om Esbo inte är din hemkommun .
du kan boka tid hos en tandläkare på Esbo tandklinikers gemensamma nummer .
Tandklinikernas tidsbeställning
tfn ( 09 ) 816.30300
du kan ringa numret på vardagar .
om du behöver besöka tandläkaren snabbt , ta kontakt med social- och hälsostationen i Kilo .
social- och hälsostationen i Kilo
Trillagatan 5
tfn ( 09 ) 816.35900
tidsbeställning på vardagar .
om du behöver akut tandläkarvård kvällstid eller under veckoslut , kan du kontakta Haartmanska sjukhuset i Helsingfors .
jourmottagningen vid Haartmanska sjukhuset har öppet vardagar kl . 14 @-@ 21 och lö @-@ sö kl . 8 @-@ 21 .
tfn ( 09 ) 310.49999 .
linkkiEsbo stad :
Mun- och tandhälsovårdenfinska _ svenska _ engelska
privat tandvård
i Esbo finns också privata tandläkare .
du kan gå till en privat tandläkare även om du inte har rätt att använda den offentliga hälsovårdens tjänster .
privat tandvård är dyrare än offentlig tandvård .
Läs mer : tandvård .
Sök tandläkarefinska
mental hälsa
om du behöver hjälp eller stöd i mental- och / eller missbruksfrågor , boka tid till en psykiatriskötare .
du kan boka tid vardagar kl . 8 @-@ 16 på numret 09.816.31300 .
linkkiEsbo stad :
information om mentalvårdstjänsternafinska _ svenska _ engelska
Psykiatriskötarna har mottagning på hälsostationerna .
mottagning för unga finns vid Nupoli .
du kan även besöka mottagningen vid kliniken för mental- och missbruksvård på servicetorget i Iso Omena utan tidsbokning måndag till fredag kl . 8.30 @-@ 10.30 och dessutom måndag till torsdag kl . 13 @-@ 14.30 .
adress : Finnviksvägen 1 , Köpcentret Iso Omena .
om du behöver krishjälp snabbt , ta kontakt med Esbo social- och krisjour ( Espoon sosiaali- ja kriisipäivystys ) .
social- och krisjouren
Åbovägen 150
tfn ( 09 ) 816.42439
öppet alla dagar dygnet runt .
linkkiEsbo stad :
social- och krisjourenfinska _ svenska _ engelska
Läs mer : mental hälsa .
linkkiFöreningen för mental hälsa i Finland :
krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
information om mentalvårdstjänsternafinska _ svenska _ engelska
sexuell hälsa
vid hälsostationernas preventivrådgivning ( ehkäisyneuvola ) får du hjälp med graviditetsprevention och familjeplanering .
ungdomar kan diskutera frågor kring sexuell hälsa med hälsovårdaren vid sin egen skola .
linkkiEsbo stad :
Preventivrådgivningsbyråerfinska _ svenska _ engelska
om du behöver en gynekologisk undersökning , ta kontakt med hälsostationen .
du kan också boka tid vid hälsostationen om du behöver ett recept för preventivmedel eller om du överväger abort .
hälsostationernas kontaktuppgifter finns på Esbo stads webbplats .
linkkiEsbo stad :
Hälsostationernafinska _ svenska _ engelska
könssjukdomar behandlas i huvudstadsregionen på polikliniken för könssjukdomar i Helsingfors .
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS :
polikliniken för könssjukdomarfinska _ svenska _ engelska
Läs mer : Sexualhälsa
när du väntar barn
kontakta rådgivningen ( neuvola ) när du upptäcker att du är gravid .
vid rådgivningen följs moderns , fostrets och hela familjens hälsotillstånd under graviditeten .
i Esbo finns flera rådgivningsbyråer på olika håll i staden .
du kan boka tid vid alla rådgivningsbyråer på samma nummer .
rådgivning och tidsbeställning vid rådgivningsbyrån
tfn ( 09 ) 816.22800
Läs mer : graviditet och förlossning .
linkkiEsbo stad :
rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
förlossning
i Esbo finns Jorv sjukhus där man kan föda barn .
om du vill kan du även föda barnet på något annat sjukhus inom samkommunen Helsingfors och Nylands sjukvårdsdistrikt ( HNS ) .
mer information hittar du på HNS webbplats .
linkkiHelsingfors och Nylands sjukvårdsdistrikt HNS :
Förlossningfinska _ svenska _ engelska
linkkiHelsingfors och Nylands sjukvårdsdistrikt :
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
handikappade personer
Esbo stad ordnar olika tjänster för handikappade , till exempel dagverksamhet och färdtjänster .
personer som har sin hemkommun i Esbo har rätt till dessa tjänster .
du kan ansöka om tjänster och stödfunktioner hos stadens socialarbetare .
mer information om tjänsterna för handikappade hittar du på Esbo stads handikappservice .
Esbo handikappservice
Kamrersvägen 2 A , vån . 4
tfn ( 09 ) 816.45285
Läs mer : handikappade personer
linkkiEsbo stad :
stödtjänster för handikappadefinska _ svenska _ engelska
ett handikappat barn
om du har ett handikappat barn kan du kontakta socialarbetaren vid handikappservicen för ditt eget område vammaispalvelut ( at ) espoo.fi .
frågor som rör skolgången för ett handikappat barn kan du ställa till skolväsendet ( opetustoimi ) samt till servicehandledaren för skolelever ( koululaisten palveluohjaaja ) .
Läs mer : ett handikappat barn
linkkiEsbo stad :
kontaktuppgifter till utbildningsväsendetfinska _ engelska
detta innehåll finns inte på det språk som du har valt .
Välj något annat språk .
finska
detta innehåll finns inte på det språk som du har valt .
Välj något annat språk .
finska
detta innehåll finns inte på det språk som du har valt .
Välj något annat språk .
finska
dagvård
förskoleundervisning
grundläggande utbildning
hemspråksundervisning för invandrare
yrkesutbildning
gymnasium
stöd och handledning för unga
Högskoleutbildning
andra studiemöjligheter
dagvård
i Esbo finns både kommunala och privata daghem .
i Esbo finns dessutom familjedagvårdare .
dagvård fås på finska och på svenska .
Ansök om dagvårdsplats minst fyra månader innan barnet ska börja i dagvården .
om du till exempel oväntat får arbete eller en studieplats kan du ansöka om vårdplats senare .
när du ansöker om vårdplats ska du fylla i en ansökningsblankett .
du kan också söka dagvårdsplats via Internet .
familjer som bor i Esbo kan också söka dagvårdsplats till sitt barn i Helsingfors , Vanda eller Grankulla .
du ska ändå lämna in din ansökan i Esbo .
mer information får du via tjänsten Helsingforsregionen.fi .
Läs mer : dagvård .
linkkiEsbo stad :
dagvårdfinska _ svenska _ engelska
linkkiEsbo stad :
ansökan om dagvårdsplatsfinska
linkkiEsbo stad :
Servicepunktfinska _ svenska _ engelska
linkkiEsbo stad :
Dagvårdens samanvändningsområdefinska _ svenska _ engelska
förskoleundervisning
i Esbo anordnas förskoleundervisningen ( esiopetus ) i daghemmen .
förskoleundervisning ges på finska och på svenska .
till förskoleundervisningen anmäler man sig via Esbo stads webbplats .
förskoleundervisningen börjar i augusti .
ansökningstiden är vanligtvis i januari .
i frågor kring barndagvård och förskoleundervisning kan du också kontakta daghemsföreståndarna eller stadens chef för småbarnsfostran ( varhaiskasvatuspäällikkö ) .
kontaktuppgifterna finns på stadens webbplats .
Läs mer : förskoleundervisning .
linkkiEsbo stad :
förskoleundervisningfinska _ svenska _ engelska
linkkiEsbo stad :
ansökan till förskoleundervisningfinska _ svenska _ engelska
grundläggande utbildning
