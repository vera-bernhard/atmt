I Esbo finns finskspråkiga och svenskspråkiga grundskolor (peruskoulu).
Undervisning kan även fås på engelska.
Skolan börjar vanligtvis det året då barnet fyller sju år.
Anmälan till grundskolan ska göras på förhand.
Anmälningstiden är vanligtvis i januari.
På stadens webbplats hittar du kontaktuppgifterna till skolorna och mer information om anmälan.
Om du har frågor om den grundläggande utbildningen kan du kontakta Resultatenheten för den finskspråkiga undervisningen (Suomenkielisen opetuksen tulosyksikkö).
Resultatenheten för den finskspråkiga undervisningen
Kamrersvägen 3 B
Tfn (09) 816 52044 och (09) 816 52043
Grundläggande utbildning.
linkkiEsbo stad:
Grundläggande utbildningfinska _ svenska _ engelska
linkkiEsbo stad:
Anmälan till skolanfinska _ svenska _ engelska
linkkiEsbo stad:
Espoo International Schoolfinska _ engelska
Internationella skolor i huvudstadsregionenfinska
linkkiExpatFinland.fi:
Internationella skolor i huvudstadsregionenengelska
linkkiEsbo stad:
Eftermiddagsverksamhetfinska _ engelska
Hemspråksundervisning för invandrare
Barn med invandrarbakgrund och barn från tvåspråkiga familjer kan få hemspråksundervisning (oman äidinkielen opetus) om tillräckligt många barn anmäler sig till gruppen för det egna språket.
Undervisning ges två timmar i veckan.
Anmälan till hemspråksundervisning görs varje år i mars.
Mer information hittar du på Esbo stads webbplats.
linkkiEsbo stad:
Förberedande undervisning för barn i förskoleåldern(pdf, 100 kb)finska _ engelska _ ryska _ estniska _ somaliska _ kinesiska _ arabiska _ kurdiska _ albanska
linkkiEsbo stad:
Förberedande undervisning för barn i förskoleåldernfinska _ engelska
linkkiEsbo stad:
Hemspråksundervisningfinska _ engelska
Yrkesutbildning
På Omnia kan man studera många olika yrken.
På Omnia ordnas för invandrare utbildning som förbereder dem på yrkesutbildning.
Den förberedande utbildningen är avsedd för unga och vuxna, som är intresserade av yrkesstudier och vill förbättra sina kunskaper i finska..
Esbobor kan också ansöka till yrkesskolorna i Helsingfors och Vanda.
Läs mer: Yrkesutbildning
Yrkesutbildningfinska _ engelska
linkkiEsbo stad:
Yrkesläroanstalterfinska _ engelska
Yrkesläroanstalterfinska _ svenska _ engelska
linkkiVanda stad:
Yrkesutbildningfinska _ svenska
Gymnasium
I Esbo finns elva finskspråkiga och ett svenskspråkigt gymnasium (lukio).
I två av gymnasierna i Esbo finns en engelskspråkig IB-linje.
Ungdomar från Esbo kan också söka till gymnasier i andra städer.
I Esbo finns ett vuxengymnasium (aikuislukio) där vuxna kan avlägga gymnasie- och studentexamen.
På gymnasiet kan man även höja vitsorden i sitt avgångsbetyg eller studera enskilda ämnen.
Invandrarungdomar kan dessutom studera finska och avlägga grundskolans lärokurs.
I gymnasiet Leppävaaran lukio ordnas för invandrare och utlänningar utbildning som förbereder dem på gymnasiet.
Utbildningen är avsedd för unga som vill studera på gymnasiet, men vars språkkunskaper inte är tillräckliga för gymnasiestudier.
Läs mer: Gymnasium
linkkiEsbo stad:
Gymnasierfinska _ svenska _ engelska
linkkiEsbo stad:
Vuxengymnasietfinska
linkkiEsbo stad:
Gymnasieförberedande utbildning för invandrarefinska _ engelska
linkkiEsbo vuxengymnasium Omnia:
Grundläggande utbildning för invandrarefinska
Om du är under 30 år gammal kan du få råd och handledning via Ohjaamo-tjänsten.
Ohjaamos personal hjälper dig om du inte har ett arbete eller en studieplats.
Du kan även fråga om andra saker, som till exempel boende eller ekonomiska frågor.
Kontaktuppgifter:
Fågelbergavägen 2 A
Puh. 040 126 7513
linkkiEsbo stad:
Ohjaamofinska _ svenska _ engelska
Högskoleutbildning
I Esbo finns tre högskolor:
yrkeshögskolan Laurea
yrkeshögskolan Metropolia.
Vid högskolorna kan du avlägga högskoleexamen.
Mer information finns på Aalto-universitetets, Laureas och Metropolias webbplatser.
Också i Helsingfors finns det universitet och yrkeshögskolor där man kan studera inom många områden.
Mer information hittar du på Helsingfors stads webbplats.
Läs mer: Högskoleutbildning
Universitet inom teknik, konst och ekonomifinska _ svenska _ engelska
Yrkeshögskolafinska _ engelska
linkkiMetropolia:
Yrkeshögskolafinska _ engelska
Högskolorfinska
Andra studiemöjligheter
Vid Esbo arbetarinstitut (Espoon työväenopisto) kan du studera till exempel språk, handarbete och matlagning eller delta i ledd motion.
Kurserna är avgiftsbelagda. Kurser anordnas både dagtid och kvällstid.
Vid arbetarinstitutet kan vem som helst studera.
Vid Esbo bildkonstskola (Espoon kuvataidekoulu) kan barn och unga studera bildkonst.
Studierna är avgiftsbelagda.
Vid Esbo musikinstitut (Espoon musiikkiopisto) kan barn och vuxna studera musik.
Läs mer: Andra studiemöjligheter
linkkiEsbo stad:
Arbetarinstitutetfinska _ svenska _ engelska
linkkiEsbo biIdkonstskola:
Bildkonst för barn och ungafinska _ svenska _ engelska
linkkiEsbo musikinstitut:
Musikundervisning för barn och vuxnafinska _ engelska
Dagvård
Förskoleundervisning
Grundläggande utbildning
Hemspråksundervisning för invandrare
Yrkesutbildning
Gymnasium
Stöd och handledning för unga
Högskoleutbildning
Andra studiemöjligheter
Dagvård
I Esbo finns både kommunala och privata daghem.
I Esbo finns dessutom familjedagvårdare.
Dagvård fås på finska och på svenska.
Ansök om dagvårdsplats minst fyra månader innan barnet ska börja i dagvården.
Om du till exempel oväntat får arbete eller en studieplats kan du ansöka om vårdplats senare.
När du ansöker om vårdplats ska du fylla i en ansökningsblankett.
Du kan också söka dagvårdsplats via Internet.
Familjer som bor i Esbo kan också söka dagvårdsplats till sitt barn i Helsingfors, Vanda eller Grankulla.
Du ska ändå lämna in din ansökan i Esbo.
Mer information får du via tjänsten Helsingforsregionen.fi.
Läs mer: Dagvård.
linkkiEsbo stad:
Dagvårdfinska _ svenska _ engelska
linkkiEsbo stad:
Ansökan om dagvårdsplatsfinska
linkkiEsbo stad:
Servicepunktfinska _ svenska _ engelska
linkkiEsbo stad:
Dagvårdens samanvändningsområdefinska _ svenska _ engelska
Förskoleundervisning
I Esbo anordnas förskoleundervisningen (esiopetus) i daghemmen.
Förskoleundervisning ges på finska och på svenska.
Till förskoleundervisningen anmäler man sig via Esbo stads webbplats.
Förskoleundervisningen börjar i augusti.
Ansökningstiden är vanligtvis i januari.
I frågor kring barndagvård och förskoleundervisning kan du också kontakta daghemsföreståndarna eller stadens chef för småbarnsfostran (varhaiskasvatuspäällikkö).
Kontaktuppgifterna finns på stadens webbplats.
Läs mer: Förskoleundervisning.
linkkiEsbo stad:
Förskoleundervisningfinska _ svenska _ engelska
linkkiEsbo stad:
Ansökan till förskoleundervisningfinska _ engelska
Grundläggande utbildning
I Esbo finns finskspråkiga och svenskspråkiga grundskolor (peruskoulu).
Undervisning kan även fås på engelska.
Skolan börjar vanligtvis det året då barnet fyller sju år.
Anmälan till grundskolan ska göras på förhand.
Anmälningstiden är vanligtvis i januari.
På stadens webbplats hittar du kontaktuppgifterna till skolorna och mer information om anmälan.
Om du har frågor om den grundläggande utbildningen kan du kontakta Resultatenheten för den finskspråkiga undervisningen (Suomenkielisen opetuksen tulosyksikkö).
Resultatenheten för den finskspråkiga undervisningen
Kamrersvägen 3 B
Tfn (09) 816 52044 och (09) 816 52043
Grundläggande utbildning.
linkkiEsbo stad:
Grundläggande utbildningfinska _ svenska _ engelska
linkkiEsbo stad:
Anmälan till skolanfinska _ svenska _ engelska
linkkiEsbo stad:
Espoo International Schoolfinska _ engelska
Internationella skolor i huvudstadsregionenfinska
linkkiExpatFinland.fi:
Internationella skolor i huvudstadsregionenengelska
linkkiEsbo stad:
Eftermiddagsverksamhetfinska _ engelska
Hemspråksundervisning för invandrare
Barn med invandrarbakgrund och barn från tvåspråkiga familjer kan få hemspråksundervisning (oman äidinkielen opetus) om tillräckligt många barn anmäler sig till gruppen för det egna språket.
Undervisning ges två timmar i veckan.
Anmälan till hemspråksundervisning görs varje år i mars.
Mer information hittar du på Esbo stads webbplats.
linkkiEsbo stad:
Förberedande undervisning för barn i förskoleåldern(pdf, 100 kb)finska _ engelska _ ryska _ estniska _ somaliska _ kinesiska _ arabiska _ kurdiska _ albanska
linkkiEsbo stad:
Förberedande undervisning för barn i förskoleåldernfinska _ engelska
linkkiEsbo stad:
Hemspråksundervisningfinska _ engelska
Yrkesutbildning
På Omnia kan man studera många olika yrken.
På Omnia ordnas för invandrare utbildning som förbereder dem på yrkesutbildning.
Den förberedande utbildningen är avsedd för unga och vuxna, som är intresserade av yrkesstudier och vill förbättra sina kunskaper i finska..
Esbobor kan också ansöka till yrkesskolorna i Helsingfors och Vanda.
Läs mer: Yrkesutbildning
Yrkesutbildningfinska _ engelska
linkkiEsbo stad:
Yrkesläroanstalterfinska _ engelska
Yrkesläroanstalterfinska _ svenska _ engelska
linkkiVanda stad:
Yrkesutbildningfinska _ svenska
Gymnasium
I Esbo finns elva finskspråkiga och ett svenskspråkigt gymnasium (lukio).
I två av gymnasierna i Esbo finns en engelskspråkig IB-linje.
Ungdomar från Esbo kan också söka till gymnasier i andra städer.
I Esbo finns ett vuxengymnasium (aikuislukio) där vuxna kan avlägga gymnasie- och studentexamen.
På gymnasiet kan man även höja vitsorden i sitt avgångsbetyg eller studera enskilda ämnen.
Invandrarungdomar kan dessutom studera finska och avlägga grundskolans lärokurs.
I gymnasiet Leppävaaran lukio ordnas för invandrare och utlänningar utbildning som förbereder dem på gymnasiet.
Utbildningen är avsedd för unga som vill studera på gymnasiet, men vars språkkunskaper inte är tillräckliga för gymnasiestudier.
Läs mer: Gymnasium
linkkiEsbo stad:
Gymnasierfinska _ svenska _ engelska
linkkiEsbo stad:
Vuxengymnasietfinska
linkkiEsbo stad:
Gymnasieförberedande utbildning för invandrarefinska _ engelska
linkkiEsbo vuxengymnasium Omnia:
Grundläggande utbildning för invandrarefinska
Om du är under 30 år gammal kan du få råd och handledning via Ohjaamo-tjänsten.
Ohjaamos personal hjälper dig om du inte har ett arbete eller en studieplats.
Du kan även fråga om andra saker, som till exempel boende eller ekonomiska frågor.
Kontaktuppgifter:
Fågelbergavägen 2 A
Puh. 040 126 7513
linkkiEsbo stad:
Ohjaamofinska _ svenska _ engelska
Högskoleutbildning
I Esbo finns tre högskolor:
yrkeshögskolan Laurea
yrkeshögskolan Metropolia.
Vid högskolorna kan du avlägga högskoleexamen.
Mer information finns på Aalto-universitetets, Laureas och Metropolias webbplatser.
Också i Helsingfors finns det universitet och yrkeshögskolor där man kan studera inom många områden.
Mer information hittar du på Helsingfors stads webbplats.
Läs mer: Högskoleutbildning
Universitet inom teknik, konst och ekonomifinska _ svenska _ engelska
Yrkeshögskolafinska _ engelska
linkkiMetropolia:
Yrkeshögskolafinska _ engelska
Högskolorfinska
Andra studiemöjligheter
Vid Esbo arbetarinstitut (Espoon työväenopisto) kan du studera till exempel språk, handarbete och matlagning eller delta i ledd motion.
Kurserna är avgiftsbelagda. Kurser anordnas både dagtid och kvällstid.
Vid arbetarinstitutet kan vem som helst studera.
Vid Esbo bildkonstskola (Espoon kuvataidekoulu) kan barn och unga studera bildkonst.
Studierna är avgiftsbelagda.
Vid Esbo musikinstitut (Espoon musiikkiopisto) kan barn och vuxna studera musik.
Läs mer: Andra studiemöjligheter
linkkiEsbo stad:
Arbetarinstitutetfinska _ svenska _ engelska
linkkiEsbo biIdkonstskola:
Bildkonst för barn och ungafinska _ svenska _ engelska
linkkiEsbo musikinstitut:
Musikundervisning för barn och vuxnafinska _ engelska
Dagvård
Förskoleundervisning
Grundläggande utbildning
Hemspråksundervisning för invandrare
Yrkesutbildning
Gymnasium
Stöd och handledning för unga
Högskoleutbildning
Andra studiemöjligheter
Dagvård
I Esbo finns både kommunala och privata daghem.
I Esbo finns dessutom familjedagvårdare.
Dagvård fås på finska och på svenska.
Ansök om dagvårdsplats minst fyra månader innan barnet ska börja i dagvården.
Om du till exempel oväntat får arbete eller en studieplats kan du ansöka om vårdplats senare.
När du ansöker om vårdplats ska du fylla i en ansökningsblankett.
Du kan också söka dagvårdsplats via Internet.
Familjer som bor i Esbo kan också söka dagvårdsplats till sitt barn i Helsingfors, Vanda eller Grankulla.
Du ska ändå lämna in din ansökan i Esbo.
Mer information får du via tjänsten Helsingforsregionen.fi.
Läs mer: Småbarnspedagogik
linkkiEsbo stad:
Dagvårdfinska _ svenska _ engelska
linkkiEsbo stad:
Ansökan om dagvårdsplatsfinska _ engelska
linkkiEsbo stad:
Servicepunktfinska _ svenska _ engelska
linkkiEsbo stad:
Dagvårdens samanvändningsområdefinska _ svenska _ engelska
Förskoleundervisning
I Esbo anordnas förskoleundervisningen (esiopetus) i daghemmen.
Förskoleundervisning ges på finska och på svenska.
Till förskoleundervisningen anmäler man sig via Esbo stads webbplats.
Förskoleundervisningen börjar i augusti.
Ansökningstiden är vanligtvis i januari.
I frågor kring barndagvård och förskoleundervisning kan du också kontakta daghemsföreståndarna eller stadens chef för småbarnsfostran (varhaiskasvatuspäällikkö).
Kontaktuppgifterna finns på stadens webbplats.
Läs mer: Förskoleundervisning.
linkkiEsbo stad:
Förskoleundervisningfinska _ svenska _ engelska
linkkiEsbo stad:
Ansökan till förskoleundervisningfinska _ engelska
Grundläggande utbildning
I Esbo finns finskspråkiga och svenskspråkiga grundskolor (peruskoulu).
Undervisning kan även fås på engelska.
Skolan börjar vanligtvis det året då barnet fyller sju år.
Anmälan till grundskolan ska göras på förhand.
Anmälningstiden är vanligtvis i januari.
På stadens webbplats hittar du kontaktuppgifterna till skolorna och mer information om anmälan.
Om du har frågor om den grundläggande utbildningen kan du kontakta Resultatenheten för den finskspråkiga undervisningen (Suomenkielisen opetuksen tulosyksikkö).
Resultatenheten för den finskspråkiga undervisningen
Kamrersvägen 3 B
Tfn (09) 816 52044 och (09) 816 52043
Grundläggande utbildning.
linkkiEsbo stad:
Grundläggande utbildningfinska _ svenska _ engelska
linkkiEsbo stad:
Anmälan till skolanfinska _ svenska _ engelska
linkkiEsbo stad:
Espoo International Schoolfinska _ engelska
Internationella skolor i huvudstadsregionenfinska
linkkiExpatFinland.fi:
Internationella skolor i huvudstadsregionenengelska
linkkiEsbo stad:
Eftermiddagsverksamhetfinska _ engelska
Hemspråksundervisning för invandrare
Barn med invandrarbakgrund och barn från tvåspråkiga familjer kan få hemspråksundervisning (oman äidinkielen opetus) om tillräckligt många barn anmäler sig till gruppen för det egna språket.
Undervisning ges två timmar i veckan.
Anmälan till hemspråksundervisning görs varje år i mars.
Mer information hittar du på Esbo stads webbplats.
linkkiEsbo stad:
Förberedande undervisning för barn i förskoleåldern(pdf, 100 kb)finska _ engelska _ ryska _ estniska _ somaliska _ kinesiska _ arabiska _ kurdiska _ albanska
linkkiEsbo stad:
Förberedande undervisning för barn i förskoleåldernfinska _ engelska
linkkiEsbo stad:
Hemspråksundervisningfinska _ engelska
Yrkesutbildning
På Omnia kan man studera många olika yrken.
På Omnia ordnas för invandrare utbildning som förbereder dem på yrkesutbildning.
Den förberedande utbildningen är avsedd för unga och vuxna, som är intresserade av yrkesstudier och vill förbättra sina kunskaper i finska..
Esbobor kan också ansöka till yrkesskolorna i Helsingfors och Vanda.
Läs mer: Yrkesutbildning
Yrkesutbildningfinska _ engelska
linkkiEsbo stad:
Yrkesläroanstalterfinska _ engelska
Yrkesläroanstalterfinska _ svenska _ engelska
linkkiVanda stad:
Yrkesutbildningfinska _ svenska
Gymnasium
I Esbo finns elva finskspråkiga och ett svenskspråkigt gymnasium (lukio).
I två av gymnasierna i Esbo finns en engelskspråkig IB-linje.
Ungdomar från Esbo kan också söka till gymnasier i andra städer.
I Esbo finns ett vuxengymnasium (aikuislukio) där vuxna kan avlägga gymnasie- och studentexamen.
På gymnasiet kan man även höja vitsorden i sitt avgångsbetyg eller studera enskilda ämnen.
Invandrarungdomar kan dessutom studera finska och avlägga grundskolans lärokurs.
I gymnasiet Leppävaaran lukio ordnas för invandrare och utlänningar utbildning som förbereder dem på gymnasiet.
Utbildningen är avsedd för unga som vill studera på gymnasiet, men vars språkkunskaper inte är tillräckliga för gymnasiestudier.
Läs mer: Gymnasium
linkkiEsbo stad:
Gymnasierfinska _ svenska _ engelska
linkkiEsbo stad:
Vuxengymnasietfinska
linkkiEsbo stad:
Gymnasieförberedande utbildning för invandrarefinska _ engelska
linkkiEsbo vuxengymnasium Omnia:
Grundläggande utbildning för invandrarefinska
Om du är under 30 år gammal kan du få råd och handledning via Ohjaamo-tjänsten.
Ohjaamos personal hjälper dig om du inte har ett arbete eller en studieplats.
Du kan även fråga om andra saker, som till exempel boende eller ekonomiska frågor.
Kontaktuppgifter:
Fågelbergavägen 2 A
Puh. 040 126 7513
linkkiEsbo stad:
Ohjaamofinska _ svenska _ engelska
Högskoleutbildning
I Esbo finns tre högskolor:
yrkeshögskolan Laurea
yrkeshögskolan Metropolia.
Vid högskolorna kan du avlägga högskoleexamen.
Mer information finns på Aalto-universitetets, Laureas och Metropolias webbplatser.
Också i Helsingfors finns det universitet och yrkeshögskolor där man kan studera inom många områden.
Mer information hittar du på Helsingfors stads webbplats.
Läs mer: Yrkeshögskolor
Universitet inom teknik, konst och ekonomifinska _ svenska _ engelska
Yrkeshögskolafinska _ engelska
linkkiMetropolia:
Yrkeshögskolafinska _ engelska
Högskolorfinska
Andra studiemöjligheter
Vid Esbo arbetarinstitut (Espoon työväenopisto) kan du studera till exempel språk, handarbete och matlagning eller delta i ledd motion.
Kurserna är avgiftsbelagda. Kurser anordnas både dagtid och kvällstid.
Vid arbetarinstitutet kan vem som helst studera.
Vid Esbo bildkonstskola (Espoon kuvataidekoulu) kan barn och unga studera bildkonst.
Studierna är avgiftsbelagda.
Vid Esbo musikinstitut (Espoon musiikkiopisto) kan barn och vuxna studera musik.
Läs mer: Studier som hobby
linkkiEsbo stad:
Arbetarinstitutetfinska _ svenska _ engelska
linkkiEsbo biIdkonstskola:
Bildkonst för barn och ungafinska _ svenska _ engelska
linkkiEsbo musikinstitut:
Musikundervisning för barn och vuxnafinska _ engelska
Hyresbostad
Ägarbostad
Bostadsrättsbostad
Delägarbostad
Tillfälligt boende
Boende i en krissituation
Stöd- och serviceboende
Bostadslöshet
Avfallshantering och återvinning
Hyresbostad
I Esbo och huvudstadsregionen är hyrorna ofta högre än i resten av Finland.
Det kan vara svårt att hitta en bostad med lämplig hyra.
Det lönar sig att avsätta tid för bostadssökandet och undersöka olika alternativ.
Privata hyresbostäder
Hos en privat hyresvärd kan det gå snabbt att få en bostad, men hyran kan vara högre än i stadens hyresbostäder.
Du kan söka privata hyresbostäder i Esbo via hyresvärdarnas webbplatser:
Sökning av hyresbostäderfinska
Sökning av hyresbostäderfinska _ engelska
Hyresbostäder för ungafinska _ engelska
Hyresbostäder för ungafinska _ engelska
Om du är studerande kan du få en hyresbostad för studerande i Esbo.
Hyresbostäder för studerande erbjuds av Helsingforsregionens studentbostadsstiftelse HOAS och Aalto-universitets studentkår AUS.
linkkiHOAS:
Hyresbostäder för studerandefinska _ svenska _ engelska
Hyresbostäder för studerandefinska _ svenska _ engelska
Stadens hyresbostäder
Stadens hyresbostäder är ofta billigare än bostäder som man hyr av företag eller privatpersoner.
Det är dock många som ansöker om stadens bostäder och endast en liten del av de sökande får en bostad.
Störst är bristen på små bostäder.
Stadens hyresbostäder förvaltas av Espoon Asunnot Oy (Espoon Asunnot Oy).
Om du vill ansöka om en hyresbostad, fyll i en ansökningsblankett för hyresbostad på Espoon Asunnot Oy:s webbplats.
Du kan även fylla i ansökningsblanketten på Espoon Asunnot Oy:s kontor.
Du kan också få blanketten hemskickad per post.
Dina möjligheter att få en bostad påverkas av ditt bostadsbehov och dina tillgångar och inkomster.
För att kunna ansöka om en hyresbostad hos staden, måste du ha uppehållstillstånd för minst ett år.
Tfn (09) 816 5800
Ansökan är giltig i tre månader.
Efter det måste du förnya din ansökan om du fortfarande letar efter bostad.
Läs mer: Hyresbostad
linkkiEsbo Bostäder Ab:
Ansökan om hyresbostad i stadenfinska _ engelska
linkkiEsbo stad:
Stadens hyresbostäderfinska _ svenska _ engelska
linkkiEsbo stad:
Seniorbostäderfinska _ svenska
Ägarbostad
På internet finns många bostadsförsäljningsannonser. Bostäderna i Esbo är tämligen dyra.
Information om köp av bostad hittar du på InfoFinlands sida Ägarbostad.
Bostadsrättsbostad
Om du ansöker om en bostadsrättsbostad, behöver du ett ordningsnummer. Du ansöker om ordningsnumret vid Esbo eller Helsingfors stad.
Läs mer: Bostadsrättsbostad.
linkkiEsbo stad:
Bostadsrättsbostäderfinska _ svenska _ engelska
Delägarbostad
Asuntosäätiö har delägarbostäder i Esbo.
Mer information hittar du på Asuntosäätiös webbplats.
Läs mer: Delägarbostad.
Delägarbostadfinska
Tillfälligt boende
I Esbo finns många olika hotell där man kan bo tillfälligt.
Läs mer: Tillfälligt boende.
linkkiVisitEspoo.fi:
Hotellfinska _ svenska _ engelska _ ryska _ kinesiska
Brand eller vattenskada
Om din bostad har skadats till exempel till följd av brand eller vattenskada kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
Kontakta ditt försäkringsbolag direkt när skadan har inträffat.
Våld i hemmet
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta tjänsten Omatila (Omatila).
Omatila ordnar vid behov boende för dig och dina barn.
Omatila-tjänsten
Kamrersvägen 6 A
Tfn 043 825 0535
Öppet
Lördag-söndag kl. 9-16
Social- och krisjouren 24 h
Tfn 09 816 42439
linkkiEsbo stad:
Hjälp till offer för familjevåldfinska _ svenska _ engelska
Om du är ung och har problem hemma, kan du kontakta Finlands Röda Kors De ungas skyddshus.
Skyddshuset finns i Alberga.
De ungas skyddshus
Tfn (09) 8195 5360
linkkiFinlands Röda Kors:
De ungas skyddshusfinska _ svenska _ engelska
Stöd- och serviceboende
En del människor, till exempel åldringar och handikappade, har svårt att klara av de dagliga sysslorna utan hjälp.
Personer som har sin hemkommun i Esbo kan få hemvårdens stödtjänster av Esbo stad, till exempel måltidstjänster eller färdtjänst.
Dessa tjänster hjälper människorna att klara sig bättre hemma.
Åldringar och handikappade som inte klarar av att bo självständigt, kan bo i ett servicehus eller på en vårdinrättning.
Läs mer: Stöd- och serviceboende
Om du har frågor kring stödtjänsterna för handikappade, kontakta handikappservicen vid Esbo stad.
Esbo stads handikappservice
Telefonrådgivning: (09) 816 45285
linkkiEsbo stad:
Stödtjänster för handikappadefinska _ svenska _ engelska
Om du har frågor kring stödtjänsterna för äldre, kontakta Esbo stads rådgivning för seniorer.
Esbo stads rådgivning för seniorer
tfn (09) 816 33333
linkkiEsbo stad:
Stödtjänster för äldrefinska _ svenska _ engelska
linkkiEsbo stad:
Information om hemvårdens stödtjänsterfinska _ svenska
linkkiEsbo stad:
Information om boende i servicehusfinska _ svenska
Bostadslöshet
Om du blir bostadslös, kontakta Esbo stads verksamhetsställe för vuxensocialarbete.
linkkiEsbo stad:
Kontaktuppgifter till vuxensocialarbetetfinska _ svenska _ engelska
Om läget är akut, kan du även kontakta social- och krisjouren i Esbo.
Social- och krisjouren
Jorvs sjukhus
Åbovägen 150
Tfn (09) 816 42439
linkkiEsbo stad:
Social- och krisjourenfinska _ svenska _ engelska
Läs mer: Bostadslöshet
Avfallshantering och återvinning
